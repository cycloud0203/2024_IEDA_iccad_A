// Benchmark "top_809568696_809776567_809698999_863110837_1234615" written by ABC on Fri Jun 14 22:42:45 2024

module top_809568696_809776567_809698999_863110837_1234615 ( 
    n74, n203, n271, n394, n411, n427, n462, n498, n650, n656, n666, n674,
    n702, n730, n737, n760, n844, n977, n1027, n1093, n1222, n1265, n1268,
    n1347, n1568, n1637, n1702, n1763, n1776, n2048, n2061, n2164, n2166,
    n2201, n2334, n2454, n2573, n2615, n2674, n2699, n2895, n3130, n3166,
    n3263, n3367, n3388, n3506, n3532, n3652, n3655, n3673, n3775, n3799,
    n3804, n3833, n3893, n3910, n3972, n4000, n4022, n4039, n4117, n4131,
    n4147, n4154, n4172, n4175, n4225, n4282, n4292, n4615, n4659, n4755,
    n4774, n4785, n4895, n4907, n5009, n5014, n5023, n5033, n5046, n5077,
    n5184, n5185, n5225, n5430, n5449, n5467, n5502, n5601, n5725, n5786,
    n5943, n5950, n5960, n6007, n6054, n6114, n6147, n6251, n6258, n6270,
    n6362, n6436, n6460, n6480, n6517, n6555, n6586, n6680, n6693, n6703,
    n6758, n6791, n6810, n6873, n6946, n6999, n7104, n7272, n7282, n7354,
    n7450, n7652, n7667, n7748, n7832, n7941, n7972, n7988, n8002, n8044,
    n8073, n8204, n8262, n8302, n8315, n8397, n8439, n8463, n8486, n8550,
    n8552, n8598, n8635, n8649, n8737, n8746, n8780, n8799, n8800, n8873,
    n8892, n8926, n8997, n9026, n9110, n9154, n9186, n9252, n9314, n9543,
    n9544, n9555, n9589, n9830, n9893, n9921, n9936, n9977, n10050, n10051,
    n10061, n10080, n10112, n10147, n10255, n10278, n10283, n10378, n10407,
    n10426, n10446, n10466, n10470, n10573, n10615, n10630, n10736, n10750,
    n10765, n10862, n10912, n10945, n11143, n11158, n11269, n11345, n11404,
    n11529, n11590, n11605, n11666, n11756, n11776, n11842, n11854, n11875,
    n11902, n11930, n11933, n11961, n12009, n12012, n12025, n12142, n12218,
    n12270, n12321, n12336, n12573, n12614, n12782, n12829, n12885, n12927,
    n12976, n13000, n13093, n13102, n13109, n13186, n13224, n13231, n13295,
    n13363, n13364, n13509, n13511, n13561, n13625, n13636, n13814, n13882,
    n13890, n13944, n13992, n14072, n14163, n14293, n14303, n14408, n14464,
    n14475, n14483,
    n8, n46, n91, n126, n278, n389, n451, n490, n543, n682, n884, n948,
    n1094, n1122, n1124, n1329, n1545, n1739, n1827, n1900, n1927, n1951,
    n2027, n2126, n2175, n2223, n2311, n2407, n2556, n2559, n2572, n2672,
    n2734, n3090, n3242, n3340, n3603, n3854, n3901, n4125, n4279, n4305,
    n4345, n4437, n4541, n4604, n4672, n4858, n4971, n5479, n5550, n5586,
    n5806, n5851, n5987, n6012, n6198, n6275, n6314, n6682, n6696, n6786,
    n6853, n6952, n6979, n7071, n7073, n7132, n7152, n7246, n7265, n7382,
    n7655, n7771, n7825, n8068, n8085, n8124, n8144, n8215, n8306, n8471,
    n8604, n8909, n9096, n9342, n9437, n9447, n9570, n9665, n9717, n10515,
    n10591, n10791, n10802, n10915, n11122, n11393, n11463, n11534, n11627,
    n11664, n11822, n11847, n12032, n12166, n12232, n12355, n12535, n12989,
    n13010, n13045, n13114, n13141, n13316, n13577, n13639, n13658, n13693,
    n13760, n13853, n13870, n13953, n13959, n14289, n14307, n14330, n14399,
    n14463  );
  input  n74, n203, n271, n394, n411, n427, n462, n498, n650, n656, n666,
    n674, n702, n730, n737, n760, n844, n977, n1027, n1093, n1222, n1265,
    n1268, n1347, n1568, n1637, n1702, n1763, n1776, n2048, n2061, n2164,
    n2166, n2201, n2334, n2454, n2573, n2615, n2674, n2699, n2895, n3130,
    n3166, n3263, n3367, n3388, n3506, n3532, n3652, n3655, n3673, n3775,
    n3799, n3804, n3833, n3893, n3910, n3972, n4000, n4022, n4039, n4117,
    n4131, n4147, n4154, n4172, n4175, n4225, n4282, n4292, n4615, n4659,
    n4755, n4774, n4785, n4895, n4907, n5009, n5014, n5023, n5033, n5046,
    n5077, n5184, n5185, n5225, n5430, n5449, n5467, n5502, n5601, n5725,
    n5786, n5943, n5950, n5960, n6007, n6054, n6114, n6147, n6251, n6258,
    n6270, n6362, n6436, n6460, n6480, n6517, n6555, n6586, n6680, n6693,
    n6703, n6758, n6791, n6810, n6873, n6946, n6999, n7104, n7272, n7282,
    n7354, n7450, n7652, n7667, n7748, n7832, n7941, n7972, n7988, n8002,
    n8044, n8073, n8204, n8262, n8302, n8315, n8397, n8439, n8463, n8486,
    n8550, n8552, n8598, n8635, n8649, n8737, n8746, n8780, n8799, n8800,
    n8873, n8892, n8926, n8997, n9026, n9110, n9154, n9186, n9252, n9314,
    n9543, n9544, n9555, n9589, n9830, n9893, n9921, n9936, n9977, n10050,
    n10051, n10061, n10080, n10112, n10147, n10255, n10278, n10283, n10378,
    n10407, n10426, n10446, n10466, n10470, n10573, n10615, n10630, n10736,
    n10750, n10765, n10862, n10912, n10945, n11143, n11158, n11269, n11345,
    n11404, n11529, n11590, n11605, n11666, n11756, n11776, n11842, n11854,
    n11875, n11902, n11930, n11933, n11961, n12009, n12012, n12025, n12142,
    n12218, n12270, n12321, n12336, n12573, n12614, n12782, n12829, n12885,
    n12927, n12976, n13000, n13093, n13102, n13109, n13186, n13224, n13231,
    n13295, n13363, n13364, n13509, n13511, n13561, n13625, n13636, n13814,
    n13882, n13890, n13944, n13992, n14072, n14163, n14293, n14303, n14408,
    n14464, n14475, n14483;
  output n8, n46, n91, n126, n278, n389, n451, n490, n543, n682, n884, n948,
    n1094, n1122, n1124, n1329, n1545, n1739, n1827, n1900, n1927, n1951,
    n2027, n2126, n2175, n2223, n2311, n2407, n2556, n2559, n2572, n2672,
    n2734, n3090, n3242, n3340, n3603, n3854, n3901, n4125, n4279, n4305,
    n4345, n4437, n4541, n4604, n4672, n4858, n4971, n5479, n5550, n5586,
    n5806, n5851, n5987, n6012, n6198, n6275, n6314, n6682, n6696, n6786,
    n6853, n6952, n6979, n7071, n7073, n7132, n7152, n7246, n7265, n7382,
    n7655, n7771, n7825, n8068, n8085, n8124, n8144, n8215, n8306, n8471,
    n8604, n8909, n9096, n9342, n9437, n9447, n9570, n9665, n9717, n10515,
    n10591, n10791, n10802, n10915, n11122, n11393, n11463, n11534, n11627,
    n11664, n11822, n11847, n12032, n12166, n12232, n12355, n12535, n12989,
    n13010, n13045, n13114, n13141, n13316, n13577, n13639, n13658, n13693,
    n13760, n13853, n13870, n13953, n13959, n14289, n14307, n14330, n14399,
    n14463;
  wire new_n386, new_n387, new_n388, new_n389_1, new_n390, new_n391,
    new_n392, new_n393, new_n394_1, new_n395, new_n396, new_n397, new_n398,
    new_n399, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411_1, new_n412,
    new_n413, new_n414, new_n415, new_n416, new_n417, new_n418, new_n419,
    new_n420, new_n421, new_n422, new_n423, new_n424, new_n425, new_n426,
    new_n427_1, new_n428, new_n429, new_n430, new_n431, new_n432, new_n433,
    new_n434, new_n435, new_n436, new_n437, new_n438, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n449, new_n450, new_n451_1, new_n452, new_n453, new_n454,
    new_n455, new_n456, new_n457, new_n458, new_n459, new_n460, new_n461,
    new_n462_1, new_n463, new_n464, new_n465, new_n466, new_n467, new_n468,
    new_n469, new_n470, new_n471, new_n472, new_n473, new_n474, new_n475,
    new_n476, new_n477, new_n478, new_n479, new_n480, new_n481, new_n482,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488, new_n489,
    new_n490_1, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498_1, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543_1, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650_1,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656_1, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666_1, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674_1, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682_1, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702_1, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730_1, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737_1, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760_1, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884_1, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948_1, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977_1, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027_1, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085,
    new_n1086, new_n1087, new_n1088, new_n1089, new_n1090, new_n1091,
    new_n1092, new_n1093_1, new_n1094_1, new_n1095, new_n1096, new_n1097,
    new_n1098, new_n1099, new_n1100, new_n1101, new_n1102, new_n1103,
    new_n1104, new_n1105, new_n1106, new_n1107, new_n1108, new_n1109,
    new_n1110, new_n1111, new_n1112, new_n1113, new_n1114, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122_1, new_n1123, new_n1124_1, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222_1, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265_1, new_n1266,
    new_n1267, new_n1268_1, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329_1, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347_1, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1502, new_n1503, new_n1504, new_n1505, new_n1506,
    new_n1507, new_n1508, new_n1509, new_n1510, new_n1511, new_n1512,
    new_n1513, new_n1514, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545_1, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564, new_n1565, new_n1566, new_n1567,
    new_n1568_1, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1626, new_n1627, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637_1, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644, new_n1645, new_n1646,
    new_n1647, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1669, new_n1670,
    new_n1671, new_n1672, new_n1673, new_n1674, new_n1675, new_n1676,
    new_n1677, new_n1678, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1690, new_n1691, new_n1692, new_n1693, new_n1694,
    new_n1695, new_n1696, new_n1697, new_n1698, new_n1699, new_n1700,
    new_n1701, new_n1702_1, new_n1703, new_n1704, new_n1705, new_n1706,
    new_n1707, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1713, new_n1714, new_n1715, new_n1716, new_n1717, new_n1718,
    new_n1719, new_n1720, new_n1721, new_n1722, new_n1723, new_n1724,
    new_n1725, new_n1726, new_n1727, new_n1728, new_n1729, new_n1730,
    new_n1731, new_n1732, new_n1733, new_n1734, new_n1735, new_n1736,
    new_n1737, new_n1738, new_n1739_1, new_n1740, new_n1741, new_n1742,
    new_n1743, new_n1744, new_n1745, new_n1746, new_n1747, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763_1, new_n1764, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1775, new_n1776_1, new_n1777, new_n1778,
    new_n1779, new_n1780, new_n1781, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1786, new_n1787, new_n1788, new_n1789, new_n1790,
    new_n1791, new_n1792, new_n1793, new_n1794, new_n1795, new_n1796,
    new_n1797, new_n1798, new_n1799, new_n1800, new_n1801, new_n1802,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1809, new_n1810, new_n1811, new_n1812, new_n1813, new_n1814,
    new_n1815, new_n1816, new_n1817, new_n1818, new_n1819, new_n1820,
    new_n1821, new_n1822, new_n1823, new_n1824, new_n1825, new_n1826,
    new_n1827_1, new_n1828, new_n1829, new_n1830, new_n1831, new_n1832,
    new_n1833, new_n1834, new_n1835, new_n1836, new_n1837, new_n1838,
    new_n1839, new_n1840, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1850,
    new_n1851, new_n1852, new_n1853, new_n1854, new_n1855, new_n1856,
    new_n1857, new_n1858, new_n1859, new_n1860, new_n1861, new_n1862,
    new_n1863, new_n1864, new_n1865, new_n1866, new_n1867, new_n1868,
    new_n1869, new_n1870, new_n1871, new_n1872, new_n1873, new_n1874,
    new_n1875, new_n1876, new_n1877, new_n1878, new_n1879, new_n1880,
    new_n1881, new_n1882, new_n1883, new_n1884, new_n1885, new_n1886,
    new_n1887, new_n1888, new_n1889, new_n1890, new_n1891, new_n1892,
    new_n1893, new_n1894, new_n1895, new_n1896, new_n1897, new_n1898,
    new_n1899, new_n1900_1, new_n1901, new_n1902, new_n1903, new_n1904,
    new_n1905, new_n1906, new_n1907, new_n1908, new_n1909, new_n1910,
    new_n1911, new_n1912, new_n1913, new_n1914, new_n1915, new_n1916,
    new_n1917, new_n1918, new_n1919, new_n1920, new_n1921, new_n1922,
    new_n1923, new_n1924, new_n1925, new_n1926, new_n1927_1, new_n1928,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1940, new_n1941,
    new_n1942, new_n1943, new_n1944, new_n1945, new_n1946, new_n1947,
    new_n1948, new_n1949, new_n1950, new_n1951_1, new_n1952, new_n1953,
    new_n1954, new_n1955, new_n1956, new_n1957, new_n1958, new_n1959,
    new_n1960, new_n1961, new_n1962, new_n1963, new_n1964, new_n1965,
    new_n1966, new_n1967, new_n1968, new_n1969, new_n1970, new_n1971,
    new_n1972, new_n1973, new_n1974, new_n1975, new_n1976, new_n1977,
    new_n1978, new_n1979, new_n1980, new_n1981, new_n1982, new_n1983,
    new_n1984, new_n1985, new_n1986, new_n1987, new_n1988, new_n1989,
    new_n1990, new_n1991, new_n1992, new_n1993, new_n1994, new_n1995,
    new_n1996, new_n1997, new_n1998, new_n1999, new_n2000, new_n2001,
    new_n2002, new_n2003, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2008, new_n2009, new_n2010, new_n2011, new_n2012, new_n2013,
    new_n2014, new_n2015, new_n2016, new_n2017, new_n2019, new_n2020,
    new_n2021, new_n2022, new_n2023, new_n2024, new_n2025, new_n2026,
    new_n2027_1, new_n2028, new_n2029, new_n2030, new_n2031, new_n2032,
    new_n2033, new_n2034, new_n2035, new_n2036, new_n2037, new_n2038,
    new_n2039, new_n2040, new_n2041, new_n2042, new_n2043, new_n2044,
    new_n2045, new_n2046, new_n2047, new_n2048_1, new_n2049, new_n2050,
    new_n2051, new_n2052, new_n2053, new_n2054, new_n2055, new_n2056,
    new_n2057, new_n2058, new_n2059, new_n2060, new_n2061_1, new_n2062,
    new_n2063, new_n2064, new_n2065, new_n2066, new_n2067, new_n2068,
    new_n2069, new_n2070, new_n2071, new_n2072, new_n2073, new_n2074,
    new_n2075, new_n2076, new_n2077, new_n2078, new_n2079, new_n2080,
    new_n2081, new_n2082, new_n2083, new_n2084, new_n2085, new_n2086,
    new_n2087, new_n2088, new_n2089, new_n2090, new_n2091, new_n2092,
    new_n2093, new_n2094, new_n2095, new_n2096, new_n2097, new_n2098,
    new_n2099, new_n2100, new_n2101, new_n2102, new_n2103, new_n2104,
    new_n2105, new_n2106, new_n2107, new_n2108, new_n2109, new_n2110,
    new_n2111, new_n2112, new_n2113, new_n2114, new_n2115, new_n2116,
    new_n2117, new_n2118, new_n2119, new_n2120, new_n2121, new_n2122,
    new_n2123, new_n2124, new_n2125, new_n2126_1, new_n2127, new_n2128,
    new_n2129, new_n2130, new_n2132, new_n2133, new_n2134, new_n2135,
    new_n2136, new_n2137, new_n2138, new_n2139, new_n2140, new_n2141,
    new_n2142, new_n2143, new_n2144, new_n2145, new_n2146, new_n2147,
    new_n2148, new_n2149, new_n2150, new_n2151, new_n2152, new_n2153,
    new_n2154, new_n2155, new_n2156, new_n2157, new_n2158, new_n2159,
    new_n2160, new_n2161, new_n2162, new_n2163, new_n2164_1, new_n2165,
    new_n2166_1, new_n2167, new_n2168, new_n2169, new_n2170, new_n2171,
    new_n2172, new_n2173, new_n2174, new_n2175_1, new_n2176, new_n2177,
    new_n2178, new_n2179, new_n2180, new_n2181, new_n2182, new_n2183,
    new_n2184, new_n2185, new_n2186, new_n2187, new_n2188, new_n2189,
    new_n2190, new_n2191, new_n2192, new_n2193, new_n2194, new_n2195,
    new_n2196, new_n2197, new_n2198, new_n2199, new_n2200, new_n2201_1,
    new_n2202, new_n2203, new_n2204, new_n2205, new_n2206, new_n2207,
    new_n2208, new_n2209, new_n2210, new_n2211, new_n2212, new_n2213,
    new_n2214, new_n2215, new_n2216, new_n2217, new_n2218, new_n2219,
    new_n2220, new_n2221, new_n2222, new_n2223_1, new_n2224, new_n2225,
    new_n2226, new_n2227, new_n2228, new_n2229, new_n2230, new_n2231,
    new_n2232, new_n2233, new_n2234, new_n2235, new_n2236, new_n2237,
    new_n2238, new_n2239, new_n2240, new_n2241, new_n2242, new_n2243,
    new_n2244, new_n2245, new_n2246, new_n2247, new_n2248, new_n2249,
    new_n2250, new_n2251, new_n2252, new_n2253, new_n2254, new_n2255,
    new_n2256, new_n2257, new_n2258, new_n2259, new_n2260, new_n2261,
    new_n2262, new_n2263, new_n2264, new_n2265, new_n2266, new_n2267,
    new_n2268, new_n2269, new_n2270, new_n2271, new_n2272, new_n2273,
    new_n2274, new_n2275, new_n2276, new_n2277, new_n2278, new_n2279,
    new_n2280, new_n2281, new_n2283, new_n2284, new_n2285, new_n2286,
    new_n2287, new_n2288, new_n2289, new_n2290, new_n2291, new_n2292,
    new_n2293, new_n2294, new_n2295, new_n2296, new_n2297, new_n2298,
    new_n2299, new_n2300, new_n2301, new_n2302, new_n2303, new_n2304,
    new_n2305, new_n2306, new_n2307, new_n2308, new_n2309, new_n2310,
    new_n2311_1, new_n2312, new_n2313, new_n2314, new_n2315, new_n2316,
    new_n2317, new_n2318, new_n2319, new_n2320, new_n2321, new_n2322,
    new_n2323, new_n2324, new_n2325, new_n2326, new_n2327, new_n2328,
    new_n2329, new_n2330, new_n2331, new_n2332, new_n2333, new_n2334_1,
    new_n2335, new_n2336, new_n2337, new_n2338, new_n2339, new_n2340,
    new_n2341, new_n2342, new_n2343, new_n2344, new_n2345, new_n2346,
    new_n2347, new_n2348, new_n2349, new_n2350, new_n2351, new_n2352,
    new_n2353, new_n2354, new_n2355, new_n2356, new_n2357, new_n2358,
    new_n2359, new_n2360, new_n2361, new_n2362, new_n2363, new_n2364,
    new_n2365, new_n2366, new_n2367, new_n2368, new_n2369, new_n2370,
    new_n2371, new_n2372, new_n2373, new_n2374, new_n2375, new_n2376,
    new_n2377, new_n2378, new_n2379, new_n2380, new_n2381, new_n2382,
    new_n2383, new_n2384, new_n2385, new_n2386, new_n2387, new_n2388,
    new_n2389, new_n2390, new_n2391, new_n2392, new_n2393, new_n2395,
    new_n2396, new_n2397, new_n2398, new_n2399, new_n2400, new_n2401,
    new_n2402, new_n2403, new_n2404, new_n2405, new_n2406, new_n2407_1,
    new_n2408, new_n2409, new_n2410, new_n2411, new_n2412, new_n2413,
    new_n2414, new_n2415, new_n2416, new_n2417, new_n2418, new_n2419,
    new_n2420, new_n2421, new_n2422, new_n2423, new_n2424, new_n2425,
    new_n2426, new_n2427, new_n2428, new_n2429, new_n2430, new_n2431,
    new_n2432, new_n2433, new_n2434, new_n2435, new_n2436, new_n2437,
    new_n2438, new_n2439, new_n2440, new_n2441, new_n2442, new_n2443,
    new_n2444, new_n2445, new_n2446, new_n2447, new_n2448, new_n2449,
    new_n2450, new_n2451, new_n2452, new_n2453, new_n2454_1, new_n2455,
    new_n2456, new_n2457, new_n2458, new_n2459, new_n2460, new_n2461,
    new_n2462, new_n2463, new_n2464, new_n2465, new_n2466, new_n2467,
    new_n2468, new_n2469, new_n2470, new_n2471, new_n2472, new_n2473,
    new_n2474, new_n2475, new_n2476, new_n2477, new_n2478, new_n2479,
    new_n2480, new_n2481, new_n2482, new_n2483, new_n2484, new_n2485,
    new_n2486, new_n2487, new_n2488, new_n2489, new_n2490, new_n2491,
    new_n2492, new_n2493, new_n2494, new_n2495, new_n2496, new_n2497,
    new_n2498, new_n2499, new_n2500, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513, new_n2514, new_n2515, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556_1, new_n2557, new_n2558,
    new_n2559_1, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572_1, new_n2573_1, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578, new_n2579, new_n2580, new_n2581, new_n2582,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2609, new_n2610, new_n2611, new_n2612, new_n2613,
    new_n2614, new_n2615_1, new_n2616, new_n2617, new_n2618, new_n2619,
    new_n2620, new_n2621, new_n2622, new_n2623, new_n2624, new_n2625,
    new_n2626, new_n2627, new_n2628, new_n2629, new_n2630, new_n2631,
    new_n2632, new_n2633, new_n2634, new_n2635, new_n2636, new_n2637,
    new_n2638, new_n2639, new_n2640, new_n2641, new_n2642, new_n2643,
    new_n2644, new_n2645, new_n2646, new_n2647, new_n2648, new_n2649,
    new_n2650, new_n2651, new_n2652, new_n2653, new_n2654, new_n2655,
    new_n2656, new_n2657, new_n2658, new_n2659, new_n2660, new_n2661,
    new_n2662, new_n2663, new_n2664, new_n2665, new_n2666, new_n2667,
    new_n2668, new_n2669, new_n2670, new_n2671, new_n2672_1, new_n2673,
    new_n2674_1, new_n2675, new_n2676, new_n2677, new_n2678, new_n2679,
    new_n2680, new_n2681, new_n2682, new_n2683, new_n2684, new_n2685,
    new_n2686, new_n2687, new_n2688, new_n2689, new_n2690, new_n2691,
    new_n2692, new_n2693, new_n2694, new_n2695, new_n2696, new_n2697,
    new_n2698, new_n2700, new_n2701, new_n2702, new_n2703, new_n2704,
    new_n2705, new_n2706, new_n2707, new_n2708, new_n2709, new_n2710,
    new_n2711, new_n2712, new_n2713, new_n2714, new_n2715, new_n2716,
    new_n2717, new_n2718, new_n2719, new_n2720, new_n2721, new_n2722,
    new_n2723, new_n2724, new_n2725, new_n2726, new_n2727, new_n2728,
    new_n2729, new_n2730, new_n2731, new_n2732, new_n2733, new_n2734_1,
    new_n2735, new_n2736, new_n2737, new_n2738, new_n2739, new_n2740,
    new_n2741, new_n2742, new_n2743, new_n2744, new_n2745, new_n2746,
    new_n2747, new_n2748, new_n2749, new_n2750, new_n2751, new_n2752,
    new_n2753, new_n2754, new_n2755, new_n2756, new_n2757, new_n2758,
    new_n2759, new_n2760, new_n2761, new_n2762, new_n2763, new_n2764,
    new_n2765, new_n2766, new_n2767, new_n2768, new_n2769, new_n2770,
    new_n2771, new_n2772, new_n2773, new_n2774, new_n2775, new_n2776,
    new_n2777, new_n2778, new_n2779, new_n2780, new_n2781, new_n2782,
    new_n2783, new_n2784, new_n2785, new_n2786, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858, new_n2859, new_n2860, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886,
    new_n2887, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895_1, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944, new_n2945, new_n2946,
    new_n2947, new_n2948, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2972, new_n2973, new_n2974, new_n2975, new_n2976, new_n2977,
    new_n2978, new_n2979, new_n2980, new_n2981, new_n2982, new_n2983,
    new_n2984, new_n2985, new_n2986, new_n2987, new_n2988, new_n2989,
    new_n2990, new_n2991, new_n2992, new_n2993, new_n2994, new_n2995,
    new_n2996, new_n2997, new_n2998, new_n2999, new_n3000, new_n3001,
    new_n3002, new_n3003, new_n3004, new_n3005, new_n3006, new_n3007,
    new_n3008, new_n3009, new_n3010, new_n3011, new_n3012, new_n3013,
    new_n3014, new_n3015, new_n3016, new_n3017, new_n3018, new_n3019,
    new_n3020, new_n3021, new_n3022, new_n3023, new_n3024, new_n3025,
    new_n3026, new_n3027, new_n3028, new_n3029, new_n3030, new_n3031,
    new_n3032, new_n3033, new_n3034, new_n3035, new_n3036, new_n3037,
    new_n3038, new_n3039, new_n3040, new_n3041, new_n3042, new_n3043,
    new_n3044, new_n3045, new_n3046, new_n3047, new_n3048, new_n3049,
    new_n3050, new_n3051, new_n3052, new_n3053, new_n3054, new_n3055,
    new_n3056, new_n3057, new_n3058, new_n3059, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090_1, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130_1, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166_1, new_n3167, new_n3168, new_n3169, new_n3171,
    new_n3172, new_n3173, new_n3174, new_n3175, new_n3176, new_n3177,
    new_n3178, new_n3179, new_n3180, new_n3181, new_n3182, new_n3183,
    new_n3184, new_n3185, new_n3186, new_n3187, new_n3188, new_n3189,
    new_n3190, new_n3191, new_n3192, new_n3193, new_n3194, new_n3195,
    new_n3196, new_n3197, new_n3198, new_n3199, new_n3200, new_n3201,
    new_n3202, new_n3203, new_n3204, new_n3205, new_n3206, new_n3207,
    new_n3208, new_n3209, new_n3210, new_n3211, new_n3212, new_n3213,
    new_n3214, new_n3215, new_n3216, new_n3217, new_n3218, new_n3219,
    new_n3220, new_n3221, new_n3222, new_n3223, new_n3224, new_n3225,
    new_n3226, new_n3227, new_n3228, new_n3229, new_n3230, new_n3231,
    new_n3232, new_n3233, new_n3234, new_n3235, new_n3236, new_n3237,
    new_n3238, new_n3239, new_n3240, new_n3241, new_n3242_1, new_n3243,
    new_n3244, new_n3245, new_n3246, new_n3247, new_n3248, new_n3249,
    new_n3250, new_n3251, new_n3252, new_n3253, new_n3254, new_n3255,
    new_n3256, new_n3257, new_n3258, new_n3260, new_n3261, new_n3262,
    new_n3263_1, new_n3264, new_n3265, new_n3266, new_n3267, new_n3268,
    new_n3269, new_n3270, new_n3271, new_n3272, new_n3273, new_n3274,
    new_n3275, new_n3276, new_n3277, new_n3278, new_n3279, new_n3280,
    new_n3281, new_n3282, new_n3283, new_n3284, new_n3285, new_n3286,
    new_n3287, new_n3288, new_n3289, new_n3290, new_n3291, new_n3292,
    new_n3293, new_n3294, new_n3295, new_n3296, new_n3297, new_n3298,
    new_n3299, new_n3300, new_n3301, new_n3302, new_n3303, new_n3304,
    new_n3305, new_n3306, new_n3307, new_n3308, new_n3309, new_n3310,
    new_n3311, new_n3312, new_n3313, new_n3314, new_n3315, new_n3316,
    new_n3317, new_n3318, new_n3319, new_n3320, new_n3321, new_n3322,
    new_n3323, new_n3324, new_n3325, new_n3326, new_n3327, new_n3328,
    new_n3329, new_n3330, new_n3331, new_n3332, new_n3333, new_n3334,
    new_n3335, new_n3336, new_n3337, new_n3338, new_n3339, new_n3340_1,
    new_n3341, new_n3342, new_n3343, new_n3344, new_n3345, new_n3346,
    new_n3348, new_n3349, new_n3350, new_n3351, new_n3352, new_n3353,
    new_n3354, new_n3355, new_n3356, new_n3357, new_n3358, new_n3359,
    new_n3360, new_n3361, new_n3362, new_n3363, new_n3364, new_n3365,
    new_n3366, new_n3367_1, new_n3368, new_n3369, new_n3370, new_n3371,
    new_n3372, new_n3373, new_n3374, new_n3375, new_n3376, new_n3377,
    new_n3378, new_n3379, new_n3380, new_n3381, new_n3382, new_n3383,
    new_n3384, new_n3385, new_n3386, new_n3387, new_n3388_1, new_n3389,
    new_n3390, new_n3391, new_n3392, new_n3393, new_n3394, new_n3395,
    new_n3396, new_n3397, new_n3398, new_n3399, new_n3400, new_n3401,
    new_n3402, new_n3403, new_n3404, new_n3405, new_n3406, new_n3407,
    new_n3408, new_n3409, new_n3410, new_n3411, new_n3412, new_n3413,
    new_n3414, new_n3415, new_n3416, new_n3417, new_n3418, new_n3419,
    new_n3420, new_n3421, new_n3422, new_n3423, new_n3424, new_n3425,
    new_n3426, new_n3427, new_n3428, new_n3429, new_n3430, new_n3431,
    new_n3432, new_n3433, new_n3434, new_n3435, new_n3436, new_n3437,
    new_n3438, new_n3439, new_n3440, new_n3441, new_n3443, new_n3444,
    new_n3445, new_n3446, new_n3447, new_n3448, new_n3449, new_n3450,
    new_n3451, new_n3452, new_n3453, new_n3454, new_n3455, new_n3456,
    new_n3457, new_n3458, new_n3459, new_n3460, new_n3461, new_n3462,
    new_n3463, new_n3464, new_n3465, new_n3466, new_n3467, new_n3468,
    new_n3469, new_n3470, new_n3471, new_n3472, new_n3473, new_n3474,
    new_n3475, new_n3476, new_n3477, new_n3478, new_n3479, new_n3480,
    new_n3481, new_n3482, new_n3483, new_n3484, new_n3485, new_n3486,
    new_n3487, new_n3488, new_n3489, new_n3490, new_n3491, new_n3492,
    new_n3493, new_n3494, new_n3495, new_n3496, new_n3497, new_n3498,
    new_n3499, new_n3500, new_n3501, new_n3502, new_n3503, new_n3504,
    new_n3505, new_n3506_1, new_n3507, new_n3508, new_n3509, new_n3510,
    new_n3511, new_n3512, new_n3513, new_n3514, new_n3515, new_n3516,
    new_n3517, new_n3518, new_n3519, new_n3520, new_n3521, new_n3522,
    new_n3523, new_n3524, new_n3525, new_n3526, new_n3527, new_n3528,
    new_n3529, new_n3530, new_n3531, new_n3533, new_n3534, new_n3535,
    new_n3536, new_n3537, new_n3538, new_n3539, new_n3540, new_n3541,
    new_n3542, new_n3543, new_n3544, new_n3545, new_n3546, new_n3547,
    new_n3548, new_n3549, new_n3550, new_n3551, new_n3552, new_n3553,
    new_n3554, new_n3555, new_n3556, new_n3557, new_n3558, new_n3559,
    new_n3560, new_n3561, new_n3562, new_n3563, new_n3564, new_n3565,
    new_n3566, new_n3567, new_n3568, new_n3569, new_n3570, new_n3571,
    new_n3572, new_n3573, new_n3574, new_n3575, new_n3576, new_n3577,
    new_n3578, new_n3579, new_n3580, new_n3581, new_n3582, new_n3583,
    new_n3584, new_n3585, new_n3586, new_n3587, new_n3588, new_n3589,
    new_n3590, new_n3591, new_n3592, new_n3593, new_n3594, new_n3595,
    new_n3596, new_n3597, new_n3598, new_n3599, new_n3600, new_n3601,
    new_n3602, new_n3603_1, new_n3604, new_n3605, new_n3606, new_n3607,
    new_n3608, new_n3609, new_n3610, new_n3611, new_n3612, new_n3613,
    new_n3614, new_n3615, new_n3616, new_n3617, new_n3618, new_n3619,
    new_n3620, new_n3621, new_n3622, new_n3623, new_n3624, new_n3625,
    new_n3626, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649, new_n3650,
    new_n3651, new_n3652_1, new_n3653, new_n3654, new_n3655_1, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673_1, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3716, new_n3717,
    new_n3718, new_n3719, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775_1, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799_1, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804_1, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3812, new_n3813, new_n3814,
    new_n3815, new_n3816, new_n3817, new_n3818, new_n3819, new_n3820,
    new_n3821, new_n3822, new_n3823, new_n3824, new_n3825, new_n3826,
    new_n3827, new_n3828, new_n3829, new_n3830, new_n3831, new_n3832,
    new_n3833_1, new_n3834, new_n3835, new_n3836, new_n3837, new_n3838,
    new_n3839, new_n3840, new_n3841, new_n3842, new_n3843, new_n3844,
    new_n3845, new_n3846, new_n3847, new_n3848, new_n3849, new_n3850,
    new_n3851, new_n3852, new_n3853, new_n3854_1, new_n3855, new_n3856,
    new_n3857, new_n3858, new_n3859, new_n3860, new_n3861, new_n3862,
    new_n3863, new_n3864, new_n3865, new_n3866, new_n3867, new_n3868,
    new_n3869, new_n3870, new_n3871, new_n3872, new_n3873, new_n3874,
    new_n3875, new_n3876, new_n3877, new_n3878, new_n3879, new_n3880,
    new_n3881, new_n3882, new_n3883, new_n3884, new_n3885, new_n3886,
    new_n3887, new_n3888, new_n3889, new_n3890, new_n3891, new_n3892,
    new_n3893_1, new_n3894, new_n3895, new_n3896, new_n3897, new_n3898,
    new_n3900, new_n3901_1, new_n3902, new_n3903, new_n3904, new_n3905,
    new_n3906, new_n3907, new_n3908, new_n3909, new_n3910_1, new_n3911,
    new_n3912, new_n3913, new_n3914, new_n3915, new_n3916, new_n3917,
    new_n3918, new_n3919, new_n3920, new_n3921, new_n3922, new_n3923,
    new_n3924, new_n3925, new_n3926, new_n3927, new_n3928, new_n3929,
    new_n3930, new_n3931, new_n3932, new_n3933, new_n3934, new_n3935,
    new_n3936, new_n3937, new_n3938, new_n3939, new_n3940, new_n3941,
    new_n3942, new_n3943, new_n3944, new_n3945, new_n3946, new_n3947,
    new_n3948, new_n3949, new_n3950, new_n3951, new_n3952, new_n3953,
    new_n3954, new_n3955, new_n3956, new_n3957, new_n3958, new_n3959,
    new_n3960, new_n3961, new_n3962, new_n3963, new_n3964, new_n3965,
    new_n3966, new_n3967, new_n3968, new_n3969, new_n3970, new_n3971,
    new_n3972_1, new_n3973, new_n3974, new_n3975, new_n3976, new_n3977,
    new_n3978, new_n3979, new_n3980, new_n3981, new_n3982, new_n3983,
    new_n3984, new_n3985, new_n3986, new_n3987, new_n3989, new_n3990,
    new_n3991, new_n3992, new_n3993, new_n3994, new_n3995, new_n3996,
    new_n3997, new_n3998, new_n3999, new_n4000_1, new_n4001, new_n4002,
    new_n4003, new_n4004, new_n4005, new_n4006, new_n4007, new_n4008,
    new_n4009, new_n4010, new_n4011, new_n4012, new_n4013, new_n4014,
    new_n4015, new_n4016, new_n4017, new_n4018, new_n4019, new_n4020,
    new_n4021, new_n4022_1, new_n4023, new_n4024, new_n4025, new_n4026,
    new_n4027, new_n4028, new_n4029, new_n4030, new_n4031, new_n4032,
    new_n4033, new_n4034, new_n4035, new_n4036, new_n4037, new_n4038,
    new_n4039_1, new_n4040, new_n4041, new_n4042, new_n4043, new_n4044,
    new_n4045, new_n4046, new_n4047, new_n4048, new_n4049, new_n4050,
    new_n4051, new_n4052, new_n4053, new_n4054, new_n4055, new_n4056,
    new_n4057, new_n4058, new_n4059, new_n4060, new_n4061, new_n4062,
    new_n4063, new_n4064, new_n4065, new_n4066, new_n4067, new_n4068,
    new_n4069, new_n4070, new_n4071, new_n4072, new_n4073, new_n4074,
    new_n4075, new_n4076, new_n4078, new_n4079, new_n4080, new_n4081,
    new_n4082, new_n4083, new_n4084, new_n4085, new_n4086, new_n4087,
    new_n4088, new_n4089, new_n4090, new_n4091, new_n4092, new_n4093,
    new_n4094, new_n4095, new_n4096, new_n4097, new_n4098, new_n4099,
    new_n4100, new_n4101, new_n4102, new_n4103, new_n4104, new_n4105,
    new_n4106, new_n4107, new_n4108, new_n4109, new_n4110, new_n4111,
    new_n4112, new_n4113, new_n4114, new_n4115, new_n4116, new_n4117_1,
    new_n4118, new_n4119, new_n4120, new_n4121, new_n4122, new_n4123,
    new_n4124, new_n4125_1, new_n4126, new_n4127, new_n4128, new_n4129,
    new_n4130, new_n4131_1, new_n4132, new_n4133, new_n4134, new_n4135,
    new_n4136, new_n4137, new_n4138, new_n4139, new_n4140, new_n4141,
    new_n4142, new_n4143, new_n4144, new_n4145, new_n4146, new_n4147_1,
    new_n4148, new_n4149, new_n4150, new_n4151, new_n4152, new_n4153,
    new_n4154_1, new_n4155, new_n4156, new_n4157, new_n4158, new_n4159,
    new_n4160, new_n4161, new_n4162, new_n4163, new_n4164, new_n4166,
    new_n4167, new_n4168, new_n4169, new_n4170, new_n4171, new_n4172_1,
    new_n4173, new_n4174, new_n4175_1, new_n4176, new_n4177, new_n4178,
    new_n4179, new_n4180, new_n4181, new_n4182, new_n4183, new_n4184,
    new_n4185, new_n4186, new_n4187, new_n4188, new_n4189, new_n4190,
    new_n4191, new_n4192, new_n4193, new_n4194, new_n4195, new_n4196,
    new_n4197, new_n4198, new_n4199, new_n4200, new_n4201, new_n4202,
    new_n4203, new_n4204, new_n4205, new_n4206, new_n4207, new_n4208,
    new_n4209, new_n4210, new_n4211, new_n4212, new_n4213, new_n4214,
    new_n4215, new_n4216, new_n4217, new_n4218, new_n4219, new_n4220,
    new_n4221, new_n4222, new_n4223, new_n4224, new_n4225_1, new_n4226,
    new_n4227, new_n4228, new_n4229, new_n4230, new_n4231, new_n4232,
    new_n4233, new_n4234, new_n4235, new_n4236, new_n4237, new_n4238,
    new_n4239, new_n4240, new_n4241, new_n4242, new_n4243, new_n4244,
    new_n4245, new_n4246, new_n4247, new_n4248, new_n4249, new_n4250,
    new_n4251, new_n4252, new_n4253, new_n4255, new_n4256, new_n4257,
    new_n4258, new_n4259, new_n4260, new_n4261, new_n4262, new_n4263,
    new_n4264, new_n4265, new_n4266, new_n4267, new_n4268, new_n4269,
    new_n4270, new_n4271, new_n4272, new_n4273, new_n4274, new_n4275,
    new_n4276, new_n4277, new_n4278, new_n4279_1, new_n4280, new_n4281,
    new_n4282_1, new_n4283, new_n4284, new_n4285, new_n4286, new_n4287,
    new_n4288, new_n4289, new_n4290, new_n4291, new_n4292_1, new_n4293,
    new_n4294, new_n4295, new_n4296, new_n4297, new_n4298, new_n4299,
    new_n4300, new_n4301, new_n4302, new_n4303, new_n4304, new_n4305_1,
    new_n4306, new_n4307, new_n4308, new_n4309, new_n4310, new_n4311,
    new_n4312, new_n4313, new_n4314, new_n4315, new_n4316, new_n4317,
    new_n4318, new_n4319, new_n4320, new_n4321, new_n4322, new_n4323,
    new_n4324, new_n4325, new_n4326, new_n4327, new_n4328, new_n4329,
    new_n4330, new_n4331, new_n4332, new_n4333, new_n4334, new_n4335,
    new_n4336, new_n4337, new_n4338, new_n4339, new_n4340, new_n4341,
    new_n4343, new_n4344, new_n4345_1, new_n4346, new_n4347, new_n4348,
    new_n4349, new_n4350, new_n4351, new_n4352, new_n4353, new_n4354,
    new_n4355, new_n4356, new_n4357, new_n4358, new_n4359, new_n4360,
    new_n4361, new_n4362, new_n4363, new_n4364, new_n4365, new_n4366,
    new_n4367, new_n4368, new_n4369, new_n4370, new_n4371, new_n4372,
    new_n4373, new_n4374, new_n4375, new_n4376, new_n4377, new_n4378,
    new_n4379, new_n4380, new_n4381, new_n4382, new_n4383, new_n4384,
    new_n4385, new_n4386, new_n4387, new_n4388, new_n4389, new_n4390,
    new_n4391, new_n4392, new_n4393, new_n4394, new_n4395, new_n4396,
    new_n4397, new_n4398, new_n4399, new_n4400, new_n4401, new_n4402,
    new_n4403, new_n4404, new_n4405, new_n4406, new_n4407, new_n4408,
    new_n4409, new_n4410, new_n4411, new_n4412, new_n4413, new_n4414,
    new_n4415, new_n4416, new_n4417, new_n4418, new_n4419, new_n4420,
    new_n4421, new_n4422, new_n4423, new_n4424, new_n4425, new_n4426,
    new_n4427, new_n4428, new_n4429, new_n4430, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436, new_n4437_1, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4522, new_n4523, new_n4524,
    new_n4525, new_n4526, new_n4527, new_n4528, new_n4529, new_n4530,
    new_n4531, new_n4532, new_n4533, new_n4534, new_n4535, new_n4536,
    new_n4537, new_n4538, new_n4539, new_n4540, new_n4541_1, new_n4542,
    new_n4543, new_n4544, new_n4545, new_n4546, new_n4547, new_n4548,
    new_n4549, new_n4550, new_n4551, new_n4552, new_n4553, new_n4554,
    new_n4555, new_n4556, new_n4557, new_n4558, new_n4559, new_n4560,
    new_n4561, new_n4562, new_n4563, new_n4564, new_n4565, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4574, new_n4575, new_n4576, new_n4577, new_n4578,
    new_n4579, new_n4580, new_n4581, new_n4582, new_n4583, new_n4584,
    new_n4585, new_n4586, new_n4587, new_n4588, new_n4589, new_n4590,
    new_n4591, new_n4592, new_n4593, new_n4594, new_n4595, new_n4596,
    new_n4597, new_n4598, new_n4599, new_n4600, new_n4601, new_n4602,
    new_n4603, new_n4604_1, new_n4605, new_n4606, new_n4607, new_n4608,
    new_n4610, new_n4611, new_n4612, new_n4613, new_n4614, new_n4615_1,
    new_n4616, new_n4617, new_n4618, new_n4619, new_n4620, new_n4621,
    new_n4622, new_n4623, new_n4624, new_n4625, new_n4626, new_n4627,
    new_n4628, new_n4629, new_n4630, new_n4631, new_n4632, new_n4633,
    new_n4634, new_n4635, new_n4636, new_n4637, new_n4638, new_n4639,
    new_n4640, new_n4641, new_n4642, new_n4643, new_n4644, new_n4645,
    new_n4646, new_n4647, new_n4648, new_n4649, new_n4650, new_n4651,
    new_n4652, new_n4653, new_n4654, new_n4655, new_n4656, new_n4657,
    new_n4658, new_n4659_1, new_n4660, new_n4661, new_n4662, new_n4663,
    new_n4664, new_n4665, new_n4666, new_n4667, new_n4668, new_n4669,
    new_n4670, new_n4671, new_n4672_1, new_n4673, new_n4674, new_n4675,
    new_n4676, new_n4677, new_n4678, new_n4679, new_n4680, new_n4681,
    new_n4682, new_n4683, new_n4684, new_n4685, new_n4686, new_n4687,
    new_n4688, new_n4689, new_n4690, new_n4691, new_n4692, new_n4693,
    new_n4694, new_n4695, new_n4696, new_n4698, new_n4699, new_n4700,
    new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706,
    new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712,
    new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718,
    new_n4719, new_n4720, new_n4721, new_n4722, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745, new_n4746, new_n4747, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755_1, new_n4756, new_n4757, new_n4758, new_n4759, new_n4760,
    new_n4761, new_n4762, new_n4763, new_n4764, new_n4765, new_n4766,
    new_n4767, new_n4768, new_n4769, new_n4770, new_n4771, new_n4772,
    new_n4773, new_n4774_1, new_n4775, new_n4776, new_n4777, new_n4778,
    new_n4779, new_n4780, new_n4781, new_n4782, new_n4783, new_n4784,
    new_n4785_1, new_n4786, new_n4787, new_n4788, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4854, new_n4855, new_n4856, new_n4857, new_n4858_1,
    new_n4859, new_n4860, new_n4861, new_n4862, new_n4863, new_n4864,
    new_n4865, new_n4866, new_n4867, new_n4868, new_n4869, new_n4870,
    new_n4871, new_n4872, new_n4873, new_n4874, new_n4875, new_n4876,
    new_n4877, new_n4878, new_n4879, new_n4880, new_n4881, new_n4882,
    new_n4883, new_n4884, new_n4885, new_n4886, new_n4887, new_n4888,
    new_n4889, new_n4890, new_n4891, new_n4892, new_n4893, new_n4894,
    new_n4895_1, new_n4896, new_n4897, new_n4898, new_n4899, new_n4900,
    new_n4901, new_n4902, new_n4903, new_n4904, new_n4905, new_n4906,
    new_n4907_1, new_n4908, new_n4909, new_n4910, new_n4911, new_n4912,
    new_n4913, new_n4914, new_n4915, new_n4916, new_n4917, new_n4918,
    new_n4919, new_n4920, new_n4921, new_n4922, new_n4923, new_n4924,
    new_n4925, new_n4926, new_n4927, new_n4928, new_n4929, new_n4930,
    new_n4931, new_n4932, new_n4933, new_n4934, new_n4935, new_n4936,
    new_n4937, new_n4938, new_n4939, new_n4940, new_n4941, new_n4942,
    new_n4943, new_n4945, new_n4946, new_n4947, new_n4948, new_n4949,
    new_n4950, new_n4951, new_n4952, new_n4953, new_n4954, new_n4955,
    new_n4956, new_n4957, new_n4958, new_n4959, new_n4960, new_n4961,
    new_n4962, new_n4963, new_n4964, new_n4965, new_n4966, new_n4967,
    new_n4968, new_n4969, new_n4970, new_n4971_1, new_n4972, new_n4973,
    new_n4974, new_n4975, new_n4976, new_n4977, new_n4978, new_n4979,
    new_n4980, new_n4981, new_n4982, new_n4983, new_n4984, new_n4985,
    new_n4986, new_n4987, new_n4988, new_n4989, new_n4990, new_n4991,
    new_n4992, new_n4993, new_n4994, new_n4995, new_n4996, new_n4997,
    new_n4998, new_n4999, new_n5000, new_n5001, new_n5002, new_n5003,
    new_n5004, new_n5005, new_n5006, new_n5007, new_n5008, new_n5009_1,
    new_n5010, new_n5011, new_n5012, new_n5013, new_n5014_1, new_n5015,
    new_n5016, new_n5017, new_n5018, new_n5019, new_n5020, new_n5021,
    new_n5022, new_n5023_1, new_n5024, new_n5025, new_n5026, new_n5027,
    new_n5028, new_n5029, new_n5030, new_n5031, new_n5033_1, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046_1,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060, new_n5061, new_n5062, new_n5063, new_n5064,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077_1, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098, new_n5099, new_n5100,
    new_n5101, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5121, new_n5122, new_n5123, new_n5124, new_n5125,
    new_n5126, new_n5127, new_n5128, new_n5129, new_n5130, new_n5131,
    new_n5132, new_n5133, new_n5134, new_n5135, new_n5136, new_n5137,
    new_n5138, new_n5139, new_n5140, new_n5141, new_n5142, new_n5143,
    new_n5144, new_n5145, new_n5146, new_n5147, new_n5148, new_n5149,
    new_n5150, new_n5151, new_n5152, new_n5153, new_n5154, new_n5155,
    new_n5156, new_n5157, new_n5158, new_n5159, new_n5160, new_n5161,
    new_n5162, new_n5163, new_n5164, new_n5165, new_n5166, new_n5167,
    new_n5168, new_n5169, new_n5170, new_n5171, new_n5172, new_n5173,
    new_n5174, new_n5175, new_n5176, new_n5177, new_n5178, new_n5179,
    new_n5180, new_n5181, new_n5182, new_n5183, new_n5184_1, new_n5185_1,
    new_n5186, new_n5187, new_n5188, new_n5189, new_n5190, new_n5191,
    new_n5192, new_n5193, new_n5194, new_n5195, new_n5196, new_n5197,
    new_n5198, new_n5199, new_n5200, new_n5201, new_n5202, new_n5203,
    new_n5204, new_n5205, new_n5206, new_n5207, new_n5208, new_n5210,
    new_n5211, new_n5212, new_n5213, new_n5214, new_n5215, new_n5216,
    new_n5217, new_n5218, new_n5219, new_n5220, new_n5221, new_n5222,
    new_n5223, new_n5224, new_n5225_1, new_n5226, new_n5227, new_n5228,
    new_n5229, new_n5230, new_n5231, new_n5232, new_n5233, new_n5234,
    new_n5235, new_n5236, new_n5237, new_n5238, new_n5239, new_n5240,
    new_n5241, new_n5242, new_n5243, new_n5244, new_n5245, new_n5246,
    new_n5247, new_n5248, new_n5249, new_n5250, new_n5251, new_n5252,
    new_n5253, new_n5254, new_n5255, new_n5256, new_n5257, new_n5258,
    new_n5259, new_n5260, new_n5261, new_n5262, new_n5263, new_n5264,
    new_n5265, new_n5266, new_n5267, new_n5268, new_n5269, new_n5270,
    new_n5271, new_n5272, new_n5273, new_n5274, new_n5275, new_n5276,
    new_n5277, new_n5278, new_n5279, new_n5280, new_n5281, new_n5282,
    new_n5283, new_n5284, new_n5285, new_n5286, new_n5287, new_n5288,
    new_n5289, new_n5290, new_n5291, new_n5292, new_n5293, new_n5294,
    new_n5295, new_n5296, new_n5297, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319,
    new_n5320, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5387, new_n5388, new_n5389, new_n5390, new_n5391, new_n5392,
    new_n5393, new_n5394, new_n5395, new_n5396, new_n5397, new_n5398,
    new_n5399, new_n5400, new_n5401, new_n5402, new_n5403, new_n5404,
    new_n5405, new_n5406, new_n5407, new_n5408, new_n5409, new_n5410,
    new_n5411, new_n5412, new_n5413, new_n5414, new_n5415, new_n5416,
    new_n5417, new_n5418, new_n5419, new_n5420, new_n5421, new_n5422,
    new_n5423, new_n5424, new_n5425, new_n5426, new_n5427, new_n5428,
    new_n5429, new_n5430_1, new_n5431, new_n5432, new_n5433, new_n5434,
    new_n5435, new_n5436, new_n5437, new_n5438, new_n5439, new_n5440,
    new_n5441, new_n5442, new_n5443, new_n5444, new_n5445, new_n5446,
    new_n5447, new_n5448, new_n5449_1, new_n5450, new_n5451, new_n5452,
    new_n5453, new_n5454, new_n5455, new_n5456, new_n5457, new_n5458,
    new_n5459, new_n5460, new_n5461, new_n5462, new_n5463, new_n5464,
    new_n5465, new_n5466, new_n5467_1, new_n5468, new_n5469, new_n5470,
    new_n5471, new_n5472, new_n5473, new_n5475, new_n5476, new_n5477,
    new_n5478, new_n5479_1, new_n5480, new_n5481, new_n5482, new_n5483,
    new_n5484, new_n5485, new_n5486, new_n5487, new_n5488, new_n5489,
    new_n5490, new_n5491, new_n5492, new_n5493, new_n5494, new_n5495,
    new_n5496, new_n5497, new_n5498, new_n5499, new_n5500, new_n5501,
    new_n5502_1, new_n5503, new_n5504, new_n5505, new_n5506, new_n5507,
    new_n5508, new_n5509, new_n5510, new_n5511, new_n5512, new_n5513,
    new_n5514, new_n5515, new_n5516, new_n5517, new_n5518, new_n5519,
    new_n5520, new_n5521, new_n5522, new_n5523, new_n5524, new_n5525,
    new_n5526, new_n5527, new_n5528, new_n5529, new_n5530, new_n5531,
    new_n5532, new_n5533, new_n5534, new_n5535, new_n5536, new_n5537,
    new_n5538, new_n5539, new_n5540, new_n5541, new_n5542, new_n5543,
    new_n5544, new_n5545, new_n5546, new_n5547, new_n5548, new_n5549,
    new_n5550_1, new_n5551, new_n5552, new_n5553, new_n5554, new_n5555,
    new_n5556, new_n5557, new_n5558, new_n5559, new_n5560, new_n5561,
    new_n5562, new_n5564, new_n5565, new_n5566, new_n5567, new_n5568,
    new_n5569, new_n5570, new_n5571, new_n5572, new_n5573, new_n5574,
    new_n5575, new_n5576, new_n5577, new_n5578, new_n5579, new_n5580,
    new_n5581, new_n5582, new_n5583, new_n5584, new_n5585, new_n5586_1,
    new_n5587, new_n5588, new_n5589, new_n5590, new_n5591, new_n5592,
    new_n5593, new_n5594, new_n5595, new_n5596, new_n5597, new_n5598,
    new_n5599, new_n5600, new_n5601_1, new_n5602, new_n5603, new_n5604,
    new_n5605, new_n5606, new_n5607, new_n5608, new_n5609, new_n5610,
    new_n5611, new_n5612, new_n5613, new_n5614, new_n5615, new_n5616,
    new_n5617, new_n5618, new_n5619, new_n5620, new_n5621, new_n5622,
    new_n5623, new_n5624, new_n5625, new_n5626, new_n5627, new_n5628,
    new_n5629, new_n5630, new_n5631, new_n5632, new_n5633, new_n5634,
    new_n5635, new_n5636, new_n5637, new_n5638, new_n5639, new_n5640,
    new_n5641, new_n5642, new_n5643, new_n5644, new_n5645, new_n5646,
    new_n5647, new_n5648, new_n5649, new_n5650, new_n5651, new_n5653,
    new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659,
    new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665,
    new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671,
    new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677,
    new_n5678, new_n5679, new_n5680, new_n5681, new_n5682, new_n5683,
    new_n5684, new_n5685, new_n5686, new_n5687, new_n5688, new_n5689,
    new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695,
    new_n5696, new_n5697, new_n5698, new_n5699, new_n5700, new_n5701,
    new_n5702, new_n5703, new_n5704, new_n5705, new_n5706, new_n5707,
    new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713,
    new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719,
    new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725_1,
    new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731,
    new_n5732, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5743, new_n5744,
    new_n5745, new_n5746, new_n5747, new_n5748, new_n5749, new_n5750,
    new_n5751, new_n5752, new_n5753, new_n5754, new_n5755, new_n5756,
    new_n5757, new_n5758, new_n5759, new_n5760, new_n5761, new_n5762,
    new_n5763, new_n5764, new_n5765, new_n5766, new_n5767, new_n5768,
    new_n5769, new_n5770, new_n5771, new_n5772, new_n5773, new_n5774,
    new_n5775, new_n5776, new_n5777, new_n5778, new_n5779, new_n5780,
    new_n5781, new_n5782, new_n5783, new_n5784, new_n5785, new_n5786_1,
    new_n5787, new_n5788, new_n5789, new_n5790, new_n5791, new_n5792,
    new_n5793, new_n5794, new_n5795, new_n5796, new_n5797, new_n5798,
    new_n5799, new_n5800, new_n5801, new_n5802, new_n5803, new_n5804,
    new_n5805, new_n5806_1, new_n5807, new_n5808, new_n5809, new_n5810,
    new_n5811, new_n5812, new_n5813, new_n5814, new_n5815, new_n5816,
    new_n5817, new_n5818, new_n5819, new_n5820, new_n5821, new_n5822,
    new_n5823, new_n5824, new_n5825, new_n5826, new_n5827, new_n5828,
    new_n5829, new_n5830, new_n5831, new_n5832, new_n5834, new_n5835,
    new_n5836, new_n5837, new_n5838, new_n5839, new_n5840, new_n5841,
    new_n5842, new_n5843, new_n5844, new_n5845, new_n5846, new_n5847,
    new_n5848, new_n5849, new_n5850, new_n5851_1, new_n5852, new_n5853,
    new_n5854, new_n5855, new_n5856, new_n5857, new_n5858, new_n5859,
    new_n5860, new_n5861, new_n5862, new_n5863, new_n5864, new_n5865,
    new_n5866, new_n5867, new_n5868, new_n5869, new_n5870, new_n5871,
    new_n5872, new_n5873, new_n5874, new_n5875, new_n5876, new_n5877,
    new_n5878, new_n5879, new_n5880, new_n5881, new_n5882, new_n5883,
    new_n5884, new_n5885, new_n5886, new_n5887, new_n5888, new_n5889,
    new_n5890, new_n5891, new_n5892, new_n5893, new_n5894, new_n5895,
    new_n5896, new_n5897, new_n5898, new_n5899, new_n5900, new_n5901,
    new_n5902, new_n5903, new_n5904, new_n5905, new_n5906, new_n5907,
    new_n5908, new_n5909, new_n5910, new_n5911, new_n5912, new_n5913,
    new_n5914, new_n5915, new_n5916, new_n5917, new_n5918, new_n5919,
    new_n5920, new_n5921, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943_1, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950_1,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960_1, new_n5961, new_n5962,
    new_n5963, new_n5964, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980,
    new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986,
    new_n5987_1, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992,
    new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998,
    new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004,
    new_n6005, new_n6006, new_n6007_1, new_n6008, new_n6009, new_n6011,
    new_n6012_1, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054_1, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6100, new_n6101, new_n6102,
    new_n6103, new_n6104, new_n6105, new_n6106, new_n6107, new_n6108,
    new_n6109, new_n6110, new_n6111, new_n6112, new_n6113, new_n6114_1,
    new_n6115, new_n6116, new_n6117, new_n6118, new_n6119, new_n6120,
    new_n6121, new_n6122, new_n6123, new_n6124, new_n6125, new_n6126,
    new_n6127, new_n6128, new_n6129, new_n6130, new_n6131, new_n6132,
    new_n6133, new_n6134, new_n6135, new_n6136, new_n6137, new_n6138,
    new_n6139, new_n6140, new_n6141, new_n6142, new_n6143, new_n6144,
    new_n6145, new_n6146, new_n6147_1, new_n6148, new_n6149, new_n6150,
    new_n6151, new_n6152, new_n6153, new_n6154, new_n6155, new_n6156,
    new_n6157, new_n6158, new_n6159, new_n6160, new_n6161, new_n6162,
    new_n6163, new_n6164, new_n6165, new_n6166, new_n6167, new_n6168,
    new_n6169, new_n6170, new_n6171, new_n6172, new_n6173, new_n6174,
    new_n6175, new_n6176, new_n6177, new_n6178, new_n6179, new_n6180,
    new_n6181, new_n6182, new_n6183, new_n6184, new_n6185, new_n6186,
    new_n6188, new_n6189, new_n6190, new_n6191, new_n6192, new_n6193,
    new_n6194, new_n6195, new_n6196, new_n6197, new_n6198_1, new_n6199,
    new_n6200, new_n6201, new_n6202, new_n6203, new_n6204, new_n6205,
    new_n6206, new_n6207, new_n6208, new_n6209, new_n6210, new_n6211,
    new_n6212, new_n6213, new_n6214, new_n6215, new_n6216, new_n6217,
    new_n6218, new_n6219, new_n6220, new_n6221, new_n6222, new_n6223,
    new_n6224, new_n6225, new_n6226, new_n6227, new_n6228, new_n6229,
    new_n6230, new_n6231, new_n6232, new_n6233, new_n6234, new_n6235,
    new_n6236, new_n6237, new_n6238, new_n6239, new_n6240, new_n6241,
    new_n6242, new_n6243, new_n6244, new_n6245, new_n6246, new_n6247,
    new_n6248, new_n6249, new_n6250, new_n6251_1, new_n6252, new_n6253,
    new_n6254, new_n6255, new_n6256, new_n6257, new_n6258_1, new_n6259,
    new_n6260, new_n6261, new_n6262, new_n6263, new_n6264, new_n6265,
    new_n6266, new_n6267, new_n6268, new_n6269, new_n6270_1, new_n6271,
    new_n6272, new_n6273, new_n6274, new_n6275_1, new_n6277, new_n6278,
    new_n6279, new_n6280, new_n6281, new_n6282, new_n6283, new_n6284,
    new_n6285, new_n6286, new_n6287, new_n6288, new_n6289, new_n6290,
    new_n6291, new_n6292, new_n6293, new_n6294, new_n6295, new_n6296,
    new_n6297, new_n6298, new_n6299, new_n6300, new_n6301, new_n6302,
    new_n6303, new_n6304, new_n6305, new_n6306, new_n6307, new_n6308,
    new_n6309, new_n6310, new_n6311, new_n6312, new_n6313, new_n6314_1,
    new_n6315, new_n6316, new_n6317, new_n6318, new_n6319, new_n6320,
    new_n6321, new_n6322, new_n6323, new_n6324, new_n6325, new_n6326,
    new_n6327, new_n6328, new_n6329, new_n6330, new_n6331, new_n6332,
    new_n6333, new_n6334, new_n6335, new_n6336, new_n6337, new_n6338,
    new_n6339, new_n6340, new_n6341, new_n6342, new_n6343, new_n6344,
    new_n6345, new_n6346, new_n6347, new_n6348, new_n6349, new_n6350,
    new_n6351, new_n6352, new_n6353, new_n6354, new_n6355, new_n6356,
    new_n6357, new_n6358, new_n6359, new_n6360, new_n6361, new_n6362_1,
    new_n6363, new_n6365, new_n6366, new_n6367, new_n6368, new_n6369,
    new_n6370, new_n6371, new_n6372, new_n6373, new_n6374, new_n6375,
    new_n6376, new_n6377, new_n6378, new_n6379, new_n6380, new_n6381,
    new_n6382, new_n6383, new_n6384, new_n6385, new_n6386, new_n6387,
    new_n6388, new_n6389, new_n6390, new_n6391, new_n6392, new_n6393,
    new_n6394, new_n6395, new_n6396, new_n6397, new_n6398, new_n6399,
    new_n6400, new_n6401, new_n6402, new_n6403, new_n6404, new_n6405,
    new_n6406, new_n6407, new_n6408, new_n6409, new_n6410, new_n6411,
    new_n6412, new_n6413, new_n6414, new_n6415, new_n6416, new_n6417,
    new_n6418, new_n6419, new_n6420, new_n6421, new_n6422, new_n6423,
    new_n6424, new_n6425, new_n6426, new_n6427, new_n6428, new_n6429,
    new_n6430, new_n6431, new_n6432, new_n6433, new_n6434, new_n6435,
    new_n6436_1, new_n6437, new_n6438, new_n6439, new_n6440, new_n6441,
    new_n6442, new_n6443, new_n6444, new_n6445, new_n6446, new_n6447,
    new_n6448, new_n6449, new_n6450, new_n6451, new_n6452, new_n6453,
    new_n6455, new_n6456, new_n6457, new_n6458, new_n6459, new_n6460_1,
    new_n6461, new_n6462, new_n6463, new_n6464, new_n6465, new_n6466,
    new_n6467, new_n6468, new_n6469, new_n6470, new_n6471, new_n6472,
    new_n6473, new_n6474, new_n6475, new_n6476, new_n6477, new_n6478,
    new_n6479, new_n6480_1, new_n6481, new_n6482, new_n6483, new_n6484,
    new_n6485, new_n6486, new_n6487, new_n6488, new_n6489, new_n6490,
    new_n6491, new_n6492, new_n6493, new_n6494, new_n6495, new_n6496,
    new_n6497, new_n6498, new_n6499, new_n6500, new_n6501, new_n6502,
    new_n6503, new_n6504, new_n6505, new_n6506, new_n6507, new_n6508,
    new_n6509, new_n6510, new_n6511, new_n6512, new_n6513, new_n6514,
    new_n6515, new_n6516, new_n6517_1, new_n6518, new_n6519, new_n6520,
    new_n6521, new_n6522, new_n6523, new_n6524, new_n6525, new_n6526,
    new_n6527, new_n6528, new_n6529, new_n6530, new_n6531, new_n6532,
    new_n6533, new_n6534, new_n6535, new_n6536, new_n6537, new_n6538,
    new_n6539, new_n6540, new_n6541, new_n6542, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555_1, new_n6556, new_n6557,
    new_n6558, new_n6559, new_n6560, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576, new_n6577, new_n6578, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6584, new_n6585, new_n6586_1, new_n6587,
    new_n6588, new_n6589, new_n6590, new_n6591, new_n6592, new_n6593,
    new_n6594, new_n6595, new_n6596, new_n6597, new_n6598, new_n6599,
    new_n6600, new_n6601, new_n6602, new_n6603, new_n6604, new_n6605,
    new_n6606, new_n6607, new_n6608, new_n6609, new_n6610, new_n6611,
    new_n6612, new_n6613, new_n6614, new_n6615, new_n6616, new_n6617,
    new_n6618, new_n6619, new_n6620, new_n6621, new_n6622, new_n6623,
    new_n6624, new_n6625, new_n6626, new_n6627, new_n6628, new_n6629,
    new_n6630, new_n6632, new_n6633, new_n6634, new_n6635, new_n6636,
    new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652, new_n6653, new_n6654,
    new_n6655, new_n6656, new_n6657, new_n6658, new_n6659, new_n6660,
    new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669, new_n6670, new_n6671, new_n6672,
    new_n6673, new_n6674, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680_1, new_n6681, new_n6682_1, new_n6683, new_n6684,
    new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690,
    new_n6691, new_n6692, new_n6693_1, new_n6694, new_n6695, new_n6696_1,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703_1, new_n6704, new_n6705, new_n6706, new_n6707, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6717, new_n6718, new_n6720, new_n6721,
    new_n6722, new_n6723, new_n6724, new_n6725, new_n6726, new_n6727,
    new_n6728, new_n6729, new_n6730, new_n6731, new_n6732, new_n6733,
    new_n6734, new_n6735, new_n6736, new_n6737, new_n6738, new_n6739,
    new_n6740, new_n6741, new_n6742, new_n6743, new_n6744, new_n6745,
    new_n6746, new_n6747, new_n6748, new_n6749, new_n6750, new_n6751,
    new_n6752, new_n6753, new_n6754, new_n6755, new_n6756, new_n6757,
    new_n6758_1, new_n6759, new_n6760, new_n6761, new_n6762, new_n6763,
    new_n6764, new_n6765, new_n6766, new_n6767, new_n6768, new_n6769,
    new_n6770, new_n6771, new_n6772, new_n6773, new_n6774, new_n6775,
    new_n6776, new_n6777, new_n6778, new_n6779, new_n6780, new_n6781,
    new_n6782, new_n6783, new_n6784, new_n6785, new_n6786_1, new_n6787,
    new_n6788, new_n6789, new_n6790, new_n6791_1, new_n6792, new_n6793,
    new_n6794, new_n6795, new_n6796, new_n6797, new_n6798, new_n6799,
    new_n6800, new_n6801, new_n6802, new_n6803, new_n6804, new_n6805,
    new_n6806, new_n6808, new_n6809, new_n6810_1, new_n6811, new_n6812,
    new_n6813, new_n6814, new_n6815, new_n6816, new_n6817, new_n6818,
    new_n6819, new_n6820, new_n6821, new_n6822, new_n6823, new_n6824,
    new_n6825, new_n6826, new_n6827, new_n6828, new_n6829, new_n6830,
    new_n6831, new_n6832, new_n6833, new_n6834, new_n6835, new_n6836,
    new_n6837, new_n6838, new_n6839, new_n6840, new_n6841, new_n6842,
    new_n6843, new_n6844, new_n6845, new_n6846, new_n6847, new_n6848,
    new_n6849, new_n6850, new_n6851, new_n6852, new_n6853_1, new_n6854,
    new_n6855, new_n6856, new_n6857, new_n6858, new_n6859, new_n6860,
    new_n6861, new_n6862, new_n6863, new_n6864, new_n6865, new_n6866,
    new_n6867, new_n6868, new_n6869, new_n6870, new_n6871, new_n6872,
    new_n6873_1, new_n6874, new_n6875, new_n6876, new_n6877, new_n6878,
    new_n6879, new_n6880, new_n6881, new_n6882, new_n6883, new_n6884,
    new_n6885, new_n6886, new_n6887, new_n6888, new_n6889, new_n6890,
    new_n6891, new_n6892, new_n6893, new_n6894, new_n6895, new_n6896,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946_1, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952_1, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979_1, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6986, new_n6987, new_n6988,
    new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994,
    new_n6995, new_n6996, new_n6997, new_n6998, new_n6999_1, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054,
    new_n7055, new_n7056, new_n7057, new_n7058, new_n7059, new_n7060,
    new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066,
    new_n7067, new_n7068, new_n7069, new_n7070, new_n7071_1, new_n7072,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104_1, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132_1, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152_1, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159, new_n7160, new_n7162, new_n7163, new_n7164,
    new_n7165, new_n7166, new_n7167, new_n7168, new_n7169, new_n7170,
    new_n7171, new_n7172, new_n7173, new_n7174, new_n7175, new_n7176,
    new_n7177, new_n7178, new_n7179, new_n7180, new_n7181, new_n7182,
    new_n7183, new_n7184, new_n7185, new_n7186, new_n7187, new_n7188,
    new_n7189, new_n7190, new_n7191, new_n7192, new_n7193, new_n7194,
    new_n7195, new_n7196, new_n7197, new_n7198, new_n7199, new_n7200,
    new_n7201, new_n7202, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229, new_n7230,
    new_n7231, new_n7232, new_n7233, new_n7234, new_n7235, new_n7236,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246_1, new_n7247, new_n7248,
    new_n7250, new_n7251, new_n7252, new_n7253, new_n7254, new_n7255,
    new_n7256, new_n7257, new_n7258, new_n7259, new_n7260, new_n7261,
    new_n7262, new_n7263, new_n7264, new_n7265_1, new_n7266, new_n7267,
    new_n7268, new_n7269, new_n7270, new_n7271, new_n7272_1, new_n7273,
    new_n7274, new_n7275, new_n7276, new_n7277, new_n7278, new_n7279,
    new_n7280, new_n7281, new_n7282_1, new_n7283, new_n7284, new_n7285,
    new_n7286, new_n7287, new_n7288, new_n7289, new_n7290, new_n7291,
    new_n7292, new_n7293, new_n7294, new_n7295, new_n7296, new_n7297,
    new_n7298, new_n7299, new_n7300, new_n7301, new_n7302, new_n7303,
    new_n7304, new_n7305, new_n7306, new_n7307, new_n7308, new_n7309,
    new_n7310, new_n7311, new_n7312, new_n7313, new_n7314, new_n7315,
    new_n7316, new_n7317, new_n7318, new_n7319, new_n7320, new_n7321,
    new_n7322, new_n7323, new_n7324, new_n7325, new_n7326, new_n7327,
    new_n7328, new_n7329, new_n7330, new_n7331, new_n7332, new_n7333,
    new_n7334, new_n7335, new_n7336, new_n7338, new_n7339, new_n7340,
    new_n7341, new_n7342, new_n7343, new_n7344, new_n7345, new_n7346,
    new_n7347, new_n7348, new_n7349, new_n7350, new_n7351, new_n7352,
    new_n7353, new_n7354_1, new_n7355, new_n7356, new_n7357, new_n7358,
    new_n7359, new_n7360, new_n7361, new_n7362, new_n7363, new_n7364,
    new_n7365, new_n7366, new_n7367, new_n7368, new_n7369, new_n7370,
    new_n7371, new_n7372, new_n7373, new_n7374, new_n7375, new_n7376,
    new_n7377, new_n7378, new_n7379, new_n7380, new_n7381, new_n7382_1,
    new_n7383, new_n7384, new_n7385, new_n7386, new_n7387, new_n7388,
    new_n7389, new_n7390, new_n7391, new_n7392, new_n7393, new_n7394,
    new_n7395, new_n7396, new_n7397, new_n7398, new_n7399, new_n7400,
    new_n7401, new_n7402, new_n7403, new_n7404, new_n7405, new_n7406,
    new_n7407, new_n7408, new_n7409, new_n7410, new_n7411, new_n7412,
    new_n7413, new_n7414, new_n7415, new_n7416, new_n7417, new_n7418,
    new_n7419, new_n7420, new_n7421, new_n7422, new_n7423, new_n7424,
    new_n7426, new_n7427, new_n7428, new_n7429, new_n7430, new_n7431,
    new_n7432, new_n7433, new_n7434, new_n7435, new_n7436, new_n7437,
    new_n7438, new_n7439, new_n7440, new_n7441, new_n7442, new_n7443,
    new_n7444, new_n7445, new_n7446, new_n7447, new_n7448, new_n7449,
    new_n7450_1, new_n7451, new_n7452, new_n7453, new_n7454, new_n7455,
    new_n7456, new_n7457, new_n7458, new_n7459, new_n7460, new_n7461,
    new_n7462, new_n7463, new_n7464, new_n7465, new_n7466, new_n7467,
    new_n7468, new_n7469, new_n7470, new_n7471, new_n7472, new_n7473,
    new_n7474, new_n7475, new_n7476, new_n7477, new_n7478, new_n7479,
    new_n7480, new_n7481, new_n7482, new_n7483, new_n7484, new_n7485,
    new_n7486, new_n7487, new_n7488, new_n7489, new_n7490, new_n7491,
    new_n7492, new_n7493, new_n7494, new_n7495, new_n7496, new_n7497,
    new_n7498, new_n7499, new_n7500, new_n7501, new_n7502, new_n7503,
    new_n7504, new_n7505, new_n7506, new_n7507, new_n7508, new_n7509,
    new_n7510, new_n7511, new_n7512, new_n7514, new_n7515, new_n7516,
    new_n7517, new_n7518, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566, new_n7567, new_n7568, new_n7569, new_n7570,
    new_n7571, new_n7572, new_n7573, new_n7574, new_n7575, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582,
    new_n7583, new_n7584, new_n7585, new_n7586, new_n7587, new_n7588,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598, new_n7599, new_n7600,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652_1, new_n7653, new_n7654, new_n7655_1,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667_1,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690, new_n7692,
    new_n7693, new_n7694, new_n7695, new_n7696, new_n7697, new_n7698,
    new_n7699, new_n7700, new_n7701, new_n7702, new_n7703, new_n7704,
    new_n7705, new_n7706, new_n7707, new_n7708, new_n7709, new_n7710,
    new_n7711, new_n7712, new_n7713, new_n7714, new_n7715, new_n7716,
    new_n7717, new_n7718, new_n7719, new_n7720, new_n7721, new_n7722,
    new_n7723, new_n7724, new_n7725, new_n7726, new_n7727, new_n7728,
    new_n7729, new_n7730, new_n7731, new_n7732, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748_1, new_n7749, new_n7750, new_n7751, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769, new_n7770,
    new_n7771_1, new_n7772, new_n7773, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7780, new_n7781, new_n7782, new_n7783,
    new_n7784, new_n7785, new_n7786, new_n7787, new_n7788, new_n7789,
    new_n7790, new_n7791, new_n7792, new_n7793, new_n7794, new_n7795,
    new_n7796, new_n7797, new_n7798, new_n7799, new_n7800, new_n7801,
    new_n7802, new_n7803, new_n7804, new_n7805, new_n7806, new_n7807,
    new_n7808, new_n7809, new_n7810, new_n7811, new_n7812, new_n7813,
    new_n7814, new_n7815, new_n7816, new_n7817, new_n7818, new_n7819,
    new_n7820, new_n7821, new_n7822, new_n7823, new_n7824, new_n7825_1,
    new_n7826, new_n7827, new_n7828, new_n7829, new_n7830, new_n7831,
    new_n7832_1, new_n7833, new_n7834, new_n7835, new_n7836, new_n7837,
    new_n7838, new_n7839, new_n7840, new_n7841, new_n7842, new_n7843,
    new_n7844, new_n7845, new_n7846, new_n7847, new_n7848, new_n7849,
    new_n7850, new_n7851, new_n7852, new_n7853, new_n7854, new_n7855,
    new_n7856, new_n7857, new_n7858, new_n7859, new_n7860, new_n7861,
    new_n7862, new_n7863, new_n7864, new_n7865, new_n7866, new_n7868,
    new_n7869, new_n7870, new_n7871, new_n7872, new_n7873, new_n7874,
    new_n7875, new_n7876, new_n7877, new_n7878, new_n7879, new_n7880,
    new_n7881, new_n7882, new_n7883, new_n7884, new_n7885, new_n7886,
    new_n7887, new_n7888, new_n7889, new_n7890, new_n7891, new_n7892,
    new_n7893, new_n7894, new_n7895, new_n7896, new_n7897, new_n7898,
    new_n7899, new_n7900, new_n7901, new_n7902, new_n7903, new_n7904,
    new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7917, new_n7918, new_n7919, new_n7920, new_n7921, new_n7922,
    new_n7923, new_n7924, new_n7925, new_n7926, new_n7927, new_n7928,
    new_n7929, new_n7930, new_n7931, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937, new_n7938, new_n7939, new_n7940,
    new_n7941_1, new_n7942, new_n7943, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949, new_n7950, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7959,
    new_n7960, new_n7961, new_n7962, new_n7963, new_n7964, new_n7965,
    new_n7966, new_n7967, new_n7968, new_n7969, new_n7970, new_n7971,
    new_n7972_1, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977,
    new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983,
    new_n7984, new_n7985, new_n7986, new_n7987, new_n7988_1, new_n7989,
    new_n7990, new_n7991, new_n7992, new_n7993, new_n7994, new_n7995,
    new_n7996, new_n7997, new_n7998, new_n7999, new_n8000, new_n8001,
    new_n8002_1, new_n8003, new_n8004, new_n8005, new_n8006, new_n8007,
    new_n8008, new_n8009, new_n8010, new_n8011, new_n8012, new_n8013,
    new_n8014, new_n8015, new_n8016, new_n8017, new_n8018, new_n8019,
    new_n8020, new_n8021, new_n8022, new_n8023, new_n8024, new_n8025,
    new_n8026, new_n8027, new_n8028, new_n8029, new_n8030, new_n8031,
    new_n8032, new_n8033, new_n8034, new_n8035, new_n8036, new_n8037,
    new_n8038, new_n8039, new_n8040, new_n8041, new_n8042, new_n8043,
    new_n8044_1, new_n8045, new_n8047, new_n8048, new_n8049, new_n8050,
    new_n8051, new_n8052, new_n8053, new_n8054, new_n8055, new_n8056,
    new_n8057, new_n8058, new_n8059, new_n8060, new_n8061, new_n8062,
    new_n8063, new_n8064, new_n8065, new_n8066, new_n8067, new_n8068_1,
    new_n8069, new_n8070, new_n8071, new_n8072, new_n8073_1, new_n8074,
    new_n8075, new_n8076, new_n8077, new_n8078, new_n8079, new_n8080,
    new_n8081, new_n8082, new_n8083, new_n8084, new_n8085_1, new_n8086,
    new_n8087, new_n8088, new_n8089, new_n8090, new_n8091, new_n8092,
    new_n8093, new_n8094, new_n8095, new_n8096, new_n8097, new_n8098,
    new_n8099, new_n8100, new_n8101, new_n8102, new_n8103, new_n8104,
    new_n8105, new_n8106, new_n8107, new_n8108, new_n8109, new_n8110,
    new_n8111, new_n8112, new_n8113, new_n8114, new_n8115, new_n8116,
    new_n8117, new_n8118, new_n8119, new_n8120, new_n8121, new_n8122,
    new_n8123, new_n8124_1, new_n8125, new_n8126, new_n8127, new_n8128,
    new_n8129, new_n8130, new_n8131, new_n8132, new_n8133, new_n8134,
    new_n8136, new_n8137, new_n8138, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144_1, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202, new_n8203, new_n8204_1, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215_1, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8224, new_n8225, new_n8226,
    new_n8227, new_n8228, new_n8229, new_n8230, new_n8231, new_n8232,
    new_n8233, new_n8234, new_n8235, new_n8236, new_n8237, new_n8238,
    new_n8239, new_n8240, new_n8241, new_n8242, new_n8243, new_n8244,
    new_n8245, new_n8246, new_n8247, new_n8248, new_n8249, new_n8250,
    new_n8251, new_n8252, new_n8253, new_n8254, new_n8255, new_n8256,
    new_n8257, new_n8258, new_n8259, new_n8260, new_n8261, new_n8262_1,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302_1, new_n8303, new_n8304,
    new_n8305, new_n8306_1, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8312, new_n8313, new_n8314, new_n8315_1, new_n8316, new_n8317,
    new_n8318, new_n8319, new_n8320, new_n8321, new_n8322, new_n8323,
    new_n8324, new_n8325, new_n8326, new_n8327, new_n8328, new_n8329,
    new_n8330, new_n8331, new_n8332, new_n8333, new_n8334, new_n8335,
    new_n8336, new_n8337, new_n8338, new_n8339, new_n8340, new_n8341,
    new_n8342, new_n8343, new_n8344, new_n8345, new_n8346, new_n8347,
    new_n8348, new_n8349, new_n8350, new_n8351, new_n8352, new_n8353,
    new_n8354, new_n8355, new_n8356, new_n8357, new_n8358, new_n8359,
    new_n8360, new_n8361, new_n8362, new_n8363, new_n8364, new_n8365,
    new_n8366, new_n8367, new_n8368, new_n8369, new_n8370, new_n8371,
    new_n8372, new_n8373, new_n8374, new_n8375, new_n8376, new_n8377,
    new_n8378, new_n8379, new_n8380, new_n8381, new_n8382, new_n8383,
    new_n8384, new_n8385, new_n8386, new_n8387, new_n8388, new_n8389,
    new_n8390, new_n8391, new_n8392, new_n8393, new_n8394, new_n8395,
    new_n8396, new_n8397_1, new_n8398, new_n8399, new_n8400, new_n8401,
    new_n8403, new_n8404, new_n8405, new_n8406, new_n8407, new_n8408,
    new_n8409, new_n8410, new_n8411, new_n8412, new_n8413, new_n8414,
    new_n8415, new_n8416, new_n8417, new_n8418, new_n8419, new_n8420,
    new_n8421, new_n8422, new_n8423, new_n8424, new_n8425, new_n8426,
    new_n8427, new_n8428, new_n8429, new_n8430, new_n8431, new_n8432,
    new_n8433, new_n8434, new_n8435, new_n8436, new_n8437, new_n8438,
    new_n8439_1, new_n8440, new_n8441, new_n8442, new_n8443, new_n8444,
    new_n8445, new_n8446, new_n8447, new_n8448, new_n8449, new_n8450,
    new_n8451, new_n8452, new_n8453, new_n8454, new_n8455, new_n8456,
    new_n8457, new_n8458, new_n8459, new_n8460, new_n8461, new_n8462,
    new_n8463_1, new_n8464, new_n8465, new_n8466, new_n8467, new_n8468,
    new_n8469, new_n8470, new_n8471_1, new_n8472, new_n8473, new_n8474,
    new_n8475, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486_1,
    new_n8487, new_n8488, new_n8489, new_n8491, new_n8492, new_n8493,
    new_n8494, new_n8495, new_n8496, new_n8497, new_n8498, new_n8499,
    new_n8500, new_n8501, new_n8502, new_n8503, new_n8504, new_n8505,
    new_n8506, new_n8507, new_n8508, new_n8509, new_n8510, new_n8511,
    new_n8512, new_n8513, new_n8514, new_n8515, new_n8516, new_n8517,
    new_n8518, new_n8519, new_n8520, new_n8521, new_n8522, new_n8523,
    new_n8524, new_n8525, new_n8526, new_n8527, new_n8528, new_n8529,
    new_n8530, new_n8531, new_n8532, new_n8533, new_n8534, new_n8535,
    new_n8536, new_n8537, new_n8538, new_n8539, new_n8540, new_n8541,
    new_n8542, new_n8543, new_n8544, new_n8545, new_n8546, new_n8547,
    new_n8548, new_n8549, new_n8550_1, new_n8551, new_n8552_1, new_n8553,
    new_n8554, new_n8555, new_n8556, new_n8557, new_n8558, new_n8559,
    new_n8560, new_n8561, new_n8562, new_n8563, new_n8564, new_n8565,
    new_n8566, new_n8567, new_n8568, new_n8569, new_n8570, new_n8571,
    new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577,
    new_n8579, new_n8580, new_n8581, new_n8582, new_n8583, new_n8584,
    new_n8585, new_n8586, new_n8587, new_n8588, new_n8589, new_n8590,
    new_n8591, new_n8592, new_n8593, new_n8594, new_n8595, new_n8596,
    new_n8597, new_n8598_1, new_n8599, new_n8600, new_n8601, new_n8602,
    new_n8603, new_n8604_1, new_n8605, new_n8606, new_n8607, new_n8608,
    new_n8609, new_n8610, new_n8611, new_n8612, new_n8613, new_n8614,
    new_n8615, new_n8616, new_n8617, new_n8618, new_n8619, new_n8620,
    new_n8621, new_n8622, new_n8623, new_n8624, new_n8625, new_n8626,
    new_n8627, new_n8628, new_n8629, new_n8630, new_n8631, new_n8632,
    new_n8633, new_n8634, new_n8635_1, new_n8636, new_n8637, new_n8638,
    new_n8639, new_n8640, new_n8641, new_n8642, new_n8643, new_n8644,
    new_n8645, new_n8646, new_n8647, new_n8648, new_n8649_1, new_n8650,
    new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656,
    new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662,
    new_n8663, new_n8664, new_n8665, new_n8666, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716, new_n8717,
    new_n8718, new_n8719, new_n8720, new_n8721, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737_1, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744, new_n8745, new_n8746_1, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8757, new_n8758, new_n8759, new_n8760,
    new_n8761, new_n8762, new_n8763, new_n8764, new_n8765, new_n8766,
    new_n8767, new_n8768, new_n8769, new_n8770, new_n8771, new_n8772,
    new_n8773, new_n8774, new_n8775, new_n8776, new_n8777, new_n8778,
    new_n8779, new_n8780_1, new_n8781, new_n8782, new_n8783, new_n8784,
    new_n8785, new_n8786, new_n8787, new_n8788, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799_1, new_n8800_1, new_n8801, new_n8802,
    new_n8803, new_n8804, new_n8805, new_n8806, new_n8807, new_n8808,
    new_n8809, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821, new_n8822, new_n8823, new_n8824, new_n8825, new_n8826,
    new_n8827, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8848, new_n8849, new_n8850, new_n8851,
    new_n8852, new_n8853, new_n8854, new_n8855, new_n8856, new_n8857,
    new_n8858, new_n8859, new_n8860, new_n8861, new_n8862, new_n8863,
    new_n8864, new_n8865, new_n8866, new_n8867, new_n8868, new_n8869,
    new_n8870, new_n8871, new_n8872, new_n8873_1, new_n8874, new_n8875,
    new_n8876, new_n8877, new_n8878, new_n8879, new_n8880, new_n8881,
    new_n8882, new_n8883, new_n8884, new_n8885, new_n8886, new_n8887,
    new_n8888, new_n8889, new_n8890, new_n8891, new_n8892_1, new_n8893,
    new_n8894, new_n8895, new_n8896, new_n8897, new_n8898, new_n8899,
    new_n8900, new_n8901, new_n8902, new_n8903, new_n8904, new_n8905,
    new_n8906, new_n8907, new_n8908, new_n8909_1, new_n8910, new_n8911,
    new_n8912, new_n8913, new_n8914, new_n8915, new_n8916, new_n8917,
    new_n8918, new_n8919, new_n8920, new_n8921, new_n8922, new_n8923,
    new_n8924, new_n8925, new_n8926_1, new_n8927, new_n8928, new_n8929,
    new_n8930, new_n8931, new_n8932, new_n8933, new_n8934, new_n8936,
    new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942,
    new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948,
    new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954,
    new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997_1, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9024, new_n9025, new_n9026_1, new_n9027,
    new_n9028, new_n9029, new_n9030, new_n9031, new_n9032, new_n9033,
    new_n9034, new_n9035, new_n9036, new_n9037, new_n9038, new_n9039,
    new_n9040, new_n9041, new_n9042, new_n9043, new_n9044, new_n9045,
    new_n9046, new_n9047, new_n9048, new_n9049, new_n9050, new_n9051,
    new_n9052, new_n9053, new_n9054, new_n9055, new_n9056, new_n9057,
    new_n9058, new_n9059, new_n9060, new_n9061, new_n9062, new_n9063,
    new_n9064, new_n9065, new_n9066, new_n9067, new_n9068, new_n9069,
    new_n9070, new_n9071, new_n9072, new_n9073, new_n9074, new_n9075,
    new_n9076, new_n9077, new_n9078, new_n9079, new_n9080, new_n9081,
    new_n9082, new_n9083, new_n9084, new_n9085, new_n9086, new_n9087,
    new_n9088, new_n9089, new_n9090, new_n9091, new_n9092, new_n9093,
    new_n9094, new_n9095, new_n9096_1, new_n9097, new_n9098, new_n9099,
    new_n9100, new_n9101, new_n9102, new_n9103, new_n9104, new_n9105,
    new_n9106, new_n9107, new_n9108, new_n9109, new_n9110_1, new_n9112,
    new_n9113, new_n9114, new_n9115, new_n9116, new_n9117, new_n9118,
    new_n9119, new_n9120, new_n9121, new_n9122, new_n9123, new_n9124,
    new_n9125, new_n9126, new_n9127, new_n9128, new_n9129, new_n9130,
    new_n9131, new_n9132, new_n9133, new_n9134, new_n9135, new_n9136,
    new_n9137, new_n9138, new_n9139, new_n9140, new_n9141, new_n9142,
    new_n9143, new_n9144, new_n9145, new_n9146, new_n9147, new_n9148,
    new_n9149, new_n9150, new_n9151, new_n9152, new_n9153, new_n9154_1,
    new_n9155, new_n9156, new_n9157, new_n9158, new_n9159, new_n9160,
    new_n9161, new_n9162, new_n9163, new_n9164, new_n9165, new_n9166,
    new_n9167, new_n9168, new_n9169, new_n9170, new_n9171, new_n9172,
    new_n9173, new_n9174, new_n9175, new_n9176, new_n9177, new_n9178,
    new_n9179, new_n9180, new_n9181, new_n9182, new_n9183, new_n9184,
    new_n9185, new_n9186_1, new_n9187, new_n9188, new_n9189, new_n9190,
    new_n9191, new_n9192, new_n9193, new_n9194, new_n9195, new_n9196,
    new_n9197, new_n9198, new_n9199, new_n9201, new_n9202, new_n9203,
    new_n9204, new_n9205, new_n9206, new_n9207, new_n9208, new_n9209,
    new_n9210, new_n9211, new_n9212, new_n9213, new_n9214, new_n9215,
    new_n9216, new_n9217, new_n9218, new_n9219, new_n9220, new_n9221,
    new_n9222, new_n9223, new_n9224, new_n9225, new_n9226, new_n9227,
    new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233,
    new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239,
    new_n9240, new_n9241, new_n9242, new_n9243, new_n9244, new_n9245,
    new_n9246, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251,
    new_n9252_1, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259, new_n9260, new_n9261, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287,
    new_n9288, new_n9289, new_n9291, new_n9292, new_n9293, new_n9294,
    new_n9295, new_n9296, new_n9297, new_n9298, new_n9299, new_n9300,
    new_n9301, new_n9302, new_n9303, new_n9304, new_n9305, new_n9306,
    new_n9307, new_n9308, new_n9309, new_n9310, new_n9311, new_n9312,
    new_n9313, new_n9314_1, new_n9315, new_n9316, new_n9317, new_n9318,
    new_n9319, new_n9320, new_n9321, new_n9322, new_n9323, new_n9324,
    new_n9325, new_n9326, new_n9327, new_n9328, new_n9329, new_n9330,
    new_n9331, new_n9332, new_n9333, new_n9334, new_n9335, new_n9336,
    new_n9337, new_n9338, new_n9339, new_n9340, new_n9341, new_n9342_1,
    new_n9343, new_n9344, new_n9345, new_n9346, new_n9347, new_n9348,
    new_n9349, new_n9350, new_n9351, new_n9352, new_n9353, new_n9354,
    new_n9355, new_n9356, new_n9357, new_n9358, new_n9359, new_n9360,
    new_n9361, new_n9362, new_n9363, new_n9364, new_n9365, new_n9366,
    new_n9367, new_n9368, new_n9369, new_n9370, new_n9371, new_n9372,
    new_n9373, new_n9374, new_n9375, new_n9376, new_n9377, new_n9378,
    new_n9379, new_n9381, new_n9382, new_n9383, new_n9384, new_n9385,
    new_n9386, new_n9387, new_n9388, new_n9389, new_n9390, new_n9391,
    new_n9392, new_n9393, new_n9394, new_n9395, new_n9396, new_n9397,
    new_n9398, new_n9399, new_n9400, new_n9401, new_n9402, new_n9403,
    new_n9404, new_n9405, new_n9406, new_n9407, new_n9408, new_n9409,
    new_n9410, new_n9411, new_n9412, new_n9413, new_n9414, new_n9415,
    new_n9416, new_n9417, new_n9418, new_n9419, new_n9420, new_n9421,
    new_n9422, new_n9423, new_n9424, new_n9425, new_n9426, new_n9427,
    new_n9428, new_n9429, new_n9430, new_n9431, new_n9432, new_n9433,
    new_n9434, new_n9435, new_n9436, new_n9437_1, new_n9438, new_n9439,
    new_n9440, new_n9441, new_n9442, new_n9443, new_n9444, new_n9445,
    new_n9446, new_n9447_1, new_n9448, new_n9449, new_n9450, new_n9451,
    new_n9452, new_n9453, new_n9454, new_n9455, new_n9456, new_n9457,
    new_n9458, new_n9459, new_n9460, new_n9461, new_n9462, new_n9463,
    new_n9464, new_n9465, new_n9466, new_n9467, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507, new_n9508, new_n9509, new_n9510, new_n9511, new_n9512,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543_1, new_n9544_1, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552, new_n9553, new_n9554,
    new_n9555_1, new_n9556, new_n9558, new_n9559, new_n9560, new_n9561,
    new_n9562, new_n9563, new_n9564, new_n9565, new_n9566, new_n9567,
    new_n9568, new_n9569, new_n9570_1, new_n9571, new_n9572, new_n9573,
    new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579,
    new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585,
    new_n9586, new_n9587, new_n9588, new_n9589_1, new_n9590, new_n9591,
    new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597,
    new_n9598, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603,
    new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609,
    new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615,
    new_n9616, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621,
    new_n9622, new_n9623, new_n9624, new_n9625, new_n9626, new_n9627,
    new_n9628, new_n9629, new_n9630, new_n9631, new_n9632, new_n9633,
    new_n9634, new_n9635, new_n9636, new_n9637, new_n9638, new_n9639,
    new_n9640, new_n9641, new_n9642, new_n9643, new_n9644, new_n9646,
    new_n9647, new_n9648, new_n9649, new_n9650, new_n9651, new_n9652,
    new_n9653, new_n9654, new_n9655, new_n9656, new_n9657, new_n9658,
    new_n9659, new_n9660, new_n9661, new_n9662, new_n9663, new_n9664,
    new_n9665_1, new_n9666, new_n9667, new_n9668, new_n9669, new_n9670,
    new_n9671, new_n9672, new_n9673, new_n9674, new_n9675, new_n9676,
    new_n9677, new_n9678, new_n9679, new_n9680, new_n9681, new_n9682,
    new_n9683, new_n9684, new_n9685, new_n9686, new_n9687, new_n9688,
    new_n9689, new_n9690, new_n9691, new_n9692, new_n9693, new_n9694,
    new_n9695, new_n9696, new_n9697, new_n9698, new_n9699, new_n9700,
    new_n9701, new_n9702, new_n9703, new_n9704, new_n9705, new_n9706,
    new_n9707, new_n9708, new_n9709, new_n9710, new_n9711, new_n9712,
    new_n9713, new_n9714, new_n9715, new_n9716, new_n9717_1, new_n9718,
    new_n9719, new_n9720, new_n9721, new_n9722, new_n9723, new_n9724,
    new_n9725, new_n9726, new_n9727, new_n9728, new_n9729, new_n9730,
    new_n9731, new_n9732, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763, new_n9764, new_n9765, new_n9766, new_n9767,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820, new_n9822,
    new_n9823, new_n9824, new_n9825, new_n9826, new_n9827, new_n9828,
    new_n9829, new_n9830_1, new_n9831, new_n9832, new_n9833, new_n9834,
    new_n9835, new_n9836, new_n9837, new_n9838, new_n9839, new_n9840,
    new_n9841, new_n9842, new_n9843, new_n9844, new_n9845, new_n9846,
    new_n9847, new_n9848, new_n9849, new_n9850, new_n9851, new_n9852,
    new_n9853, new_n9854, new_n9855, new_n9856, new_n9857, new_n9858,
    new_n9859, new_n9860, new_n9861, new_n9862, new_n9863, new_n9864,
    new_n9865, new_n9866, new_n9867, new_n9868, new_n9869, new_n9870,
    new_n9871, new_n9872, new_n9873, new_n9874, new_n9875, new_n9876,
    new_n9877, new_n9878, new_n9879, new_n9880, new_n9881, new_n9882,
    new_n9883, new_n9884, new_n9885, new_n9886, new_n9887, new_n9888,
    new_n9889, new_n9890, new_n9891, new_n9892, new_n9893_1, new_n9894,
    new_n9895, new_n9896, new_n9897, new_n9898, new_n9899, new_n9900,
    new_n9901, new_n9902, new_n9903, new_n9904, new_n9905, new_n9906,
    new_n9907, new_n9908, new_n9910, new_n9911, new_n9912, new_n9913,
    new_n9914, new_n9915, new_n9916, new_n9917, new_n9918, new_n9919,
    new_n9920, new_n9921_1, new_n9922, new_n9923, new_n9924, new_n9925,
    new_n9926, new_n9927, new_n9928, new_n9929, new_n9930, new_n9931,
    new_n9932, new_n9933, new_n9934, new_n9935, new_n9936_1, new_n9937,
    new_n9938, new_n9939, new_n9940, new_n9941, new_n9942, new_n9943,
    new_n9944, new_n9945, new_n9946, new_n9947, new_n9948, new_n9949,
    new_n9950, new_n9951, new_n9952, new_n9953, new_n9954, new_n9955,
    new_n9956, new_n9957, new_n9958, new_n9959, new_n9960, new_n9961,
    new_n9962, new_n9963, new_n9964, new_n9965, new_n9966, new_n9967,
    new_n9968, new_n9969, new_n9970, new_n9971, new_n9972, new_n9973,
    new_n9974, new_n9975, new_n9976, new_n9977_1, new_n9978, new_n9979,
    new_n9980, new_n9981, new_n9982, new_n9983, new_n9984, new_n9985,
    new_n9986, new_n9987, new_n9988, new_n9989, new_n9990, new_n9991,
    new_n9992, new_n9993, new_n9994, new_n9995, new_n9996, new_n9998,
    new_n9999, new_n10000, new_n10001, new_n10002, new_n10003, new_n10004,
    new_n10005, new_n10006, new_n10007, new_n10008, new_n10009, new_n10010,
    new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017, new_n10018, new_n10019, new_n10020, new_n10021, new_n10022,
    new_n10023, new_n10024, new_n10025, new_n10026, new_n10027, new_n10028,
    new_n10029, new_n10030, new_n10031, new_n10032, new_n10033, new_n10034,
    new_n10035, new_n10036, new_n10037, new_n10038, new_n10039, new_n10040,
    new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046,
    new_n10047, new_n10048, new_n10049, new_n10050_1, new_n10051_1,
    new_n10052, new_n10053, new_n10054, new_n10055, new_n10056, new_n10057,
    new_n10058, new_n10059, new_n10060, new_n10061_1, new_n10062,
    new_n10063, new_n10064, new_n10065, new_n10066, new_n10067, new_n10068,
    new_n10069, new_n10070, new_n10071, new_n10072, new_n10073, new_n10074,
    new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080_1, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096, new_n10097,
    new_n10098, new_n10099, new_n10100, new_n10101, new_n10102, new_n10103,
    new_n10104, new_n10105, new_n10106, new_n10107, new_n10108, new_n10109,
    new_n10110, new_n10111, new_n10112_1, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147_1, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158, new_n10159, new_n10160, new_n10161,
    new_n10162, new_n10163, new_n10164, new_n10165, new_n10166, new_n10167,
    new_n10168, new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174, new_n10176, new_n10177, new_n10178, new_n10179, new_n10180,
    new_n10181, new_n10182, new_n10183, new_n10184, new_n10185, new_n10186,
    new_n10187, new_n10188, new_n10189, new_n10190, new_n10191, new_n10192,
    new_n10193, new_n10194, new_n10195, new_n10196, new_n10197, new_n10198,
    new_n10199, new_n10200, new_n10201, new_n10202, new_n10203, new_n10204,
    new_n10205, new_n10206, new_n10207, new_n10208, new_n10209, new_n10210,
    new_n10211, new_n10212, new_n10213, new_n10214, new_n10215, new_n10216,
    new_n10217, new_n10218, new_n10219, new_n10220, new_n10221, new_n10222,
    new_n10223, new_n10224, new_n10225, new_n10226, new_n10227, new_n10228,
    new_n10229, new_n10230, new_n10231, new_n10232, new_n10233, new_n10234,
    new_n10235, new_n10236, new_n10237, new_n10238, new_n10239, new_n10240,
    new_n10241, new_n10242, new_n10243, new_n10244, new_n10245, new_n10246,
    new_n10247, new_n10248, new_n10249, new_n10250, new_n10251, new_n10252,
    new_n10253, new_n10254, new_n10255_1, new_n10256, new_n10257,
    new_n10258, new_n10259, new_n10260, new_n10261, new_n10262, new_n10264,
    new_n10265, new_n10266, new_n10267, new_n10268, new_n10269, new_n10270,
    new_n10271, new_n10272, new_n10273, new_n10274, new_n10275, new_n10276,
    new_n10277, new_n10278_1, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283_1, new_n10284, new_n10285, new_n10286,
    new_n10287, new_n10288, new_n10289, new_n10290, new_n10291, new_n10292,
    new_n10293, new_n10294, new_n10295, new_n10296, new_n10297, new_n10298,
    new_n10299, new_n10300, new_n10301, new_n10302, new_n10303, new_n10304,
    new_n10305, new_n10306, new_n10307, new_n10308, new_n10309, new_n10310,
    new_n10311, new_n10312, new_n10313, new_n10314, new_n10315, new_n10316,
    new_n10317, new_n10318, new_n10319, new_n10320, new_n10321, new_n10322,
    new_n10323, new_n10324, new_n10325, new_n10326, new_n10327, new_n10328,
    new_n10329, new_n10330, new_n10331, new_n10332, new_n10333, new_n10334,
    new_n10335, new_n10336, new_n10337, new_n10338, new_n10339, new_n10340,
    new_n10341, new_n10342, new_n10343, new_n10344, new_n10345, new_n10346,
    new_n10347, new_n10348, new_n10349, new_n10350, new_n10352, new_n10353,
    new_n10354, new_n10355, new_n10356, new_n10357, new_n10358, new_n10359,
    new_n10360, new_n10361, new_n10362, new_n10363, new_n10364, new_n10365,
    new_n10366, new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372, new_n10373, new_n10374, new_n10375, new_n10376, new_n10377,
    new_n10378_1, new_n10379, new_n10380, new_n10381, new_n10382,
    new_n10383, new_n10384, new_n10385, new_n10386, new_n10387, new_n10388,
    new_n10389, new_n10390, new_n10391, new_n10392, new_n10393, new_n10394,
    new_n10395, new_n10396, new_n10397, new_n10398, new_n10399, new_n10400,
    new_n10401, new_n10402, new_n10403, new_n10404, new_n10405, new_n10406,
    new_n10407_1, new_n10408, new_n10409, new_n10410, new_n10411,
    new_n10412, new_n10413, new_n10414, new_n10415, new_n10416, new_n10417,
    new_n10418, new_n10419, new_n10420, new_n10421, new_n10422, new_n10423,
    new_n10424, new_n10425, new_n10426_1, new_n10427, new_n10428,
    new_n10429, new_n10430, new_n10431, new_n10432, new_n10433, new_n10434,
    new_n10435, new_n10436, new_n10437, new_n10438, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446_1,
    new_n10447, new_n10448, new_n10449, new_n10450, new_n10451, new_n10452,
    new_n10453, new_n10454, new_n10455, new_n10456, new_n10457, new_n10458,
    new_n10459, new_n10460, new_n10461, new_n10462, new_n10463, new_n10464,
    new_n10465, new_n10466_1, new_n10467, new_n10468, new_n10469,
    new_n10470_1, new_n10471, new_n10472, new_n10473, new_n10474,
    new_n10475, new_n10476, new_n10477, new_n10478, new_n10479, new_n10480,
    new_n10481, new_n10482, new_n10483, new_n10484, new_n10485, new_n10486,
    new_n10487, new_n10488, new_n10489, new_n10490, new_n10491, new_n10492,
    new_n10493, new_n10494, new_n10495, new_n10496, new_n10497, new_n10498,
    new_n10499, new_n10500, new_n10501, new_n10502, new_n10503, new_n10504,
    new_n10505, new_n10506, new_n10507, new_n10508, new_n10509, new_n10510,
    new_n10511, new_n10512, new_n10513, new_n10514, new_n10515_1,
    new_n10516, new_n10517, new_n10518, new_n10519, new_n10520, new_n10521,
    new_n10522, new_n10523, new_n10524, new_n10525, new_n10526, new_n10528,
    new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534,
    new_n10535, new_n10536, new_n10537, new_n10538, new_n10539, new_n10540,
    new_n10541, new_n10542, new_n10543, new_n10544, new_n10545, new_n10546,
    new_n10547, new_n10548, new_n10549, new_n10550, new_n10551, new_n10552,
    new_n10553, new_n10554, new_n10555, new_n10556, new_n10557, new_n10558,
    new_n10559, new_n10560, new_n10561, new_n10562, new_n10563, new_n10564,
    new_n10565, new_n10566, new_n10567, new_n10568, new_n10569, new_n10570,
    new_n10571, new_n10572, new_n10573_1, new_n10574, new_n10575,
    new_n10576, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588, new_n10589, new_n10590, new_n10591_1, new_n10592,
    new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611, new_n10612, new_n10613, new_n10614, new_n10616, new_n10617,
    new_n10618, new_n10619, new_n10620, new_n10621, new_n10622, new_n10623,
    new_n10624, new_n10625, new_n10626, new_n10627, new_n10628, new_n10629,
    new_n10630_1, new_n10631, new_n10632, new_n10633, new_n10634,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644, new_n10645, new_n10646,
    new_n10647, new_n10648, new_n10649, new_n10650, new_n10651, new_n10652,
    new_n10653, new_n10654, new_n10655, new_n10656, new_n10657, new_n10658,
    new_n10659, new_n10660, new_n10661, new_n10662, new_n10663, new_n10664,
    new_n10665, new_n10666, new_n10667, new_n10668, new_n10669, new_n10670,
    new_n10671, new_n10672, new_n10673, new_n10674, new_n10675, new_n10676,
    new_n10677, new_n10678, new_n10679, new_n10680, new_n10681, new_n10682,
    new_n10683, new_n10684, new_n10685, new_n10686, new_n10687, new_n10688,
    new_n10689, new_n10690, new_n10691, new_n10692, new_n10693, new_n10694,
    new_n10695, new_n10696, new_n10697, new_n10698, new_n10699, new_n10700,
    new_n10701, new_n10702, new_n10703, new_n10705, new_n10706, new_n10707,
    new_n10708, new_n10709, new_n10710, new_n10711, new_n10712, new_n10713,
    new_n10714, new_n10715, new_n10716, new_n10717, new_n10718, new_n10719,
    new_n10720, new_n10721, new_n10722, new_n10723, new_n10724, new_n10725,
    new_n10726, new_n10727, new_n10728, new_n10729, new_n10730, new_n10731,
    new_n10732, new_n10733, new_n10734, new_n10735, new_n10736_1,
    new_n10737, new_n10738, new_n10739, new_n10740, new_n10741, new_n10742,
    new_n10743, new_n10744, new_n10745, new_n10746, new_n10747, new_n10748,
    new_n10749, new_n10750_1, new_n10751, new_n10752, new_n10753,
    new_n10754, new_n10755, new_n10756, new_n10757, new_n10758, new_n10759,
    new_n10760, new_n10761, new_n10762, new_n10763, new_n10764,
    new_n10765_1, new_n10766, new_n10767, new_n10768, new_n10769,
    new_n10770, new_n10771, new_n10772, new_n10773, new_n10774, new_n10775,
    new_n10776, new_n10777, new_n10778, new_n10779, new_n10780, new_n10781,
    new_n10782, new_n10783, new_n10784, new_n10785, new_n10786, new_n10787,
    new_n10788, new_n10789, new_n10790, new_n10791_1, new_n10792,
    new_n10794, new_n10795, new_n10796, new_n10797, new_n10798, new_n10799,
    new_n10800, new_n10801, new_n10802_1, new_n10803, new_n10804,
    new_n10805, new_n10806, new_n10807, new_n10808, new_n10809, new_n10810,
    new_n10811, new_n10812, new_n10813, new_n10814, new_n10815, new_n10816,
    new_n10817, new_n10818, new_n10819, new_n10820, new_n10821, new_n10822,
    new_n10823, new_n10824, new_n10825, new_n10826, new_n10827, new_n10828,
    new_n10829, new_n10830, new_n10831, new_n10832, new_n10833, new_n10834,
    new_n10835, new_n10836, new_n10837, new_n10838, new_n10839, new_n10840,
    new_n10841, new_n10842, new_n10843, new_n10844, new_n10845, new_n10846,
    new_n10847, new_n10848, new_n10849, new_n10850, new_n10851, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862_1, new_n10863,
    new_n10864, new_n10865, new_n10866, new_n10867, new_n10868, new_n10869,
    new_n10870, new_n10871, new_n10872, new_n10873, new_n10874, new_n10875,
    new_n10876, new_n10877, new_n10878, new_n10879, new_n10880, new_n10881,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911,
    new_n10912_1, new_n10913, new_n10914, new_n10915_1, new_n10916,
    new_n10917, new_n10918, new_n10919, new_n10920, new_n10921, new_n10922,
    new_n10923, new_n10924, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943, new_n10944, new_n10945_1,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961, new_n10962, new_n10963,
    new_n10964, new_n10965, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10971, new_n10972, new_n10973, new_n10974, new_n10975, new_n10976,
    new_n10977, new_n10978, new_n10979, new_n10980, new_n10981, new_n10982,
    new_n10983, new_n10984, new_n10985, new_n10986, new_n10987, new_n10988,
    new_n10989, new_n10990, new_n10991, new_n10992, new_n10993, new_n10994,
    new_n10995, new_n10996, new_n10997, new_n10998, new_n10999, new_n11000,
    new_n11001, new_n11002, new_n11003, new_n11004, new_n11005, new_n11006,
    new_n11007, new_n11008, new_n11009, new_n11010, new_n11011, new_n11012,
    new_n11013, new_n11014, new_n11015, new_n11016, new_n11017, new_n11018,
    new_n11019, new_n11020, new_n11021, new_n11022, new_n11023, new_n11024,
    new_n11025, new_n11026, new_n11027, new_n11028, new_n11029, new_n11030,
    new_n11031, new_n11032, new_n11033, new_n11034, new_n11035, new_n11036,
    new_n11037, new_n11038, new_n11039, new_n11040, new_n11041, new_n11042,
    new_n11043, new_n11044, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056, new_n11057, new_n11059, new_n11060, new_n11061,
    new_n11062, new_n11063, new_n11064, new_n11065, new_n11066, new_n11067,
    new_n11068, new_n11069, new_n11070, new_n11071, new_n11072, new_n11073,
    new_n11074, new_n11075, new_n11076, new_n11077, new_n11078, new_n11079,
    new_n11080, new_n11081, new_n11082, new_n11083, new_n11084, new_n11085,
    new_n11086, new_n11087, new_n11088, new_n11089, new_n11090, new_n11091,
    new_n11092, new_n11093, new_n11094, new_n11095, new_n11096, new_n11097,
    new_n11098, new_n11099, new_n11100, new_n11101, new_n11102, new_n11103,
    new_n11104, new_n11105, new_n11106, new_n11107, new_n11108, new_n11109,
    new_n11110, new_n11111, new_n11112, new_n11113, new_n11114, new_n11115,
    new_n11116, new_n11117, new_n11118, new_n11119, new_n11120, new_n11121,
    new_n11122_1, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143_1,
    new_n11144, new_n11145, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156,
    new_n11157, new_n11158_1, new_n11159, new_n11160, new_n11161,
    new_n11162, new_n11163, new_n11164, new_n11165, new_n11166, new_n11167,
    new_n11168, new_n11169, new_n11170, new_n11171, new_n11172, new_n11173,
    new_n11174, new_n11175, new_n11176, new_n11177, new_n11178, new_n11179,
    new_n11180, new_n11181, new_n11182, new_n11183, new_n11184, new_n11185,
    new_n11186, new_n11187, new_n11188, new_n11189, new_n11190, new_n11191,
    new_n11192, new_n11193, new_n11194, new_n11195, new_n11196, new_n11197,
    new_n11198, new_n11199, new_n11200, new_n11201, new_n11202, new_n11203,
    new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209,
    new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215,
    new_n11216, new_n11217, new_n11218, new_n11219, new_n11220, new_n11221,
    new_n11222, new_n11223, new_n11224, new_n11225, new_n11226, new_n11227,
    new_n11228, new_n11229, new_n11230, new_n11231, new_n11232, new_n11233,
    new_n11235, new_n11236, new_n11237, new_n11238, new_n11239, new_n11240,
    new_n11241, new_n11242, new_n11243, new_n11244, new_n11245, new_n11246,
    new_n11247, new_n11248, new_n11249, new_n11250, new_n11251, new_n11252,
    new_n11253, new_n11254, new_n11255, new_n11256, new_n11257, new_n11258,
    new_n11259, new_n11260, new_n11261, new_n11262, new_n11263, new_n11264,
    new_n11265, new_n11266, new_n11267, new_n11268, new_n11269_1,
    new_n11270, new_n11271, new_n11272, new_n11273, new_n11274, new_n11275,
    new_n11276, new_n11277, new_n11278, new_n11279, new_n11280, new_n11281,
    new_n11282, new_n11283, new_n11284, new_n11285, new_n11286, new_n11287,
    new_n11288, new_n11289, new_n11290, new_n11291, new_n11292, new_n11293,
    new_n11294, new_n11295, new_n11296, new_n11297, new_n11298, new_n11299,
    new_n11300, new_n11301, new_n11302, new_n11303, new_n11304, new_n11305,
    new_n11306, new_n11307, new_n11308, new_n11309, new_n11310, new_n11311,
    new_n11312, new_n11313, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11323, new_n11324,
    new_n11325, new_n11326, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345_1, new_n11346, new_n11347,
    new_n11348, new_n11349, new_n11350, new_n11351, new_n11352, new_n11353,
    new_n11354, new_n11355, new_n11356, new_n11357, new_n11358, new_n11359,
    new_n11360, new_n11361, new_n11362, new_n11363, new_n11364, new_n11365,
    new_n11366, new_n11367, new_n11368, new_n11369, new_n11370, new_n11371,
    new_n11372, new_n11373, new_n11374, new_n11375, new_n11376, new_n11377,
    new_n11378, new_n11379, new_n11380, new_n11381, new_n11382, new_n11383,
    new_n11384, new_n11385, new_n11386, new_n11387, new_n11388, new_n11389,
    new_n11390, new_n11391, new_n11392, new_n11393_1, new_n11394,
    new_n11395, new_n11396, new_n11397, new_n11398, new_n11399, new_n11400,
    new_n11401, new_n11402, new_n11403, new_n11404_1, new_n11405,
    new_n11406, new_n11407, new_n11408, new_n11409, new_n11410, new_n11412,
    new_n11413, new_n11414, new_n11415, new_n11416, new_n11417, new_n11418,
    new_n11419, new_n11420, new_n11421, new_n11422, new_n11423, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463_1, new_n11464, new_n11465,
    new_n11466, new_n11467, new_n11468, new_n11469, new_n11470, new_n11471,
    new_n11472, new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478, new_n11479, new_n11480, new_n11481, new_n11482, new_n11483,
    new_n11484, new_n11485, new_n11486, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496, new_n11497, new_n11498, new_n11500, new_n11501, new_n11502,
    new_n11503, new_n11504, new_n11505, new_n11506, new_n11507, new_n11508,
    new_n11509, new_n11510, new_n11511, new_n11512, new_n11513, new_n11514,
    new_n11515, new_n11516, new_n11517, new_n11518, new_n11519, new_n11520,
    new_n11521, new_n11522, new_n11523, new_n11524, new_n11525, new_n11526,
    new_n11527, new_n11528, new_n11529_1, new_n11530, new_n11531,
    new_n11532, new_n11533, new_n11534_1, new_n11535, new_n11536,
    new_n11537, new_n11538, new_n11539, new_n11540, new_n11541, new_n11542,
    new_n11543, new_n11544, new_n11545, new_n11546, new_n11547, new_n11548,
    new_n11549, new_n11550, new_n11551, new_n11552, new_n11553, new_n11554,
    new_n11555, new_n11556, new_n11557, new_n11558, new_n11559, new_n11560,
    new_n11561, new_n11562, new_n11563, new_n11564, new_n11565, new_n11566,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579, new_n11580, new_n11581, new_n11582, new_n11583, new_n11584,
    new_n11585, new_n11586, new_n11588, new_n11589, new_n11590_1,
    new_n11591, new_n11592, new_n11593, new_n11594, new_n11595, new_n11596,
    new_n11597, new_n11598, new_n11599, new_n11600, new_n11601, new_n11602,
    new_n11603, new_n11604, new_n11605_1, new_n11606, new_n11607,
    new_n11608, new_n11609, new_n11610, new_n11611, new_n11612, new_n11613,
    new_n11614, new_n11615, new_n11616, new_n11617, new_n11618, new_n11619,
    new_n11620, new_n11621, new_n11622, new_n11623, new_n11624, new_n11625,
    new_n11626, new_n11627_1, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662, new_n11663, new_n11664_1, new_n11665,
    new_n11666_1, new_n11667, new_n11668, new_n11669, new_n11670,
    new_n11671, new_n11672, new_n11673, new_n11674, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706, new_n11707,
    new_n11708, new_n11709, new_n11710, new_n11711, new_n11712, new_n11713,
    new_n11714, new_n11715, new_n11716, new_n11717, new_n11718, new_n11719,
    new_n11720, new_n11721, new_n11722, new_n11723, new_n11724, new_n11725,
    new_n11726, new_n11727, new_n11728, new_n11729, new_n11730, new_n11731,
    new_n11732, new_n11733, new_n11734, new_n11735, new_n11736, new_n11737,
    new_n11738, new_n11739, new_n11740, new_n11741, new_n11742, new_n11743,
    new_n11744, new_n11745, new_n11746, new_n11747, new_n11748, new_n11749,
    new_n11750, new_n11751, new_n11752, new_n11753, new_n11754, new_n11755,
    new_n11756_1, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11764, new_n11765, new_n11766, new_n11767,
    new_n11768, new_n11769, new_n11770, new_n11771, new_n11772, new_n11773,
    new_n11774, new_n11775, new_n11776_1, new_n11777, new_n11778,
    new_n11779, new_n11780, new_n11781, new_n11782, new_n11783, new_n11784,
    new_n11785, new_n11786, new_n11787, new_n11788, new_n11789, new_n11790,
    new_n11791, new_n11792, new_n11793, new_n11794, new_n11795, new_n11796,
    new_n11797, new_n11798, new_n11799, new_n11800, new_n11801, new_n11802,
    new_n11803, new_n11804, new_n11805, new_n11806, new_n11807, new_n11808,
    new_n11809, new_n11810, new_n11811, new_n11812, new_n11813, new_n11814,
    new_n11815, new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821, new_n11822_1, new_n11823, new_n11824, new_n11825,
    new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831,
    new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837,
    new_n11838, new_n11839, new_n11840, new_n11841, new_n11842_1,
    new_n11843, new_n11844, new_n11845, new_n11846, new_n11847_1,
    new_n11848, new_n11849, new_n11850, new_n11852, new_n11853,
    new_n11854_1, new_n11855, new_n11856, new_n11857, new_n11858,
    new_n11859, new_n11860, new_n11861, new_n11862, new_n11863, new_n11864,
    new_n11865, new_n11866, new_n11867, new_n11868, new_n11869, new_n11870,
    new_n11871, new_n11872, new_n11873, new_n11874, new_n11875_1,
    new_n11876, new_n11877, new_n11878, new_n11879, new_n11880, new_n11881,
    new_n11882, new_n11883, new_n11884, new_n11885, new_n11886, new_n11887,
    new_n11888, new_n11889, new_n11890, new_n11891, new_n11892, new_n11893,
    new_n11894, new_n11895, new_n11896, new_n11897, new_n11898, new_n11899,
    new_n11900, new_n11901, new_n11902_1, new_n11903, new_n11904,
    new_n11905, new_n11906, new_n11907, new_n11908, new_n11909, new_n11910,
    new_n11911, new_n11912, new_n11913, new_n11914, new_n11915, new_n11916,
    new_n11917, new_n11918, new_n11919, new_n11920, new_n11921, new_n11922,
    new_n11923, new_n11924, new_n11925, new_n11926, new_n11927, new_n11928,
    new_n11929, new_n11930_1, new_n11931, new_n11932, new_n11933_1,
    new_n11934, new_n11935, new_n11936, new_n11937, new_n11938, new_n11939,
    new_n11940, new_n11942, new_n11943, new_n11944, new_n11945, new_n11946,
    new_n11947, new_n11948, new_n11949, new_n11950, new_n11951, new_n11952,
    new_n11953, new_n11954, new_n11955, new_n11956, new_n11957, new_n11958,
    new_n11959, new_n11960, new_n11961_1, new_n11962, new_n11963,
    new_n11964, new_n11965, new_n11966, new_n11967, new_n11968, new_n11969,
    new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975,
    new_n11976, new_n11977, new_n11978, new_n11979, new_n11980, new_n11981,
    new_n11982, new_n11983, new_n11984, new_n11985, new_n11986, new_n11987,
    new_n11988, new_n11989, new_n11990, new_n11991, new_n11992, new_n11993,
    new_n11994, new_n11995, new_n11996, new_n11997, new_n11998, new_n11999,
    new_n12000, new_n12001, new_n12002, new_n12003, new_n12004, new_n12005,
    new_n12006, new_n12007, new_n12008, new_n12009_1, new_n12010,
    new_n12011, new_n12012_1, new_n12013, new_n12014, new_n12015,
    new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021,
    new_n12022, new_n12023, new_n12024, new_n12025_1, new_n12026,
    new_n12027, new_n12028, new_n12030, new_n12031, new_n12032_1,
    new_n12033, new_n12034, new_n12035, new_n12036, new_n12037, new_n12038,
    new_n12039, new_n12040, new_n12041, new_n12042, new_n12043, new_n12044,
    new_n12045, new_n12046, new_n12047, new_n12048, new_n12049, new_n12050,
    new_n12051, new_n12052, new_n12053, new_n12054, new_n12055, new_n12056,
    new_n12057, new_n12058, new_n12059, new_n12060, new_n12061, new_n12062,
    new_n12063, new_n12064, new_n12065, new_n12066, new_n12067, new_n12068,
    new_n12069, new_n12070, new_n12071, new_n12072, new_n12073, new_n12074,
    new_n12075, new_n12076, new_n12077, new_n12078, new_n12079, new_n12080,
    new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086,
    new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092,
    new_n12093, new_n12094, new_n12095, new_n12096, new_n12097, new_n12098,
    new_n12099, new_n12100, new_n12101, new_n12102, new_n12103, new_n12104,
    new_n12105, new_n12106, new_n12107, new_n12108, new_n12109, new_n12110,
    new_n12111, new_n12112, new_n12113, new_n12114, new_n12115, new_n12116,
    new_n12118, new_n12119, new_n12120, new_n12121, new_n12122, new_n12123,
    new_n12124, new_n12125, new_n12126, new_n12127, new_n12128, new_n12129,
    new_n12130, new_n12131, new_n12132, new_n12133, new_n12134, new_n12135,
    new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141,
    new_n12142_1, new_n12143, new_n12144, new_n12145, new_n12146,
    new_n12147, new_n12148, new_n12149, new_n12150, new_n12151, new_n12152,
    new_n12153, new_n12154, new_n12155, new_n12156, new_n12157, new_n12158,
    new_n12159, new_n12160, new_n12161, new_n12162, new_n12163, new_n12164,
    new_n12165, new_n12166_1, new_n12167, new_n12168, new_n12169,
    new_n12170, new_n12171, new_n12172, new_n12173, new_n12174, new_n12175,
    new_n12176, new_n12177, new_n12178, new_n12179, new_n12180, new_n12181,
    new_n12182, new_n12183, new_n12184, new_n12185, new_n12186, new_n12187,
    new_n12188, new_n12189, new_n12190, new_n12191, new_n12192, new_n12193,
    new_n12194, new_n12195, new_n12196, new_n12197, new_n12198, new_n12199,
    new_n12200, new_n12201, new_n12202, new_n12203, new_n12204, new_n12205,
    new_n12206, new_n12207, new_n12209, new_n12210, new_n12211, new_n12212,
    new_n12213, new_n12214, new_n12215, new_n12216, new_n12217,
    new_n12218_1, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223, new_n12224, new_n12225, new_n12226, new_n12227, new_n12228,
    new_n12229, new_n12230, new_n12231, new_n12232_1, new_n12233,
    new_n12234, new_n12235, new_n12236, new_n12237, new_n12238, new_n12239,
    new_n12240, new_n12241, new_n12242, new_n12243, new_n12244, new_n12245,
    new_n12246, new_n12247, new_n12248, new_n12249, new_n12250, new_n12251,
    new_n12252, new_n12253, new_n12254, new_n12255, new_n12256, new_n12257,
    new_n12258, new_n12259, new_n12260, new_n12261, new_n12262, new_n12263,
    new_n12264, new_n12265, new_n12266, new_n12267, new_n12268, new_n12269,
    new_n12270_1, new_n12271, new_n12272, new_n12273, new_n12274,
    new_n12275, new_n12276, new_n12277, new_n12278, new_n12279, new_n12280,
    new_n12281, new_n12282, new_n12283, new_n12284, new_n12285, new_n12286,
    new_n12287, new_n12288, new_n12289, new_n12290, new_n12291, new_n12292,
    new_n12293, new_n12294, new_n12295, new_n12296, new_n12298, new_n12299,
    new_n12300, new_n12301, new_n12302, new_n12303, new_n12304, new_n12305,
    new_n12306, new_n12307, new_n12308, new_n12309, new_n12310, new_n12311,
    new_n12312, new_n12313, new_n12314, new_n12315, new_n12316, new_n12317,
    new_n12318, new_n12319, new_n12320, new_n12321_1, new_n12322,
    new_n12323, new_n12324, new_n12325, new_n12326, new_n12327, new_n12328,
    new_n12329, new_n12330, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336_1, new_n12337, new_n12338, new_n12339,
    new_n12340, new_n12341, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346, new_n12347, new_n12348, new_n12349, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12354, new_n12355_1, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364, new_n12365, new_n12366, new_n12367, new_n12368,
    new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374,
    new_n12375, new_n12376, new_n12377, new_n12378, new_n12379, new_n12380,
    new_n12381, new_n12382, new_n12383, new_n12384, new_n12386, new_n12387,
    new_n12388, new_n12389, new_n12390, new_n12391, new_n12392, new_n12393,
    new_n12394, new_n12395, new_n12396, new_n12397, new_n12398, new_n12399,
    new_n12400, new_n12401, new_n12402, new_n12403, new_n12404, new_n12405,
    new_n12406, new_n12407, new_n12408, new_n12409, new_n12410, new_n12411,
    new_n12412, new_n12413, new_n12414, new_n12415, new_n12416, new_n12417,
    new_n12418, new_n12419, new_n12420, new_n12421, new_n12422, new_n12423,
    new_n12424, new_n12425, new_n12426, new_n12427, new_n12428, new_n12429,
    new_n12430, new_n12431, new_n12432, new_n12433, new_n12434, new_n12435,
    new_n12436, new_n12437, new_n12438, new_n12439, new_n12440, new_n12441,
    new_n12442, new_n12443, new_n12444, new_n12445, new_n12446, new_n12447,
    new_n12448, new_n12449, new_n12450, new_n12451, new_n12452, new_n12453,
    new_n12454, new_n12455, new_n12456, new_n12457, new_n12458, new_n12459,
    new_n12460, new_n12461, new_n12462, new_n12463, new_n12464, new_n12465,
    new_n12466, new_n12467, new_n12468, new_n12469, new_n12470, new_n12471,
    new_n12472, new_n12473, new_n12474, new_n12475, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489, new_n12490,
    new_n12491, new_n12492, new_n12493, new_n12494, new_n12495, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507, new_n12508,
    new_n12509, new_n12510, new_n12511, new_n12512, new_n12513, new_n12514,
    new_n12515, new_n12516, new_n12517, new_n12518, new_n12519, new_n12520,
    new_n12521, new_n12522, new_n12523, new_n12524, new_n12525, new_n12526,
    new_n12527, new_n12528, new_n12529, new_n12530, new_n12531, new_n12532,
    new_n12533, new_n12534, new_n12535_1, new_n12536, new_n12537,
    new_n12538, new_n12539, new_n12540, new_n12541, new_n12542, new_n12543,
    new_n12544, new_n12545, new_n12546, new_n12547, new_n12548, new_n12549,
    new_n12550, new_n12551, new_n12552, new_n12553, new_n12554, new_n12555,
    new_n12556, new_n12557, new_n12558, new_n12559, new_n12560, new_n12561,
    new_n12562, new_n12563, new_n12565, new_n12566, new_n12567, new_n12568,
    new_n12569, new_n12570, new_n12571, new_n12572, new_n12573_1,
    new_n12574, new_n12575, new_n12576, new_n12577, new_n12578, new_n12579,
    new_n12580, new_n12581, new_n12582, new_n12583, new_n12584, new_n12585,
    new_n12586, new_n12587, new_n12588, new_n12589, new_n12590, new_n12591,
    new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597,
    new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603,
    new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614_1,
    new_n12615, new_n12616, new_n12617, new_n12618, new_n12619, new_n12620,
    new_n12621, new_n12622, new_n12623, new_n12624, new_n12625, new_n12626,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649, new_n12650,
    new_n12651, new_n12653, new_n12654, new_n12655, new_n12656, new_n12657,
    new_n12658, new_n12659, new_n12660, new_n12661, new_n12662, new_n12663,
    new_n12664, new_n12665, new_n12666, new_n12667, new_n12668, new_n12669,
    new_n12670, new_n12671, new_n12672, new_n12673, new_n12674, new_n12675,
    new_n12676, new_n12677, new_n12678, new_n12679, new_n12680, new_n12681,
    new_n12682, new_n12683, new_n12684, new_n12685, new_n12686, new_n12687,
    new_n12688, new_n12689, new_n12690, new_n12691, new_n12692, new_n12693,
    new_n12694, new_n12695, new_n12696, new_n12697, new_n12698, new_n12699,
    new_n12700, new_n12701, new_n12702, new_n12703, new_n12704, new_n12705,
    new_n12706, new_n12707, new_n12708, new_n12709, new_n12710, new_n12711,
    new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717,
    new_n12718, new_n12719, new_n12720, new_n12721, new_n12722, new_n12723,
    new_n12724, new_n12725, new_n12726, new_n12727, new_n12728, new_n12729,
    new_n12730, new_n12731, new_n12732, new_n12733, new_n12734, new_n12735,
    new_n12736, new_n12737, new_n12738, new_n12739, new_n12740, new_n12742,
    new_n12743, new_n12744, new_n12745, new_n12746, new_n12747, new_n12748,
    new_n12749, new_n12750, new_n12751, new_n12752, new_n12753, new_n12754,
    new_n12755, new_n12756, new_n12757, new_n12758, new_n12759, new_n12760,
    new_n12761, new_n12762, new_n12763, new_n12764, new_n12765, new_n12766,
    new_n12767, new_n12768, new_n12769, new_n12770, new_n12771, new_n12772,
    new_n12773, new_n12774, new_n12775, new_n12776, new_n12777, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782_1, new_n12783,
    new_n12784, new_n12785, new_n12786, new_n12787, new_n12788, new_n12789,
    new_n12790, new_n12791, new_n12792, new_n12793, new_n12794, new_n12795,
    new_n12796, new_n12797, new_n12798, new_n12799, new_n12800, new_n12801,
    new_n12802, new_n12803, new_n12804, new_n12805, new_n12806, new_n12807,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12830, new_n12831, new_n12832,
    new_n12833, new_n12834, new_n12835, new_n12836, new_n12837, new_n12838,
    new_n12839, new_n12840, new_n12841, new_n12842, new_n12843, new_n12844,
    new_n12845, new_n12846, new_n12847, new_n12848, new_n12849, new_n12850,
    new_n12851, new_n12852, new_n12853, new_n12854, new_n12855, new_n12856,
    new_n12857, new_n12858, new_n12859, new_n12860, new_n12861, new_n12862,
    new_n12863, new_n12864, new_n12865, new_n12866, new_n12867, new_n12868,
    new_n12869, new_n12870, new_n12871, new_n12872, new_n12873, new_n12874,
    new_n12875, new_n12876, new_n12877, new_n12878, new_n12879, new_n12880,
    new_n12881, new_n12882, new_n12883, new_n12884, new_n12885_1,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892, new_n12893, new_n12894, new_n12895, new_n12896, new_n12897,
    new_n12898, new_n12899, new_n12900, new_n12901, new_n12902, new_n12903,
    new_n12904, new_n12905, new_n12906, new_n12907, new_n12908, new_n12909,
    new_n12910, new_n12911, new_n12912, new_n12913, new_n12914, new_n12915,
    new_n12916, new_n12918, new_n12919, new_n12920, new_n12921, new_n12922,
    new_n12923, new_n12924, new_n12925, new_n12926, new_n12927_1,
    new_n12928, new_n12929, new_n12930, new_n12931, new_n12932, new_n12933,
    new_n12934, new_n12935, new_n12936, new_n12937, new_n12938, new_n12939,
    new_n12940, new_n12941, new_n12942, new_n12943, new_n12944, new_n12945,
    new_n12946, new_n12947, new_n12948, new_n12949, new_n12950, new_n12951,
    new_n12952, new_n12953, new_n12954, new_n12955, new_n12956, new_n12957,
    new_n12958, new_n12959, new_n12960, new_n12961, new_n12962, new_n12963,
    new_n12964, new_n12965, new_n12966, new_n12967, new_n12968, new_n12969,
    new_n12970, new_n12971, new_n12972, new_n12973, new_n12974, new_n12975,
    new_n12976_1, new_n12977, new_n12978, new_n12979, new_n12980,
    new_n12981, new_n12982, new_n12983, new_n12984, new_n12985, new_n12986,
    new_n12987, new_n12988, new_n12989_1, new_n12990, new_n12991,
    new_n12992, new_n12993, new_n12994, new_n12995, new_n12996, new_n12997,
    new_n12998, new_n12999, new_n13000_1, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13006, new_n13007, new_n13008, new_n13009,
    new_n13010_1, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045_1, new_n13046, new_n13047, new_n13048, new_n13049,
    new_n13050, new_n13051, new_n13052, new_n13053, new_n13054, new_n13055,
    new_n13056, new_n13057, new_n13058, new_n13059, new_n13060, new_n13061,
    new_n13062, new_n13063, new_n13064, new_n13065, new_n13066, new_n13067,
    new_n13068, new_n13069, new_n13070, new_n13071, new_n13072, new_n13073,
    new_n13074, new_n13075, new_n13076, new_n13077, new_n13078, new_n13079,
    new_n13080, new_n13081, new_n13082, new_n13083, new_n13084, new_n13085,
    new_n13086, new_n13087, new_n13088, new_n13089, new_n13090, new_n13091,
    new_n13092, new_n13093_1;
not_3  g00000(new_n386, n2674);
nor_4  g00001(new_n387, n10426, new_n386);
not_3  g00002(new_n388, n4895);
nor_4  g00003(new_n389_1, n8598, new_n388);
not_3  g00004(new_n390, n8780);
not_3  g00005(new_n391, n12270);
nand_4 g00006(new_n392, new_n391, new_n390);
nor_4  g00007(new_n393, new_n392, new_n389_1);
not_3  g00008(new_n394_1, n1268);
nor_4  g00009(new_n395, new_n394_1, n1265);
nor_4  g00010(new_n396, n8892, n1265);
nor_4  g00011(new_n397, new_n396, new_n395);
nor_4  g00012(new_n398, new_n397, n8598);
not_3  g00013(new_n399, n5046);
nor_4  g00014(new_n400, n6362, new_n399);
nor_4  g00015(new_n401, n1268, n394);
not_3  g00016(new_n402, new_n401);
nor_4  g00017(new_n403, new_n402, new_n400);
not_3  g00018(new_n404, n8649);
nor_4  g00019(new_n405, new_n404, n5950);
nor_4  g00020(new_n406, n12927, n10050);
not_3  g00021(new_n407, new_n406);
nor_4  g00022(new_n408, new_n407, new_n405);
not_3  g00023(new_n409, n8439);
nor_4  g00024(new_n410, new_n409, n702);
nor_4  g00025(new_n411_1, n3910, n844);
not_3  g00026(new_n412, new_n411_1);
nor_4  g00027(new_n413, new_n412, new_n410);
not_3  g00028(new_n414, n2061);
nor_4  g00029(new_n415, n9026, new_n414);
not_3  g00030(new_n416, n9186);
not_3  g00031(new_n417, n12336);
nand_4 g00032(new_n418, new_n417, new_n416);
nor_4  g00033(new_n419, new_n418, new_n415);
not_3  g00034(new_n420, n10147);
nor_4  g00035(new_n421, new_n420, n8397);
nor_4  g00036(new_n422, n14464, n12976);
not_3  g00037(new_n423, new_n422);
nor_4  g00038(new_n424, new_n423, new_n421);
not_3  g00039(new_n425, n7667);
nor_4  g00040(new_n426, n11930, new_n425);
nor_4  g00041(new_n427_1, n13636, n11930);
nor_4  g00042(new_n428, new_n427_1, new_n426);
nor_4  g00043(new_n429, new_n428, n8397);
not_3  g00044(new_n430, n14408);
nor_4  g00045(new_n431, n14483, new_n430);
nor_4  g00046(new_n432, n14303, n7667);
not_3  g00047(new_n433, new_n432);
nor_4  g00048(new_n434, new_n433, new_n431);
not_3  g00049(new_n435, n12025);
nor_4  g00050(new_n436, new_n435, n6460);
nor_4  g00051(new_n437, n5023, n3673);
not_3  g00052(new_n438, new_n437);
nor_4  g00053(new_n439, new_n438, new_n436);
not_3  g00054(new_n440, n3130);
nor_4  g00055(new_n441, n13000, new_n440);
nor_4  g00056(new_n442, n13000, n10446);
nor_4  g00057(new_n443, new_n442, new_n441);
nor_4  g00058(new_n444, new_n443, n6460);
not_3  g00059(new_n445, n5786);
nor_4  g00060(new_n446, n8486, new_n445);
nor_4  g00061(new_n447, n9589, n8552);
not_3  g00062(new_n448, new_n447);
nor_4  g00063(new_n449, new_n448, new_n446);
nor_4  g00064(new_n450, n8997, n3532);
not_3  g00065(new_n451_1, n3532);
nand_4 g00066(new_n452, n11345, new_n451_1);
not_3  g00067(new_n453, new_n452);
nor_4  g00068(new_n454, new_n453, new_n450);
nor_4  g00069(new_n455, new_n454, n8486);
not_3  g00070(new_n456, n6480);
nor_4  g00071(new_n457, n6791, new_n456);
nor_4  g00072(new_n458, n11345, n3263);
not_3  g00073(new_n459, new_n458);
nor_4  g00074(new_n460, new_n459, new_n457);
not_3  g00075(new_n461, n4615);
nor_4  g00076(new_n462_1, n4785, new_n461);
nor_4  g00077(new_n463, n9921, n730);
not_3  g00078(new_n464, new_n463);
nor_4  g00079(new_n465, new_n464, new_n462_1);
not_3  g00080(new_n466, n427);
nor_4  g00081(new_n467, n9893, new_n466);
nor_4  g00082(new_n468, n6999, n6517);
not_3  g00083(new_n469, new_n468);
nor_4  g00084(new_n470, new_n469, new_n467);
not_3  g00085(new_n471, new_n470);
not_3  g00086(new_n472, n12321);
nor_4  g00087(new_n473, new_n472, n5502);
nor_4  g00088(new_n474, n14072, n9544);
not_3  g00089(new_n475, new_n474);
nor_4  g00090(new_n476, new_n475, new_n473);
not_3  g00091(new_n477, new_n476);
not_3  g00092(new_n478, n6555);
nor_4  g00093(new_n479, n9555, new_n478);
nor_4  g00094(new_n480, n10736, n7972);
not_3  g00095(new_n481, new_n480);
nor_4  g00096(new_n482, new_n481, new_n479);
not_3  g00097(new_n483, new_n482);
not_3  g00098(new_n484, n4659);
nor_4  g00099(new_n485, new_n484, n4131);
nor_4  g00100(new_n486, n12573, n10470);
not_3  g00101(new_n487, new_n486);
nor_4  g00102(new_n488, new_n487, new_n485);
not_3  g00103(new_n489, new_n488);
not_3  g00104(new_n490_1, n11590);
nor_4  g00105(new_n491, new_n490_1, n5014);
nor_4  g00106(new_n492, n11158, n10407);
not_3  g00107(new_n493, new_n492);
nor_4  g00108(new_n494, new_n493, new_n491);
not_3  g00109(new_n495, new_n494);
not_3  g00110(new_n496, n9154);
nor_4  g00111(new_n497, n11933, new_n496);
nor_4  g00112(new_n498_1, n6436, n3833);
not_3  g00113(new_n499, new_n498_1);
nor_4  g00114(new_n500, new_n499, new_n497);
not_3  g00115(new_n501, new_n500);
not_3  g00116(new_n502, n11875);
nor_4  g00117(new_n503, new_n502, n8262);
nor_4  g00118(new_n504, n10061, n4117);
not_3  g00119(new_n505, new_n504);
nor_4  g00120(new_n506, new_n505, new_n503);
not_3  g00121(new_n507, n4022);
not_3  g00122(new_n508, n1568);
nand_4 g00123(new_n509, n8635, new_n508);
nand_4 g00124(new_n510, new_n509, new_n507);
nor_4  g00125(new_n511, new_n510, n13814);
not_3  g00126(new_n512, n8800);
nor_4  g00127(new_n513, new_n512, n8463);
not_3  g00128(new_n514, n203);
not_3  g00129(new_n515, n5184);
nand_4 g00130(new_n516, new_n515, new_n514);
nor_4  g00131(new_n517, new_n516, new_n513);
not_3  g00132(new_n518, n4154);
nor_4  g00133(new_n519, new_n518, n4000);
not_3  g00134(new_n520, n3506);
not_3  g00135(new_n521, n6703);
nand_4 g00136(new_n522, new_n521, new_n520);
nor_4  g00137(new_n523, new_n522, new_n519);
not_3  g00138(new_n524, n7652);
nor_4  g00139(new_n525, n8073, new_n524);
not_3  g00140(new_n526, n650);
not_3  g00141(new_n527, n13093);
nand_4 g00142(new_n528, new_n527, new_n526);
nor_4  g00143(new_n529, new_n528, new_n525);
not_3  g00144(new_n530, n3804);
nor_4  g00145(new_n531, n10112, new_n530);
nor_4  g00146(new_n532, n10466, n10112);
nor_4  g00147(new_n533, new_n532, new_n531);
nor_4  g00148(new_n534, new_n533, n8073);
not_3  g00149(new_n535, n13882);
nor_4  g00150(new_n536, new_n535, n5943);
nor_4  g00151(new_n537, n6680, n3804);
not_3  g00152(new_n538, new_n537);
nor_4  g00153(new_n539, new_n538, new_n536);
not_3  g00154(new_n540, n8746);
nor_4  g00155(new_n541, new_n540, n5430);
nor_4  g00156(new_n542, n8550, n5725);
not_3  g00157(new_n543_1, new_n542);
nor_4  g00158(new_n544, new_n543_1, new_n541);
nor_4  g00159(new_n545, n5430, n760);
not_3  g00160(new_n546, new_n545);
not_3  g00161(new_n547, n13295);
nor_4  g00162(new_n548, new_n547, n3799);
nor_4  g00163(new_n549, new_n548, new_n546);
not_3  g00164(new_n550, n3367);
nor_4  g00165(new_n551, n9543, new_n550);
nor_4  g00166(new_n552, n11776, n6873);
not_3  g00167(new_n553, new_n552);
nor_4  g00168(new_n554, new_n553, new_n551);
not_3  g00169(new_n555, n271);
nor_4  g00170(new_n556, n6007, new_n555);
nor_4  g00171(new_n557, n6007, n5960);
nor_4  g00172(new_n558, new_n557, new_n556);
nor_4  g00173(new_n559, new_n558, n9543);
not_3  g00174(new_n560, n13224);
nor_4  g00175(new_n561, new_n560, n11605);
nor_4  g00176(new_n562, n9977, n5225);
not_3  g00177(new_n563, new_n562);
nor_4  g00178(new_n564, new_n563, new_n561);
not_3  g00179(new_n565, n74);
nor_4  g00180(new_n566, n9314, new_n565);
not_3  g00181(new_n567, n9110);
not_3  g00182(new_n568, n13109);
nand_4 g00183(new_n569, new_n568, new_n567);
nor_4  g00184(new_n570, new_n569, new_n566);
not_3  g00185(new_n571, n1763);
nor_4  g00186(new_n572, n12009, new_n571);
nor_4  g00187(new_n573, n5033, n4172);
not_3  g00188(new_n574, new_n573);
nor_4  g00189(new_n575, new_n574, new_n572);
not_3  g00190(new_n576, n1222);
nor_4  g00191(new_n577, n11961, new_n576);
nor_4  g00192(new_n578, n7832, n1776);
not_3  g00193(new_n579, new_n578);
nor_4  g00194(new_n580, new_n579, new_n577);
not_3  g00195(new_n581, n11842);
nor_4  g00196(new_n582, new_n581, n1027);
nor_4  g00197(new_n583, n2048, n1027);
nor_4  g00198(new_n584, new_n583, new_n582);
nor_4  g00199(new_n585, new_n584, n11961);
not_3  g00200(new_n586, n2166);
not_3  g00201(new_n587, n8002);
nand_4 g00202(new_n588, new_n587, new_n586);
not_3  g00203(new_n589, n6147);
nand_4 g00204(new_n590, n2201, new_n586);
nand_4 g00205(new_n591, new_n590, new_n589);
nor_4  g00206(new_n592, new_n591, n11842);
nand_4 g00207(new_n593, new_n592, new_n588);
nand_4 g00208(new_n594, new_n593, new_n585);
nand_4 g00209(new_n595, new_n594, new_n580);
not_3  g00210(new_n596, n1776);
nor_4  g00211(new_n597, n14475, new_n596);
nor_4  g00212(new_n598, n14475, n13625);
nor_4  g00213(new_n599, new_n598, new_n597);
nor_4  g00214(new_n600, new_n599, n10573);
nand_4 g00215(new_n601, new_n600, new_n595);
not_3  g00216(new_n602, n13102);
nor_4  g00217(new_n603, new_n602, n10573);
nor_4  g00218(new_n604, n13363, n7354);
not_3  g00219(new_n605, new_n604);
nor_4  g00220(new_n606, new_n605, new_n603);
nand_4 g00221(new_n607, new_n606, new_n601);
not_3  g00222(new_n608, n13363);
nor_4  g00223(new_n609, new_n608, n6054);
nor_4  g00224(new_n610, n6054, n2573);
nor_4  g00225(new_n611, new_n610, new_n609);
nor_4  g00226(new_n612, new_n611, n12009);
nand_4 g00227(new_n613, new_n612, new_n607);
nand_4 g00228(new_n614, new_n613, new_n575);
not_3  g00229(new_n615, n4172);
nor_4  g00230(new_n616, n4774, new_n615);
nor_4  g00231(new_n617, n4774, n4755);
nor_4  g00232(new_n618, new_n617, new_n616);
nor_4  g00233(new_n619, new_n618, n9314);
nand_4 g00234(new_n620, new_n619, new_n614);
nand_4 g00235(new_n621, new_n620, new_n570);
nor_4  g00236(new_n622, new_n567, n7104);
nor_4  g00237(new_n623, n13231, n7104);
nor_4  g00238(new_n624, new_n623, new_n622);
nor_4  g00239(new_n625, new_n624, n11605);
nand_4 g00240(new_n626, new_n625, new_n621);
nand_4 g00241(new_n627, new_n626, new_n564);
not_3  g00242(new_n628, n9977);
nor_4  g00243(new_n629, new_n628, n1347);
nor_4  g00244(new_n630, n8315, n1347);
nor_4  g00245(new_n631, new_n630, new_n629);
nor_4  g00246(new_n632, new_n631, n6258);
nand_4 g00247(new_n633, new_n632, new_n627);
not_3  g00248(new_n634, n13890);
nor_4  g00249(new_n635, new_n634, n6258);
not_3  g00250(new_n636, n2334);
nand_4 g00251(new_n637, new_n636, new_n555);
nor_4  g00252(new_n638, new_n637, new_n635);
nand_4 g00253(new_n639, new_n638, new_n633);
nand_4 g00254(new_n640, new_n639, new_n559);
nand_4 g00255(new_n641, new_n640, new_n554);
not_3  g00256(new_n642, n6873);
nor_4  g00257(new_n643, n7988, new_n642);
nor_4  g00258(new_n644, n10912, n7988);
nor_4  g00259(new_n645, new_n644, new_n643);
nor_4  g00260(new_n646, new_n645, n10630);
nand_4 g00261(new_n647, new_n646, new_n641);
not_3  g00262(new_n648, n5185);
nor_4  g00263(new_n649, n10630, new_n648);
nor_4  g00264(new_n650_1, n3799, n3652);
not_3  g00265(new_n651, new_n650_1);
nor_4  g00266(new_n652, new_n651, new_n649);
nand_4 g00267(new_n653, new_n652, new_n647);
nand_4 g00268(new_n654, new_n653, new_n549);
nand_4 g00269(new_n655, new_n654, new_n544);
not_3  g00270(new_n656_1, n5725);
nor_4  g00271(new_n657, new_n656_1, n2164);
nor_4  g00272(new_n658, n14163, n2164);
nor_4  g00273(new_n659, new_n658, new_n657);
nor_4  g00274(new_n660, new_n659, n5943);
nand_4 g00275(new_n661, new_n660, new_n655);
nand_4 g00276(new_n662, new_n661, new_n539);
nand_4 g00277(new_n663, new_n662, new_n534);
nand_4 g00278(new_n664, new_n663, new_n529);
nor_4  g00279(new_n665, n9252, new_n526);
nor_4  g00280(new_n666_1, n11902, n9252);
nor_4  g00281(new_n667, new_n666_1, new_n665);
nor_4  g00282(new_n668, new_n667, n411);
nand_4 g00283(new_n669, new_n668, new_n664);
not_3  g00284(new_n670, n8799);
nor_4  g00285(new_n671, new_n670, n411);
nor_4  g00286(new_n672, n12614, n10765);
not_3  g00287(new_n673, new_n672);
nor_4  g00288(new_n674_1, new_n673, new_n671);
nand_4 g00289(new_n675, new_n674_1, new_n669);
not_3  g00290(new_n676, n3388);
not_3  g00291(new_n677, n4000);
nand_4 g00292(new_n678, new_n677, new_n676);
not_3  g00293(new_n679, n12142);
nor_4  g00294(new_n680, new_n679, n10765);
nor_4  g00295(new_n681, new_n680, new_n678);
nand_4 g00296(new_n682_1, new_n681, new_n675);
nand_4 g00297(new_n683, new_n682_1, new_n523);
nor_4  g00298(new_n684, n11269, new_n521);
nor_4  g00299(new_n685, n11269, n462);
nor_4  g00300(new_n686, new_n685, new_n684);
nor_4  g00301(new_n687, new_n686, n8926);
nand_4 g00302(new_n688, new_n687, new_n683);
not_3  g00303(new_n689, n3893);
nor_4  g00304(new_n690, n8926, new_n689);
nor_4  g00305(new_n691, n8044, n2454);
not_3  g00306(new_n692, new_n691);
nor_4  g00307(new_n693, new_n692, new_n690);
nand_4 g00308(new_n694, new_n693, new_n688);
not_3  g00309(new_n695, n8044);
nor_4  g00310(new_n696, n8204, new_n695);
nor_4  g00311(new_n697, n14293, n8204);
nor_4  g00312(new_n698, new_n697, new_n696);
nor_4  g00313(new_n699, new_n698, n8463);
nand_4 g00314(new_n700, new_n699, new_n694);
nand_4 g00315(new_n701, new_n700, new_n517);
nor_4  g00316(new_n702_1, new_n515, n2895);
nor_4  g00317(new_n703, n2895, n737);
nor_4  g00318(new_n704, new_n703, new_n702_1);
nor_4  g00319(new_n705, new_n704, n1568);
nand_4 g00320(new_n706, new_n705, new_n701);
nand_4 g00321(new_n707, new_n706, new_n511);
nor_4  g00322(new_n708, n10255, new_n507);
nor_4  g00323(new_n709, n10255, n5449);
nor_4  g00324(new_n710, new_n709, new_n708);
nor_4  g00325(new_n711, new_n710, n8262);
nand_4 g00326(new_n712, new_n711, new_n707);
nand_4 g00327(new_n713, new_n712, new_n506);
not_3  g00328(new_n714, new_n713);
not_3  g00329(new_n715, n10061);
nor_4  g00330(new_n716, n12885, new_n715);
nor_4  g00331(new_n717, n12885, n11666);
nor_4  g00332(new_n718, new_n717, new_n716);
nor_4  g00333(new_n719, new_n718, n11933);
not_3  g00334(new_n720, new_n719);
nor_4  g00335(new_n721, new_n720, new_n714);
nor_4  g00336(new_n722, new_n721, new_n501);
nor_4  g00337(new_n723, n11143, n5014);
not_3  g00338(new_n724, new_n723);
not_3  g00339(new_n725, n2699);
nor_4  g00340(new_n726, n6436, new_n725);
nor_4  g00341(new_n727, new_n726, new_n724);
not_3  g00342(new_n728, new_n727);
nor_4  g00343(new_n729, new_n728, new_n722);
nor_4  g00344(new_n730_1, new_n729, new_n495);
nor_4  g00345(new_n731, n10051, n4131);
not_3  g00346(new_n732, new_n731);
not_3  g00347(new_n733, n13992);
nor_4  g00348(new_n734, new_n733, n10407);
nor_4  g00349(new_n735, new_n734, new_n732);
not_3  g00350(new_n736, new_n735);
nor_4  g00351(new_n737_1, new_n736, new_n730_1);
nor_4  g00352(new_n738, new_n737_1, new_n489);
not_3  g00353(new_n739, n10470);
nor_4  g00354(new_n740, new_n739, n6693);
nor_4  g00355(new_n741, n12829, n6693);
nor_4  g00356(new_n742, new_n741, new_n740);
nor_4  g00357(new_n743, new_n742, n9555);
not_3  g00358(new_n744, new_n743);
nor_4  g00359(new_n745, new_n744, new_n738);
nor_4  g00360(new_n746, new_n745, new_n483);
not_3  g00361(new_n747, n7972);
nor_4  g00362(new_n748, new_n747, n3972);
nor_4  g00363(new_n749, n10945, n3972);
nor_4  g00364(new_n750, new_n749, new_n748);
nor_4  g00365(new_n751, new_n750, n7450);
not_3  g00366(new_n752, new_n751);
nor_4  g00367(new_n753, new_n752, new_n746);
not_3  g00368(new_n754, n10615);
nor_4  g00369(new_n755, new_n754, n7450);
nor_4  g00370(new_n756, n9830, n8302);
not_3  g00371(new_n757, new_n756);
nor_4  g00372(new_n758, new_n757, new_n755);
not_3  g00373(new_n759, new_n758);
nor_4  g00374(new_n760_1, new_n759, new_n753);
not_3  g00375(new_n761, n8302);
nor_4  g00376(new_n762, new_n761, n3166);
nor_4  g00377(new_n763, n6270, n3166);
nor_4  g00378(new_n764, new_n763, new_n762);
nor_4  g00379(new_n765, new_n764, n5502);
not_3  g00380(new_n766, new_n765);
nor_4  g00381(new_n767, new_n766, new_n760_1);
nor_4  g00382(new_n768, new_n767, new_n477);
not_3  g00383(new_n769, n14072);
nor_4  g00384(new_n770, new_n769, n6251);
nor_4  g00385(new_n771, n6251, n1702);
nor_4  g00386(new_n772, new_n771, new_n770);
nor_4  g00387(new_n773, new_n772, n6758);
not_3  g00388(new_n774, new_n773);
nor_4  g00389(new_n775, new_n774, new_n768);
not_3  g00390(new_n776, n4147);
nor_4  g00391(new_n777, n6758, new_n776);
nor_4  g00392(new_n778, n10378, n10080);
not_3  g00393(new_n779, new_n778);
nor_4  g00394(new_n780, new_n779, new_n777);
not_3  g00395(new_n781, new_n780);
nor_4  g00396(new_n782, new_n781, new_n775);
not_3  g00397(new_n783, n10080);
nor_4  g00398(new_n784, new_n783, n977);
nor_4  g00399(new_n785, n4282, n977);
nor_4  g00400(new_n786, new_n785, new_n784);
nor_4  g00401(new_n787, new_n786, n9893);
not_3  g00402(new_n788, new_n787);
nor_4  g00403(new_n789, new_n788, new_n782);
nor_4  g00404(new_n790, new_n789, new_n471);
not_3  g00405(new_n791, n6999);
nor_4  g00406(new_n792, n10862, new_n791);
nor_4  g00407(new_n793, n12218, n10862);
nor_4  g00408(new_n794, new_n793, new_n792);
nor_4  g00409(new_n795, new_n794, n9936);
not_3  g00410(new_n796, new_n795);
nor_4  g00411(new_n797, new_n796, new_n790);
not_3  g00412(new_n798, n1093);
nor_4  g00413(new_n799, n9936, new_n798);
not_3  g00414(new_n800, n2615);
not_3  g00415(new_n801, n8737);
nand_4 g00416(new_n802, new_n801, new_n800);
nor_4  g00417(new_n803, new_n802, new_n799);
not_3  g00418(new_n804, new_n803);
nor_4  g00419(new_n805, new_n804, new_n797);
nor_4  g00420(new_n806, n13561, new_n801);
nor_4  g00421(new_n807, n13561, n656);
nor_4  g00422(new_n808, new_n807, new_n806);
nor_4  g00423(new_n809, new_n808, n4785);
not_3  g00424(new_n810, new_n809);
nor_4  g00425(new_n811, new_n810, new_n805);
not_3  g00426(new_n812, new_n811);
nand_4 g00427(new_n813, new_n812, new_n465);
not_3  g00428(new_n814, n9921);
nor_4  g00429(new_n815, n10283, new_n814);
nor_4  g00430(new_n816, n10283, n3775);
nor_4  g00431(new_n817, new_n816, new_n815);
nor_4  g00432(new_n818, new_n817, n6791);
nand_4 g00433(new_n819, new_n818, new_n813);
nand_4 g00434(new_n820, new_n819, new_n460);
nand_4 g00435(new_n821, new_n820, new_n455);
nand_4 g00436(new_n822, new_n821, new_n449);
not_3  g00437(new_n823, n9589);
nor_4  g00438(new_n824, n10750, new_n823);
nor_4  g00439(new_n825, n10750, n1637);
nor_4  g00440(new_n826, new_n825, new_n824);
nor_4  g00441(new_n827, new_n826, n498);
nand_4 g00442(new_n828, new_n827, new_n822);
not_3  g00443(new_n829, n11404);
nor_4  g00444(new_n830, new_n829, n498);
nor_4  g00445(new_n831, n4175, n3130);
not_3  g00446(new_n832, new_n831);
nor_4  g00447(new_n833, new_n832, new_n830);
nand_4 g00448(new_n834, new_n833, new_n828);
nand_4 g00449(new_n835, new_n834, new_n444);
nand_4 g00450(new_n836, new_n835, new_n439);
not_3  g00451(new_n837, n5023);
nor_4  g00452(new_n838, new_n837, n4225);
nor_4  g00453(new_n839, n6586, n4225);
nor_4  g00454(new_n840, new_n839, new_n838);
nor_4  g00455(new_n841, new_n840, n14483);
nand_4 g00456(new_n842, new_n841, new_n836);
nand_4 g00457(new_n843, new_n842, new_n434);
nand_4 g00458(new_n844_1, new_n843, new_n429);
nand_4 g00459(new_n845, new_n844_1, new_n424);
not_3  g00460(new_n846, n12976);
nor_4  g00461(new_n847, new_n846, n6810);
nor_4  g00462(new_n848, n12012, n6810);
nor_4  g00463(new_n849, new_n848, new_n847);
nor_4  g00464(new_n850, new_n849, n11756);
nand_4 g00465(new_n851, new_n850, new_n845);
not_3  g00466(new_n852, n666);
nor_4  g00467(new_n853, n11756, new_n852);
nor_4  g00468(new_n854, n13511, n13364);
not_3  g00469(new_n855, new_n854);
nor_4  g00470(new_n856, new_n855, new_n853);
nand_4 g00471(new_n857, new_n856, new_n851);
not_3  g00472(new_n858, n3655);
not_3  g00473(new_n859, n9026);
nand_4 g00474(new_n860, new_n859, new_n858);
not_3  g00475(new_n861, n4907);
nor_4  g00476(new_n862, n13364, new_n861);
nor_4  g00477(new_n863, new_n862, new_n860);
nand_4 g00478(new_n864, new_n863, new_n857);
nand_4 g00479(new_n865, new_n864, new_n419);
nor_4  g00480(new_n866, new_n417, n4292);
nor_4  g00481(new_n867, n6114, n4292);
nor_4  g00482(new_n868, new_n867, new_n866);
nor_4  g00483(new_n869, new_n868, n7272);
nand_4 g00484(new_n870, new_n869, new_n865);
not_3  g00485(new_n871, n7748);
not_3  g00486(new_n872, n7272);
nand_4 g00487(new_n873, n12782, new_n872);
nand_4 g00488(new_n874, new_n873, new_n871);
nor_4  g00489(new_n875, new_n874, n13186);
nand_4 g00490(new_n876, new_n875, new_n870);
not_3  g00491(new_n877, n11854);
not_3  g00492(new_n878, n13186);
nand_4 g00493(new_n879, new_n878, n10278);
nand_4 g00494(new_n880, new_n879, new_n877);
nor_4  g00495(new_n881, new_n880, n702);
nand_4 g00496(new_n882, new_n881, new_n876);
nand_4 g00497(new_n883, new_n882, new_n413);
not_3  g00498(new_n884_1, n674);
not_3  g00499(new_n885, n5077);
nand_4 g00500(new_n886, new_n885, new_n884_1);
not_3  g00501(new_n887, n8873);
nor_4  g00502(new_n888, new_n887, n3910);
nor_4  g00503(new_n889, new_n888, new_n886);
nand_4 g00504(new_n890, new_n889, new_n883);
not_3  g00505(new_n891, n5467);
nor_4  g00506(new_n892, new_n891, n5077);
not_3  g00507(new_n893, n7282);
not_3  g00508(new_n894, n13944);
nand_4 g00509(new_n895, new_n894, new_n893);
nor_4  g00510(new_n896, new_n895, new_n892);
nand_4 g00511(new_n897, new_n896, new_n890);
nor_4  g00512(new_n898, new_n894, n7941);
nor_4  g00513(new_n899, n7941, n6946);
nor_4  g00514(new_n900, new_n899, new_n898);
nor_4  g00515(new_n901, new_n900, n5950);
nand_4 g00516(new_n902, new_n901, new_n897);
nand_4 g00517(new_n903, new_n902, new_n408);
not_3  g00518(new_n904, n10050);
nor_4  g00519(new_n905, new_n904, n4039);
nor_4  g00520(new_n906, n11529, n4039);
nor_4  g00521(new_n907, new_n906, new_n905);
nor_4  g00522(new_n908, new_n907, n6362);
nand_4 g00523(new_n909, new_n908, new_n903);
nand_4 g00524(new_n910, new_n909, new_n403);
nand_4 g00525(new_n911, new_n910, new_n398);
nand_4 g00526(new_n912, new_n911, new_n393);
nor_4  g00527(new_n913, new_n391, n5601);
nor_4  g00528(new_n914, n5601, n5009);
nor_4  g00529(new_n915, new_n914, new_n913);
nor_4  g00530(new_n916, new_n915, n10426);
nand_4 g00531(new_n917, new_n916, new_n912);
nand_4 g00532(new_n918, new_n917, n13509);
nor_4  g00533(n8, new_n918, new_n387);
not_3  g00534(new_n920, n10378);
nor_4  g00535(new_n921, new_n920, n4282);
not_3  g00536(new_n922, n6758);
nand_4 g00537(new_n923, n6251, new_n776);
nand_4 g00538(new_n924, new_n923, new_n922);
nor_4  g00539(new_n925, new_n924, n4282);
not_3  g00540(new_n926, n1702);
nand_4 g00541(new_n927, n9544, new_n926);
nand_4 g00542(new_n928, new_n927, new_n776);
nor_4  g00543(new_n929, new_n928, n14072);
not_3  g00544(new_n930, n5502);
nand_4 g00545(new_n931, new_n930, new_n926);
not_3  g00546(new_n932, n3166);
nor_4  g00547(new_n933, n12321, new_n932);
nor_4  g00548(new_n934, new_n933, new_n931);
not_3  g00549(new_n935, n9830);
nor_4  g00550(new_n936, new_n935, n6270);
nand_4 g00551(new_n937, new_n472, new_n761);
nor_4  g00552(new_n938, new_n937, new_n936);
nor_4  g00553(new_n939, n7450, n6270);
not_3  g00554(new_n940, new_n939);
not_3  g00555(new_n941, n3972);
nor_4  g00556(new_n942, n10615, new_n941);
nor_4  g00557(new_n943, new_n942, new_n940);
not_3  g00558(new_n944, n10736);
nor_4  g00559(new_n945, n10945, new_n944);
nor_4  g00560(new_n946, n10615, n7972);
not_3  g00561(new_n947, new_n946);
nor_4  g00562(new_n948_1, new_n947, new_n945);
not_3  g00563(new_n949, n9555);
nand_4 g00564(new_n950, n6693, new_n478);
nand_4 g00565(new_n951, new_n950, new_n949);
nor_4  g00566(new_n952, new_n951, n10945);
not_3  g00567(new_n953, new_n952);
not_3  g00568(new_n954, n12573);
nor_4  g00569(new_n955, n12829, new_n954);
nand_4 g00570(new_n956, new_n739, new_n478);
nor_4  g00571(new_n957, new_n956, new_n955);
not_3  g00572(new_n958, new_n957);
nor_4  g00573(new_n959, new_n731, new_n485);
nor_4  g00574(new_n960, new_n959, n12829);
not_3  g00575(new_n961, new_n960);
nand_4 g00576(new_n962, new_n733, n11158);
nand_4 g00577(new_n963, new_n962, new_n484);
nor_4  g00578(new_n964, new_n963, n10407);
not_3  g00579(new_n965, new_n964);
nor_4  g00580(new_n966, new_n723, new_n491);
nor_4  g00581(new_n967, new_n966, n13992);
not_3  g00582(new_n968, new_n967);
not_3  g00583(new_n969, n3833);
nor_4  g00584(new_n970, new_n969, n2699);
nor_4  g00585(new_n971, n11590, n6436);
not_3  g00586(new_n972, new_n971);
nor_4  g00587(new_n973, new_n972, new_n970);
not_3  g00588(new_n974, new_n973);
not_3  g00589(new_n975, n11933);
nand_4 g00590(new_n976, n12885, new_n496);
nand_4 g00591(new_n977_1, new_n976, new_n975);
nor_4  g00592(new_n978, new_n977_1, n2699);
not_3  g00593(new_n979, new_n978);
not_3  g00594(new_n980, n4117);
nor_4  g00595(new_n981, n11666, new_n980);
nor_4  g00596(new_n982, n10061, n9154);
not_3  g00597(new_n983, new_n982);
nor_4  g00598(new_n984, new_n983, new_n981);
not_3  g00599(new_n985, new_n984);
not_3  g00600(new_n986, n8262);
nand_4 g00601(new_n987, new_n502, n10255);
nand_4 g00602(new_n988, new_n987, new_n986);
nor_4  g00603(new_n989, new_n988, n11666);
not_3  g00604(new_n990, new_n989);
not_3  g00605(new_n991, n13814);
nor_4  g00606(new_n992, new_n991, n5449);
nand_4 g00607(new_n993, new_n502, new_n507);
nor_4  g00608(new_n994, new_n993, new_n992);
not_3  g00609(new_n995, new_n994);
not_3  g00610(new_n996, n5449);
nand_4 g00611(new_n997, new_n996, new_n508);
not_3  g00612(new_n998, n2895);
nor_4  g00613(new_n999, n8635, new_n998);
nor_4  g00614(new_n1000, new_n999, new_n997);
not_3  g00615(new_n1001, new_n1000);
nor_4  g00616(new_n1002, n737, new_n514);
nor_4  g00617(new_n1003, n8635, n5184);
not_3  g00618(new_n1004, new_n1003);
nor_4  g00619(new_n1005, new_n1004, new_n1002);
not_3  g00620(new_n1006, new_n1005);
not_3  g00621(new_n1007, n2454);
nor_4  g00622(new_n1008, n14293, new_n1007);
nand_4 g00623(new_n1009, new_n512, new_n695);
nor_4  g00624(new_n1010, new_n1009, new_n1008);
not_3  g00625(new_n1011, new_n1010);
not_3  g00626(new_n1012, n8926);
nand_4 g00627(new_n1013, n11269, new_n689);
nand_4 g00628(new_n1014, new_n1013, new_n1012);
nor_4  g00629(new_n1015, new_n1014, n14293);
not_3  g00630(new_n1016, new_n1015);
nor_4  g00631(new_n1017, new_n520, n462);
nor_4  g00632(new_n1018, n6703, n3893);
not_3  g00633(new_n1019, new_n1018);
nor_4  g00634(new_n1020, new_n1019, new_n1017);
not_3  g00635(new_n1021, new_n1020);
nor_4  g00636(new_n1022, n4000, n462);
not_3  g00637(new_n1023, new_n1022);
nor_4  g00638(new_n1024, n4154, new_n676);
nor_4  g00639(new_n1025, new_n1024, new_n1023);
not_3  g00640(new_n1026, new_n1025);
not_3  g00641(new_n1027_1, n12614);
nor_4  g00642(new_n1028, new_n1027_1, n12142);
not_3  g00643(new_n1029, n10765);
nand_4 g00644(new_n1030, new_n1029, new_n518);
nor_4  g00645(new_n1031, new_n1030, new_n1028);
not_3  g00646(new_n1032, new_n1031);
not_3  g00647(new_n1033, n411);
nand_4 g00648(new_n1034, n9252, new_n670);
nand_4 g00649(new_n1035, new_n1034, new_n1033);
nor_4  g00650(new_n1036, new_n1035, n12142);
not_3  g00651(new_n1037, new_n1036);
nor_4  g00652(new_n1038, new_n527, n11902);
nor_4  g00653(new_n1039, n8799, n650);
not_3  g00654(new_n1040, new_n1039);
nor_4  g00655(new_n1041, new_n1040, new_n1038);
not_3  g00656(new_n1042, new_n1041);
nor_4  g00657(new_n1043, n10112, n8073);
nor_4  g00658(new_n1044, new_n1043, new_n525);
nor_4  g00659(new_n1045, new_n1044, n11902);
not_3  g00660(new_n1046, new_n1045);
not_3  g00661(new_n1047, n6680);
nor_4  g00662(new_n1048, n10466, new_n1047);
nand_4 g00663(new_n1049, new_n524, new_n530);
nor_4  g00664(new_n1050, new_n1049, new_n1048);
not_3  g00665(new_n1051, new_n1050);
not_3  g00666(new_n1052, n5943);
nand_4 g00667(new_n1053, new_n535, n2164);
nand_4 g00668(new_n1054, new_n1053, new_n1052);
nor_4  g00669(new_n1055, new_n1054, n10466);
not_3  g00670(new_n1056, new_n1055);
not_3  g00671(new_n1057, n8550);
nor_4  g00672(new_n1058, n14163, new_n1057);
nor_4  g00673(new_n1059, n13882, n5725);
not_3  g00674(new_n1060, new_n1059);
nor_4  g00675(new_n1061, new_n1060, new_n1058);
not_3  g00676(new_n1062, new_n1061);
nor_4  g00677(new_n1063, new_n545, new_n541);
nor_4  g00678(new_n1064, new_n1063, n14163);
not_3  g00679(new_n1065, new_n1064);
not_3  g00680(new_n1066, n3652);
nor_4  g00681(new_n1067, n13295, new_n1066);
not_3  g00682(new_n1068, n3799);
nand_4 g00683(new_n1069, new_n540, new_n1068);
nor_4  g00684(new_n1070, new_n1069, new_n1067);
not_3  g00685(new_n1071, new_n1070);
nor_4  g00686(new_n1072, n10630, n7988);
nor_4  g00687(new_n1073, new_n1072, new_n649);
nor_4  g00688(new_n1074, new_n1073, n13295);
not_3  g00689(new_n1075, new_n1074);
not_3  g00690(new_n1076, n10912);
nand_4 g00691(new_n1077, n11776, new_n1076);
nand_4 g00692(new_n1078, new_n1077, new_n648);
nor_4  g00693(new_n1079, new_n1078, n6873);
nor_4  g00694(new_n1080, n10912, n9543);
not_3  g00695(new_n1081, new_n1080);
not_3  g00696(new_n1082, n6007);
nor_4  g00697(new_n1083, new_n1082, n3367);
nor_4  g00698(new_n1084, new_n1083, new_n1081);
nor_4  g00699(new_n1085, n5960, new_n636);
nor_4  g00700(new_n1086, n3367, n271);
not_3  g00701(new_n1087, new_n1086);
nor_4  g00702(new_n1088, new_n1087, new_n1085);
nor_4  g00703(new_n1089, n6258, n1347);
nor_4  g00704(new_n1090, new_n1089, new_n635);
nor_4  g00705(new_n1091, new_n1090, n5960);
not_3  g00706(new_n1092, n8315);
nand_4 g00707(new_n1093_1, new_n1092, n5225);
nand_4 g00708(new_n1094_1, new_n1093_1, new_n628);
nor_4  g00709(new_n1095, new_n1094_1, n13890);
nor_4  g00710(new_n1096, n13231, new_n568);
nor_4  g00711(new_n1097, n13224, n9110);
not_3  g00712(new_n1098, new_n1097);
nor_4  g00713(new_n1099, new_n1098, new_n1096);
nor_4  g00714(new_n1100, n9314, n4774);
nor_4  g00715(new_n1101, new_n1100, new_n566);
nor_4  g00716(new_n1102, new_n1101, n13231);
not_3  g00717(new_n1103, n7354);
nor_4  g00718(new_n1104, new_n1103, n2573);
nand_4 g00719(new_n1105, new_n608, new_n571);
nor_4  g00720(new_n1106, new_n1105, new_n1104);
nor_4  g00721(new_n1107, n10573, n2573);
not_3  g00722(new_n1108, new_n1107);
not_3  g00723(new_n1109, n14475);
nor_4  g00724(new_n1110, new_n1109, n13102);
nor_4  g00725(new_n1111, new_n1110, new_n1108);
not_3  g00726(new_n1112, n7832);
nor_4  g00727(new_n1113, n13625, new_n1112);
nor_4  g00728(new_n1114, n13102, n1776);
not_3  g00729(new_n1115, new_n1114);
nor_4  g00730(new_n1116, new_n1115, new_n1113);
nor_4  g00731(new_n1117, new_n589, n2048);
nor_4  g00732(new_n1118, n11842, n1222);
not_3  g00733(new_n1119, new_n1118);
nor_4  g00734(new_n1120, new_n1119, new_n1117);
nor_4  g00735(new_n1121, n13509, n2201);
not_3  g00736(new_n1122_1, new_n1121);
nor_4  g00737(new_n1123, new_n1122_1, new_n387);
nor_4  g00738(new_n1124_1, n9893, n977);
nor_4  g00739(new_n1125, new_n1124_1, new_n467);
nand_4 g00740(new_n1126, new_n1125, new_n468);
nand_4 g00741(new_n1127, new_n1126, new_n795);
nand_4 g00742(new_n1128, new_n1127, new_n803);
nand_4 g00743(new_n1129, new_n1128, new_n809);
nand_4 g00744(new_n1130, new_n1129, new_n465);
nand_4 g00745(new_n1131, new_n1130, new_n818);
nand_4 g00746(new_n1132, new_n1131, new_n460);
nand_4 g00747(new_n1133, new_n1132, new_n455);
nand_4 g00748(new_n1134, new_n1133, new_n449);
nand_4 g00749(new_n1135, new_n1134, new_n827);
nand_4 g00750(new_n1136, new_n1135, new_n833);
nand_4 g00751(new_n1137, new_n1136, new_n444);
nand_4 g00752(new_n1138, new_n1137, new_n439);
nand_4 g00753(new_n1139, new_n1138, new_n841);
nand_4 g00754(new_n1140, new_n1139, new_n434);
nand_4 g00755(new_n1141, new_n1140, new_n429);
nand_4 g00756(new_n1142, new_n1141, new_n424);
nand_4 g00757(new_n1143, new_n1142, new_n850);
nand_4 g00758(new_n1144, new_n1143, new_n856);
nand_4 g00759(new_n1145, new_n1144, new_n863);
nand_4 g00760(new_n1146, new_n1145, new_n419);
nand_4 g00761(new_n1147, new_n1146, new_n869);
nand_4 g00762(new_n1148, new_n1147, new_n875);
nand_4 g00763(new_n1149, new_n1148, new_n881);
nand_4 g00764(new_n1150, new_n1149, new_n413);
nand_4 g00765(new_n1151, new_n1150, new_n889);
nand_4 g00766(new_n1152, new_n1151, new_n896);
nand_4 g00767(new_n1153, new_n1152, new_n901);
nand_4 g00768(new_n1154, new_n1153, new_n408);
nand_4 g00769(new_n1155, new_n1154, new_n908);
nand_4 g00770(new_n1156, new_n1155, new_n403);
nand_4 g00771(new_n1157, new_n1156, new_n398);
nand_4 g00772(new_n1158, new_n1157, new_n393);
nand_4 g00773(new_n1159, new_n1158, new_n916);
nand_4 g00774(new_n1160, new_n1159, new_n1123);
nor_4  g00775(new_n1161, n2166, n2048);
not_3  g00776(new_n1162, new_n1161);
nor_4  g00777(new_n1163, new_n587, n2201);
nor_4  g00778(new_n1164, new_n1163, new_n1162);
nand_4 g00779(new_n1165, new_n1164, new_n1160);
nand_4 g00780(new_n1166, new_n1165, new_n1120);
nor_4  g00781(new_n1167, n11961, n1027);
nor_4  g00782(new_n1168, new_n1167, new_n577);
nor_4  g00783(new_n1169, new_n1168, n13625);
nand_4 g00784(new_n1170, new_n1169, new_n1166);
nand_4 g00785(new_n1171, new_n1170, new_n1116);
nand_4 g00786(new_n1172, new_n1171, new_n1111);
nand_4 g00787(new_n1173, new_n1172, new_n1106);
nor_4  g00788(new_n1174, n12009, n4755);
not_3  g00789(new_n1175, new_n1174);
not_3  g00790(new_n1176, n6054);
nor_4  g00791(new_n1177, new_n1176, n1763);
nor_4  g00792(new_n1178, new_n1177, new_n1175);
nand_4 g00793(new_n1179, new_n1178, new_n1173);
not_3  g00794(new_n1180, n4755);
nand_4 g00795(new_n1181, n5033, new_n1180);
nand_4 g00796(new_n1182, new_n1181, new_n565);
nor_4  g00797(new_n1183, new_n1182, n4172);
nand_4 g00798(new_n1184, new_n1183, new_n1179);
nand_4 g00799(new_n1185, new_n1184, new_n1102);
nand_4 g00800(new_n1186, new_n1185, new_n1099);
not_3  g00801(new_n1187, n11605);
nand_4 g00802(new_n1188, new_n1187, new_n1092);
not_3  g00803(new_n1189, n7104);
nor_4  g00804(new_n1190, n13224, new_n1189);
nor_4  g00805(new_n1191, new_n1190, new_n1188);
nand_4 g00806(new_n1192, new_n1191, new_n1186);
nand_4 g00807(new_n1193, new_n1192, new_n1095);
nand_4 g00808(new_n1194, new_n1193, new_n1091);
nand_4 g00809(new_n1195, new_n1194, new_n1088);
nand_4 g00810(new_n1196, new_n1195, new_n1084);
nand_4 g00811(new_n1197, new_n1196, new_n1079);
not_3  g00812(new_n1198, new_n1197);
nor_4  g00813(new_n1199, new_n1198, new_n1075);
nor_4  g00814(new_n1200, new_n1199, new_n1071);
nor_4  g00815(new_n1201, new_n1200, new_n1065);
nor_4  g00816(new_n1202, new_n1201, new_n1062);
nor_4  g00817(new_n1203, new_n1202, new_n1056);
nor_4  g00818(new_n1204, new_n1203, new_n1051);
nor_4  g00819(new_n1205, new_n1204, new_n1046);
nor_4  g00820(new_n1206, new_n1205, new_n1042);
nor_4  g00821(new_n1207, new_n1206, new_n1037);
nor_4  g00822(new_n1208, new_n1207, new_n1032);
nor_4  g00823(new_n1209, new_n1208, new_n1026);
nor_4  g00824(new_n1210, new_n1209, new_n1021);
nor_4  g00825(new_n1211, new_n1210, new_n1016);
nor_4  g00826(new_n1212, new_n1211, new_n1011);
nor_4  g00827(new_n1213, n8463, n8204);
nor_4  g00828(new_n1214, new_n1213, new_n513);
nor_4  g00829(new_n1215, new_n1214, n737);
not_3  g00830(new_n1216, new_n1215);
nor_4  g00831(new_n1217, new_n1216, new_n1212);
nor_4  g00832(new_n1218, new_n1217, new_n1006);
nor_4  g00833(new_n1219, new_n1218, new_n1001);
nor_4  g00834(new_n1220, new_n1219, new_n995);
nor_4  g00835(new_n1221, new_n1220, new_n990);
nor_4  g00836(new_n1222_1, new_n1221, new_n985);
nor_4  g00837(new_n1223, new_n1222_1, new_n979);
nor_4  g00838(new_n1224, new_n1223, new_n974);
nor_4  g00839(new_n1225, new_n1224, new_n968);
nor_4  g00840(new_n1226, new_n1225, new_n965);
nor_4  g00841(new_n1227, new_n1226, new_n961);
nor_4  g00842(new_n1228, new_n1227, new_n958);
nor_4  g00843(new_n1229, new_n1228, new_n953);
not_3  g00844(new_n1230, new_n1229);
nand_4 g00845(new_n1231, new_n1230, new_n948_1);
nand_4 g00846(new_n1232, new_n1231, new_n943);
nand_4 g00847(new_n1233, new_n1232, new_n938);
nand_4 g00848(new_n1234, new_n1233, new_n934);
nand_4 g00849(new_n1235, new_n1234, new_n929);
nand_4 g00850(new_n1236, new_n1235, new_n925);
nand_4 g00851(new_n1237, new_n1236, n10080);
nor_4  g00852(n46, new_n1237, new_n921);
not_3  g00853(new_n1239, new_n612);
not_3  g00854(new_n1240, new_n606);
not_3  g00855(new_n1241, new_n600);
not_3  g00856(new_n1242, new_n580);
not_3  g00857(new_n1243, new_n585);
not_3  g00858(new_n1244, new_n592);
not_3  g00859(new_n1245, n13509);
nand_4 g00860(new_n1246, new_n1245, new_n386);
nor_4  g00861(new_n1247, new_n1246, new_n913);
not_3  g00862(new_n1248, new_n1247);
nor_4  g00863(new_n1249, n5046, n394);
not_3  g00864(new_n1250, new_n1249);
nor_4  g00865(new_n1251, new_n1250, new_n905);
not_3  g00866(new_n1252, new_n1251);
not_3  g00867(new_n1253, new_n906);
not_3  g00868(new_n1254, n5950);
nor_4  g00869(new_n1255, n12927, new_n1254);
nor_4  g00870(new_n1256, new_n1255, new_n1253);
not_3  g00871(new_n1257, new_n1256);
nor_4  g00872(new_n1258, n12927, n8649);
not_3  g00873(new_n1259, new_n1258);
nor_4  g00874(new_n1260, new_n1259, new_n898);
not_3  g00875(new_n1261, new_n1260);
nor_4  g00876(new_n1262, new_n893, n6946);
nor_4  g00877(new_n1263, n6946, n5077);
nor_4  g00878(new_n1264, new_n1263, new_n1262);
nor_4  g00879(new_n1265_1, new_n1264, n7941);
not_3  g00880(new_n1266, new_n1265_1);
not_3  g00881(new_n1267, n3910);
nor_4  g00882(new_n1268_1, new_n1267, n674);
nand_4 g00883(new_n1269, new_n893, new_n891);
nor_4  g00884(new_n1270, new_n1269, new_n1268_1);
not_3  g00885(new_n1271, new_n1270);
nor_4  g00886(new_n1272, new_n878, n11854);
nor_4  g00887(new_n1273, n8439, n844);
not_3  g00888(new_n1274, new_n1273);
nor_4  g00889(new_n1275, new_n1274, new_n1272);
not_3  g00890(new_n1276, new_n1275);
nor_4  g00891(new_n1277, n10278, new_n871);
nor_4  g00892(new_n1278, n10278, n7272);
nor_4  g00893(new_n1279, new_n1278, new_n1277);
nor_4  g00894(new_n1280, new_n1279, n11854);
not_3  g00895(new_n1281, new_n1280);
nor_4  g00896(new_n1282, n12782, n7748);
not_3  g00897(new_n1283, new_n1282);
nor_4  g00898(new_n1284, new_n1283, new_n866);
nor_4  g00899(new_n1285, new_n416, n6114);
nor_4  g00900(new_n1286, n9026, n6114);
nor_4  g00901(new_n1287, new_n1286, new_n1285);
nor_4  g00902(new_n1288, new_n1287, n4292);
nand_4 g00903(new_n1289, n13364, new_n858);
nand_4 g00904(new_n1290, new_n1289, new_n414);
nor_4  g00905(new_n1291, new_n1290, n9186);
nand_4 g00906(new_n1292, new_n861, new_n858);
not_3  g00907(new_n1293, n11756);
nor_4  g00908(new_n1294, n13511, new_n1293);
nor_4  g00909(new_n1295, new_n1294, new_n1292);
nor_4  g00910(new_n1296, n13511, n666);
not_3  g00911(new_n1297, new_n1296);
nor_4  g00912(new_n1298, new_n1297, new_n847);
not_3  g00913(new_n1299, new_n848);
not_3  g00914(new_n1300, n8397);
nor_4  g00915(new_n1301, n14464, new_n1300);
nor_4  g00916(new_n1302, new_n1301, new_n1299);
nor_4  g00917(new_n1303, n14408, n14303);
not_3  g00918(new_n1304, new_n1303);
nor_4  g00919(new_n1305, new_n1304, new_n838);
not_3  g00920(new_n1306, n3673);
nor_4  g00921(new_n1307, n6586, new_n1306);
nor_4  g00922(new_n1308, n6586, n6460);
nor_4  g00923(new_n1309, new_n1308, new_n1307);
nor_4  g00924(new_n1310, new_n1309, n4225);
not_3  g00925(new_n1311, n10446);
not_3  g00926(new_n1312, n4175);
nand_4 g00927(new_n1313, new_n1312, n498);
nand_4 g00928(new_n1314, new_n1313, new_n1311);
nor_4  g00929(new_n1315, new_n1314, n13000);
nand_4 g00930(new_n1316, new_n829, new_n1312);
nor_4  g00931(new_n1317, new_n1316, new_n824);
not_3  g00932(new_n1318, n1637);
not_3  g00933(new_n1319, n8552);
nand_4 g00934(new_n1320, new_n1319, n8486);
nand_4 g00935(new_n1321, new_n1320, new_n1318);
nor_4  g00936(new_n1322, new_n1321, n10750);
nor_4  g00937(new_n1323, n6480, n3263);
not_3  g00938(new_n1324, new_n1323);
nor_4  g00939(new_n1325, new_n1324, new_n815);
nor_4  g00940(new_n1326, n4615, n730);
not_3  g00941(new_n1327, new_n1326);
nor_4  g00942(new_n1328, new_n1327, new_n806);
not_3  g00943(new_n1329_1, new_n807);
not_3  g00944(new_n1330, n9936);
nor_4  g00945(new_n1331, new_n1330, n2615);
nor_4  g00946(new_n1332, new_n1331, new_n1329_1);
nor_4  g00947(new_n1333, n2615, n1093);
not_3  g00948(new_n1334, new_n1333);
nor_4  g00949(new_n1335, new_n1334, new_n792);
nor_4  g00950(new_n1336, n6517, n427);
not_3  g00951(new_n1337, new_n1336);
nor_4  g00952(new_n1338, new_n1337, new_n784);
nor_4  g00953(new_n1339, n6758, n4282);
nor_4  g00954(new_n1340, new_n1339, new_n921);
nor_4  g00955(new_n1341, new_n1340, n977);
nor_4  g00956(new_n1342, n10378, n4147);
not_3  g00957(new_n1343, new_n1342);
nor_4  g00958(new_n1344, new_n1343, new_n770);
not_3  g00959(new_n1345, new_n771);
nor_4  g00960(new_n1346, n9544, new_n930);
nor_4  g00961(new_n1347_1, new_n1346, new_n1345);
nor_4  g00962(new_n1348, n12321, n9544);
not_3  g00963(new_n1349, new_n1348);
nor_4  g00964(new_n1350, new_n1349, new_n762);
nor_4  g00965(new_n1351, new_n939, new_n936);
nor_4  g00966(new_n1352, new_n1351, n3166);
nand_4 g00967(new_n1353, new_n754, new_n935);
nor_4  g00968(new_n1354, new_n1353, new_n748);
nor_4  g00969(new_n1355, n10945, n9555);
nor_4  g00970(new_n1356, new_n1355, new_n945);
nor_4  g00971(new_n1357, new_n1356, n3972);
nor_4  g00972(new_n1358, n10736, n6555);
not_3  g00973(new_n1359, new_n1358);
nor_4  g00974(new_n1360, new_n1359, new_n740);
nor_4  g00975(new_n1361, n12829, n4131);
nor_4  g00976(new_n1362, new_n1361, new_n955);
nor_4  g00977(new_n1363, new_n1362, n6693);
not_3  g00978(new_n1364, n10407);
nor_4  g00979(new_n1365, new_n1364, n10051);
nand_4 g00980(new_n1366, new_n954, new_n484);
nor_4  g00981(new_n1367, new_n1366, new_n1365);
not_3  g00982(new_n1368, n10051);
nand_4 g00983(new_n1369, new_n733, new_n1368);
not_3  g00984(new_n1370, n5014);
nor_4  g00985(new_n1371, n11158, new_n1370);
nor_4  g00986(new_n1372, new_n1371, new_n1369);
not_3  g00987(new_n1373, n11143);
nand_4 g00988(new_n1374, new_n1373, new_n725);
not_3  g00989(new_n1375, n11158);
nand_4 g00990(new_n1376, new_n1373, n6436);
nand_4 g00991(new_n1377, new_n1376, new_n1375);
nor_4  g00992(new_n1378, new_n1377, n11590);
nand_4 g00993(new_n1379, new_n1378, new_n1374);
nand_4 g00994(new_n1380, new_n1379, new_n1372);
nand_4 g00995(new_n1381, new_n1380, new_n1367);
nand_4 g00996(new_n1382, new_n1381, new_n1363);
nand_4 g00997(new_n1383, new_n1382, new_n1360);
nand_4 g00998(new_n1384, new_n1383, new_n1357);
nand_4 g00999(new_n1385, new_n1384, new_n1354);
nand_4 g01000(new_n1386, new_n1385, new_n1352);
nand_4 g01001(new_n1387, new_n1386, new_n1350);
nand_4 g01002(new_n1388, new_n1387, new_n1347_1);
nand_4 g01003(new_n1389, new_n1388, new_n1344);
nand_4 g01004(new_n1390, new_n1389, new_n1341);
nand_4 g01005(new_n1391, new_n1390, new_n1338);
not_3  g01006(new_n1392, new_n793);
not_3  g01007(new_n1393, n9893);
nor_4  g01008(new_n1394, new_n1393, n6517);
nor_4  g01009(new_n1395, new_n1394, new_n1392);
nand_4 g01010(new_n1396, new_n1395, new_n1391);
nand_4 g01011(new_n1397, new_n1396, new_n1335);
nand_4 g01012(new_n1398, new_n1397, new_n1332);
nand_4 g01013(new_n1399, new_n1398, new_n1328);
not_3  g01014(new_n1400, new_n816);
not_3  g01015(new_n1401, n4785);
nor_4  g01016(new_n1402, new_n1401, n730);
nor_4  g01017(new_n1403, new_n1402, new_n1400);
nand_4 g01018(new_n1404, new_n1403, new_n1399);
nand_4 g01019(new_n1405, new_n1404, new_n1325);
not_3  g01020(new_n1406, n3263);
nor_4  g01021(new_n1407, n8997, new_n1406);
nor_4  g01022(new_n1408, n8997, n6791);
nor_4  g01023(new_n1409, new_n1408, new_n1407);
nor_4  g01024(new_n1410, new_n1409, n3532);
nand_4 g01025(new_n1411, new_n1410, new_n1405);
nand_4 g01026(new_n1412, new_n452, new_n445);
nor_4  g01027(new_n1413, new_n1412, n8552);
nand_4 g01028(new_n1414, new_n1413, new_n1411);
nand_4 g01029(new_n1415, new_n1414, new_n1322);
nand_4 g01030(new_n1416, new_n1415, new_n1317);
nand_4 g01031(new_n1417, new_n1416, new_n1315);
nand_4 g01032(new_n1418, new_n435, new_n1306);
nor_4  g01033(new_n1419, new_n1418, new_n441);
nand_4 g01034(new_n1420, new_n1419, new_n1417);
nand_4 g01035(new_n1421, new_n1420, new_n1310);
nand_4 g01036(new_n1422, new_n1421, new_n1305);
not_3  g01037(new_n1423, n13636);
not_3  g01038(new_n1424, n14303);
nand_4 g01039(new_n1425, n14483, new_n1424);
nand_4 g01040(new_n1426, new_n1425, new_n1423);
nor_4  g01041(new_n1427, new_n1426, n11930);
nand_4 g01042(new_n1428, new_n1427, new_n1422);
not_3  g01043(new_n1429, n14464);
nand_4 g01044(new_n1430, new_n1429, new_n420);
nor_4  g01045(new_n1431, new_n1430, new_n426);
nand_4 g01046(new_n1432, new_n1431, new_n1428);
nand_4 g01047(new_n1433, new_n1432, new_n1302);
nand_4 g01048(new_n1434, new_n1433, new_n1298);
nand_4 g01049(new_n1435, new_n1434, new_n1295);
nand_4 g01050(new_n1436, new_n1435, new_n1291);
nand_4 g01051(new_n1437, new_n1436, new_n1288);
nand_4 g01052(new_n1438, new_n1437, new_n1284);
not_3  g01053(new_n1439, new_n1438);
nor_4  g01054(new_n1440, new_n1439, new_n1281);
nor_4  g01055(new_n1441, new_n1440, new_n1276);
nand_4 g01056(new_n1442, new_n887, new_n884_1);
not_3  g01057(new_n1443, n702);
nor_4  g01058(new_n1444, n844, new_n1443);
nor_4  g01059(new_n1445, new_n1444, new_n1442);
not_3  g01060(new_n1446, new_n1445);
nor_4  g01061(new_n1447, new_n1446, new_n1441);
nor_4  g01062(new_n1448, new_n1447, new_n1271);
nor_4  g01063(new_n1449, new_n1448, new_n1266);
nor_4  g01064(new_n1450, new_n1449, new_n1261);
nor_4  g01065(new_n1451, new_n1450, new_n1257);
nor_4  g01066(new_n1452, new_n1451, new_n1252);
not_3  g01067(new_n1453, n394);
nor_4  g01068(new_n1454, n8892, new_n1453);
nor_4  g01069(new_n1455, n8892, n6362);
nor_4  g01070(new_n1456, new_n1455, new_n1454);
nor_4  g01071(new_n1457, new_n1456, n1265);
not_3  g01072(new_n1458, new_n1457);
nor_4  g01073(new_n1459, new_n1458, new_n1452);
nor_4  g01074(new_n1460, n8780, n4895);
not_3  g01075(new_n1461, new_n1460);
nor_4  g01076(new_n1462, new_n1461, new_n395);
not_3  g01077(new_n1463, new_n1462);
nor_4  g01078(new_n1464, new_n1463, new_n1459);
nor_4  g01079(new_n1465, new_n390, n5009);
nor_4  g01080(new_n1466, n8598, n5009);
nor_4  g01081(new_n1467, new_n1466, new_n1465);
nor_4  g01082(new_n1468, new_n1467, n5601);
not_3  g01083(new_n1469, new_n1468);
nor_4  g01084(new_n1470, new_n1469, new_n1464);
nor_4  g01085(new_n1471, new_n1470, new_n1248);
not_3  g01086(new_n1472, n10426);
nor_4  g01087(new_n1473, n13509, new_n1472);
nor_4  g01088(new_n1474, new_n1473, new_n588);
not_3  g01089(new_n1475, new_n1474);
nor_4  g01090(new_n1476, new_n1475, new_n1471);
nor_4  g01091(new_n1477, new_n1476, new_n1244);
nor_4  g01092(new_n1478, new_n1477, new_n1243);
nor_4  g01093(new_n1479, new_n1478, new_n1242);
nor_4  g01094(new_n1480, new_n1479, new_n1241);
nor_4  g01095(new_n1481, new_n1480, new_n1240);
nor_4  g01096(new_n1482, new_n1481, new_n1239);
not_3  g01097(new_n1483, new_n1482);
nand_4 g01098(new_n1484, new_n1483, new_n575);
nand_4 g01099(new_n1485, new_n1484, new_n619);
nand_4 g01100(new_n1486, new_n1485, new_n570);
nand_4 g01101(new_n1487, new_n1486, new_n625);
nand_4 g01102(new_n1488, new_n1487, new_n564);
nand_4 g01103(new_n1489, new_n1488, new_n632);
nand_4 g01104(new_n1490, new_n1489, new_n638);
nand_4 g01105(new_n1491, new_n1490, new_n559);
nand_4 g01106(new_n1492, new_n1491, new_n554);
nand_4 g01107(new_n1493, new_n1492, new_n646);
nand_4 g01108(new_n1494, new_n1493, new_n652);
nand_4 g01109(new_n1495, new_n1494, new_n549);
nand_4 g01110(new_n1496, new_n1495, new_n544);
nand_4 g01111(new_n1497, new_n1496, new_n660);
nand_4 g01112(new_n1498, new_n1497, new_n539);
nand_4 g01113(new_n1499, new_n1498, new_n534);
nand_4 g01114(new_n1500, new_n1499, new_n529);
nand_4 g01115(new_n1501, new_n1500, new_n668);
nand_4 g01116(new_n1502, new_n1501, new_n674_1);
nand_4 g01117(new_n1503, new_n1502, new_n681);
nand_4 g01118(new_n1504, new_n1503, new_n523);
nand_4 g01119(new_n1505, new_n1504, new_n687);
nand_4 g01120(new_n1506, new_n1505, new_n693);
nand_4 g01121(new_n1507, new_n1506, new_n699);
nand_4 g01122(new_n1508, new_n1507, new_n517);
nand_4 g01123(new_n1509, new_n1508, new_n705);
nand_4 g01124(new_n1510, new_n1509, new_n511);
nand_4 g01125(new_n1511, new_n1510, new_n711);
nand_4 g01126(new_n1512, new_n1511, new_n506);
nand_4 g01127(new_n1513, new_n1512, new_n719);
nand_4 g01128(new_n1514, new_n1513, n3833);
nor_4  g01129(n91, new_n1514, new_n497);
not_3  g01130(new_n1516, new_n1079);
not_3  g01131(new_n1517, new_n1084);
not_3  g01132(new_n1518, new_n1088);
not_3  g01133(new_n1519, new_n1091);
not_3  g01134(new_n1520, new_n1095);
not_3  g01135(new_n1521, new_n1191);
not_3  g01136(new_n1522, new_n1099);
not_3  g01137(new_n1523, new_n1102);
not_3  g01138(new_n1524, new_n1183);
not_3  g01139(new_n1525, new_n1178);
not_3  g01140(new_n1526, new_n1106);
not_3  g01141(new_n1527, new_n1111);
not_3  g01142(new_n1528, new_n1116);
not_3  g01143(new_n1529, new_n1169);
not_3  g01144(new_n1530, new_n1120);
not_3  g01145(new_n1531, new_n1164);
not_3  g01146(new_n1532, new_n1123);
not_3  g01147(new_n1533, new_n916);
not_3  g01148(new_n1534, new_n393);
not_3  g01149(new_n1535, new_n398);
not_3  g01150(new_n1536, new_n403);
not_3  g01151(new_n1537, new_n908);
nand_4 g01152(new_n1538, new_n988, new_n504);
nand_4 g01153(new_n1539, new_n1538, new_n719);
nand_4 g01154(new_n1540, new_n1539, new_n500);
nand_4 g01155(new_n1541, new_n1540, new_n727);
nand_4 g01156(new_n1542, new_n1541, new_n494);
nand_4 g01157(new_n1543, new_n1542, new_n735);
nand_4 g01158(new_n1544, new_n1543, new_n488);
nand_4 g01159(new_n1545_1, new_n1544, new_n743);
nand_4 g01160(new_n1546, new_n1545_1, new_n482);
nand_4 g01161(new_n1547, new_n1546, new_n751);
nand_4 g01162(new_n1548, new_n1547, new_n758);
nand_4 g01163(new_n1549, new_n1548, new_n765);
nand_4 g01164(new_n1550, new_n1549, new_n476);
nand_4 g01165(new_n1551, new_n1550, new_n773);
nand_4 g01166(new_n1552, new_n1551, new_n780);
nand_4 g01167(new_n1553, new_n1552, new_n787);
nand_4 g01168(new_n1554, new_n1553, new_n470);
nand_4 g01169(new_n1555, new_n1554, new_n795);
nand_4 g01170(new_n1556, new_n1555, new_n803);
nand_4 g01171(new_n1557, new_n1556, new_n809);
nand_4 g01172(new_n1558, new_n1557, new_n465);
nand_4 g01173(new_n1559, new_n1558, new_n818);
nand_4 g01174(new_n1560, new_n1559, new_n460);
nand_4 g01175(new_n1561, new_n1560, new_n455);
nand_4 g01176(new_n1562, new_n1561, new_n449);
nand_4 g01177(new_n1563, new_n1562, new_n827);
nand_4 g01178(new_n1564, new_n1563, new_n833);
nand_4 g01179(new_n1565, new_n1564, new_n444);
nand_4 g01180(new_n1566, new_n1565, new_n439);
nand_4 g01181(new_n1567, new_n1566, new_n841);
nand_4 g01182(new_n1568_1, new_n1567, new_n434);
nand_4 g01183(new_n1569, new_n1568_1, new_n429);
nand_4 g01184(new_n1570, new_n1569, new_n424);
nand_4 g01185(new_n1571, new_n1570, new_n850);
nand_4 g01186(new_n1572, new_n1571, new_n856);
nand_4 g01187(new_n1573, new_n1572, new_n863);
nand_4 g01188(new_n1574, new_n1573, new_n419);
nand_4 g01189(new_n1575, new_n1574, new_n869);
nand_4 g01190(new_n1576, new_n1575, new_n875);
nand_4 g01191(new_n1577, new_n1576, new_n881);
nand_4 g01192(new_n1578, new_n1577, new_n413);
nand_4 g01193(new_n1579, new_n1578, new_n889);
nand_4 g01194(new_n1580, new_n1579, new_n896);
nand_4 g01195(new_n1581, new_n1580, new_n901);
nand_4 g01196(new_n1582, new_n1581, new_n408);
not_3  g01197(new_n1583, new_n1582);
nor_4  g01198(new_n1584, new_n1583, new_n1537);
nor_4  g01199(new_n1585, new_n1584, new_n1536);
nor_4  g01200(new_n1586, new_n1585, new_n1535);
nor_4  g01201(new_n1587, new_n1586, new_n1534);
nor_4  g01202(new_n1588, new_n1587, new_n1533);
nor_4  g01203(new_n1589, new_n1588, new_n1532);
nor_4  g01204(new_n1590, new_n1589, new_n1531);
nor_4  g01205(new_n1591, new_n1590, new_n1530);
nor_4  g01206(new_n1592, new_n1591, new_n1529);
nor_4  g01207(new_n1593, new_n1592, new_n1528);
nor_4  g01208(new_n1594, new_n1593, new_n1527);
nor_4  g01209(new_n1595, new_n1594, new_n1526);
nor_4  g01210(new_n1596, new_n1595, new_n1525);
nor_4  g01211(new_n1597, new_n1596, new_n1524);
nor_4  g01212(new_n1598, new_n1597, new_n1523);
nor_4  g01213(new_n1599, new_n1598, new_n1522);
nor_4  g01214(new_n1600, new_n1599, new_n1521);
nor_4  g01215(new_n1601, new_n1600, new_n1520);
nor_4  g01216(new_n1602, new_n1601, new_n1519);
nor_4  g01217(new_n1603, new_n1602, new_n1518);
nor_4  g01218(new_n1604, new_n1603, new_n1517);
nor_4  g01219(new_n1605, new_n1604, new_n1516);
nor_4  g01220(new_n1606, new_n1605, new_n1075);
nor_4  g01221(new_n1607, new_n1606, new_n1071);
not_3  g01222(new_n1608, new_n1607);
nand_4 g01223(new_n1609, new_n1608, new_n1064);
nand_4 g01224(new_n1610, new_n1609, new_n1061);
nand_4 g01225(new_n1611, new_n1610, new_n1055);
nand_4 g01226(new_n1612, new_n1611, new_n1050);
nand_4 g01227(new_n1613, new_n1612, new_n1045);
nand_4 g01228(new_n1614, new_n1613, new_n1041);
nand_4 g01229(new_n1615, new_n1614, new_n1036);
nand_4 g01230(new_n1616, new_n1615, new_n1031);
nand_4 g01231(new_n1617, new_n1616, new_n1025);
nand_4 g01232(new_n1618, new_n1617, new_n1020);
nand_4 g01233(new_n1619, new_n1618, new_n1015);
nand_4 g01234(new_n1620, new_n1619, new_n1010);
nand_4 g01235(new_n1621, new_n1620, new_n1215);
nand_4 g01236(new_n1622, new_n1621, new_n1005);
nand_4 g01237(new_n1623, new_n1622, new_n1000);
nand_4 g01238(new_n1624, new_n1623, n4022);
nor_4  g01239(n126, new_n1624, new_n992);
not_3  g01240(new_n1626, new_n1363);
not_3  g01241(new_n1627, new_n1367);
not_3  g01242(new_n1628, new_n1372);
not_3  g01243(new_n1629, new_n1378);
nor_4  g01244(new_n1630, n11933, n2699);
nor_4  g01245(new_n1631, new_n1630, new_n970);
nor_4  g01246(new_n1632, new_n1631, n11143);
not_3  g01247(new_n1633, new_n1632);
nor_4  g01248(new_n1634, n9154, n3833);
not_3  g01249(new_n1635, new_n1634);
nor_4  g01250(new_n1636, new_n1635, new_n716);
not_3  g01251(new_n1637_1, new_n1636);
nor_4  g01252(new_n1638, n11666, n8262);
nor_4  g01253(new_n1639, new_n1638, new_n981);
nor_4  g01254(new_n1640, new_n1639, n12885);
not_3  g01255(new_n1641, new_n1640);
nor_4  g01256(new_n1642, n11875, n4117);
not_3  g01257(new_n1643, new_n1642);
nor_4  g01258(new_n1644, new_n1643, new_n708);
not_3  g01259(new_n1645, new_n1644);
not_3  g01260(new_n1646, new_n709);
nor_4  g01261(new_n1647, n13814, new_n508);
nor_4  g01262(new_n1648, new_n1647, new_n1646);
not_3  g01263(new_n1649, new_n1648);
not_3  g01264(new_n1650, n8635);
nand_4 g01265(new_n1651, new_n991, new_n1650);
nor_4  g01266(new_n1652, new_n1651, new_n702_1);
not_3  g01267(new_n1653, new_n1652);
not_3  g01268(new_n1654, n737);
nand_4 g01269(new_n1655, n8463, new_n514);
nand_4 g01270(new_n1656, new_n1655, new_n1654);
nor_4  g01271(new_n1657, new_n1656, n2895);
not_3  g01272(new_n1658, new_n1657);
nor_4  g01273(new_n1659, n8800, n203);
not_3  g01274(new_n1660, new_n1659);
nor_4  g01275(new_n1661, new_n1660, new_n696);
not_3  g01276(new_n1662, new_n1661);
nor_4  g01277(new_n1663, n14293, n8926);
nor_4  g01278(new_n1664, new_n1663, new_n1008);
nor_4  g01279(new_n1665, new_n1664, n8204);
not_3  g01280(new_n1666, new_n1665);
nor_4  g01281(new_n1667, n3893, n2454);
not_3  g01282(new_n1668, new_n1667);
nor_4  g01283(new_n1669, new_n1668, new_n684);
not_3  g01284(new_n1670, new_n1669);
nor_4  g01285(new_n1671, new_n1029, n3388);
nor_4  g01286(new_n1672, n4154, n3506);
not_3  g01287(new_n1673, new_n1672);
nor_4  g01288(new_n1674, new_n1673, new_n1671);
not_3  g01289(new_n1675, new_n1674);
nor_4  g01290(new_n1676, n12142, n411);
nor_4  g01291(new_n1677, new_n1676, new_n1028);
nor_4  g01292(new_n1678, new_n1677, n3388);
not_3  g01293(new_n1679, new_n1678);
nor_4  g01294(new_n1680, n12614, n8799);
not_3  g01295(new_n1681, new_n1680);
nor_4  g01296(new_n1682, new_n1681, new_n665);
not_3  g01297(new_n1683, new_n1682);
nor_4  g01298(new_n1684, n11902, n8073);
nor_4  g01299(new_n1685, new_n1684, new_n1038);
nor_4  g01300(new_n1686, new_n1685, n9252);
not_3  g01301(new_n1687, new_n1686);
nor_4  g01302(new_n1688, n13882, n6680);
not_3  g01303(new_n1689, new_n1688);
nor_4  g01304(new_n1690, new_n1689, new_n657);
not_3  g01305(new_n1691, new_n1690);
nor_4  g01306(new_n1692, n14163, n5430);
nor_4  g01307(new_n1693, new_n1692, new_n1058);
nor_4  g01308(new_n1694, new_n1693, n2164);
nor_4  g01309(new_n1695, n13295, n10630);
nor_4  g01310(new_n1696, new_n1695, new_n1067);
nor_4  g01311(new_n1697, new_n1696, n760);
nand_4 g01312(new_n1698, new_n648, new_n1066);
nor_4  g01313(new_n1699, new_n1698, new_n643);
not_3  g01314(new_n1700, n5960);
nand_4 g01315(new_n1701, n6258, new_n636);
nand_4 g01316(new_n1702_1, new_n1701, new_n1700);
nor_4  g01317(new_n1703, new_n1702_1, n6007);
nand_4 g01318(new_n1704, new_n634, new_n636);
nor_4  g01319(new_n1705, new_n1704, new_n629);
not_3  g01320(new_n1706, new_n630);
nor_4  g01321(new_n1707, new_n1187, n5225);
nor_4  g01322(new_n1708, new_n1707, new_n1706);
not_3  g01323(new_n1709, n5225);
nand_4 g01324(new_n1710, new_n560, new_n1709);
nor_4  g01325(new_n1711, new_n1710, new_n622);
not_3  g01326(new_n1712, new_n623);
not_3  g01327(new_n1713, n9314);
nor_4  g01328(new_n1714, n13109, new_n1713);
nor_4  g01329(new_n1715, new_n1714, new_n1712);
nor_4  g01330(new_n1716, n13109, n74);
not_3  g01331(new_n1717, new_n1716);
nor_4  g01332(new_n1718, new_n1717, new_n616);
not_3  g01333(new_n1719, new_n1181);
nor_4  g01334(new_n1720, new_n1719, new_n1174);
nor_4  g01335(new_n1721, new_n1720, n4774);
nor_4  g01336(new_n1722, n5033, n1763);
not_3  g01337(new_n1723, new_n1722);
nor_4  g01338(new_n1724, new_n1723, new_n609);
nor_4  g01339(new_n1725, new_n1107, new_n1104);
nor_4  g01340(new_n1726, new_n1725, n6054);
nor_4  g01341(new_n1727, n13102, n7354);
not_3  g01342(new_n1728, new_n1727);
nor_4  g01343(new_n1729, new_n1728, new_n597);
nor_4  g01344(new_n1730, n13625, n11961);
nor_4  g01345(new_n1731, new_n1730, new_n1113);
nor_4  g01346(new_n1732, new_n1731, n14475);
not_3  g01347(new_n1733, n1027);
nand_4 g01348(new_n1734, n11842, new_n1733);
nand_4 g01349(new_n1735, new_n1734, new_n576);
nor_4  g01350(new_n1736, new_n1735, n7832);
nor_4  g01351(new_n1737, new_n1161, new_n1117);
nor_4  g01352(new_n1738, new_n1737, n1027);
nor_4  g01353(new_n1739_1, new_n1245, n8002);
not_3  g01354(new_n1740, n2201);
nand_4 g01355(new_n1741, new_n589, new_n1740);
nor_4  g01356(new_n1742, new_n1741, new_n1739_1);
nand_4 g01357(new_n1743, new_n1472, new_n587);
not_3  g01358(new_n1744, n5601);
nor_4  g01359(new_n1745, new_n1744, n2674);
nor_4  g01360(new_n1746, new_n1745, new_n1743);
nand_4 g01361(new_n1747, new_n391, new_n386);
nor_4  g01362(new_n1748, new_n1747, new_n1465);
nor_4  g01363(new_n1749, n8598, n1265);
nor_4  g01364(new_n1750, new_n1749, new_n389_1);
nor_4  g01365(new_n1751, new_n1750, n5009);
nor_4  g01366(new_n1752, n4895, n1268);
not_3  g01367(new_n1753, new_n1752);
nor_4  g01368(new_n1754, new_n1753, new_n1454);
not_3  g01369(new_n1755, new_n1455);
not_3  g01370(new_n1756, n4039);
nor_4  g01371(new_n1757, n5046, new_n1756);
nor_4  g01372(new_n1758, new_n1757, new_n1755);
not_3  g01373(new_n1759, n11529);
nand_4 g01374(new_n1760, n12927, new_n1759);
nand_4 g01375(new_n1761, new_n1760, new_n399);
nor_4  g01376(new_n1762, new_n1761, n10050);
nand_4 g01377(new_n1763_1, new_n1759, new_n1254);
not_3  g01378(new_n1764, n7941);
nor_4  g01379(new_n1765, n8649, new_n1764);
nor_4  g01380(new_n1766, new_n1765, new_n1763_1);
nor_4  g01381(new_n1767, n13944, n8649);
not_3  g01382(new_n1768, new_n1767);
nor_4  g01383(new_n1769, new_n1768, new_n1262);
not_3  g01384(new_n1770, n844);
nor_4  g01385(new_n1771, n8873, new_n1770);
nor_4  g01386(new_n1772, n5467, n3910);
not_3  g01387(new_n1773, new_n1772);
nor_4  g01388(new_n1774, new_n1773, new_n1771);
nor_4  g01389(new_n1775, n11854, n702);
nor_4  g01390(new_n1776_1, new_n1775, new_n410);
nor_4  g01391(new_n1777, new_n1776_1, n8873);
nor_4  g01392(new_n1778, n13186, n8439);
not_3  g01393(new_n1779, new_n1778);
nor_4  g01394(new_n1780, new_n1779, new_n1277);
not_3  g01395(new_n1781, n12782);
nor_4  g01396(new_n1782, new_n1781, n7272);
nor_4  g01397(new_n1783, n7272, n4292);
nor_4  g01398(new_n1784, new_n1783, new_n1782);
nor_4  g01399(new_n1785, new_n1784, n10278);
not_3  g01400(new_n1786, n6114);
nand_4 g01401(new_n1787, n9186, new_n1786);
nand_4 g01402(new_n1788, new_n1787, new_n417);
nor_4  g01403(new_n1789, new_n1788, n12782);
not_3  g01404(new_n1790, n13511);
nor_4  g01405(new_n1791, new_n1790, n4907);
not_3  g01406(new_n1792, n13364);
nand_4 g01407(new_n1793, new_n1792, new_n414);
nor_4  g01408(new_n1794, new_n1793, new_n1791);
not_3  g01409(new_n1795, n12012);
nand_4 g01410(new_n1796, n14464, new_n1795);
nand_4 g01411(new_n1797, new_n1796, new_n852);
nor_4  g01412(new_n1798, new_n1797, n12976);
nand_4 g01413(new_n1799, new_n1795, new_n1300);
not_3  g01414(new_n1800, n11930);
nor_4  g01415(new_n1801, new_n1800, n10147);
nor_4  g01416(new_n1802, new_n1801, new_n1799);
nor_4  g01417(new_n1803, new_n1424, n13636);
nor_4  g01418(new_n1804, n10147, n7667);
not_3  g01419(new_n1805, new_n1804);
nor_4  g01420(new_n1806, new_n1805, new_n1803);
not_3  g01421(new_n1807, n14483);
nand_4 g01422(new_n1808, new_n430, n4225);
nand_4 g01423(new_n1809, new_n1808, new_n1807);
nor_4  g01424(new_n1810, new_n1809, n13636);
nor_4  g01425(new_n1811, n14408, n5023);
nand_4 g01426(new_n1812, new_n1811, new_n1309);
nand_4 g01427(new_n1813, new_n1812, new_n1810);
nand_4 g01428(new_n1814, new_n1813, new_n1806);
nand_4 g01429(new_n1815, new_n1814, new_n1802);
nand_4 g01430(new_n1816, new_n1815, new_n1798);
nand_4 g01431(new_n1817, new_n1293, new_n861);
not_3  g01432(new_n1818, n6810);
nor_4  g01433(new_n1819, new_n1818, n666);
nor_4  g01434(new_n1820, new_n1819, new_n1817);
nand_4 g01435(new_n1821, new_n1820, new_n1816);
nand_4 g01436(new_n1822, new_n1821, new_n1794);
not_3  g01437(new_n1823, new_n1286);
nor_4  g01438(new_n1824, new_n858, n2061);
nor_4  g01439(new_n1825, new_n1824, new_n1823);
nand_4 g01440(new_n1826, new_n1825, new_n1822);
nand_4 g01441(new_n1827_1, new_n1826, new_n1789);
nand_4 g01442(new_n1828, new_n1827_1, new_n1785);
nand_4 g01443(new_n1829, new_n1828, new_n1780);
nand_4 g01444(new_n1830, new_n1829, new_n1777);
nand_4 g01445(new_n1831, new_n1830, new_n1774);
not_3  g01446(new_n1832, new_n1263);
nor_4  g01447(new_n1833, n5467, new_n884_1);
nor_4  g01448(new_n1834, new_n1833, new_n1832);
nand_4 g01449(new_n1835, new_n1834, new_n1831);
nand_4 g01450(new_n1836, new_n1835, new_n1769);
nand_4 g01451(new_n1837, new_n1836, new_n1766);
nand_4 g01452(new_n1838, new_n1837, new_n1762);
nand_4 g01453(new_n1839, new_n1838, new_n1758);
nand_4 g01454(new_n1840, new_n1839, new_n1754);
nand_4 g01455(new_n1841, new_n1840, new_n1751);
nand_4 g01456(new_n1842, new_n1841, new_n1748);
nand_4 g01457(new_n1843, new_n1842, new_n1746);
nand_4 g01458(new_n1844, new_n1843, new_n1742);
nand_4 g01459(new_n1845, new_n1844, new_n1738);
nand_4 g01460(new_n1846, new_n1845, new_n1736);
nand_4 g01461(new_n1847, new_n1846, new_n1732);
nand_4 g01462(new_n1848, new_n1847, new_n1729);
nand_4 g01463(new_n1849, new_n1848, new_n1726);
nand_4 g01464(new_n1850, new_n1849, new_n1724);
nand_4 g01465(new_n1851, new_n1850, new_n1721);
nand_4 g01466(new_n1852, new_n1851, new_n1718);
nand_4 g01467(new_n1853, new_n1852, new_n1715);
nand_4 g01468(new_n1854, new_n1853, new_n1711);
nand_4 g01469(new_n1855, new_n1854, new_n1708);
nand_4 g01470(new_n1856, new_n1855, new_n1705);
nand_4 g01471(new_n1857, new_n1856, new_n1703);
nor_4  g01472(new_n1858, n11776, n3367);
not_3  g01473(new_n1859, new_n1858);
nor_4  g01474(new_n1860, new_n1859, new_n556);
nand_4 g01475(new_n1861, new_n1860, new_n1857);
not_3  g01476(new_n1862, new_n1077);
nor_4  g01477(new_n1863, new_n1080, new_n1862);
nor_4  g01478(new_n1864, new_n1863, n7988);
nand_4 g01479(new_n1865, new_n1864, new_n1861);
nand_4 g01480(new_n1866, new_n1865, new_n1699);
nand_4 g01481(new_n1867, new_n1866, new_n1697);
not_3  g01482(new_n1868, n760);
nand_4 g01483(new_n1869, n3799, new_n1868);
nand_4 g01484(new_n1870, new_n1869, new_n1057);
nor_4  g01485(new_n1871, new_n1870, n8746);
nand_4 g01486(new_n1872, new_n1871, new_n1867);
nand_4 g01487(new_n1873, new_n1872, new_n1694);
not_3  g01488(new_n1874, new_n1873);
nor_4  g01489(new_n1875, new_n1874, new_n1691);
nor_4  g01490(new_n1876, n10466, n5943);
nor_4  g01491(new_n1877, new_n1876, new_n1048);
nor_4  g01492(new_n1878, new_n1877, n10112);
not_3  g01493(new_n1879, new_n1878);
nor_4  g01494(new_n1880, new_n1879, new_n1875);
nand_4 g01495(new_n1881, new_n527, new_n524);
nor_4  g01496(new_n1882, new_n1881, new_n531);
not_3  g01497(new_n1883, new_n1882);
nor_4  g01498(new_n1884, new_n1883, new_n1880);
nor_4  g01499(new_n1885, new_n1884, new_n1687);
nor_4  g01500(new_n1886, new_n1885, new_n1683);
nor_4  g01501(new_n1887, new_n1886, new_n1679);
nor_4  g01502(new_n1888, new_n1887, new_n1675);
nor_4  g01503(new_n1889, new_n1022, new_n1017);
nor_4  g01504(new_n1890, new_n1889, n11269);
not_3  g01505(new_n1891, new_n1890);
nor_4  g01506(new_n1892, new_n1891, new_n1888);
nor_4  g01507(new_n1893, new_n1892, new_n1670);
nor_4  g01508(new_n1894, new_n1893, new_n1666);
nor_4  g01509(new_n1895, new_n1894, new_n1662);
nor_4  g01510(new_n1896, new_n1895, new_n1658);
nor_4  g01511(new_n1897, new_n1896, new_n1653);
nor_4  g01512(new_n1898, new_n1897, new_n1649);
nor_4  g01513(new_n1899, new_n1898, new_n1645);
nor_4  g01514(new_n1900_1, new_n1899, new_n1641);
nor_4  g01515(new_n1901, new_n1900_1, new_n1637_1);
nor_4  g01516(new_n1902, new_n1901, new_n1633);
nor_4  g01517(new_n1903, new_n1902, new_n1629);
nor_4  g01518(new_n1904, new_n1903, new_n1628);
nor_4  g01519(new_n1905, new_n1904, new_n1627);
nor_4  g01520(new_n1906, new_n1905, new_n1626);
not_3  g01521(new_n1907, new_n1906);
nand_4 g01522(new_n1908, new_n1907, new_n1360);
nand_4 g01523(new_n1909, new_n1908, new_n1357);
nand_4 g01524(new_n1910, new_n1909, new_n1354);
nand_4 g01525(new_n1911, new_n1910, new_n1352);
nand_4 g01526(new_n1912, new_n1911, new_n1350);
nand_4 g01527(new_n1913, new_n1912, new_n1347_1);
nand_4 g01528(new_n1914, new_n1913, new_n1344);
nand_4 g01529(new_n1915, new_n1914, new_n1341);
nand_4 g01530(new_n1916, new_n1915, new_n1338);
nand_4 g01531(new_n1917, new_n1916, new_n1395);
nand_4 g01532(new_n1918, new_n1917, new_n1335);
nand_4 g01533(new_n1919, new_n1918, new_n1332);
nand_4 g01534(new_n1920, new_n1919, new_n1328);
nand_4 g01535(new_n1921, new_n1920, new_n1403);
nand_4 g01536(new_n1922, new_n1921, new_n1325);
nand_4 g01537(new_n1923, new_n1922, new_n1410);
nand_4 g01538(new_n1924, new_n1923, new_n1413);
nand_4 g01539(new_n1925, new_n1924, new_n1322);
nand_4 g01540(new_n1926, new_n1925, new_n1317);
nand_4 g01541(new_n1927_1, new_n1926, new_n1315);
nand_4 g01542(new_n1928, new_n1927_1, n12025);
nor_4  g01543(n278, new_n1928, new_n441);
not_3  g01544(new_n1930, new_n1289);
nand_4 g01545(new_n1931, new_n1789, new_n1823);
nand_4 g01546(new_n1932, new_n1931, new_n1785);
nand_4 g01547(new_n1933, new_n1932, new_n1780);
nand_4 g01548(new_n1934, new_n1933, new_n1777);
nand_4 g01549(new_n1935, new_n1934, new_n1774);
nand_4 g01550(new_n1936, new_n1935, new_n1834);
nand_4 g01551(new_n1937, new_n1936, new_n1769);
nand_4 g01552(new_n1938, new_n1937, new_n1766);
nand_4 g01553(new_n1939, new_n1938, new_n1762);
nand_4 g01554(new_n1940, new_n1939, new_n1758);
nand_4 g01555(new_n1941, new_n1940, new_n1754);
nand_4 g01556(new_n1942, new_n1941, new_n1751);
nand_4 g01557(new_n1943, new_n1942, new_n1748);
nand_4 g01558(new_n1944, new_n1943, new_n1746);
nand_4 g01559(new_n1945, new_n1944, new_n1742);
nand_4 g01560(new_n1946, new_n1945, new_n1738);
nand_4 g01561(new_n1947, new_n1946, new_n1736);
nand_4 g01562(new_n1948, new_n1947, new_n1732);
nand_4 g01563(new_n1949, new_n1948, new_n1729);
nand_4 g01564(new_n1950, new_n1949, new_n1726);
nand_4 g01565(new_n1951_1, new_n1950, new_n1724);
nand_4 g01566(new_n1952, new_n1951_1, new_n1721);
nand_4 g01567(new_n1953, new_n1952, new_n1718);
nand_4 g01568(new_n1954, new_n1953, new_n1715);
nand_4 g01569(new_n1955, new_n1954, new_n1711);
nand_4 g01570(new_n1956, new_n1955, new_n1708);
nand_4 g01571(new_n1957, new_n1956, new_n1705);
nand_4 g01572(new_n1958, new_n1957, new_n1703);
nand_4 g01573(new_n1959, new_n1958, new_n1860);
nand_4 g01574(new_n1960, new_n1959, new_n1864);
nand_4 g01575(new_n1961, new_n1960, new_n1699);
nand_4 g01576(new_n1962, new_n1961, new_n1697);
nand_4 g01577(new_n1963, new_n1962, new_n1871);
nand_4 g01578(new_n1964, new_n1963, new_n1694);
nand_4 g01579(new_n1965, new_n1964, new_n1690);
not_3  g01580(new_n1966, new_n1965);
nor_4  g01581(new_n1967, new_n1966, new_n1879);
nor_4  g01582(new_n1968, new_n1967, new_n1883);
nor_4  g01583(new_n1969, new_n1968, new_n1687);
nor_4  g01584(new_n1970, new_n1969, new_n1683);
nor_4  g01585(new_n1971, new_n1970, new_n1679);
nor_4  g01586(new_n1972, new_n1971, new_n1675);
nor_4  g01587(new_n1973, new_n1972, new_n1891);
nor_4  g01588(new_n1974, new_n1973, new_n1670);
nor_4  g01589(new_n1975, new_n1974, new_n1666);
nor_4  g01590(new_n1976, new_n1975, new_n1662);
nor_4  g01591(new_n1977, new_n1976, new_n1658);
nor_4  g01592(new_n1978, new_n1977, new_n1653);
nor_4  g01593(new_n1979, new_n1978, new_n1649);
nor_4  g01594(new_n1980, new_n1979, new_n1645);
nor_4  g01595(new_n1981, new_n1980, new_n1641);
nor_4  g01596(new_n1982, new_n1981, new_n1637_1);
nor_4  g01597(new_n1983, new_n1982, new_n1633);
nor_4  g01598(new_n1984, new_n1983, new_n1629);
nor_4  g01599(new_n1985, new_n1984, new_n1628);
not_3  g01600(new_n1986, new_n1985);
nand_4 g01601(new_n1987, new_n1986, new_n1367);
nand_4 g01602(new_n1988, new_n1987, new_n1363);
nand_4 g01603(new_n1989, new_n1988, new_n1360);
nand_4 g01604(new_n1990, new_n1989, new_n1357);
nand_4 g01605(new_n1991, new_n1990, new_n1354);
nand_4 g01606(new_n1992, new_n1991, new_n1352);
nand_4 g01607(new_n1993, new_n1992, new_n1350);
nand_4 g01608(new_n1994, new_n1993, new_n1347_1);
nand_4 g01609(new_n1995, new_n1994, new_n1344);
nand_4 g01610(new_n1996, new_n1995, new_n1341);
nand_4 g01611(new_n1997, new_n1996, new_n1338);
nand_4 g01612(new_n1998, new_n1997, new_n1395);
nand_4 g01613(new_n1999, new_n1998, new_n1335);
nand_4 g01614(new_n2000, new_n1999, new_n1332);
nand_4 g01615(new_n2001, new_n2000, new_n1328);
nand_4 g01616(new_n2002, new_n2001, new_n1403);
nand_4 g01617(new_n2003, new_n2002, new_n1325);
nand_4 g01618(new_n2004, new_n2003, new_n1410);
nand_4 g01619(new_n2005, new_n2004, new_n1413);
nand_4 g01620(new_n2006, new_n2005, new_n1322);
nand_4 g01621(new_n2007, new_n2006, new_n1317);
nand_4 g01622(new_n2008, new_n2007, new_n1315);
nand_4 g01623(new_n2009, new_n2008, new_n1419);
nand_4 g01624(new_n2010, new_n2009, new_n1310);
nand_4 g01625(new_n2011, new_n2010, new_n1305);
nand_4 g01626(new_n2012, new_n2011, new_n1427);
nand_4 g01627(new_n2013, new_n2012, new_n1431);
nand_4 g01628(new_n2014, new_n2013, new_n1302);
nand_4 g01629(new_n2015, new_n2014, new_n1298);
nand_4 g01630(new_n2016, new_n2015, new_n1295);
nand_4 g01631(new_n2017, new_n2016, n2061);
nor_4  g01632(n389, new_n2017, new_n1930);
not_3  g01633(new_n2019, new_n408);
not_3  g01634(new_n2020, new_n901);
not_3  g01635(new_n2021, new_n896);
not_3  g01636(new_n2022, new_n889);
not_3  g01637(new_n2023, new_n413);
not_3  g01638(new_n2024, new_n881);
not_3  g01639(new_n2025, new_n875);
not_3  g01640(new_n2026, new_n869);
not_3  g01641(new_n2027_1, new_n419);
not_3  g01642(new_n2028, new_n863);
not_3  g01643(new_n2029, new_n856);
not_3  g01644(new_n2030, new_n850);
not_3  g01645(new_n2031, new_n424);
not_3  g01646(new_n2032, new_n429);
not_3  g01647(new_n2033, new_n434);
not_3  g01648(new_n2034, new_n841);
not_3  g01649(new_n2035, new_n439);
not_3  g01650(new_n2036, new_n444);
not_3  g01651(new_n2037, new_n833);
not_3  g01652(new_n2038, new_n827);
not_3  g01653(new_n2039, new_n449);
not_3  g01654(new_n2040, new_n455);
not_3  g01655(new_n2041, new_n460);
not_3  g01656(new_n2042, new_n818);
not_3  g01657(new_n2043, new_n465);
nand_4 g01658(new_n2044, new_n1168, new_n578);
nand_4 g01659(new_n2045, new_n2044, new_n600);
nand_4 g01660(new_n2046, new_n2045, new_n606);
nand_4 g01661(new_n2047, new_n2046, new_n612);
nand_4 g01662(new_n2048_1, new_n2047, new_n575);
nand_4 g01663(new_n2049, new_n2048_1, new_n619);
nand_4 g01664(new_n2050, new_n2049, new_n570);
nand_4 g01665(new_n2051, new_n2050, new_n625);
nand_4 g01666(new_n2052, new_n2051, new_n564);
nand_4 g01667(new_n2053, new_n2052, new_n632);
nand_4 g01668(new_n2054, new_n2053, new_n638);
nand_4 g01669(new_n2055, new_n2054, new_n559);
nand_4 g01670(new_n2056, new_n2055, new_n554);
nand_4 g01671(new_n2057, new_n2056, new_n646);
nand_4 g01672(new_n2058, new_n2057, new_n652);
nand_4 g01673(new_n2059, new_n2058, new_n549);
nand_4 g01674(new_n2060, new_n2059, new_n544);
nand_4 g01675(new_n2061_1, new_n2060, new_n660);
nand_4 g01676(new_n2062, new_n2061_1, new_n539);
nand_4 g01677(new_n2063, new_n2062, new_n534);
nand_4 g01678(new_n2064, new_n2063, new_n529);
nand_4 g01679(new_n2065, new_n2064, new_n668);
nand_4 g01680(new_n2066, new_n2065, new_n674_1);
nand_4 g01681(new_n2067, new_n2066, new_n681);
nand_4 g01682(new_n2068, new_n2067, new_n523);
nand_4 g01683(new_n2069, new_n2068, new_n687);
nand_4 g01684(new_n2070, new_n2069, new_n693);
nand_4 g01685(new_n2071, new_n2070, new_n699);
nand_4 g01686(new_n2072, new_n2071, new_n517);
nand_4 g01687(new_n2073, new_n2072, new_n705);
nand_4 g01688(new_n2074, new_n2073, new_n511);
nand_4 g01689(new_n2075, new_n2074, new_n711);
nand_4 g01690(new_n2076, new_n2075, new_n506);
nand_4 g01691(new_n2077, new_n2076, new_n719);
nand_4 g01692(new_n2078, new_n2077, new_n500);
nand_4 g01693(new_n2079, new_n2078, new_n727);
nand_4 g01694(new_n2080, new_n2079, new_n494);
nand_4 g01695(new_n2081, new_n2080, new_n735);
nand_4 g01696(new_n2082, new_n2081, new_n488);
nand_4 g01697(new_n2083, new_n2082, new_n743);
nand_4 g01698(new_n2084, new_n2083, new_n482);
nand_4 g01699(new_n2085, new_n2084, new_n751);
nand_4 g01700(new_n2086, new_n2085, new_n758);
nand_4 g01701(new_n2087, new_n2086, new_n765);
nand_4 g01702(new_n2088, new_n2087, new_n476);
nand_4 g01703(new_n2089, new_n2088, new_n773);
nand_4 g01704(new_n2090, new_n2089, new_n780);
nand_4 g01705(new_n2091, new_n2090, new_n787);
nand_4 g01706(new_n2092, new_n2091, new_n470);
nand_4 g01707(new_n2093, new_n2092, new_n795);
nand_4 g01708(new_n2094, new_n2093, new_n803);
not_3  g01709(new_n2095, new_n2094);
nor_4  g01710(new_n2096, new_n2095, new_n810);
nor_4  g01711(new_n2097, new_n2096, new_n2043);
nor_4  g01712(new_n2098, new_n2097, new_n2042);
nor_4  g01713(new_n2099, new_n2098, new_n2041);
nor_4  g01714(new_n2100, new_n2099, new_n2040);
nor_4  g01715(new_n2101, new_n2100, new_n2039);
nor_4  g01716(new_n2102, new_n2101, new_n2038);
nor_4  g01717(new_n2103, new_n2102, new_n2037);
nor_4  g01718(new_n2104, new_n2103, new_n2036);
nor_4  g01719(new_n2105, new_n2104, new_n2035);
nor_4  g01720(new_n2106, new_n2105, new_n2034);
nor_4  g01721(new_n2107, new_n2106, new_n2033);
nor_4  g01722(new_n2108, new_n2107, new_n2032);
nor_4  g01723(new_n2109, new_n2108, new_n2031);
nor_4  g01724(new_n2110, new_n2109, new_n2030);
nor_4  g01725(new_n2111, new_n2110, new_n2029);
nor_4  g01726(new_n2112, new_n2111, new_n2028);
nor_4  g01727(new_n2113, new_n2112, new_n2027_1);
nor_4  g01728(new_n2114, new_n2113, new_n2026);
nor_4  g01729(new_n2115, new_n2114, new_n2025);
nor_4  g01730(new_n2116, new_n2115, new_n2024);
nor_4  g01731(new_n2117, new_n2116, new_n2023);
nor_4  g01732(new_n2118, new_n2117, new_n2022);
nor_4  g01733(new_n2119, new_n2118, new_n2021);
nor_4  g01734(new_n2120, new_n2119, new_n2020);
nor_4  g01735(new_n2121, new_n2120, new_n2019);
nor_4  g01736(new_n2122, new_n2121, new_n1537);
not_3  g01737(new_n2123, new_n2122);
nand_4 g01738(new_n2124, new_n2123, new_n403);
nand_4 g01739(new_n2125, new_n2124, new_n398);
nand_4 g01740(new_n2126_1, new_n2125, new_n393);
nand_4 g01741(new_n2127, new_n2126_1, new_n916);
nand_4 g01742(new_n2128, new_n2127, new_n1123);
nand_4 g01743(new_n2129, new_n2128, new_n1164);
nand_4 g01744(new_n2130, new_n2129, n11842);
nor_4  g01745(n451, new_n2130, new_n1117);
not_3  g01746(new_n2132, new_n1694);
not_3  g01747(new_n2133, new_n1871);
not_3  g01748(new_n2134, new_n1697);
not_3  g01749(new_n2135, new_n1699);
not_3  g01750(new_n2136, new_n1864);
not_3  g01751(new_n2137, new_n1860);
not_3  g01752(new_n2138, new_n1703);
not_3  g01753(new_n2139, new_n1705);
not_3  g01754(new_n2140, new_n1708);
not_3  g01755(new_n2141, new_n1711);
not_3  g01756(new_n2142, new_n1715);
not_3  g01757(new_n2143, new_n1718);
not_3  g01758(new_n2144, new_n1721);
not_3  g01759(new_n2145, new_n1724);
not_3  g01760(new_n2146, new_n1811);
nor_4  g01761(new_n2147, new_n2146, new_n1307);
not_3  g01762(new_n2148, new_n1308);
not_3  g01763(new_n2149, n13000);
nor_4  g01764(new_n2150, new_n2149, n12025);
nor_4  g01765(new_n2151, new_n2150, new_n2148);
nor_4  g01766(new_n2152, n10446, new_n1312);
nor_4  g01767(new_n2153, n12025, n3130);
not_3  g01768(new_n2154, new_n2153);
nor_4  g01769(new_n2155, new_n2154, new_n2152);
nor_4  g01770(new_n2156, n10750, n498);
nor_4  g01771(new_n2157, new_n2156, new_n830);
nor_4  g01772(new_n2158, new_n2157, n10446);
nor_4  g01773(new_n2159, new_n1319, n1637);
nor_4  g01774(new_n2160, n11404, n9589);
not_3  g01775(new_n2161, new_n2160);
nor_4  g01776(new_n2162, new_n2161, new_n2159);
nor_4  g01777(new_n2163, n8486, n3532);
nor_4  g01778(new_n2164_1, new_n2163, new_n446);
nor_4  g01779(new_n2165, new_n2164_1, n1637);
nor_4  g01780(new_n2166_1, n11345, n5786);
not_3  g01781(new_n2167, new_n2166_1);
nor_4  g01782(new_n2168, new_n2167, new_n1407);
nor_4  g01783(new_n2169, n10283, n6791);
nor_4  g01784(new_n2170, new_n2169, new_n457);
nor_4  g01785(new_n2171, new_n2170, n8997);
not_3  g01786(new_n2172, n3775);
nand_4 g01787(new_n2173, new_n2172, n730);
nand_4 g01788(new_n2174, new_n2173, new_n456);
nor_4  g01789(new_n2175_1, new_n2174, n9921);
nand_4 g01790(new_n2176, new_n1401, new_n2172);
not_3  g01791(new_n2177, n13561);
nor_4  g01792(new_n2178, new_n2177, n4615);
nor_4  g01793(new_n2179, new_n2178, new_n2176);
nor_4  g01794(new_n2180, new_n800, n656);
nor_4  g01795(new_n2181, n8737, n4615);
not_3  g01796(new_n2182, new_n2181);
nor_4  g01797(new_n2183, new_n2182, new_n2180);
nor_4  g01798(new_n2184, n10862, n9936);
nor_4  g01799(new_n2185, new_n2184, new_n799);
nor_4  g01800(new_n2186, new_n2185, n656);
not_3  g01801(new_n2187, n12218);
nand_4 g01802(new_n2188, new_n2187, n6517);
nand_4 g01803(new_n2189, new_n2188, new_n798);
nor_4  g01804(new_n2190, new_n2189, n6999);
nor_4  g01805(new_n2191, new_n1125, n12218);
nor_4  g01806(new_n2192, n10080, n427);
not_3  g01807(new_n2193, new_n2192);
nor_4  g01808(new_n2194, new_n2193, new_n921);
nand_4 g01809(new_n2195, new_n940, new_n938);
nand_4 g01810(new_n2196, new_n2195, new_n934);
nand_4 g01811(new_n2197, new_n2196, new_n929);
nand_4 g01812(new_n2198, new_n2197, new_n925);
nand_4 g01813(new_n2199, new_n2198, new_n2194);
nand_4 g01814(new_n2200, new_n2199, new_n2191);
nand_4 g01815(new_n2201_1, new_n2200, new_n2190);
nand_4 g01816(new_n2202, new_n2201_1, new_n2186);
nand_4 g01817(new_n2203, new_n2202, new_n2183);
nand_4 g01818(new_n2204, new_n2203, new_n2179);
nand_4 g01819(new_n2205, new_n2204, new_n2175_1);
nand_4 g01820(new_n2206, new_n2205, new_n2171);
nand_4 g01821(new_n2207, new_n2206, new_n2168);
nand_4 g01822(new_n2208, new_n2207, new_n2165);
nand_4 g01823(new_n2209, new_n2208, new_n2162);
nand_4 g01824(new_n2210, new_n2209, new_n2158);
nand_4 g01825(new_n2211, new_n2210, new_n2155);
nand_4 g01826(new_n2212, new_n2211, new_n2151);
nand_4 g01827(new_n2213, new_n2212, new_n2147);
nand_4 g01828(new_n2214, new_n2213, new_n1810);
nand_4 g01829(new_n2215, new_n2214, new_n1806);
nand_4 g01830(new_n2216, new_n2215, new_n1802);
nand_4 g01831(new_n2217, new_n2216, new_n1798);
nand_4 g01832(new_n2218, new_n2217, new_n1820);
nand_4 g01833(new_n2219, new_n2218, new_n1794);
nand_4 g01834(new_n2220, new_n2219, new_n1825);
nand_4 g01835(new_n2221, new_n2220, new_n1789);
nand_4 g01836(new_n2222, new_n2221, new_n1785);
nand_4 g01837(new_n2223_1, new_n2222, new_n1780);
nand_4 g01838(new_n2224, new_n2223_1, new_n1777);
nand_4 g01839(new_n2225, new_n2224, new_n1774);
nand_4 g01840(new_n2226, new_n2225, new_n1834);
nand_4 g01841(new_n2227, new_n2226, new_n1769);
nand_4 g01842(new_n2228, new_n2227, new_n1766);
nand_4 g01843(new_n2229, new_n2228, new_n1762);
nand_4 g01844(new_n2230, new_n2229, new_n1758);
nand_4 g01845(new_n2231, new_n2230, new_n1754);
nand_4 g01846(new_n2232, new_n2231, new_n1751);
nand_4 g01847(new_n2233, new_n2232, new_n1748);
nand_4 g01848(new_n2234, new_n2233, new_n1746);
nand_4 g01849(new_n2235, new_n2234, new_n1742);
nand_4 g01850(new_n2236, new_n2235, new_n1738);
nand_4 g01851(new_n2237, new_n2236, new_n1736);
nand_4 g01852(new_n2238, new_n2237, new_n1732);
nand_4 g01853(new_n2239, new_n2238, new_n1729);
nand_4 g01854(new_n2240, new_n2239, new_n1726);
not_3  g01855(new_n2241, new_n2240);
nor_4  g01856(new_n2242, new_n2241, new_n2145);
nor_4  g01857(new_n2243, new_n2242, new_n2144);
nor_4  g01858(new_n2244, new_n2243, new_n2143);
nor_4  g01859(new_n2245, new_n2244, new_n2142);
nor_4  g01860(new_n2246, new_n2245, new_n2141);
nor_4  g01861(new_n2247, new_n2246, new_n2140);
nor_4  g01862(new_n2248, new_n2247, new_n2139);
nor_4  g01863(new_n2249, new_n2248, new_n2138);
nor_4  g01864(new_n2250, new_n2249, new_n2137);
nor_4  g01865(new_n2251, new_n2250, new_n2136);
nor_4  g01866(new_n2252, new_n2251, new_n2135);
nor_4  g01867(new_n2253, new_n2252, new_n2134);
nor_4  g01868(new_n2254, new_n2253, new_n2133);
nor_4  g01869(new_n2255, new_n2254, new_n2132);
nor_4  g01870(new_n2256, new_n2255, new_n1691);
nor_4  g01871(new_n2257, new_n2256, new_n1879);
nor_4  g01872(new_n2258, new_n2257, new_n1883);
nor_4  g01873(new_n2259, new_n2258, new_n1687);
nor_4  g01874(new_n2260, new_n2259, new_n1683);
nor_4  g01875(new_n2261, new_n2260, new_n1679);
nor_4  g01876(new_n2262, new_n2261, new_n1675);
nor_4  g01877(new_n2263, new_n2262, new_n1891);
nor_4  g01878(new_n2264, new_n2263, new_n1670);
nor_4  g01879(new_n2265, new_n2264, new_n1666);
not_3  g01880(new_n2266, new_n2265);
nand_4 g01881(new_n2267, new_n2266, new_n1661);
nand_4 g01882(new_n2268, new_n2267, new_n1657);
nand_4 g01883(new_n2269, new_n2268, new_n1652);
nand_4 g01884(new_n2270, new_n2269, new_n1648);
nand_4 g01885(new_n2271, new_n2270, new_n1644);
nand_4 g01886(new_n2272, new_n2271, new_n1640);
nand_4 g01887(new_n2273, new_n2272, new_n1636);
nand_4 g01888(new_n2274, new_n2273, new_n1632);
nand_4 g01889(new_n2275, new_n2274, new_n1378);
nand_4 g01890(new_n2276, new_n2275, new_n1372);
nand_4 g01891(new_n2277, new_n2276, new_n1367);
nand_4 g01892(new_n2278, new_n2277, new_n1363);
nand_4 g01893(new_n2279, new_n2278, new_n1360);
nand_4 g01894(new_n2280, new_n2279, new_n1357);
nand_4 g01895(new_n2281, new_n2280, n10615);
nor_4  g01896(n490, new_n2281, new_n748);
not_3  g01897(new_n2283, new_n1726);
not_3  g01898(new_n2284, new_n1729);
not_3  g01899(new_n2285, new_n1732);
not_3  g01900(new_n2286, new_n1736);
not_3  g01901(new_n2287, new_n1738);
not_3  g01902(new_n2288, new_n1742);
not_3  g01903(new_n2289, new_n1746);
not_3  g01904(new_n2290, new_n1748);
not_3  g01905(new_n2291, new_n1751);
not_3  g01906(new_n2292, new_n1754);
not_3  g01907(new_n2293, new_n1758);
not_3  g01908(new_n2294, new_n1762);
not_3  g01909(new_n2295, new_n1766);
not_3  g01910(new_n2296, new_n1769);
not_3  g01911(new_n2297, new_n1834);
not_3  g01912(new_n2298, new_n1774);
not_3  g01913(new_n2299, new_n1777);
not_3  g01914(new_n2300, new_n1780);
not_3  g01915(new_n2301, new_n1785);
not_3  g01916(new_n2302, new_n1789);
not_3  g01917(new_n2303, new_n1825);
not_3  g01918(new_n2304, new_n1794);
not_3  g01919(new_n2305, new_n1820);
not_3  g01920(new_n2306, new_n1695);
nand_4 g01921(new_n2307, new_n2306, new_n1070);
nand_4 g01922(new_n2308, new_n2307, new_n1064);
nand_4 g01923(new_n2309, new_n2308, new_n1061);
nand_4 g01924(new_n2310, new_n2309, new_n1055);
nand_4 g01925(new_n2311_1, new_n2310, new_n1050);
nand_4 g01926(new_n2312, new_n2311_1, new_n1045);
nand_4 g01927(new_n2313, new_n2312, new_n1041);
nand_4 g01928(new_n2314, new_n2313, new_n1036);
nand_4 g01929(new_n2315, new_n2314, new_n1031);
nand_4 g01930(new_n2316, new_n2315, new_n1025);
nand_4 g01931(new_n2317, new_n2316, new_n1020);
nand_4 g01932(new_n2318, new_n2317, new_n1015);
nand_4 g01933(new_n2319, new_n2318, new_n1010);
nand_4 g01934(new_n2320, new_n2319, new_n1215);
nand_4 g01935(new_n2321, new_n2320, new_n1005);
nand_4 g01936(new_n2322, new_n2321, new_n1000);
nand_4 g01937(new_n2323, new_n2322, new_n994);
nand_4 g01938(new_n2324, new_n2323, new_n989);
nand_4 g01939(new_n2325, new_n2324, new_n984);
nand_4 g01940(new_n2326, new_n2325, new_n978);
nand_4 g01941(new_n2327, new_n2326, new_n973);
nand_4 g01942(new_n2328, new_n2327, new_n967);
nand_4 g01943(new_n2329, new_n2328, new_n964);
nand_4 g01944(new_n2330, new_n2329, new_n960);
nand_4 g01945(new_n2331, new_n2330, new_n957);
nand_4 g01946(new_n2332, new_n2331, new_n952);
nand_4 g01947(new_n2333, new_n2332, new_n948_1);
nand_4 g01948(new_n2334_1, new_n2333, new_n943);
nand_4 g01949(new_n2335, new_n2334_1, new_n938);
nand_4 g01950(new_n2336, new_n2335, new_n934);
nand_4 g01951(new_n2337, new_n2336, new_n929);
nand_4 g01952(new_n2338, new_n2337, new_n925);
nand_4 g01953(new_n2339, new_n2338, new_n2194);
nand_4 g01954(new_n2340, new_n2339, new_n2191);
nand_4 g01955(new_n2341, new_n2340, new_n2190);
nand_4 g01956(new_n2342, new_n2341, new_n2186);
nand_4 g01957(new_n2343, new_n2342, new_n2183);
nand_4 g01958(new_n2344, new_n2343, new_n2179);
nand_4 g01959(new_n2345, new_n2344, new_n2175_1);
nand_4 g01960(new_n2346, new_n2345, new_n2171);
nand_4 g01961(new_n2347, new_n2346, new_n2168);
nand_4 g01962(new_n2348, new_n2347, new_n2165);
nand_4 g01963(new_n2349, new_n2348, new_n2162);
nand_4 g01964(new_n2350, new_n2349, new_n2158);
nand_4 g01965(new_n2351, new_n2350, new_n2155);
nand_4 g01966(new_n2352, new_n2351, new_n2151);
nand_4 g01967(new_n2353, new_n2352, new_n2147);
nand_4 g01968(new_n2354, new_n2353, new_n1810);
nand_4 g01969(new_n2355, new_n2354, new_n1806);
nand_4 g01970(new_n2356, new_n2355, new_n1802);
nand_4 g01971(new_n2357, new_n2356, new_n1798);
not_3  g01972(new_n2358, new_n2357);
nor_4  g01973(new_n2359, new_n2358, new_n2305);
nor_4  g01974(new_n2360, new_n2359, new_n2304);
nor_4  g01975(new_n2361, new_n2360, new_n2303);
nor_4  g01976(new_n2362, new_n2361, new_n2302);
nor_4  g01977(new_n2363, new_n2362, new_n2301);
nor_4  g01978(new_n2364, new_n2363, new_n2300);
nor_4  g01979(new_n2365, new_n2364, new_n2299);
nor_4  g01980(new_n2366, new_n2365, new_n2298);
nor_4  g01981(new_n2367, new_n2366, new_n2297);
nor_4  g01982(new_n2368, new_n2367, new_n2296);
nor_4  g01983(new_n2369, new_n2368, new_n2295);
nor_4  g01984(new_n2370, new_n2369, new_n2294);
nor_4  g01985(new_n2371, new_n2370, new_n2293);
nor_4  g01986(new_n2372, new_n2371, new_n2292);
nor_4  g01987(new_n2373, new_n2372, new_n2291);
nor_4  g01988(new_n2374, new_n2373, new_n2290);
nor_4  g01989(new_n2375, new_n2374, new_n2289);
nor_4  g01990(new_n2376, new_n2375, new_n2288);
nor_4  g01991(new_n2377, new_n2376, new_n2287);
nor_4  g01992(new_n2378, new_n2377, new_n2286);
nor_4  g01993(new_n2379, new_n2378, new_n2285);
nor_4  g01994(new_n2380, new_n2379, new_n2284);
nor_4  g01995(new_n2381, new_n2380, new_n2283);
nor_4  g01996(new_n2382, new_n2381, new_n2145);
nor_4  g01997(new_n2383, new_n2382, new_n2144);
nor_4  g01998(new_n2384, new_n2383, new_n2143);
nor_4  g01999(new_n2385, new_n2384, new_n2142);
not_3  g02000(new_n2386, new_n2385);
nand_4 g02001(new_n2387, new_n2386, new_n1711);
nand_4 g02002(new_n2388, new_n2387, new_n1708);
nand_4 g02003(new_n2389, new_n2388, new_n1705);
nand_4 g02004(new_n2390, new_n2389, new_n1703);
nand_4 g02005(new_n2391, new_n2390, new_n1860);
nand_4 g02006(new_n2392, new_n2391, new_n1864);
nand_4 g02007(new_n2393, new_n2392, n5185);
nor_4  g02008(n543, new_n2393, new_n643);
not_3  g02009(new_n2395, new_n1284);
not_3  g02010(new_n2396, new_n1288);
not_3  g02011(new_n2397, new_n1291);
not_3  g02012(new_n2398, new_n1295);
not_3  g02013(new_n2399, new_n1298);
not_3  g02014(new_n2400, new_n1302);
not_3  g02015(new_n2401, new_n1431);
not_3  g02016(new_n2402, new_n1427);
not_3  g02017(new_n2403, new_n1305);
not_3  g02018(new_n2404, new_n1310);
not_3  g02019(new_n2405, new_n1419);
not_3  g02020(new_n2406, new_n1315);
not_3  g02021(new_n2407_1, new_n1317);
not_3  g02022(new_n2408, new_n1322);
not_3  g02023(new_n2409, new_n1413);
not_3  g02024(new_n2410, new_n1410);
not_3  g02025(new_n2411, new_n1325);
not_3  g02026(new_n2412, new_n1403);
not_3  g02027(new_n2413, new_n1328);
nand_4 g02028(new_n2414, new_n1716, new_n618);
nand_4 g02029(new_n2415, new_n2414, new_n1715);
nand_4 g02030(new_n2416, new_n2415, new_n1711);
nand_4 g02031(new_n2417, new_n2416, new_n1708);
nand_4 g02032(new_n2418, new_n2417, new_n1705);
nand_4 g02033(new_n2419, new_n2418, new_n1703);
nand_4 g02034(new_n2420, new_n2419, new_n1860);
nand_4 g02035(new_n2421, new_n2420, new_n1864);
nand_4 g02036(new_n2422, new_n2421, new_n1699);
nand_4 g02037(new_n2423, new_n2422, new_n1697);
nand_4 g02038(new_n2424, new_n2423, new_n1871);
nand_4 g02039(new_n2425, new_n2424, new_n1694);
nand_4 g02040(new_n2426, new_n2425, new_n1690);
nand_4 g02041(new_n2427, new_n2426, new_n1878);
nand_4 g02042(new_n2428, new_n2427, new_n1882);
nand_4 g02043(new_n2429, new_n2428, new_n1686);
nand_4 g02044(new_n2430, new_n2429, new_n1682);
nand_4 g02045(new_n2431, new_n2430, new_n1678);
nand_4 g02046(new_n2432, new_n2431, new_n1674);
nand_4 g02047(new_n2433, new_n2432, new_n1890);
nand_4 g02048(new_n2434, new_n2433, new_n1669);
nand_4 g02049(new_n2435, new_n2434, new_n1665);
nand_4 g02050(new_n2436, new_n2435, new_n1661);
nand_4 g02051(new_n2437, new_n2436, new_n1657);
nand_4 g02052(new_n2438, new_n2437, new_n1652);
nand_4 g02053(new_n2439, new_n2438, new_n1648);
nand_4 g02054(new_n2440, new_n2439, new_n1644);
nand_4 g02055(new_n2441, new_n2440, new_n1640);
nand_4 g02056(new_n2442, new_n2441, new_n1636);
nand_4 g02057(new_n2443, new_n2442, new_n1632);
nand_4 g02058(new_n2444, new_n2443, new_n1378);
nand_4 g02059(new_n2445, new_n2444, new_n1372);
nand_4 g02060(new_n2446, new_n2445, new_n1367);
nand_4 g02061(new_n2447, new_n2446, new_n1363);
nand_4 g02062(new_n2448, new_n2447, new_n1360);
nand_4 g02063(new_n2449, new_n2448, new_n1357);
nand_4 g02064(new_n2450, new_n2449, new_n1354);
nand_4 g02065(new_n2451, new_n2450, new_n1352);
nand_4 g02066(new_n2452, new_n2451, new_n1350);
nand_4 g02067(new_n2453, new_n2452, new_n1347_1);
nand_4 g02068(new_n2454_1, new_n2453, new_n1344);
nand_4 g02069(new_n2455, new_n2454_1, new_n1341);
nand_4 g02070(new_n2456, new_n2455, new_n1338);
nand_4 g02071(new_n2457, new_n2456, new_n1395);
nand_4 g02072(new_n2458, new_n2457, new_n1335);
nand_4 g02073(new_n2459, new_n2458, new_n1332);
not_3  g02074(new_n2460, new_n2459);
nor_4  g02075(new_n2461, new_n2460, new_n2413);
nor_4  g02076(new_n2462, new_n2461, new_n2412);
nor_4  g02077(new_n2463, new_n2462, new_n2411);
nor_4  g02078(new_n2464, new_n2463, new_n2410);
nor_4  g02079(new_n2465, new_n2464, new_n2409);
nor_4  g02080(new_n2466, new_n2465, new_n2408);
nor_4  g02081(new_n2467, new_n2466, new_n2407_1);
nor_4  g02082(new_n2468, new_n2467, new_n2406);
nor_4  g02083(new_n2469, new_n2468, new_n2405);
nor_4  g02084(new_n2470, new_n2469, new_n2404);
nor_4  g02085(new_n2471, new_n2470, new_n2403);
nor_4  g02086(new_n2472, new_n2471, new_n2402);
nor_4  g02087(new_n2473, new_n2472, new_n2401);
nor_4  g02088(new_n2474, new_n2473, new_n2400);
nor_4  g02089(new_n2475, new_n2474, new_n2399);
nor_4  g02090(new_n2476, new_n2475, new_n2398);
nor_4  g02091(new_n2477, new_n2476, new_n2397);
nor_4  g02092(new_n2478, new_n2477, new_n2396);
nor_4  g02093(new_n2479, new_n2478, new_n2395);
nor_4  g02094(new_n2480, new_n2479, new_n1281);
nor_4  g02095(new_n2481, new_n2480, new_n1276);
nor_4  g02096(new_n2482, new_n2481, new_n1446);
nor_4  g02097(new_n2483, new_n2482, new_n1271);
nor_4  g02098(new_n2484, new_n2483, new_n1266);
not_3  g02099(new_n2485, new_n2484);
nand_4 g02100(new_n2486, new_n2485, new_n1260);
nand_4 g02101(new_n2487, new_n2486, new_n1256);
nand_4 g02102(new_n2488, new_n2487, new_n1251);
nand_4 g02103(new_n2489, new_n2488, new_n1457);
nand_4 g02104(new_n2490, new_n2489, new_n1462);
nand_4 g02105(new_n2491, new_n2490, new_n1468);
nand_4 g02106(new_n2492, new_n2491, new_n1247);
nand_4 g02107(new_n2493, new_n2492, new_n1474);
nand_4 g02108(new_n2494, new_n2493, new_n592);
nand_4 g02109(new_n2495, new_n2494, new_n585);
nand_4 g02110(new_n2496, new_n2495, new_n580);
nand_4 g02111(new_n2497, new_n2496, new_n600);
nand_4 g02112(new_n2498, new_n2497, new_n606);
nand_4 g02113(new_n2499, new_n2498, new_n612);
nand_4 g02114(new_n2500, new_n2499, n5033);
nor_4  g02115(n682, new_n2500, new_n572);
not_3  g02116(new_n2502, new_n1810);
not_3  g02117(new_n2503, new_n2147);
not_3  g02118(new_n2504, new_n2151);
not_3  g02119(new_n2505, new_n2155);
not_3  g02120(new_n2506, new_n2158);
not_3  g02121(new_n2507, new_n2162);
not_3  g02122(new_n2508, new_n2165);
not_3  g02123(new_n2509, new_n2168);
not_3  g02124(new_n2510, new_n2171);
not_3  g02125(new_n2511, new_n2175_1);
not_3  g02126(new_n2512, new_n2179);
not_3  g02127(new_n2513, new_n2183);
not_3  g02128(new_n2514, new_n2186);
not_3  g02129(new_n2515, new_n2190);
not_3  g02130(new_n2516, new_n2191);
not_3  g02131(new_n2517, new_n2194);
not_3  g02132(new_n2518, new_n925);
not_3  g02133(new_n2519, new_n929);
not_3  g02134(new_n2520, new_n934);
nand_4 g02135(new_n2521, new_n1188, new_n1095);
nand_4 g02136(new_n2522, new_n2521, new_n1091);
nand_4 g02137(new_n2523, new_n2522, new_n1088);
nand_4 g02138(new_n2524, new_n2523, new_n1084);
nand_4 g02139(new_n2525, new_n2524, new_n1079);
nand_4 g02140(new_n2526, new_n2525, new_n1074);
nand_4 g02141(new_n2527, new_n2526, new_n1070);
nand_4 g02142(new_n2528, new_n2527, new_n1064);
nand_4 g02143(new_n2529, new_n2528, new_n1061);
nand_4 g02144(new_n2530, new_n2529, new_n1055);
nand_4 g02145(new_n2531, new_n2530, new_n1050);
nand_4 g02146(new_n2532, new_n2531, new_n1045);
nand_4 g02147(new_n2533, new_n2532, new_n1041);
nand_4 g02148(new_n2534, new_n2533, new_n1036);
nand_4 g02149(new_n2535, new_n2534, new_n1031);
nand_4 g02150(new_n2536, new_n2535, new_n1025);
nand_4 g02151(new_n2537, new_n2536, new_n1020);
nand_4 g02152(new_n2538, new_n2537, new_n1015);
nand_4 g02153(new_n2539, new_n2538, new_n1010);
nand_4 g02154(new_n2540, new_n2539, new_n1215);
nand_4 g02155(new_n2541, new_n2540, new_n1005);
nand_4 g02156(new_n2542, new_n2541, new_n1000);
nand_4 g02157(new_n2543, new_n2542, new_n994);
nand_4 g02158(new_n2544, new_n2543, new_n989);
nand_4 g02159(new_n2545, new_n2544, new_n984);
nand_4 g02160(new_n2546, new_n2545, new_n978);
nand_4 g02161(new_n2547, new_n2546, new_n973);
nand_4 g02162(new_n2548, new_n2547, new_n967);
nand_4 g02163(new_n2549, new_n2548, new_n964);
nand_4 g02164(new_n2550, new_n2549, new_n960);
nand_4 g02165(new_n2551, new_n2550, new_n957);
nand_4 g02166(new_n2552, new_n2551, new_n952);
nand_4 g02167(new_n2553, new_n2552, new_n948_1);
nand_4 g02168(new_n2554, new_n2553, new_n943);
nand_4 g02169(new_n2555, new_n2554, new_n938);
not_3  g02170(new_n2556_1, new_n2555);
nor_4  g02171(new_n2557, new_n2556_1, new_n2520);
nor_4  g02172(new_n2558, new_n2557, new_n2519);
nor_4  g02173(new_n2559_1, new_n2558, new_n2518);
nor_4  g02174(new_n2560, new_n2559_1, new_n2517);
nor_4  g02175(new_n2561, new_n2560, new_n2516);
nor_4  g02176(new_n2562, new_n2561, new_n2515);
nor_4  g02177(new_n2563, new_n2562, new_n2514);
nor_4  g02178(new_n2564, new_n2563, new_n2513);
nor_4  g02179(new_n2565, new_n2564, new_n2512);
nor_4  g02180(new_n2566, new_n2565, new_n2511);
nor_4  g02181(new_n2567, new_n2566, new_n2510);
nor_4  g02182(new_n2568, new_n2567, new_n2509);
nor_4  g02183(new_n2569, new_n2568, new_n2508);
nor_4  g02184(new_n2570, new_n2569, new_n2507);
nor_4  g02185(new_n2571, new_n2570, new_n2506);
nor_4  g02186(new_n2572_1, new_n2571, new_n2505);
nor_4  g02187(new_n2573_1, new_n2572_1, new_n2504);
nor_4  g02188(new_n2574, new_n2573_1, new_n2503);
nor_4  g02189(new_n2575, new_n2574, new_n2502);
not_3  g02190(new_n2576, new_n2575);
nand_4 g02191(new_n2577, new_n2576, new_n1806);
nand_4 g02192(new_n2578, new_n2577, new_n1802);
nand_4 g02193(new_n2579, new_n2578, new_n1798);
nand_4 g02194(new_n2580, new_n2579, new_n1820);
nand_4 g02195(new_n2581, new_n2580, new_n1794);
nand_4 g02196(new_n2582, new_n2581, new_n1825);
nand_4 g02197(new_n2583, new_n2582, new_n1789);
nand_4 g02198(new_n2584, new_n2583, new_n1785);
nand_4 g02199(new_n2585, new_n2584, new_n1780);
nand_4 g02200(new_n2586, new_n2585, new_n1777);
nand_4 g02201(new_n2587, new_n2586, new_n1774);
nand_4 g02202(new_n2588, new_n2587, new_n1834);
nand_4 g02203(new_n2589, new_n2588, new_n1769);
nand_4 g02204(new_n2590, new_n2589, new_n1766);
nand_4 g02205(new_n2591, new_n2590, new_n1762);
nand_4 g02206(new_n2592, new_n2591, new_n1758);
nand_4 g02207(new_n2593, new_n2592, new_n1754);
nand_4 g02208(new_n2594, new_n2593, new_n1751);
nand_4 g02209(new_n2595, new_n2594, new_n1748);
nand_4 g02210(new_n2596, new_n2595, new_n1746);
nand_4 g02211(new_n2597, new_n2596, new_n1742);
nand_4 g02212(new_n2598, new_n2597, new_n1738);
nand_4 g02213(new_n2599, new_n2598, new_n1736);
nand_4 g02214(new_n2600, new_n2599, new_n1732);
nand_4 g02215(new_n2601, new_n2600, new_n1729);
nand_4 g02216(new_n2602, new_n2601, new_n1726);
nand_4 g02217(new_n2603, new_n2602, new_n1724);
nand_4 g02218(new_n2604, new_n2603, new_n1721);
nand_4 g02219(new_n2605, new_n2604, new_n1718);
nand_4 g02220(new_n2606, new_n2605, new_n1715);
nand_4 g02221(new_n2607, new_n2606, n13224);
nor_4  g02222(n884, new_n2607, new_n622);
not_3  g02223(new_n2609, new_n1332);
not_3  g02224(new_n2610, new_n1335);
not_3  g02225(new_n2611, new_n1395);
nand_4 g02226(new_n2612, new_n1743, new_n1742);
nand_4 g02227(new_n2613, new_n2612, new_n1738);
nand_4 g02228(new_n2614, new_n2613, new_n1736);
nand_4 g02229(new_n2615_1, new_n2614, new_n1732);
nand_4 g02230(new_n2616, new_n2615_1, new_n1729);
nand_4 g02231(new_n2617, new_n2616, new_n1726);
nand_4 g02232(new_n2618, new_n2617, new_n1724);
nand_4 g02233(new_n2619, new_n2618, new_n1721);
nand_4 g02234(new_n2620, new_n2619, new_n1718);
nand_4 g02235(new_n2621, new_n2620, new_n1715);
nand_4 g02236(new_n2622, new_n2621, new_n1711);
nand_4 g02237(new_n2623, new_n2622, new_n1708);
nand_4 g02238(new_n2624, new_n2623, new_n1705);
nand_4 g02239(new_n2625, new_n2624, new_n1703);
nand_4 g02240(new_n2626, new_n2625, new_n1860);
nand_4 g02241(new_n2627, new_n2626, new_n1864);
nand_4 g02242(new_n2628, new_n2627, new_n1699);
nand_4 g02243(new_n2629, new_n2628, new_n1697);
nand_4 g02244(new_n2630, new_n2629, new_n1871);
nand_4 g02245(new_n2631, new_n2630, new_n1694);
nand_4 g02246(new_n2632, new_n2631, new_n1690);
nand_4 g02247(new_n2633, new_n2632, new_n1878);
nand_4 g02248(new_n2634, new_n2633, new_n1882);
nand_4 g02249(new_n2635, new_n2634, new_n1686);
nand_4 g02250(new_n2636, new_n2635, new_n1682);
nand_4 g02251(new_n2637, new_n2636, new_n1678);
nand_4 g02252(new_n2638, new_n2637, new_n1674);
nand_4 g02253(new_n2639, new_n2638, new_n1890);
nand_4 g02254(new_n2640, new_n2639, new_n1669);
nand_4 g02255(new_n2641, new_n2640, new_n1665);
nand_4 g02256(new_n2642, new_n2641, new_n1661);
nand_4 g02257(new_n2643, new_n2642, new_n1657);
nand_4 g02258(new_n2644, new_n2643, new_n1652);
nand_4 g02259(new_n2645, new_n2644, new_n1648);
nand_4 g02260(new_n2646, new_n2645, new_n1644);
nand_4 g02261(new_n2647, new_n2646, new_n1640);
nand_4 g02262(new_n2648, new_n2647, new_n1636);
nand_4 g02263(new_n2649, new_n2648, new_n1632);
nand_4 g02264(new_n2650, new_n2649, new_n1378);
nand_4 g02265(new_n2651, new_n2650, new_n1372);
nand_4 g02266(new_n2652, new_n2651, new_n1367);
nand_4 g02267(new_n2653, new_n2652, new_n1363);
nand_4 g02268(new_n2654, new_n2653, new_n1360);
nand_4 g02269(new_n2655, new_n2654, new_n1357);
nand_4 g02270(new_n2656, new_n2655, new_n1354);
nand_4 g02271(new_n2657, new_n2656, new_n1352);
nand_4 g02272(new_n2658, new_n2657, new_n1350);
nand_4 g02273(new_n2659, new_n2658, new_n1347_1);
nand_4 g02274(new_n2660, new_n2659, new_n1344);
nand_4 g02275(new_n2661, new_n2660, new_n1341);
nand_4 g02276(new_n2662, new_n2661, new_n1338);
not_3  g02277(new_n2663, new_n2662);
nor_4  g02278(new_n2664, new_n2663, new_n2611);
nor_4  g02279(new_n2665, new_n2664, new_n2610);
nor_4  g02280(new_n2666, new_n2665, new_n2609);
nor_4  g02281(new_n2667, new_n2666, new_n2413);
nor_4  g02282(new_n2668, new_n2667, new_n2412);
nor_4  g02283(new_n2669, new_n2668, new_n2411);
nor_4  g02284(new_n2670, new_n2669, new_n2410);
nor_4  g02285(new_n2671, new_n2670, new_n2409);
nor_4  g02286(new_n2672_1, new_n2671, new_n2408);
nor_4  g02287(new_n2673, new_n2672_1, new_n2407_1);
nor_4  g02288(new_n2674_1, new_n2673, new_n2406);
nor_4  g02289(new_n2675, new_n2674_1, new_n2405);
nor_4  g02290(new_n2676, new_n2675, new_n2404);
nor_4  g02291(new_n2677, new_n2676, new_n2403);
nor_4  g02292(new_n2678, new_n2677, new_n2402);
nor_4  g02293(new_n2679, new_n2678, new_n2401);
nor_4  g02294(new_n2680, new_n2679, new_n2400);
nor_4  g02295(new_n2681, new_n2680, new_n2399);
nor_4  g02296(new_n2682, new_n2681, new_n2398);
nor_4  g02297(new_n2683, new_n2682, new_n2397);
nor_4  g02298(new_n2684, new_n2683, new_n2396);
nor_4  g02299(new_n2685, new_n2684, new_n2395);
nor_4  g02300(new_n2686, new_n2685, new_n1281);
nor_4  g02301(new_n2687, new_n2686, new_n1276);
nor_4  g02302(new_n2688, new_n2687, new_n1446);
nor_4  g02303(new_n2689, new_n2688, new_n1271);
nor_4  g02304(new_n2690, new_n2689, new_n1266);
not_3  g02305(new_n2691, new_n2690);
nand_4 g02306(new_n2692, new_n2691, new_n1260);
nand_4 g02307(new_n2693, new_n2692, new_n1256);
nand_4 g02308(new_n2694, new_n2693, new_n1251);
nand_4 g02309(new_n2695, new_n2694, new_n1457);
nand_4 g02310(new_n2696, new_n2695, new_n1462);
nand_4 g02311(new_n2697, new_n2696, new_n1468);
nand_4 g02312(new_n2698, new_n2697, n2674);
nor_4  g02313(n948, new_n2698, new_n913);
nand_4 g02314(new_n2700, new_n1356, new_n946);
nand_4 g02315(new_n2701, new_n2700, new_n943);
nand_4 g02316(new_n2702, new_n2701, new_n938);
nand_4 g02317(new_n2703, new_n2702, new_n934);
nand_4 g02318(new_n2704, new_n2703, new_n929);
nand_4 g02319(new_n2705, new_n2704, new_n925);
nand_4 g02320(new_n2706, new_n2705, new_n2194);
nand_4 g02321(new_n2707, new_n2706, new_n2191);
nand_4 g02322(new_n2708, new_n2707, new_n2190);
nand_4 g02323(new_n2709, new_n2708, new_n2186);
nand_4 g02324(new_n2710, new_n2709, new_n2183);
nand_4 g02325(new_n2711, new_n2710, new_n2179);
nand_4 g02326(new_n2712, new_n2711, new_n2175_1);
nand_4 g02327(new_n2713, new_n2712, new_n2171);
nand_4 g02328(new_n2714, new_n2713, new_n2168);
nand_4 g02329(new_n2715, new_n2714, new_n2165);
nand_4 g02330(new_n2716, new_n2715, new_n2162);
nand_4 g02331(new_n2717, new_n2716, new_n2158);
nand_4 g02332(new_n2718, new_n2717, new_n2155);
nand_4 g02333(new_n2719, new_n2718, new_n2151);
nand_4 g02334(new_n2720, new_n2719, new_n2147);
nand_4 g02335(new_n2721, new_n2720, new_n1810);
nand_4 g02336(new_n2722, new_n2721, new_n1806);
nand_4 g02337(new_n2723, new_n2722, new_n1802);
nand_4 g02338(new_n2724, new_n2723, new_n1798);
nand_4 g02339(new_n2725, new_n2724, new_n1820);
nand_4 g02340(new_n2726, new_n2725, new_n1794);
nand_4 g02341(new_n2727, new_n2726, new_n1825);
nand_4 g02342(new_n2728, new_n2727, new_n1789);
nand_4 g02343(new_n2729, new_n2728, new_n1785);
nand_4 g02344(new_n2730, new_n2729, new_n1780);
nand_4 g02345(new_n2731, new_n2730, new_n1777);
nand_4 g02346(new_n2732, new_n2731, new_n1774);
nand_4 g02347(new_n2733, new_n2732, new_n1834);
nand_4 g02348(new_n2734_1, new_n2733, new_n1769);
nand_4 g02349(new_n2735, new_n2734_1, new_n1766);
nand_4 g02350(new_n2736, new_n2735, new_n1762);
nand_4 g02351(new_n2737, new_n2736, new_n1758);
nand_4 g02352(new_n2738, new_n2737, new_n1754);
nand_4 g02353(new_n2739, new_n2738, new_n1751);
nand_4 g02354(new_n2740, new_n2739, new_n1748);
nand_4 g02355(new_n2741, new_n2740, new_n1746);
nand_4 g02356(new_n2742, new_n2741, new_n1742);
nand_4 g02357(new_n2743, new_n2742, new_n1738);
nand_4 g02358(new_n2744, new_n2743, new_n1736);
nand_4 g02359(new_n2745, new_n2744, new_n1732);
not_3  g02360(new_n2746, new_n2745);
nor_4  g02361(new_n2747, new_n2746, new_n2284);
nor_4  g02362(new_n2748, new_n2747, new_n2283);
nor_4  g02363(new_n2749, new_n2748, new_n2145);
nor_4  g02364(new_n2750, new_n2749, new_n2144);
nor_4  g02365(new_n2751, new_n2750, new_n2143);
nor_4  g02366(new_n2752, new_n2751, new_n2142);
nor_4  g02367(new_n2753, new_n2752, new_n2141);
nor_4  g02368(new_n2754, new_n2753, new_n2140);
nor_4  g02369(new_n2755, new_n2754, new_n2139);
nor_4  g02370(new_n2756, new_n2755, new_n2138);
nor_4  g02371(new_n2757, new_n2756, new_n2137);
nor_4  g02372(new_n2758, new_n2757, new_n2136);
nor_4  g02373(new_n2759, new_n2758, new_n2135);
nor_4  g02374(new_n2760, new_n2759, new_n2134);
nor_4  g02375(new_n2761, new_n2760, new_n2133);
nor_4  g02376(new_n2762, new_n2761, new_n2132);
nor_4  g02377(new_n2763, new_n2762, new_n1691);
nor_4  g02378(new_n2764, new_n2763, new_n1879);
nor_4  g02379(new_n2765, new_n2764, new_n1883);
nor_4  g02380(new_n2766, new_n2765, new_n1687);
nor_4  g02381(new_n2767, new_n2766, new_n1683);
nor_4  g02382(new_n2768, new_n2767, new_n1679);
nor_4  g02383(new_n2769, new_n2768, new_n1675);
nor_4  g02384(new_n2770, new_n2769, new_n1891);
not_3  g02385(new_n2771, new_n2770);
nand_4 g02386(new_n2772, new_n2771, new_n1669);
nand_4 g02387(new_n2773, new_n2772, new_n1665);
nand_4 g02388(new_n2774, new_n2773, new_n1661);
nand_4 g02389(new_n2775, new_n2774, new_n1657);
nand_4 g02390(new_n2776, new_n2775, new_n1652);
nand_4 g02391(new_n2777, new_n2776, new_n1648);
nand_4 g02392(new_n2778, new_n2777, new_n1644);
nand_4 g02393(new_n2779, new_n2778, new_n1640);
nand_4 g02394(new_n2780, new_n2779, new_n1636);
nand_4 g02395(new_n2781, new_n2780, new_n1632);
nand_4 g02396(new_n2782, new_n2781, new_n1378);
nand_4 g02397(new_n2783, new_n2782, new_n1372);
nand_4 g02398(new_n2784, new_n2783, new_n1367);
nand_4 g02399(new_n2785, new_n2784, new_n1363);
nand_4 g02400(new_n2786, new_n2785, n6555);
nor_4  g02401(n1094, new_n2786, new_n740);
not_3  g02402(new_n2788, new_n1798);
not_3  g02403(new_n2789, new_n1802);
not_3  g02404(new_n2790, new_n1806);
not_3  g02405(new_n2791, new_n1745);
nand_4 g02406(new_n2792, new_n2791, new_n1472);
nand_4 g02407(new_n2793, new_n2792, new_n1121);
nand_4 g02408(new_n2794, new_n2793, new_n1164);
nand_4 g02409(new_n2795, new_n2794, new_n1120);
nand_4 g02410(new_n2796, new_n2795, new_n1169);
nand_4 g02411(new_n2797, new_n2796, new_n1116);
nand_4 g02412(new_n2798, new_n2797, new_n1111);
nand_4 g02413(new_n2799, new_n2798, new_n1106);
nand_4 g02414(new_n2800, new_n2799, new_n1178);
nand_4 g02415(new_n2801, new_n2800, new_n1183);
nand_4 g02416(new_n2802, new_n2801, new_n1102);
nand_4 g02417(new_n2803, new_n2802, new_n1099);
nand_4 g02418(new_n2804, new_n2803, new_n1191);
nand_4 g02419(new_n2805, new_n2804, new_n1095);
nand_4 g02420(new_n2806, new_n2805, new_n1091);
nand_4 g02421(new_n2807, new_n2806, new_n1088);
nand_4 g02422(new_n2808, new_n2807, new_n1084);
nand_4 g02423(new_n2809, new_n2808, new_n1079);
nand_4 g02424(new_n2810, new_n2809, new_n1074);
nand_4 g02425(new_n2811, new_n2810, new_n1070);
nand_4 g02426(new_n2812, new_n2811, new_n1064);
nand_4 g02427(new_n2813, new_n2812, new_n1061);
nand_4 g02428(new_n2814, new_n2813, new_n1055);
nand_4 g02429(new_n2815, new_n2814, new_n1050);
nand_4 g02430(new_n2816, new_n2815, new_n1045);
nand_4 g02431(new_n2817, new_n2816, new_n1041);
nand_4 g02432(new_n2818, new_n2817, new_n1036);
nand_4 g02433(new_n2819, new_n2818, new_n1031);
nand_4 g02434(new_n2820, new_n2819, new_n1025);
nand_4 g02435(new_n2821, new_n2820, new_n1020);
nand_4 g02436(new_n2822, new_n2821, new_n1015);
nand_4 g02437(new_n2823, new_n2822, new_n1010);
nand_4 g02438(new_n2824, new_n2823, new_n1215);
nand_4 g02439(new_n2825, new_n2824, new_n1005);
nand_4 g02440(new_n2826, new_n2825, new_n1000);
nand_4 g02441(new_n2827, new_n2826, new_n994);
nand_4 g02442(new_n2828, new_n2827, new_n989);
nand_4 g02443(new_n2829, new_n2828, new_n984);
nand_4 g02444(new_n2830, new_n2829, new_n978);
nand_4 g02445(new_n2831, new_n2830, new_n973);
nand_4 g02446(new_n2832, new_n2831, new_n967);
nand_4 g02447(new_n2833, new_n2832, new_n964);
nand_4 g02448(new_n2834, new_n2833, new_n960);
nand_4 g02449(new_n2835, new_n2834, new_n957);
nand_4 g02450(new_n2836, new_n2835, new_n952);
nand_4 g02451(new_n2837, new_n2836, new_n948_1);
nand_4 g02452(new_n2838, new_n2837, new_n943);
nand_4 g02453(new_n2839, new_n2838, new_n938);
nand_4 g02454(new_n2840, new_n2839, new_n934);
nand_4 g02455(new_n2841, new_n2840, new_n929);
nand_4 g02456(new_n2842, new_n2841, new_n925);
not_3  g02457(new_n2843, new_n2842);
nor_4  g02458(new_n2844, new_n2843, new_n2517);
nor_4  g02459(new_n2845, new_n2844, new_n2516);
nor_4  g02460(new_n2846, new_n2845, new_n2515);
nor_4  g02461(new_n2847, new_n2846, new_n2514);
nor_4  g02462(new_n2848, new_n2847, new_n2513);
nor_4  g02463(new_n2849, new_n2848, new_n2512);
nor_4  g02464(new_n2850, new_n2849, new_n2511);
nor_4  g02465(new_n2851, new_n2850, new_n2510);
nor_4  g02466(new_n2852, new_n2851, new_n2509);
nor_4  g02467(new_n2853, new_n2852, new_n2508);
nor_4  g02468(new_n2854, new_n2853, new_n2507);
nor_4  g02469(new_n2855, new_n2854, new_n2506);
nor_4  g02470(new_n2856, new_n2855, new_n2505);
nor_4  g02471(new_n2857, new_n2856, new_n2504);
nor_4  g02472(new_n2858, new_n2857, new_n2503);
nor_4  g02473(new_n2859, new_n2858, new_n2502);
nor_4  g02474(new_n2860, new_n2859, new_n2790);
nor_4  g02475(new_n2861, new_n2860, new_n2789);
nor_4  g02476(new_n2862, new_n2861, new_n2788);
nor_4  g02477(new_n2863, new_n2862, new_n2305);
nor_4  g02478(new_n2864, new_n2863, new_n2304);
nor_4  g02479(new_n2865, new_n2864, new_n2303);
nor_4  g02480(new_n2866, new_n2865, new_n2302);
nor_4  g02481(new_n2867, new_n2866, new_n2301);
nor_4  g02482(new_n2868, new_n2867, new_n2300);
not_3  g02483(new_n2869, new_n2868);
nand_4 g02484(new_n2870, new_n2869, new_n1777);
nand_4 g02485(new_n2871, new_n2870, new_n1774);
nand_4 g02486(new_n2872, new_n2871, new_n1834);
nand_4 g02487(new_n2873, new_n2872, new_n1769);
nand_4 g02488(new_n2874, new_n2873, new_n1766);
nand_4 g02489(new_n2875, new_n2874, new_n1762);
nand_4 g02490(new_n2876, new_n2875, new_n1758);
nand_4 g02491(new_n2877, new_n2876, new_n1754);
nand_4 g02492(new_n2878, new_n2877, new_n1751);
nand_4 g02493(new_n2879, new_n2878, n12270);
nor_4  g02494(n1122, new_n2879, new_n1465);
not_3  g02495(new_n2881, n9543);
not_3  g02496(new_n2882, new_n1083);
nand_4 g02497(new_n2883, new_n2882, new_n2881);
nand_4 g02498(new_n2884, new_n2883, new_n552);
nand_4 g02499(new_n2885, new_n2884, new_n646);
nand_4 g02500(new_n2886, new_n2885, new_n652);
nand_4 g02501(new_n2887, new_n2886, new_n549);
nand_4 g02502(new_n2888, new_n2887, new_n544);
nand_4 g02503(new_n2889, new_n2888, new_n660);
nand_4 g02504(new_n2890, new_n2889, new_n539);
nand_4 g02505(new_n2891, new_n2890, new_n534);
nand_4 g02506(new_n2892, new_n2891, new_n529);
nand_4 g02507(new_n2893, new_n2892, new_n668);
nand_4 g02508(new_n2894, new_n2893, new_n674_1);
nand_4 g02509(new_n2895_1, new_n2894, new_n681);
nand_4 g02510(new_n2896, new_n2895_1, new_n523);
nand_4 g02511(new_n2897, new_n2896, new_n687);
nand_4 g02512(new_n2898, new_n2897, new_n693);
nand_4 g02513(new_n2899, new_n2898, new_n699);
nand_4 g02514(new_n2900, new_n2899, new_n517);
nand_4 g02515(new_n2901, new_n2900, new_n705);
nand_4 g02516(new_n2902, new_n2901, new_n511);
nand_4 g02517(new_n2903, new_n2902, new_n711);
nand_4 g02518(new_n2904, new_n2903, new_n506);
nand_4 g02519(new_n2905, new_n2904, new_n719);
nand_4 g02520(new_n2906, new_n2905, new_n500);
nand_4 g02521(new_n2907, new_n2906, new_n727);
nand_4 g02522(new_n2908, new_n2907, new_n494);
nand_4 g02523(new_n2909, new_n2908, new_n735);
nand_4 g02524(new_n2910, new_n2909, new_n488);
nand_4 g02525(new_n2911, new_n2910, new_n743);
nand_4 g02526(new_n2912, new_n2911, new_n482);
nand_4 g02527(new_n2913, new_n2912, new_n751);
nand_4 g02528(new_n2914, new_n2913, new_n758);
nand_4 g02529(new_n2915, new_n2914, new_n765);
nand_4 g02530(new_n2916, new_n2915, new_n476);
nand_4 g02531(new_n2917, new_n2916, new_n773);
nand_4 g02532(new_n2918, new_n2917, new_n780);
nand_4 g02533(new_n2919, new_n2918, new_n787);
nand_4 g02534(new_n2920, new_n2919, new_n470);
nand_4 g02535(new_n2921, new_n2920, new_n795);
nand_4 g02536(new_n2922, new_n2921, new_n803);
nand_4 g02537(new_n2923, new_n2922, new_n809);
nand_4 g02538(new_n2924, new_n2923, new_n465);
nand_4 g02539(new_n2925, new_n2924, new_n818);
nand_4 g02540(new_n2926, new_n2925, new_n460);
nand_4 g02541(new_n2927, new_n2926, new_n455);
nand_4 g02542(new_n2928, new_n2927, new_n449);
not_3  g02543(new_n2929, new_n2928);
nor_4  g02544(new_n2930, new_n2929, new_n2038);
nor_4  g02545(new_n2931, new_n2930, new_n2037);
nor_4  g02546(new_n2932, new_n2931, new_n2036);
nor_4  g02547(new_n2933, new_n2932, new_n2035);
nor_4  g02548(new_n2934, new_n2933, new_n2034);
nor_4  g02549(new_n2935, new_n2934, new_n2033);
nor_4  g02550(new_n2936, new_n2935, new_n2032);
nor_4  g02551(new_n2937, new_n2936, new_n2031);
nor_4  g02552(new_n2938, new_n2937, new_n2030);
nor_4  g02553(new_n2939, new_n2938, new_n2029);
nor_4  g02554(new_n2940, new_n2939, new_n2028);
nor_4  g02555(new_n2941, new_n2940, new_n2027_1);
nor_4  g02556(new_n2942, new_n2941, new_n2026);
nor_4  g02557(new_n2943, new_n2942, new_n2025);
nor_4  g02558(new_n2944, new_n2943, new_n2024);
nor_4  g02559(new_n2945, new_n2944, new_n2023);
nor_4  g02560(new_n2946, new_n2945, new_n2022);
nor_4  g02561(new_n2947, new_n2946, new_n2021);
nor_4  g02562(new_n2948, new_n2947, new_n2020);
nor_4  g02563(new_n2949, new_n2948, new_n2019);
nor_4  g02564(new_n2950, new_n2949, new_n1537);
nor_4  g02565(new_n2951, new_n2950, new_n1536);
nor_4  g02566(new_n2952, new_n2951, new_n1535);
nor_4  g02567(new_n2953, new_n2952, new_n1534);
not_3  g02568(new_n2954, new_n2953);
nand_4 g02569(new_n2955, new_n2954, new_n916);
nand_4 g02570(new_n2956, new_n2955, new_n1123);
nand_4 g02571(new_n2957, new_n2956, new_n1164);
nand_4 g02572(new_n2958, new_n2957, new_n1120);
nand_4 g02573(new_n2959, new_n2958, new_n1169);
nand_4 g02574(new_n2960, new_n2959, new_n1116);
nand_4 g02575(new_n2961, new_n2960, new_n1111);
nand_4 g02576(new_n2962, new_n2961, new_n1106);
nand_4 g02577(new_n2963, new_n2962, new_n1178);
nand_4 g02578(new_n2964, new_n2963, new_n1183);
nand_4 g02579(new_n2965, new_n2964, new_n1102);
nand_4 g02580(new_n2966, new_n2965, new_n1099);
nand_4 g02581(new_n2967, new_n2966, new_n1191);
nand_4 g02582(new_n2968, new_n2967, new_n1095);
nand_4 g02583(new_n2969, new_n2968, new_n1091);
nand_4 g02584(new_n2970, new_n2969, n271);
nor_4  g02585(n1124, new_n2970, new_n1085);
not_3  g02586(new_n2972, new_n1749);
nand_4 g02587(new_n2973, new_n2972, new_n393);
nand_4 g02588(new_n2974, new_n2973, new_n916);
nand_4 g02589(new_n2975, new_n2974, new_n1123);
nand_4 g02590(new_n2976, new_n2975, new_n1164);
nand_4 g02591(new_n2977, new_n2976, new_n1120);
nand_4 g02592(new_n2978, new_n2977, new_n1169);
nand_4 g02593(new_n2979, new_n2978, new_n1116);
nand_4 g02594(new_n2980, new_n2979, new_n1111);
nand_4 g02595(new_n2981, new_n2980, new_n1106);
nand_4 g02596(new_n2982, new_n2981, new_n1178);
nand_4 g02597(new_n2983, new_n2982, new_n1183);
nand_4 g02598(new_n2984, new_n2983, new_n1102);
nand_4 g02599(new_n2985, new_n2984, new_n1099);
nand_4 g02600(new_n2986, new_n2985, new_n1191);
nand_4 g02601(new_n2987, new_n2986, new_n1095);
nand_4 g02602(new_n2988, new_n2987, new_n1091);
nand_4 g02603(new_n2989, new_n2988, new_n1088);
nand_4 g02604(new_n2990, new_n2989, new_n1084);
nand_4 g02605(new_n2991, new_n2990, new_n1079);
nand_4 g02606(new_n2992, new_n2991, new_n1074);
nand_4 g02607(new_n2993, new_n2992, new_n1070);
nand_4 g02608(new_n2994, new_n2993, new_n1064);
nand_4 g02609(new_n2995, new_n2994, new_n1061);
nand_4 g02610(new_n2996, new_n2995, new_n1055);
nand_4 g02611(new_n2997, new_n2996, new_n1050);
nand_4 g02612(new_n2998, new_n2997, new_n1045);
nand_4 g02613(new_n2999, new_n2998, new_n1041);
nand_4 g02614(new_n3000, new_n2999, new_n1036);
nand_4 g02615(new_n3001, new_n3000, new_n1031);
nand_4 g02616(new_n3002, new_n3001, new_n1025);
nand_4 g02617(new_n3003, new_n3002, new_n1020);
nand_4 g02618(new_n3004, new_n3003, new_n1015);
nand_4 g02619(new_n3005, new_n3004, new_n1010);
nand_4 g02620(new_n3006, new_n3005, new_n1215);
nand_4 g02621(new_n3007, new_n3006, new_n1005);
nand_4 g02622(new_n3008, new_n3007, new_n1000);
nand_4 g02623(new_n3009, new_n3008, new_n994);
nand_4 g02624(new_n3010, new_n3009, new_n989);
nand_4 g02625(new_n3011, new_n3010, new_n984);
nand_4 g02626(new_n3012, new_n3011, new_n978);
nand_4 g02627(new_n3013, new_n3012, new_n973);
nand_4 g02628(new_n3014, new_n3013, new_n967);
nand_4 g02629(new_n3015, new_n3014, new_n964);
nand_4 g02630(new_n3016, new_n3015, new_n960);
nand_4 g02631(new_n3017, new_n3016, new_n957);
nand_4 g02632(new_n3018, new_n3017, new_n952);
nand_4 g02633(new_n3019, new_n3018, new_n948_1);
nand_4 g02634(new_n3020, new_n3019, new_n943);
nand_4 g02635(new_n3021, new_n3020, new_n938);
nand_4 g02636(new_n3022, new_n3021, new_n934);
nand_4 g02637(new_n3023, new_n3022, new_n929);
not_3  g02638(new_n3024, new_n3023);
nor_4  g02639(new_n3025, new_n3024, new_n2518);
nor_4  g02640(new_n3026, new_n3025, new_n2517);
nor_4  g02641(new_n3027, new_n3026, new_n2516);
nor_4  g02642(new_n3028, new_n3027, new_n2515);
nor_4  g02643(new_n3029, new_n3028, new_n2514);
nor_4  g02644(new_n3030, new_n3029, new_n2513);
nor_4  g02645(new_n3031, new_n3030, new_n2512);
nor_4  g02646(new_n3032, new_n3031, new_n2511);
nor_4  g02647(new_n3033, new_n3032, new_n2510);
nor_4  g02648(new_n3034, new_n3033, new_n2509);
nor_4  g02649(new_n3035, new_n3034, new_n2508);
nor_4  g02650(new_n3036, new_n3035, new_n2507);
nor_4  g02651(new_n3037, new_n3036, new_n2506);
nor_4  g02652(new_n3038, new_n3037, new_n2505);
nor_4  g02653(new_n3039, new_n3038, new_n2504);
nor_4  g02654(new_n3040, new_n3039, new_n2503);
nor_4  g02655(new_n3041, new_n3040, new_n2502);
nor_4  g02656(new_n3042, new_n3041, new_n2790);
nor_4  g02657(new_n3043, new_n3042, new_n2789);
nor_4  g02658(new_n3044, new_n3043, new_n2788);
nor_4  g02659(new_n3045, new_n3044, new_n2305);
nor_4  g02660(new_n3046, new_n3045, new_n2304);
nor_4  g02661(new_n3047, new_n3046, new_n2303);
nor_4  g02662(new_n3048, new_n3047, new_n2302);
nor_4  g02663(new_n3049, new_n3048, new_n2301);
nor_4  g02664(new_n3050, new_n3049, new_n2300);
nor_4  g02665(new_n3051, new_n3050, new_n2299);
not_3  g02666(new_n3052, new_n3051);
nand_4 g02667(new_n3053, new_n3052, new_n1774);
nand_4 g02668(new_n3054, new_n3053, new_n1834);
nand_4 g02669(new_n3055, new_n3054, new_n1769);
nand_4 g02670(new_n3056, new_n3055, new_n1766);
nand_4 g02671(new_n3057, new_n3056, new_n1762);
nand_4 g02672(new_n3058, new_n3057, new_n1758);
nand_4 g02673(new_n3059, new_n3058, n1268);
nor_4  g02674(n1329, new_n3059, new_n1454);
not_3  g02675(new_n3061, new_n687);
not_3  g02676(new_n3062, new_n523);
not_3  g02677(new_n3063, new_n681);
not_3  g02678(new_n3064, new_n674_1);
not_3  g02679(new_n3065, new_n668);
not_3  g02680(new_n3066, new_n529);
not_3  g02681(new_n3067, new_n534);
not_3  g02682(new_n3068, new_n539);
not_3  g02683(new_n3069, new_n660);
not_3  g02684(new_n3070, new_n544);
not_3  g02685(new_n3071, new_n549);
not_3  g02686(new_n3072, new_n652);
not_3  g02687(new_n3073, new_n646);
not_3  g02688(new_n3074, new_n554);
not_3  g02689(new_n3075, new_n559);
not_3  g02690(new_n3076, new_n638);
not_3  g02691(new_n3077, new_n632);
not_3  g02692(new_n3078, new_n564);
not_3  g02693(new_n3079, new_n625);
not_3  g02694(new_n3080, new_n570);
not_3  g02695(new_n3081, new_n619);
not_3  g02696(new_n3082, new_n575);
nand_4 g02697(new_n3083, new_n1634, new_n718);
nand_4 g02698(new_n3084, new_n3083, new_n1632);
nand_4 g02699(new_n3085, new_n3084, new_n1378);
nand_4 g02700(new_n3086, new_n3085, new_n1372);
nand_4 g02701(new_n3087, new_n3086, new_n1367);
nand_4 g02702(new_n3088, new_n3087, new_n1363);
nand_4 g02703(new_n3089, new_n3088, new_n1360);
nand_4 g02704(new_n3090_1, new_n3089, new_n1357);
nand_4 g02705(new_n3091, new_n3090_1, new_n1354);
nand_4 g02706(new_n3092, new_n3091, new_n1352);
nand_4 g02707(new_n3093, new_n3092, new_n1350);
nand_4 g02708(new_n3094, new_n3093, new_n1347_1);
nand_4 g02709(new_n3095, new_n3094, new_n1344);
nand_4 g02710(new_n3096, new_n3095, new_n1341);
nand_4 g02711(new_n3097, new_n3096, new_n1338);
nand_4 g02712(new_n3098, new_n3097, new_n1395);
nand_4 g02713(new_n3099, new_n3098, new_n1335);
nand_4 g02714(new_n3100, new_n3099, new_n1332);
nand_4 g02715(new_n3101, new_n3100, new_n1328);
nand_4 g02716(new_n3102, new_n3101, new_n1403);
nand_4 g02717(new_n3103, new_n3102, new_n1325);
nand_4 g02718(new_n3104, new_n3103, new_n1410);
nand_4 g02719(new_n3105, new_n3104, new_n1413);
nand_4 g02720(new_n3106, new_n3105, new_n1322);
nand_4 g02721(new_n3107, new_n3106, new_n1317);
nand_4 g02722(new_n3108, new_n3107, new_n1315);
nand_4 g02723(new_n3109, new_n3108, new_n1419);
nand_4 g02724(new_n3110, new_n3109, new_n1310);
nand_4 g02725(new_n3111, new_n3110, new_n1305);
nand_4 g02726(new_n3112, new_n3111, new_n1427);
nand_4 g02727(new_n3113, new_n3112, new_n1431);
nand_4 g02728(new_n3114, new_n3113, new_n1302);
nand_4 g02729(new_n3115, new_n3114, new_n1298);
nand_4 g02730(new_n3116, new_n3115, new_n1295);
nand_4 g02731(new_n3117, new_n3116, new_n1291);
nand_4 g02732(new_n3118, new_n3117, new_n1288);
nand_4 g02733(new_n3119, new_n3118, new_n1284);
nand_4 g02734(new_n3120, new_n3119, new_n1280);
nand_4 g02735(new_n3121, new_n3120, new_n1275);
nand_4 g02736(new_n3122, new_n3121, new_n1445);
nand_4 g02737(new_n3123, new_n3122, new_n1270);
nand_4 g02738(new_n3124, new_n3123, new_n1265_1);
nand_4 g02739(new_n3125, new_n3124, new_n1260);
nand_4 g02740(new_n3126, new_n3125, new_n1256);
nand_4 g02741(new_n3127, new_n3126, new_n1251);
nand_4 g02742(new_n3128, new_n3127, new_n1457);
nand_4 g02743(new_n3129, new_n3128, new_n1462);
nand_4 g02744(new_n3130_1, new_n3129, new_n1468);
nand_4 g02745(new_n3131, new_n3130_1, new_n1247);
nand_4 g02746(new_n3132, new_n3131, new_n1474);
nand_4 g02747(new_n3133, new_n3132, new_n592);
not_3  g02748(new_n3134, new_n3133);
nor_4  g02749(new_n3135, new_n3134, new_n1243);
nor_4  g02750(new_n3136, new_n3135, new_n1242);
nor_4  g02751(new_n3137, new_n3136, new_n1241);
nor_4  g02752(new_n3138, new_n3137, new_n1240);
nor_4  g02753(new_n3139, new_n3138, new_n1239);
nor_4  g02754(new_n3140, new_n3139, new_n3082);
nor_4  g02755(new_n3141, new_n3140, new_n3081);
nor_4  g02756(new_n3142, new_n3141, new_n3080);
nor_4  g02757(new_n3143, new_n3142, new_n3079);
nor_4  g02758(new_n3144, new_n3143, new_n3078);
nor_4  g02759(new_n3145, new_n3144, new_n3077);
nor_4  g02760(new_n3146, new_n3145, new_n3076);
nor_4  g02761(new_n3147, new_n3146, new_n3075);
nor_4  g02762(new_n3148, new_n3147, new_n3074);
nor_4  g02763(new_n3149, new_n3148, new_n3073);
nor_4  g02764(new_n3150, new_n3149, new_n3072);
nor_4  g02765(new_n3151, new_n3150, new_n3071);
nor_4  g02766(new_n3152, new_n3151, new_n3070);
nor_4  g02767(new_n3153, new_n3152, new_n3069);
nor_4  g02768(new_n3154, new_n3153, new_n3068);
nor_4  g02769(new_n3155, new_n3154, new_n3067);
nor_4  g02770(new_n3156, new_n3155, new_n3066);
nor_4  g02771(new_n3157, new_n3156, new_n3065);
nor_4  g02772(new_n3158, new_n3157, new_n3064);
nor_4  g02773(new_n3159, new_n3158, new_n3063);
nor_4  g02774(new_n3160, new_n3159, new_n3062);
nor_4  g02775(new_n3161, new_n3160, new_n3061);
not_3  g02776(new_n3162, new_n3161);
nand_4 g02777(new_n3163, new_n3162, new_n693);
nand_4 g02778(new_n3164, new_n3163, new_n699);
nand_4 g02779(new_n3165, new_n3164, new_n517);
nand_4 g02780(new_n3166_1, new_n3165, new_n705);
nand_4 g02781(new_n3167, new_n3166_1, new_n511);
nand_4 g02782(new_n3168, new_n3167, new_n711);
nand_4 g02783(new_n3169, new_n3168, n4117);
nor_4  g02784(n1545, new_n3169, new_n503);
not_3  g02785(new_n3171, new_n1783);
nand_4 g02786(new_n3172, new_n3171, new_n875);
nand_4 g02787(new_n3173, new_n3172, new_n881);
nand_4 g02788(new_n3174, new_n3173, new_n413);
nand_4 g02789(new_n3175, new_n3174, new_n889);
nand_4 g02790(new_n3176, new_n3175, new_n896);
nand_4 g02791(new_n3177, new_n3176, new_n901);
nand_4 g02792(new_n3178, new_n3177, new_n408);
nand_4 g02793(new_n3179, new_n3178, new_n908);
nand_4 g02794(new_n3180, new_n3179, new_n403);
nand_4 g02795(new_n3181, new_n3180, new_n398);
nand_4 g02796(new_n3182, new_n3181, new_n393);
nand_4 g02797(new_n3183, new_n3182, new_n916);
nand_4 g02798(new_n3184, new_n3183, new_n1123);
nand_4 g02799(new_n3185, new_n3184, new_n1164);
nand_4 g02800(new_n3186, new_n3185, new_n1120);
nand_4 g02801(new_n3187, new_n3186, new_n1169);
nand_4 g02802(new_n3188, new_n3187, new_n1116);
nand_4 g02803(new_n3189, new_n3188, new_n1111);
nand_4 g02804(new_n3190, new_n3189, new_n1106);
nand_4 g02805(new_n3191, new_n3190, new_n1178);
nand_4 g02806(new_n3192, new_n3191, new_n1183);
nand_4 g02807(new_n3193, new_n3192, new_n1102);
nand_4 g02808(new_n3194, new_n3193, new_n1099);
nand_4 g02809(new_n3195, new_n3194, new_n1191);
nand_4 g02810(new_n3196, new_n3195, new_n1095);
nand_4 g02811(new_n3197, new_n3196, new_n1091);
nand_4 g02812(new_n3198, new_n3197, new_n1088);
nand_4 g02813(new_n3199, new_n3198, new_n1084);
nand_4 g02814(new_n3200, new_n3199, new_n1079);
nand_4 g02815(new_n3201, new_n3200, new_n1074);
nand_4 g02816(new_n3202, new_n3201, new_n1070);
nand_4 g02817(new_n3203, new_n3202, new_n1064);
nand_4 g02818(new_n3204, new_n3203, new_n1061);
nand_4 g02819(new_n3205, new_n3204, new_n1055);
nand_4 g02820(new_n3206, new_n3205, new_n1050);
not_3  g02821(new_n3207, new_n3206);
nor_4  g02822(new_n3208, new_n3207, new_n1046);
nor_4  g02823(new_n3209, new_n3208, new_n1042);
nor_4  g02824(new_n3210, new_n3209, new_n1037);
nor_4  g02825(new_n3211, new_n3210, new_n1032);
nor_4  g02826(new_n3212, new_n3211, new_n1026);
nor_4  g02827(new_n3213, new_n3212, new_n1021);
nor_4  g02828(new_n3214, new_n3213, new_n1016);
nor_4  g02829(new_n3215, new_n3214, new_n1011);
nor_4  g02830(new_n3216, new_n3215, new_n1216);
nor_4  g02831(new_n3217, new_n3216, new_n1006);
nor_4  g02832(new_n3218, new_n3217, new_n1001);
nor_4  g02833(new_n3219, new_n3218, new_n995);
nor_4  g02834(new_n3220, new_n3219, new_n990);
nor_4  g02835(new_n3221, new_n3220, new_n985);
nor_4  g02836(new_n3222, new_n3221, new_n979);
nor_4  g02837(new_n3223, new_n3222, new_n974);
nor_4  g02838(new_n3224, new_n3223, new_n968);
nor_4  g02839(new_n3225, new_n3224, new_n965);
nor_4  g02840(new_n3226, new_n3225, new_n961);
not_3  g02841(new_n3227, new_n3226);
nand_4 g02842(new_n3228, new_n3227, new_n957);
nand_4 g02843(new_n3229, new_n3228, new_n952);
nand_4 g02844(new_n3230, new_n3229, new_n948_1);
nand_4 g02845(new_n3231, new_n3230, new_n943);
nand_4 g02846(new_n3232, new_n3231, new_n938);
nand_4 g02847(new_n3233, new_n3232, new_n934);
nand_4 g02848(new_n3234, new_n3233, new_n929);
nand_4 g02849(new_n3235, new_n3234, new_n925);
nand_4 g02850(new_n3236, new_n3235, new_n2194);
nand_4 g02851(new_n3237, new_n3236, new_n2191);
nand_4 g02852(new_n3238, new_n3237, new_n2190);
nand_4 g02853(new_n3239, new_n3238, new_n2186);
nand_4 g02854(new_n3240, new_n3239, new_n2183);
nand_4 g02855(new_n3241, new_n3240, new_n2179);
nand_4 g02856(new_n3242_1, new_n3241, new_n2175_1);
nand_4 g02857(new_n3243, new_n3242_1, new_n2171);
nand_4 g02858(new_n3244, new_n3243, new_n2168);
nand_4 g02859(new_n3245, new_n3244, new_n2165);
nand_4 g02860(new_n3246, new_n3245, new_n2162);
nand_4 g02861(new_n3247, new_n3246, new_n2158);
nand_4 g02862(new_n3248, new_n3247, new_n2155);
nand_4 g02863(new_n3249, new_n3248, new_n2151);
nand_4 g02864(new_n3250, new_n3249, new_n2147);
nand_4 g02865(new_n3251, new_n3250, new_n1810);
nand_4 g02866(new_n3252, new_n3251, new_n1806);
nand_4 g02867(new_n3253, new_n3252, new_n1802);
nand_4 g02868(new_n3254, new_n3253, new_n1798);
nand_4 g02869(new_n3255, new_n3254, new_n1820);
nand_4 g02870(new_n3256, new_n3255, new_n1794);
nand_4 g02871(new_n3257, new_n3256, new_n1825);
nand_4 g02872(new_n3258, new_n3257, n12336);
nor_4  g02873(n1739, new_n3258, new_n1285);
nand_4 g02874(new_n3260, new_n1460, new_n397);
nand_4 g02875(new_n3261, new_n3260, new_n1468);
nand_4 g02876(new_n3262, new_n3261, new_n1247);
nand_4 g02877(new_n3263_1, new_n3262, new_n1474);
nand_4 g02878(new_n3264, new_n3263_1, new_n592);
nand_4 g02879(new_n3265, new_n3264, new_n585);
nand_4 g02880(new_n3266, new_n3265, new_n580);
nand_4 g02881(new_n3267, new_n3266, new_n600);
nand_4 g02882(new_n3268, new_n3267, new_n606);
nand_4 g02883(new_n3269, new_n3268, new_n612);
nand_4 g02884(new_n3270, new_n3269, new_n575);
nand_4 g02885(new_n3271, new_n3270, new_n619);
nand_4 g02886(new_n3272, new_n3271, new_n570);
nand_4 g02887(new_n3273, new_n3272, new_n625);
nand_4 g02888(new_n3274, new_n3273, new_n564);
nand_4 g02889(new_n3275, new_n3274, new_n632);
nand_4 g02890(new_n3276, new_n3275, new_n638);
nand_4 g02891(new_n3277, new_n3276, new_n559);
nand_4 g02892(new_n3278, new_n3277, new_n554);
nand_4 g02893(new_n3279, new_n3278, new_n646);
nand_4 g02894(new_n3280, new_n3279, new_n652);
nand_4 g02895(new_n3281, new_n3280, new_n549);
nand_4 g02896(new_n3282, new_n3281, new_n544);
nand_4 g02897(new_n3283, new_n3282, new_n660);
nand_4 g02898(new_n3284, new_n3283, new_n539);
nand_4 g02899(new_n3285, new_n3284, new_n534);
nand_4 g02900(new_n3286, new_n3285, new_n529);
nand_4 g02901(new_n3287, new_n3286, new_n668);
nand_4 g02902(new_n3288, new_n3287, new_n674_1);
nand_4 g02903(new_n3289, new_n3288, new_n681);
nand_4 g02904(new_n3290, new_n3289, new_n523);
nand_4 g02905(new_n3291, new_n3290, new_n687);
nand_4 g02906(new_n3292, new_n3291, new_n693);
nand_4 g02907(new_n3293, new_n3292, new_n699);
nand_4 g02908(new_n3294, new_n3293, new_n517);
nand_4 g02909(new_n3295, new_n3294, new_n705);
nand_4 g02910(new_n3296, new_n3295, new_n511);
nand_4 g02911(new_n3297, new_n3296, new_n711);
nand_4 g02912(new_n3298, new_n3297, new_n506);
nand_4 g02913(new_n3299, new_n3298, new_n719);
nand_4 g02914(new_n3300, new_n3299, new_n500);
nand_4 g02915(new_n3301, new_n3300, new_n727);
nand_4 g02916(new_n3302, new_n3301, new_n494);
nand_4 g02917(new_n3303, new_n3302, new_n735);
nand_4 g02918(new_n3304, new_n3303, new_n488);
nand_4 g02919(new_n3305, new_n3304, new_n743);
nand_4 g02920(new_n3306, new_n3305, new_n482);
nand_4 g02921(new_n3307, new_n3306, new_n751);
nand_4 g02922(new_n3308, new_n3307, new_n758);
nand_4 g02923(new_n3309, new_n3308, new_n765);
nand_4 g02924(new_n3310, new_n3309, new_n476);
not_3  g02925(new_n3311, new_n3310);
nor_4  g02926(new_n3312, new_n3311, new_n774);
nor_4  g02927(new_n3313, new_n3312, new_n781);
nor_4  g02928(new_n3314, new_n3313, new_n788);
nor_4  g02929(new_n3315, new_n3314, new_n471);
nor_4  g02930(new_n3316, new_n3315, new_n796);
nor_4  g02931(new_n3317, new_n3316, new_n804);
nor_4  g02932(new_n3318, new_n3317, new_n810);
nor_4  g02933(new_n3319, new_n3318, new_n2043);
nor_4  g02934(new_n3320, new_n3319, new_n2042);
nor_4  g02935(new_n3321, new_n3320, new_n2041);
nor_4  g02936(new_n3322, new_n3321, new_n2040);
nor_4  g02937(new_n3323, new_n3322, new_n2039);
nor_4  g02938(new_n3324, new_n3323, new_n2038);
nor_4  g02939(new_n3325, new_n3324, new_n2037);
nor_4  g02940(new_n3326, new_n3325, new_n2036);
nor_4  g02941(new_n3327, new_n3326, new_n2035);
nor_4  g02942(new_n3328, new_n3327, new_n2034);
nor_4  g02943(new_n3329, new_n3328, new_n2033);
nor_4  g02944(new_n3330, new_n3329, new_n2032);
nor_4  g02945(new_n3331, new_n3330, new_n2031);
nor_4  g02946(new_n3332, new_n3331, new_n2030);
nor_4  g02947(new_n3333, new_n3332, new_n2029);
nor_4  g02948(new_n3334, new_n3333, new_n2028);
nor_4  g02949(new_n3335, new_n3334, new_n2027_1);
nor_4  g02950(new_n3336, new_n3335, new_n2026);
nor_4  g02951(new_n3337, new_n3336, new_n2025);
nor_4  g02952(new_n3338, new_n3337, new_n2024);
not_3  g02953(new_n3339, new_n3338);
nand_4 g02954(new_n3340_1, new_n3339, new_n413);
nand_4 g02955(new_n3341, new_n3340_1, new_n889);
nand_4 g02956(new_n3342, new_n3341, new_n896);
nand_4 g02957(new_n3343, new_n3342, new_n901);
nand_4 g02958(new_n3344, new_n3343, new_n408);
nand_4 g02959(new_n3345, new_n3344, new_n908);
nand_4 g02960(new_n3346, new_n3345, n394);
nor_4  g02961(n1827, new_n3346, new_n400);
not_3  g02962(new_n3348, new_n506);
not_3  g02963(new_n3349, new_n711);
not_3  g02964(new_n3350, new_n511);
not_3  g02965(new_n3351, new_n705);
not_3  g02966(new_n3352, new_n517);
not_3  g02967(new_n3353, new_n699);
not_3  g02968(new_n3354, new_n693);
nand_4 g02969(new_n3355, new_n1323, new_n817);
nand_4 g02970(new_n3356, new_n3355, new_n1410);
nand_4 g02971(new_n3357, new_n3356, new_n1413);
nand_4 g02972(new_n3358, new_n3357, new_n1322);
nand_4 g02973(new_n3359, new_n3358, new_n1317);
nand_4 g02974(new_n3360, new_n3359, new_n1315);
nand_4 g02975(new_n3361, new_n3360, new_n1419);
nand_4 g02976(new_n3362, new_n3361, new_n1310);
nand_4 g02977(new_n3363, new_n3362, new_n1305);
nand_4 g02978(new_n3364, new_n3363, new_n1427);
nand_4 g02979(new_n3365, new_n3364, new_n1431);
nand_4 g02980(new_n3366, new_n3365, new_n1302);
nand_4 g02981(new_n3367_1, new_n3366, new_n1298);
nand_4 g02982(new_n3368, new_n3367_1, new_n1295);
nand_4 g02983(new_n3369, new_n3368, new_n1291);
nand_4 g02984(new_n3370, new_n3369, new_n1288);
nand_4 g02985(new_n3371, new_n3370, new_n1284);
nand_4 g02986(new_n3372, new_n3371, new_n1280);
nand_4 g02987(new_n3373, new_n3372, new_n1275);
nand_4 g02988(new_n3374, new_n3373, new_n1445);
nand_4 g02989(new_n3375, new_n3374, new_n1270);
nand_4 g02990(new_n3376, new_n3375, new_n1265_1);
nand_4 g02991(new_n3377, new_n3376, new_n1260);
nand_4 g02992(new_n3378, new_n3377, new_n1256);
nand_4 g02993(new_n3379, new_n3378, new_n1251);
nand_4 g02994(new_n3380, new_n3379, new_n1457);
nand_4 g02995(new_n3381, new_n3380, new_n1462);
nand_4 g02996(new_n3382, new_n3381, new_n1468);
nand_4 g02997(new_n3383, new_n3382, new_n1247);
nand_4 g02998(new_n3384, new_n3383, new_n1474);
nand_4 g02999(new_n3385, new_n3384, new_n592);
nand_4 g03000(new_n3386, new_n3385, new_n585);
nand_4 g03001(new_n3387, new_n3386, new_n580);
nand_4 g03002(new_n3388_1, new_n3387, new_n600);
nand_4 g03003(new_n3389, new_n3388_1, new_n606);
nand_4 g03004(new_n3390, new_n3389, new_n612);
nand_4 g03005(new_n3391, new_n3390, new_n575);
nand_4 g03006(new_n3392, new_n3391, new_n619);
nand_4 g03007(new_n3393, new_n3392, new_n570);
nand_4 g03008(new_n3394, new_n3393, new_n625);
nand_4 g03009(new_n3395, new_n3394, new_n564);
nand_4 g03010(new_n3396, new_n3395, new_n632);
nand_4 g03011(new_n3397, new_n3396, new_n638);
nand_4 g03012(new_n3398, new_n3397, new_n559);
nand_4 g03013(new_n3399, new_n3398, new_n554);
nand_4 g03014(new_n3400, new_n3399, new_n646);
nand_4 g03015(new_n3401, new_n3400, new_n652);
nand_4 g03016(new_n3402, new_n3401, new_n549);
nand_4 g03017(new_n3403, new_n3402, new_n544);
nand_4 g03018(new_n3404, new_n3403, new_n660);
nand_4 g03019(new_n3405, new_n3404, new_n539);
not_3  g03020(new_n3406, new_n3405);
nor_4  g03021(new_n3407, new_n3406, new_n3067);
nor_4  g03022(new_n3408, new_n3407, new_n3066);
nor_4  g03023(new_n3409, new_n3408, new_n3065);
nor_4  g03024(new_n3410, new_n3409, new_n3064);
nor_4  g03025(new_n3411, new_n3410, new_n3063);
nor_4  g03026(new_n3412, new_n3411, new_n3062);
nor_4  g03027(new_n3413, new_n3412, new_n3061);
nor_4  g03028(new_n3414, new_n3413, new_n3354);
nor_4  g03029(new_n3415, new_n3414, new_n3353);
nor_4  g03030(new_n3416, new_n3415, new_n3352);
nor_4  g03031(new_n3417, new_n3416, new_n3351);
nor_4  g03032(new_n3418, new_n3417, new_n3350);
nor_4  g03033(new_n3419, new_n3418, new_n3349);
nor_4  g03034(new_n3420, new_n3419, new_n3348);
nor_4  g03035(new_n3421, new_n3420, new_n720);
nor_4  g03036(new_n3422, new_n3421, new_n501);
nor_4  g03037(new_n3423, new_n3422, new_n728);
nor_4  g03038(new_n3424, new_n3423, new_n495);
nor_4  g03039(new_n3425, new_n3424, new_n736);
nor_4  g03040(new_n3426, new_n3425, new_n489);
nor_4  g03041(new_n3427, new_n3426, new_n744);
nor_4  g03042(new_n3428, new_n3427, new_n483);
nor_4  g03043(new_n3429, new_n3428, new_n752);
nor_4  g03044(new_n3430, new_n3429, new_n759);
nor_4  g03045(new_n3431, new_n3430, new_n766);
nor_4  g03046(new_n3432, new_n3431, new_n477);
nor_4  g03047(new_n3433, new_n3432, new_n774);
not_3  g03048(new_n3434, new_n3433);
nand_4 g03049(new_n3435, new_n3434, new_n780);
nand_4 g03050(new_n3436, new_n3435, new_n787);
nand_4 g03051(new_n3437, new_n3436, new_n470);
nand_4 g03052(new_n3438, new_n3437, new_n795);
nand_4 g03053(new_n3439, new_n3438, new_n803);
nand_4 g03054(new_n3440, new_n3439, new_n809);
nand_4 g03055(new_n3441, new_n3440, n730);
nor_4  g03056(n1900, new_n3441, new_n462_1);
not_3  g03057(new_n3443, new_n2178);
nand_4 g03058(new_n3444, new_n3443, new_n1401);
nand_4 g03059(new_n3445, new_n3444, new_n463);
nand_4 g03060(new_n3446, new_n3445, new_n818);
nand_4 g03061(new_n3447, new_n3446, new_n460);
nand_4 g03062(new_n3448, new_n3447, new_n455);
nand_4 g03063(new_n3449, new_n3448, new_n449);
nand_4 g03064(new_n3450, new_n3449, new_n827);
nand_4 g03065(new_n3451, new_n3450, new_n833);
nand_4 g03066(new_n3452, new_n3451, new_n444);
nand_4 g03067(new_n3453, new_n3452, new_n439);
nand_4 g03068(new_n3454, new_n3453, new_n841);
nand_4 g03069(new_n3455, new_n3454, new_n434);
nand_4 g03070(new_n3456, new_n3455, new_n429);
nand_4 g03071(new_n3457, new_n3456, new_n424);
nand_4 g03072(new_n3458, new_n3457, new_n850);
nand_4 g03073(new_n3459, new_n3458, new_n856);
nand_4 g03074(new_n3460, new_n3459, new_n863);
nand_4 g03075(new_n3461, new_n3460, new_n419);
nand_4 g03076(new_n3462, new_n3461, new_n869);
nand_4 g03077(new_n3463, new_n3462, new_n875);
nand_4 g03078(new_n3464, new_n3463, new_n881);
nand_4 g03079(new_n3465, new_n3464, new_n413);
nand_4 g03080(new_n3466, new_n3465, new_n889);
nand_4 g03081(new_n3467, new_n3466, new_n896);
nand_4 g03082(new_n3468, new_n3467, new_n901);
nand_4 g03083(new_n3469, new_n3468, new_n408);
nand_4 g03084(new_n3470, new_n3469, new_n908);
nand_4 g03085(new_n3471, new_n3470, new_n403);
nand_4 g03086(new_n3472, new_n3471, new_n398);
nand_4 g03087(new_n3473, new_n3472, new_n393);
nand_4 g03088(new_n3474, new_n3473, new_n916);
nand_4 g03089(new_n3475, new_n3474, new_n1123);
nand_4 g03090(new_n3476, new_n3475, new_n1164);
nand_4 g03091(new_n3477, new_n3476, new_n1120);
nand_4 g03092(new_n3478, new_n3477, new_n1169);
nand_4 g03093(new_n3479, new_n3478, new_n1116);
nand_4 g03094(new_n3480, new_n3479, new_n1111);
nand_4 g03095(new_n3481, new_n3480, new_n1106);
nand_4 g03096(new_n3482, new_n3481, new_n1178);
nand_4 g03097(new_n3483, new_n3482, new_n1183);
nand_4 g03098(new_n3484, new_n3483, new_n1102);
nand_4 g03099(new_n3485, new_n3484, new_n1099);
nand_4 g03100(new_n3486, new_n3485, new_n1191);
nand_4 g03101(new_n3487, new_n3486, new_n1095);
nand_4 g03102(new_n3488, new_n3487, new_n1091);
nand_4 g03103(new_n3489, new_n3488, new_n1088);
not_3  g03104(new_n3490, new_n3489);
nor_4  g03105(new_n3491, new_n3490, new_n1517);
nor_4  g03106(new_n3492, new_n3491, new_n1516);
nor_4  g03107(new_n3493, new_n3492, new_n1075);
nor_4  g03108(new_n3494, new_n3493, new_n1071);
nor_4  g03109(new_n3495, new_n3494, new_n1065);
nor_4  g03110(new_n3496, new_n3495, new_n1062);
nor_4  g03111(new_n3497, new_n3496, new_n1056);
nor_4  g03112(new_n3498, new_n3497, new_n1051);
nor_4  g03113(new_n3499, new_n3498, new_n1046);
nor_4  g03114(new_n3500, new_n3499, new_n1042);
nor_4  g03115(new_n3501, new_n3500, new_n1037);
nor_4  g03116(new_n3502, new_n3501, new_n1032);
nor_4  g03117(new_n3503, new_n3502, new_n1026);
nor_4  g03118(new_n3504, new_n3503, new_n1021);
nor_4  g03119(new_n3505, new_n3504, new_n1016);
nor_4  g03120(new_n3506_1, new_n3505, new_n1011);
nor_4  g03121(new_n3507, new_n3506_1, new_n1216);
nor_4  g03122(new_n3508, new_n3507, new_n1006);
nor_4  g03123(new_n3509, new_n3508, new_n1001);
nor_4  g03124(new_n3510, new_n3509, new_n995);
nor_4  g03125(new_n3511, new_n3510, new_n990);
nor_4  g03126(new_n3512, new_n3511, new_n985);
nor_4  g03127(new_n3513, new_n3512, new_n979);
nor_4  g03128(new_n3514, new_n3513, new_n974);
not_3  g03129(new_n3515, new_n3514);
nand_4 g03130(new_n3516, new_n3515, new_n967);
nand_4 g03131(new_n3517, new_n3516, new_n964);
nand_4 g03132(new_n3518, new_n3517, new_n960);
nand_4 g03133(new_n3519, new_n3518, new_n957);
nand_4 g03134(new_n3520, new_n3519, new_n952);
nand_4 g03135(new_n3521, new_n3520, new_n948_1);
nand_4 g03136(new_n3522, new_n3521, new_n943);
nand_4 g03137(new_n3523, new_n3522, new_n938);
nand_4 g03138(new_n3524, new_n3523, new_n934);
nand_4 g03139(new_n3525, new_n3524, new_n929);
nand_4 g03140(new_n3526, new_n3525, new_n925);
nand_4 g03141(new_n3527, new_n3526, new_n2194);
nand_4 g03142(new_n3528, new_n3527, new_n2191);
nand_4 g03143(new_n3529, new_n3528, new_n2190);
nand_4 g03144(new_n3530, new_n3529, new_n2186);
nand_4 g03145(new_n3531, new_n3530, n8737);
nor_4  g03146(n1927, new_n3531, new_n2180);
not_3  g03147(new_n3533, new_n1760);
not_3  g03148(new_n3534, new_n938);
not_3  g03149(new_n3535, new_n943);
not_3  g03150(new_n3536, new_n948_1);
not_3  g03151(new_n3537, n6362);
not_3  g03152(new_n3538, new_n1757);
nand_4 g03153(new_n3539, new_n3538, new_n3537);
nand_4 g03154(new_n3540, new_n3539, new_n401);
nand_4 g03155(new_n3541, new_n3540, new_n398);
nand_4 g03156(new_n3542, new_n3541, new_n393);
nand_4 g03157(new_n3543, new_n3542, new_n916);
nand_4 g03158(new_n3544, new_n3543, new_n1123);
nand_4 g03159(new_n3545, new_n3544, new_n1164);
nand_4 g03160(new_n3546, new_n3545, new_n1120);
nand_4 g03161(new_n3547, new_n3546, new_n1169);
nand_4 g03162(new_n3548, new_n3547, new_n1116);
nand_4 g03163(new_n3549, new_n3548, new_n1111);
nand_4 g03164(new_n3550, new_n3549, new_n1106);
nand_4 g03165(new_n3551, new_n3550, new_n1178);
nand_4 g03166(new_n3552, new_n3551, new_n1183);
nand_4 g03167(new_n3553, new_n3552, new_n1102);
nand_4 g03168(new_n3554, new_n3553, new_n1099);
nand_4 g03169(new_n3555, new_n3554, new_n1191);
nand_4 g03170(new_n3556, new_n3555, new_n1095);
nand_4 g03171(new_n3557, new_n3556, new_n1091);
nand_4 g03172(new_n3558, new_n3557, new_n1088);
nand_4 g03173(new_n3559, new_n3558, new_n1084);
nand_4 g03174(new_n3560, new_n3559, new_n1079);
nand_4 g03175(new_n3561, new_n3560, new_n1074);
nand_4 g03176(new_n3562, new_n3561, new_n1070);
nand_4 g03177(new_n3563, new_n3562, new_n1064);
nand_4 g03178(new_n3564, new_n3563, new_n1061);
nand_4 g03179(new_n3565, new_n3564, new_n1055);
nand_4 g03180(new_n3566, new_n3565, new_n1050);
nand_4 g03181(new_n3567, new_n3566, new_n1045);
nand_4 g03182(new_n3568, new_n3567, new_n1041);
nand_4 g03183(new_n3569, new_n3568, new_n1036);
nand_4 g03184(new_n3570, new_n3569, new_n1031);
nand_4 g03185(new_n3571, new_n3570, new_n1025);
nand_4 g03186(new_n3572, new_n3571, new_n1020);
nand_4 g03187(new_n3573, new_n3572, new_n1015);
nand_4 g03188(new_n3574, new_n3573, new_n1010);
nand_4 g03189(new_n3575, new_n3574, new_n1215);
nand_4 g03190(new_n3576, new_n3575, new_n1005);
nand_4 g03191(new_n3577, new_n3576, new_n1000);
nand_4 g03192(new_n3578, new_n3577, new_n994);
nand_4 g03193(new_n3579, new_n3578, new_n989);
nand_4 g03194(new_n3580, new_n3579, new_n984);
nand_4 g03195(new_n3581, new_n3580, new_n978);
nand_4 g03196(new_n3582, new_n3581, new_n973);
nand_4 g03197(new_n3583, new_n3582, new_n967);
nand_4 g03198(new_n3584, new_n3583, new_n964);
not_3  g03199(new_n3585, new_n3584);
nor_4  g03200(new_n3586, new_n3585, new_n961);
nor_4  g03201(new_n3587, new_n3586, new_n958);
nor_4  g03202(new_n3588, new_n3587, new_n953);
nor_4  g03203(new_n3589, new_n3588, new_n3536);
nor_4  g03204(new_n3590, new_n3589, new_n3535);
nor_4  g03205(new_n3591, new_n3590, new_n3534);
nor_4  g03206(new_n3592, new_n3591, new_n2520);
nor_4  g03207(new_n3593, new_n3592, new_n2519);
nor_4  g03208(new_n3594, new_n3593, new_n2518);
nor_4  g03209(new_n3595, new_n3594, new_n2517);
nor_4  g03210(new_n3596, new_n3595, new_n2516);
nor_4  g03211(new_n3597, new_n3596, new_n2515);
nor_4  g03212(new_n3598, new_n3597, new_n2514);
nor_4  g03213(new_n3599, new_n3598, new_n2513);
nor_4  g03214(new_n3600, new_n3599, new_n2512);
nor_4  g03215(new_n3601, new_n3600, new_n2511);
nor_4  g03216(new_n3602, new_n3601, new_n2510);
nor_4  g03217(new_n3603_1, new_n3602, new_n2509);
nor_4  g03218(new_n3604, new_n3603_1, new_n2508);
nor_4  g03219(new_n3605, new_n3604, new_n2507);
nor_4  g03220(new_n3606, new_n3605, new_n2506);
nor_4  g03221(new_n3607, new_n3606, new_n2505);
nor_4  g03222(new_n3608, new_n3607, new_n2504);
nor_4  g03223(new_n3609, new_n3608, new_n2503);
not_3  g03224(new_n3610, new_n3609);
nand_4 g03225(new_n3611, new_n3610, new_n1810);
nand_4 g03226(new_n3612, new_n3611, new_n1806);
nand_4 g03227(new_n3613, new_n3612, new_n1802);
nand_4 g03228(new_n3614, new_n3613, new_n1798);
nand_4 g03229(new_n3615, new_n3614, new_n1820);
nand_4 g03230(new_n3616, new_n3615, new_n1794);
nand_4 g03231(new_n3617, new_n3616, new_n1825);
nand_4 g03232(new_n3618, new_n3617, new_n1789);
nand_4 g03233(new_n3619, new_n3618, new_n1785);
nand_4 g03234(new_n3620, new_n3619, new_n1780);
nand_4 g03235(new_n3621, new_n3620, new_n1777);
nand_4 g03236(new_n3622, new_n3621, new_n1774);
nand_4 g03237(new_n3623, new_n3622, new_n1834);
nand_4 g03238(new_n3624, new_n3623, new_n1769);
nand_4 g03239(new_n3625, new_n3624, new_n1766);
nand_4 g03240(new_n3626, new_n3625, n10050);
nor_4  g03241(n1951, new_n3626, new_n3533);
nand_4 g03242(new_n3628, new_n2176, new_n2175_1);
nand_4 g03243(new_n3629, new_n3628, new_n2171);
nand_4 g03244(new_n3630, new_n3629, new_n2168);
nand_4 g03245(new_n3631, new_n3630, new_n2165);
nand_4 g03246(new_n3632, new_n3631, new_n2162);
nand_4 g03247(new_n3633, new_n3632, new_n2158);
nand_4 g03248(new_n3634, new_n3633, new_n2155);
nand_4 g03249(new_n3635, new_n3634, new_n2151);
nand_4 g03250(new_n3636, new_n3635, new_n2147);
nand_4 g03251(new_n3637, new_n3636, new_n1810);
nand_4 g03252(new_n3638, new_n3637, new_n1806);
nand_4 g03253(new_n3639, new_n3638, new_n1802);
nand_4 g03254(new_n3640, new_n3639, new_n1798);
nand_4 g03255(new_n3641, new_n3640, new_n1820);
nand_4 g03256(new_n3642, new_n3641, new_n1794);
nand_4 g03257(new_n3643, new_n3642, new_n1825);
nand_4 g03258(new_n3644, new_n3643, new_n1789);
nand_4 g03259(new_n3645, new_n3644, new_n1785);
nand_4 g03260(new_n3646, new_n3645, new_n1780);
nand_4 g03261(new_n3647, new_n3646, new_n1777);
nand_4 g03262(new_n3648, new_n3647, new_n1774);
nand_4 g03263(new_n3649, new_n3648, new_n1834);
nand_4 g03264(new_n3650, new_n3649, new_n1769);
nand_4 g03265(new_n3651, new_n3650, new_n1766);
nand_4 g03266(new_n3652_1, new_n3651, new_n1762);
nand_4 g03267(new_n3653, new_n3652_1, new_n1758);
nand_4 g03268(new_n3654, new_n3653, new_n1754);
nand_4 g03269(new_n3655_1, new_n3654, new_n1751);
nand_4 g03270(new_n3656, new_n3655_1, new_n1748);
nand_4 g03271(new_n3657, new_n3656, new_n1746);
nand_4 g03272(new_n3658, new_n3657, new_n1742);
nand_4 g03273(new_n3659, new_n3658, new_n1738);
nand_4 g03274(new_n3660, new_n3659, new_n1736);
nand_4 g03275(new_n3661, new_n3660, new_n1732);
nand_4 g03276(new_n3662, new_n3661, new_n1729);
not_3  g03277(new_n3663, new_n3662);
nor_4  g03278(new_n3664, new_n3663, new_n2283);
nor_4  g03279(new_n3665, new_n3664, new_n2145);
nor_4  g03280(new_n3666, new_n3665, new_n2144);
nor_4  g03281(new_n3667, new_n3666, new_n2143);
nor_4  g03282(new_n3668, new_n3667, new_n2142);
nor_4  g03283(new_n3669, new_n3668, new_n2141);
nor_4  g03284(new_n3670, new_n3669, new_n2140);
nor_4  g03285(new_n3671, new_n3670, new_n2139);
nor_4  g03286(new_n3672, new_n3671, new_n2138);
nor_4  g03287(new_n3673_1, new_n3672, new_n2137);
nor_4  g03288(new_n3674, new_n3673_1, new_n2136);
nor_4  g03289(new_n3675, new_n3674, new_n2135);
nor_4  g03290(new_n3676, new_n3675, new_n2134);
nor_4  g03291(new_n3677, new_n3676, new_n2133);
nor_4  g03292(new_n3678, new_n3677, new_n2132);
nor_4  g03293(new_n3679, new_n3678, new_n1691);
nor_4  g03294(new_n3680, new_n3679, new_n1879);
nor_4  g03295(new_n3681, new_n3680, new_n1883);
nor_4  g03296(new_n3682, new_n3681, new_n1687);
not_3  g03297(new_n3683, new_n3682);
nand_4 g03298(new_n3684, new_n3683, new_n1682);
nand_4 g03299(new_n3685, new_n3684, new_n1678);
nand_4 g03300(new_n3686, new_n3685, new_n1674);
nand_4 g03301(new_n3687, new_n3686, new_n1890);
nand_4 g03302(new_n3688, new_n3687, new_n1669);
nand_4 g03303(new_n3689, new_n3688, new_n1665);
nand_4 g03304(new_n3690, new_n3689, new_n1661);
nand_4 g03305(new_n3691, new_n3690, new_n1657);
nand_4 g03306(new_n3692, new_n3691, new_n1652);
nand_4 g03307(new_n3693, new_n3692, new_n1648);
nand_4 g03308(new_n3694, new_n3693, new_n1644);
nand_4 g03309(new_n3695, new_n3694, new_n1640);
nand_4 g03310(new_n3696, new_n3695, new_n1636);
nand_4 g03311(new_n3697, new_n3696, new_n1632);
nand_4 g03312(new_n3698, new_n3697, new_n1378);
nand_4 g03313(new_n3699, new_n3698, new_n1372);
nand_4 g03314(new_n3700, new_n3699, new_n1367);
nand_4 g03315(new_n3701, new_n3700, new_n1363);
nand_4 g03316(new_n3702, new_n3701, new_n1360);
nand_4 g03317(new_n3703, new_n3702, new_n1357);
nand_4 g03318(new_n3704, new_n3703, new_n1354);
nand_4 g03319(new_n3705, new_n3704, new_n1352);
nand_4 g03320(new_n3706, new_n3705, new_n1350);
nand_4 g03321(new_n3707, new_n3706, new_n1347_1);
nand_4 g03322(new_n3708, new_n3707, new_n1344);
nand_4 g03323(new_n3709, new_n3708, new_n1341);
nand_4 g03324(new_n3710, new_n3709, new_n1338);
nand_4 g03325(new_n3711, new_n3710, new_n1395);
nand_4 g03326(new_n3712, new_n3711, new_n1335);
nand_4 g03327(new_n3713, new_n3712, new_n1332);
nand_4 g03328(new_n3714, new_n3713, n4615);
nor_4  g03329(n2027, new_n3714, new_n806);
not_3  g03330(new_n3716, new_n1338);
not_3  g03331(new_n3717, new_n1341);
not_3  g03332(new_n3718, new_n1344);
not_3  g03333(new_n3719, new_n1347_1);
not_3  g03334(new_n3720, new_n1350);
not_3  g03335(new_n3721, new_n1352);
not_3  g03336(new_n3722, new_n1354);
not_3  g03337(new_n3723, new_n1466);
nand_4 g03338(new_n3724, new_n1748, new_n3723);
nand_4 g03339(new_n3725, new_n3724, new_n1746);
nand_4 g03340(new_n3726, new_n3725, new_n1742);
nand_4 g03341(new_n3727, new_n3726, new_n1738);
nand_4 g03342(new_n3728, new_n3727, new_n1736);
nand_4 g03343(new_n3729, new_n3728, new_n1732);
nand_4 g03344(new_n3730, new_n3729, new_n1729);
nand_4 g03345(new_n3731, new_n3730, new_n1726);
nand_4 g03346(new_n3732, new_n3731, new_n1724);
nand_4 g03347(new_n3733, new_n3732, new_n1721);
nand_4 g03348(new_n3734, new_n3733, new_n1718);
nand_4 g03349(new_n3735, new_n3734, new_n1715);
nand_4 g03350(new_n3736, new_n3735, new_n1711);
nand_4 g03351(new_n3737, new_n3736, new_n1708);
nand_4 g03352(new_n3738, new_n3737, new_n1705);
nand_4 g03353(new_n3739, new_n3738, new_n1703);
nand_4 g03354(new_n3740, new_n3739, new_n1860);
nand_4 g03355(new_n3741, new_n3740, new_n1864);
nand_4 g03356(new_n3742, new_n3741, new_n1699);
nand_4 g03357(new_n3743, new_n3742, new_n1697);
nand_4 g03358(new_n3744, new_n3743, new_n1871);
nand_4 g03359(new_n3745, new_n3744, new_n1694);
nand_4 g03360(new_n3746, new_n3745, new_n1690);
nand_4 g03361(new_n3747, new_n3746, new_n1878);
nand_4 g03362(new_n3748, new_n3747, new_n1882);
nand_4 g03363(new_n3749, new_n3748, new_n1686);
nand_4 g03364(new_n3750, new_n3749, new_n1682);
nand_4 g03365(new_n3751, new_n3750, new_n1678);
nand_4 g03366(new_n3752, new_n3751, new_n1674);
nand_4 g03367(new_n3753, new_n3752, new_n1890);
nand_4 g03368(new_n3754, new_n3753, new_n1669);
nand_4 g03369(new_n3755, new_n3754, new_n1665);
nand_4 g03370(new_n3756, new_n3755, new_n1661);
nand_4 g03371(new_n3757, new_n3756, new_n1657);
nand_4 g03372(new_n3758, new_n3757, new_n1652);
nand_4 g03373(new_n3759, new_n3758, new_n1648);
nand_4 g03374(new_n3760, new_n3759, new_n1644);
nand_4 g03375(new_n3761, new_n3760, new_n1640);
nand_4 g03376(new_n3762, new_n3761, new_n1636);
nand_4 g03377(new_n3763, new_n3762, new_n1632);
nand_4 g03378(new_n3764, new_n3763, new_n1378);
nand_4 g03379(new_n3765, new_n3764, new_n1372);
nand_4 g03380(new_n3766, new_n3765, new_n1367);
nand_4 g03381(new_n3767, new_n3766, new_n1363);
nand_4 g03382(new_n3768, new_n3767, new_n1360);
nand_4 g03383(new_n3769, new_n3768, new_n1357);
not_3  g03384(new_n3770, new_n3769);
nor_4  g03385(new_n3771, new_n3770, new_n3722);
nor_4  g03386(new_n3772, new_n3771, new_n3721);
nor_4  g03387(new_n3773, new_n3772, new_n3720);
nor_4  g03388(new_n3774, new_n3773, new_n3719);
nor_4  g03389(new_n3775_1, new_n3774, new_n3718);
nor_4  g03390(new_n3776, new_n3775_1, new_n3717);
nor_4  g03391(new_n3777, new_n3776, new_n3716);
nor_4  g03392(new_n3778, new_n3777, new_n2611);
nor_4  g03393(new_n3779, new_n3778, new_n2610);
nor_4  g03394(new_n3780, new_n3779, new_n2609);
nor_4  g03395(new_n3781, new_n3780, new_n2413);
nor_4  g03396(new_n3782, new_n3781, new_n2412);
nor_4  g03397(new_n3783, new_n3782, new_n2411);
nor_4  g03398(new_n3784, new_n3783, new_n2410);
nor_4  g03399(new_n3785, new_n3784, new_n2409);
nor_4  g03400(new_n3786, new_n3785, new_n2408);
nor_4  g03401(new_n3787, new_n3786, new_n2407_1);
nor_4  g03402(new_n3788, new_n3787, new_n2406);
nor_4  g03403(new_n3789, new_n3788, new_n2405);
nor_4  g03404(new_n3790, new_n3789, new_n2404);
nor_4  g03405(new_n3791, new_n3790, new_n2403);
nor_4  g03406(new_n3792, new_n3791, new_n2402);
nor_4  g03407(new_n3793, new_n3792, new_n2401);
nor_4  g03408(new_n3794, new_n3793, new_n2400);
not_3  g03409(new_n3795, new_n3794);
nand_4 g03410(new_n3796, new_n3795, new_n1298);
nand_4 g03411(new_n3797, new_n3796, new_n1295);
nand_4 g03412(new_n3798, new_n3797, new_n1291);
nand_4 g03413(new_n3799_1, new_n3798, new_n1288);
nand_4 g03414(new_n3800, new_n3799_1, new_n1284);
nand_4 g03415(new_n3801, new_n3800, new_n1280);
nand_4 g03416(new_n3802, new_n3801, new_n1275);
nand_4 g03417(new_n3803, new_n3802, new_n1445);
nand_4 g03418(new_n3804_1, new_n3803, new_n1270);
nand_4 g03419(new_n3805, new_n3804_1, new_n1265_1);
nand_4 g03420(new_n3806, new_n3805, new_n1260);
nand_4 g03421(new_n3807, new_n3806, new_n1256);
nand_4 g03422(new_n3808, new_n3807, new_n1251);
nand_4 g03423(new_n3809, new_n3808, new_n1457);
nand_4 g03424(new_n3810, new_n3809, n4895);
nor_4  g03425(n2126, new_n3810, new_n395);
nand_4 g03426(new_n3812, new_n1702_1, new_n1086);
nand_4 g03427(new_n3813, new_n3812, new_n1084);
nand_4 g03428(new_n3814, new_n3813, new_n1079);
nand_4 g03429(new_n3815, new_n3814, new_n1074);
nand_4 g03430(new_n3816, new_n3815, new_n1070);
nand_4 g03431(new_n3817, new_n3816, new_n1064);
nand_4 g03432(new_n3818, new_n3817, new_n1061);
nand_4 g03433(new_n3819, new_n3818, new_n1055);
nand_4 g03434(new_n3820, new_n3819, new_n1050);
nand_4 g03435(new_n3821, new_n3820, new_n1045);
nand_4 g03436(new_n3822, new_n3821, new_n1041);
nand_4 g03437(new_n3823, new_n3822, new_n1036);
nand_4 g03438(new_n3824, new_n3823, new_n1031);
nand_4 g03439(new_n3825, new_n3824, new_n1025);
nand_4 g03440(new_n3826, new_n3825, new_n1020);
nand_4 g03441(new_n3827, new_n3826, new_n1015);
nand_4 g03442(new_n3828, new_n3827, new_n1010);
nand_4 g03443(new_n3829, new_n3828, new_n1215);
nand_4 g03444(new_n3830, new_n3829, new_n1005);
nand_4 g03445(new_n3831, new_n3830, new_n1000);
nand_4 g03446(new_n3832, new_n3831, new_n994);
nand_4 g03447(new_n3833_1, new_n3832, new_n989);
nand_4 g03448(new_n3834, new_n3833_1, new_n984);
nand_4 g03449(new_n3835, new_n3834, new_n978);
nand_4 g03450(new_n3836, new_n3835, new_n973);
nand_4 g03451(new_n3837, new_n3836, new_n967);
nand_4 g03452(new_n3838, new_n3837, new_n964);
nand_4 g03453(new_n3839, new_n3838, new_n960);
nand_4 g03454(new_n3840, new_n3839, new_n957);
nand_4 g03455(new_n3841, new_n3840, new_n952);
nand_4 g03456(new_n3842, new_n3841, new_n948_1);
nand_4 g03457(new_n3843, new_n3842, new_n943);
nand_4 g03458(new_n3844, new_n3843, new_n938);
nand_4 g03459(new_n3845, new_n3844, new_n934);
nand_4 g03460(new_n3846, new_n3845, new_n929);
nand_4 g03461(new_n3847, new_n3846, new_n925);
nand_4 g03462(new_n3848, new_n3847, new_n2194);
nand_4 g03463(new_n3849, new_n3848, new_n2191);
nand_4 g03464(new_n3850, new_n3849, new_n2190);
nand_4 g03465(new_n3851, new_n3850, new_n2186);
nand_4 g03466(new_n3852, new_n3851, new_n2183);
nand_4 g03467(new_n3853, new_n3852, new_n2179);
nand_4 g03468(new_n3854_1, new_n3853, new_n2175_1);
nand_4 g03469(new_n3855, new_n3854_1, new_n2171);
nand_4 g03470(new_n3856, new_n3855, new_n2168);
nand_4 g03471(new_n3857, new_n3856, new_n2165);
nand_4 g03472(new_n3858, new_n3857, new_n2162);
nand_4 g03473(new_n3859, new_n3858, new_n2158);
nand_4 g03474(new_n3860, new_n3859, new_n2155);
nand_4 g03475(new_n3861, new_n3860, new_n2151);
not_3  g03476(new_n3862, new_n3861);
nor_4  g03477(new_n3863, new_n3862, new_n2503);
nor_4  g03478(new_n3864, new_n3863, new_n2502);
nor_4  g03479(new_n3865, new_n3864, new_n2790);
nor_4  g03480(new_n3866, new_n3865, new_n2789);
nor_4  g03481(new_n3867, new_n3866, new_n2788);
nor_4  g03482(new_n3868, new_n3867, new_n2305);
nor_4  g03483(new_n3869, new_n3868, new_n2304);
nor_4  g03484(new_n3870, new_n3869, new_n2303);
nor_4  g03485(new_n3871, new_n3870, new_n2302);
nor_4  g03486(new_n3872, new_n3871, new_n2301);
nor_4  g03487(new_n3873, new_n3872, new_n2300);
nor_4  g03488(new_n3874, new_n3873, new_n2299);
nor_4  g03489(new_n3875, new_n3874, new_n2298);
nor_4  g03490(new_n3876, new_n3875, new_n2297);
nor_4  g03491(new_n3877, new_n3876, new_n2296);
nor_4  g03492(new_n3878, new_n3877, new_n2295);
nor_4  g03493(new_n3879, new_n3878, new_n2294);
nor_4  g03494(new_n3880, new_n3879, new_n2293);
nor_4  g03495(new_n3881, new_n3880, new_n2292);
nor_4  g03496(new_n3882, new_n3881, new_n2291);
nor_4  g03497(new_n3883, new_n3882, new_n2290);
nor_4  g03498(new_n3884, new_n3883, new_n2289);
nor_4  g03499(new_n3885, new_n3884, new_n2288);
nor_4  g03500(new_n3886, new_n3885, new_n2287);
nor_4  g03501(new_n3887, new_n3886, new_n2286);
not_3  g03502(new_n3888, new_n3887);
nand_4 g03503(new_n3889, new_n3888, new_n1732);
nand_4 g03504(new_n3890, new_n3889, new_n1729);
nand_4 g03505(new_n3891, new_n3890, new_n1726);
nand_4 g03506(new_n3892, new_n3891, new_n1724);
nand_4 g03507(new_n3893_1, new_n3892, new_n1721);
nand_4 g03508(new_n3894, new_n3893_1, new_n1718);
nand_4 g03509(new_n3895, new_n3894, new_n1715);
nand_4 g03510(new_n3896, new_n3895, new_n1711);
nand_4 g03511(new_n3897, new_n3896, new_n1708);
nand_4 g03512(new_n3898, new_n3897, n13890);
nor_4  g03513(n2175, new_n3898, new_n629);
not_3  g03514(new_n3900, new_n442);
nand_4 g03515(new_n3901_1, new_n1419, new_n3900);
nand_4 g03516(new_n3902, new_n3901_1, new_n1310);
nand_4 g03517(new_n3903, new_n3902, new_n1305);
nand_4 g03518(new_n3904, new_n3903, new_n1427);
nand_4 g03519(new_n3905, new_n3904, new_n1431);
nand_4 g03520(new_n3906, new_n3905, new_n1302);
nand_4 g03521(new_n3907, new_n3906, new_n1298);
nand_4 g03522(new_n3908, new_n3907, new_n1295);
nand_4 g03523(new_n3909, new_n3908, new_n1291);
nand_4 g03524(new_n3910_1, new_n3909, new_n1288);
nand_4 g03525(new_n3911, new_n3910_1, new_n1284);
nand_4 g03526(new_n3912, new_n3911, new_n1280);
nand_4 g03527(new_n3913, new_n3912, new_n1275);
nand_4 g03528(new_n3914, new_n3913, new_n1445);
nand_4 g03529(new_n3915, new_n3914, new_n1270);
nand_4 g03530(new_n3916, new_n3915, new_n1265_1);
nand_4 g03531(new_n3917, new_n3916, new_n1260);
nand_4 g03532(new_n3918, new_n3917, new_n1256);
nand_4 g03533(new_n3919, new_n3918, new_n1251);
nand_4 g03534(new_n3920, new_n3919, new_n1457);
nand_4 g03535(new_n3921, new_n3920, new_n1462);
nand_4 g03536(new_n3922, new_n3921, new_n1468);
nand_4 g03537(new_n3923, new_n3922, new_n1247);
nand_4 g03538(new_n3924, new_n3923, new_n1474);
nand_4 g03539(new_n3925, new_n3924, new_n592);
nand_4 g03540(new_n3926, new_n3925, new_n585);
nand_4 g03541(new_n3927, new_n3926, new_n580);
nand_4 g03542(new_n3928, new_n3927, new_n600);
nand_4 g03543(new_n3929, new_n3928, new_n606);
nand_4 g03544(new_n3930, new_n3929, new_n612);
nand_4 g03545(new_n3931, new_n3930, new_n575);
nand_4 g03546(new_n3932, new_n3931, new_n619);
nand_4 g03547(new_n3933, new_n3932, new_n570);
nand_4 g03548(new_n3934, new_n3933, new_n625);
nand_4 g03549(new_n3935, new_n3934, new_n564);
nand_4 g03550(new_n3936, new_n3935, new_n632);
nand_4 g03551(new_n3937, new_n3936, new_n638);
nand_4 g03552(new_n3938, new_n3937, new_n559);
nand_4 g03553(new_n3939, new_n3938, new_n554);
nand_4 g03554(new_n3940, new_n3939, new_n646);
nand_4 g03555(new_n3941, new_n3940, new_n652);
nand_4 g03556(new_n3942, new_n3941, new_n549);
nand_4 g03557(new_n3943, new_n3942, new_n544);
nand_4 g03558(new_n3944, new_n3943, new_n660);
nand_4 g03559(new_n3945, new_n3944, new_n539);
nand_4 g03560(new_n3946, new_n3945, new_n534);
nand_4 g03561(new_n3947, new_n3946, new_n529);
nand_4 g03562(new_n3948, new_n3947, new_n668);
nand_4 g03563(new_n3949, new_n3948, new_n674_1);
nand_4 g03564(new_n3950, new_n3949, new_n681);
nand_4 g03565(new_n3951, new_n3950, new_n523);
not_3  g03566(new_n3952, new_n3951);
nor_4  g03567(new_n3953, new_n3952, new_n3061);
nor_4  g03568(new_n3954, new_n3953, new_n3354);
nor_4  g03569(new_n3955, new_n3954, new_n3353);
nor_4  g03570(new_n3956, new_n3955, new_n3352);
nor_4  g03571(new_n3957, new_n3956, new_n3351);
nor_4  g03572(new_n3958, new_n3957, new_n3350);
nor_4  g03573(new_n3959, new_n3958, new_n3349);
nor_4  g03574(new_n3960, new_n3959, new_n3348);
nor_4  g03575(new_n3961, new_n3960, new_n720);
nor_4  g03576(new_n3962, new_n3961, new_n501);
nor_4  g03577(new_n3963, new_n3962, new_n728);
nor_4  g03578(new_n3964, new_n3963, new_n495);
nor_4  g03579(new_n3965, new_n3964, new_n736);
nor_4  g03580(new_n3966, new_n3965, new_n489);
nor_4  g03581(new_n3967, new_n3966, new_n744);
nor_4  g03582(new_n3968, new_n3967, new_n483);
nor_4  g03583(new_n3969, new_n3968, new_n752);
nor_4  g03584(new_n3970, new_n3969, new_n759);
nor_4  g03585(new_n3971, new_n3970, new_n766);
nor_4  g03586(new_n3972_1, new_n3971, new_n477);
nor_4  g03587(new_n3973, new_n3972_1, new_n774);
nor_4  g03588(new_n3974, new_n3973, new_n781);
nor_4  g03589(new_n3975, new_n3974, new_n788);
nor_4  g03590(new_n3976, new_n3975, new_n471);
nor_4  g03591(new_n3977, new_n3976, new_n796);
nor_4  g03592(new_n3978, new_n3977, new_n804);
nor_4  g03593(new_n3979, new_n3978, new_n810);
not_3  g03594(new_n3980, new_n3979);
nand_4 g03595(new_n3981, new_n3980, new_n465);
nand_4 g03596(new_n3982, new_n3981, new_n818);
nand_4 g03597(new_n3983, new_n3982, new_n460);
nand_4 g03598(new_n3984, new_n3983, new_n455);
nand_4 g03599(new_n3985, new_n3984, new_n449);
nand_4 g03600(new_n3986, new_n3985, new_n827);
nand_4 g03601(new_n3987, new_n3986, n4175);
nor_4  g03602(n2223, new_n3987, new_n830);
not_3  g03603(new_n3989, new_n1043);
nand_4 g03604(new_n3990, new_n3989, new_n529);
nand_4 g03605(new_n3991, new_n3990, new_n668);
nand_4 g03606(new_n3992, new_n3991, new_n674_1);
nand_4 g03607(new_n3993, new_n3992, new_n681);
nand_4 g03608(new_n3994, new_n3993, new_n523);
nand_4 g03609(new_n3995, new_n3994, new_n687);
nand_4 g03610(new_n3996, new_n3995, new_n693);
nand_4 g03611(new_n3997, new_n3996, new_n699);
nand_4 g03612(new_n3998, new_n3997, new_n517);
nand_4 g03613(new_n3999, new_n3998, new_n705);
nand_4 g03614(new_n4000_1, new_n3999, new_n511);
nand_4 g03615(new_n4001, new_n4000_1, new_n711);
nand_4 g03616(new_n4002, new_n4001, new_n506);
nand_4 g03617(new_n4003, new_n4002, new_n719);
nand_4 g03618(new_n4004, new_n4003, new_n500);
nand_4 g03619(new_n4005, new_n4004, new_n727);
nand_4 g03620(new_n4006, new_n4005, new_n494);
nand_4 g03621(new_n4007, new_n4006, new_n735);
nand_4 g03622(new_n4008, new_n4007, new_n488);
nand_4 g03623(new_n4009, new_n4008, new_n743);
nand_4 g03624(new_n4010, new_n4009, new_n482);
nand_4 g03625(new_n4011, new_n4010, new_n751);
nand_4 g03626(new_n4012, new_n4011, new_n758);
nand_4 g03627(new_n4013, new_n4012, new_n765);
nand_4 g03628(new_n4014, new_n4013, new_n476);
nand_4 g03629(new_n4015, new_n4014, new_n773);
nand_4 g03630(new_n4016, new_n4015, new_n780);
nand_4 g03631(new_n4017, new_n4016, new_n787);
nand_4 g03632(new_n4018, new_n4017, new_n470);
nand_4 g03633(new_n4019, new_n4018, new_n795);
nand_4 g03634(new_n4020, new_n4019, new_n803);
nand_4 g03635(new_n4021, new_n4020, new_n809);
nand_4 g03636(new_n4022_1, new_n4021, new_n465);
nand_4 g03637(new_n4023, new_n4022_1, new_n818);
nand_4 g03638(new_n4024, new_n4023, new_n460);
nand_4 g03639(new_n4025, new_n4024, new_n455);
nand_4 g03640(new_n4026, new_n4025, new_n449);
nand_4 g03641(new_n4027, new_n4026, new_n827);
nand_4 g03642(new_n4028, new_n4027, new_n833);
nand_4 g03643(new_n4029, new_n4028, new_n444);
nand_4 g03644(new_n4030, new_n4029, new_n439);
nand_4 g03645(new_n4031, new_n4030, new_n841);
nand_4 g03646(new_n4032, new_n4031, new_n434);
nand_4 g03647(new_n4033, new_n4032, new_n429);
nand_4 g03648(new_n4034, new_n4033, new_n424);
nand_4 g03649(new_n4035, new_n4034, new_n850);
nand_4 g03650(new_n4036, new_n4035, new_n856);
nand_4 g03651(new_n4037, new_n4036, new_n863);
nand_4 g03652(new_n4038, new_n4037, new_n419);
nand_4 g03653(new_n4039_1, new_n4038, new_n869);
nand_4 g03654(new_n4040, new_n4039_1, new_n875);
not_3  g03655(new_n4041, new_n4040);
nor_4  g03656(new_n4042, new_n4041, new_n2024);
nor_4  g03657(new_n4043, new_n4042, new_n2023);
nor_4  g03658(new_n4044, new_n4043, new_n2022);
nor_4  g03659(new_n4045, new_n4044, new_n2021);
nor_4  g03660(new_n4046, new_n4045, new_n2020);
nor_4  g03661(new_n4047, new_n4046, new_n2019);
nor_4  g03662(new_n4048, new_n4047, new_n1537);
nor_4  g03663(new_n4049, new_n4048, new_n1536);
nor_4  g03664(new_n4050, new_n4049, new_n1535);
nor_4  g03665(new_n4051, new_n4050, new_n1534);
nor_4  g03666(new_n4052, new_n4051, new_n1533);
nor_4  g03667(new_n4053, new_n4052, new_n1532);
nor_4  g03668(new_n4054, new_n4053, new_n1531);
nor_4  g03669(new_n4055, new_n4054, new_n1530);
nor_4  g03670(new_n4056, new_n4055, new_n1529);
nor_4  g03671(new_n4057, new_n4056, new_n1528);
nor_4  g03672(new_n4058, new_n4057, new_n1527);
nor_4  g03673(new_n4059, new_n4058, new_n1526);
nor_4  g03674(new_n4060, new_n4059, new_n1525);
nor_4  g03675(new_n4061, new_n4060, new_n1524);
nor_4  g03676(new_n4062, new_n4061, new_n1523);
nor_4  g03677(new_n4063, new_n4062, new_n1522);
nor_4  g03678(new_n4064, new_n4063, new_n1521);
nor_4  g03679(new_n4065, new_n4064, new_n1520);
nor_4  g03680(new_n4066, new_n4065, new_n1519);
nor_4  g03681(new_n4067, new_n4066, new_n1518);
nor_4  g03682(new_n4068, new_n4067, new_n1517);
not_3  g03683(new_n4069, new_n4068);
nand_4 g03684(new_n4070, new_n4069, new_n1079);
nand_4 g03685(new_n4071, new_n4070, new_n1074);
nand_4 g03686(new_n4072, new_n4071, new_n1070);
nand_4 g03687(new_n4073, new_n4072, new_n1064);
nand_4 g03688(new_n4074, new_n4073, new_n1061);
nand_4 g03689(new_n4075, new_n4074, new_n1055);
nand_4 g03690(new_n4076, new_n4075, n3804);
nor_4  g03691(n2311, new_n4076, new_n1048);
nand_4 g03692(new_n4078, new_n1799, new_n1798);
nand_4 g03693(new_n4079, new_n4078, new_n1820);
nand_4 g03694(new_n4080, new_n4079, new_n1794);
nand_4 g03695(new_n4081, new_n4080, new_n1825);
nand_4 g03696(new_n4082, new_n4081, new_n1789);
nand_4 g03697(new_n4083, new_n4082, new_n1785);
nand_4 g03698(new_n4084, new_n4083, new_n1780);
nand_4 g03699(new_n4085, new_n4084, new_n1777);
nand_4 g03700(new_n4086, new_n4085, new_n1774);
nand_4 g03701(new_n4087, new_n4086, new_n1834);
nand_4 g03702(new_n4088, new_n4087, new_n1769);
nand_4 g03703(new_n4089, new_n4088, new_n1766);
nand_4 g03704(new_n4090, new_n4089, new_n1762);
nand_4 g03705(new_n4091, new_n4090, new_n1758);
nand_4 g03706(new_n4092, new_n4091, new_n1754);
nand_4 g03707(new_n4093, new_n4092, new_n1751);
nand_4 g03708(new_n4094, new_n4093, new_n1748);
nand_4 g03709(new_n4095, new_n4094, new_n1746);
nand_4 g03710(new_n4096, new_n4095, new_n1742);
nand_4 g03711(new_n4097, new_n4096, new_n1738);
nand_4 g03712(new_n4098, new_n4097, new_n1736);
nand_4 g03713(new_n4099, new_n4098, new_n1732);
nand_4 g03714(new_n4100, new_n4099, new_n1729);
nand_4 g03715(new_n4101, new_n4100, new_n1726);
nand_4 g03716(new_n4102, new_n4101, new_n1724);
nand_4 g03717(new_n4103, new_n4102, new_n1721);
nand_4 g03718(new_n4104, new_n4103, new_n1718);
nand_4 g03719(new_n4105, new_n4104, new_n1715);
nand_4 g03720(new_n4106, new_n4105, new_n1711);
nand_4 g03721(new_n4107, new_n4106, new_n1708);
nand_4 g03722(new_n4108, new_n4107, new_n1705);
nand_4 g03723(new_n4109, new_n4108, new_n1703);
nand_4 g03724(new_n4110, new_n4109, new_n1860);
nand_4 g03725(new_n4111, new_n4110, new_n1864);
nand_4 g03726(new_n4112, new_n4111, new_n1699);
not_3  g03727(new_n4113, new_n4112);
nor_4  g03728(new_n4114, new_n4113, new_n2134);
nor_4  g03729(new_n4115, new_n4114, new_n2133);
nor_4  g03730(new_n4116, new_n4115, new_n2132);
nor_4  g03731(new_n4117_1, new_n4116, new_n1691);
nor_4  g03732(new_n4118, new_n4117_1, new_n1879);
nor_4  g03733(new_n4119, new_n4118, new_n1883);
nor_4  g03734(new_n4120, new_n4119, new_n1687);
nor_4  g03735(new_n4121, new_n4120, new_n1683);
nor_4  g03736(new_n4122, new_n4121, new_n1679);
nor_4  g03737(new_n4123, new_n4122, new_n1675);
nor_4  g03738(new_n4124, new_n4123, new_n1891);
nor_4  g03739(new_n4125_1, new_n4124, new_n1670);
nor_4  g03740(new_n4126, new_n4125_1, new_n1666);
nor_4  g03741(new_n4127, new_n4126, new_n1662);
nor_4  g03742(new_n4128, new_n4127, new_n1658);
nor_4  g03743(new_n4129, new_n4128, new_n1653);
nor_4  g03744(new_n4130, new_n4129, new_n1649);
nor_4  g03745(new_n4131_1, new_n4130, new_n1645);
nor_4  g03746(new_n4132, new_n4131_1, new_n1641);
not_3  g03747(new_n4133, new_n4132);
nand_4 g03748(new_n4134, new_n4133, new_n1636);
nand_4 g03749(new_n4135, new_n4134, new_n1632);
nand_4 g03750(new_n4136, new_n4135, new_n1378);
nand_4 g03751(new_n4137, new_n4136, new_n1372);
nand_4 g03752(new_n4138, new_n4137, new_n1367);
nand_4 g03753(new_n4139, new_n4138, new_n1363);
nand_4 g03754(new_n4140, new_n4139, new_n1360);
nand_4 g03755(new_n4141, new_n4140, new_n1357);
nand_4 g03756(new_n4142, new_n4141, new_n1354);
nand_4 g03757(new_n4143, new_n4142, new_n1352);
nand_4 g03758(new_n4144, new_n4143, new_n1350);
nand_4 g03759(new_n4145, new_n4144, new_n1347_1);
nand_4 g03760(new_n4146, new_n4145, new_n1344);
nand_4 g03761(new_n4147_1, new_n4146, new_n1341);
nand_4 g03762(new_n4148, new_n4147_1, new_n1338);
nand_4 g03763(new_n4149, new_n4148, new_n1395);
nand_4 g03764(new_n4150, new_n4149, new_n1335);
nand_4 g03765(new_n4151, new_n4150, new_n1332);
nand_4 g03766(new_n4152, new_n4151, new_n1328);
nand_4 g03767(new_n4153, new_n4152, new_n1403);
nand_4 g03768(new_n4154_1, new_n4153, new_n1325);
nand_4 g03769(new_n4155, new_n4154_1, new_n1410);
nand_4 g03770(new_n4156, new_n4155, new_n1413);
nand_4 g03771(new_n4157, new_n4156, new_n1322);
nand_4 g03772(new_n4158, new_n4157, new_n1317);
nand_4 g03773(new_n4159, new_n4158, new_n1315);
nand_4 g03774(new_n4160, new_n4159, new_n1419);
nand_4 g03775(new_n4161, new_n4160, new_n1310);
nand_4 g03776(new_n4162, new_n4161, new_n1305);
nand_4 g03777(new_n4163, new_n4162, new_n1427);
nand_4 g03778(new_n4164, new_n4163, n10147);
nor_4  g03779(n2407, new_n4164, new_n426);
not_3  g03780(new_n4166, new_n1676);
nand_4 g03781(new_n4167, new_n4166, new_n1031);
nand_4 g03782(new_n4168, new_n4167, new_n1025);
nand_4 g03783(new_n4169, new_n4168, new_n1020);
nand_4 g03784(new_n4170, new_n4169, new_n1015);
nand_4 g03785(new_n4171, new_n4170, new_n1010);
nand_4 g03786(new_n4172_1, new_n4171, new_n1215);
nand_4 g03787(new_n4173, new_n4172_1, new_n1005);
nand_4 g03788(new_n4174, new_n4173, new_n1000);
nand_4 g03789(new_n4175_1, new_n4174, new_n994);
nand_4 g03790(new_n4176, new_n4175_1, new_n989);
nand_4 g03791(new_n4177, new_n4176, new_n984);
nand_4 g03792(new_n4178, new_n4177, new_n978);
nand_4 g03793(new_n4179, new_n4178, new_n973);
nand_4 g03794(new_n4180, new_n4179, new_n967);
nand_4 g03795(new_n4181, new_n4180, new_n964);
nand_4 g03796(new_n4182, new_n4181, new_n960);
nand_4 g03797(new_n4183, new_n4182, new_n957);
nand_4 g03798(new_n4184, new_n4183, new_n952);
nand_4 g03799(new_n4185, new_n4184, new_n948_1);
nand_4 g03800(new_n4186, new_n4185, new_n943);
nand_4 g03801(new_n4187, new_n4186, new_n938);
nand_4 g03802(new_n4188, new_n4187, new_n934);
nand_4 g03803(new_n4189, new_n4188, new_n929);
nand_4 g03804(new_n4190, new_n4189, new_n925);
nand_4 g03805(new_n4191, new_n4190, new_n2194);
nand_4 g03806(new_n4192, new_n4191, new_n2191);
nand_4 g03807(new_n4193, new_n4192, new_n2190);
nand_4 g03808(new_n4194, new_n4193, new_n2186);
nand_4 g03809(new_n4195, new_n4194, new_n2183);
nand_4 g03810(new_n4196, new_n4195, new_n2179);
nand_4 g03811(new_n4197, new_n4196, new_n2175_1);
nand_4 g03812(new_n4198, new_n4197, new_n2171);
nand_4 g03813(new_n4199, new_n4198, new_n2168);
nand_4 g03814(new_n4200, new_n4199, new_n2165);
nand_4 g03815(new_n4201, new_n4200, new_n2162);
nand_4 g03816(new_n4202, new_n4201, new_n2158);
nand_4 g03817(new_n4203, new_n4202, new_n2155);
nand_4 g03818(new_n4204, new_n4203, new_n2151);
nand_4 g03819(new_n4205, new_n4204, new_n2147);
nand_4 g03820(new_n4206, new_n4205, new_n1810);
nand_4 g03821(new_n4207, new_n4206, new_n1806);
nand_4 g03822(new_n4208, new_n4207, new_n1802);
nand_4 g03823(new_n4209, new_n4208, new_n1798);
nand_4 g03824(new_n4210, new_n4209, new_n1820);
nand_4 g03825(new_n4211, new_n4210, new_n1794);
nand_4 g03826(new_n4212, new_n4211, new_n1825);
not_3  g03827(new_n4213, new_n4212);
nor_4  g03828(new_n4214, new_n4213, new_n2302);
nor_4  g03829(new_n4215, new_n4214, new_n2301);
nor_4  g03830(new_n4216, new_n4215, new_n2300);
nor_4  g03831(new_n4217, new_n4216, new_n2299);
nor_4  g03832(new_n4218, new_n4217, new_n2298);
nor_4  g03833(new_n4219, new_n4218, new_n2297);
nor_4  g03834(new_n4220, new_n4219, new_n2296);
nor_4  g03835(new_n4221, new_n4220, new_n2295);
nor_4  g03836(new_n4222, new_n4221, new_n2294);
nor_4  g03837(new_n4223, new_n4222, new_n2293);
nor_4  g03838(new_n4224, new_n4223, new_n2292);
nor_4  g03839(new_n4225_1, new_n4224, new_n2291);
nor_4  g03840(new_n4226, new_n4225_1, new_n2290);
nor_4  g03841(new_n4227, new_n4226, new_n2289);
nor_4  g03842(new_n4228, new_n4227, new_n2288);
nor_4  g03843(new_n4229, new_n4228, new_n2287);
nor_4  g03844(new_n4230, new_n4229, new_n2286);
nor_4  g03845(new_n4231, new_n4230, new_n2285);
nor_4  g03846(new_n4232, new_n4231, new_n2284);
nor_4  g03847(new_n4233, new_n4232, new_n2283);
nor_4  g03848(new_n4234, new_n4233, new_n2145);
nor_4  g03849(new_n4235, new_n4234, new_n2144);
nor_4  g03850(new_n4236, new_n4235, new_n2143);
nor_4  g03851(new_n4237, new_n4236, new_n2142);
not_3  g03852(new_n4238, new_n4237);
nand_4 g03853(new_n4239, new_n4238, new_n1711);
nand_4 g03854(new_n4240, new_n4239, new_n1708);
nand_4 g03855(new_n4241, new_n4240, new_n1705);
nand_4 g03856(new_n4242, new_n4241, new_n1703);
nand_4 g03857(new_n4243, new_n4242, new_n1860);
nand_4 g03858(new_n4244, new_n4243, new_n1864);
nand_4 g03859(new_n4245, new_n4244, new_n1699);
nand_4 g03860(new_n4246, new_n4245, new_n1697);
nand_4 g03861(new_n4247, new_n4246, new_n1871);
nand_4 g03862(new_n4248, new_n4247, new_n1694);
nand_4 g03863(new_n4249, new_n4248, new_n1690);
nand_4 g03864(new_n4250, new_n4249, new_n1878);
nand_4 g03865(new_n4251, new_n4250, new_n1882);
nand_4 g03866(new_n4252, new_n4251, new_n1686);
nand_4 g03867(new_n4253, new_n4252, n8799);
nor_4  g03868(n2556, new_n4253, new_n665);
nand_4 g03869(new_n4255, new_n1727, new_n599);
nand_4 g03870(new_n4256, new_n4255, new_n1726);
nand_4 g03871(new_n4257, new_n4256, new_n1724);
nand_4 g03872(new_n4258, new_n4257, new_n1721);
nand_4 g03873(new_n4259, new_n4258, new_n1718);
nand_4 g03874(new_n4260, new_n4259, new_n1715);
nand_4 g03875(new_n4261, new_n4260, new_n1711);
nand_4 g03876(new_n4262, new_n4261, new_n1708);
nand_4 g03877(new_n4263, new_n4262, new_n1705);
nand_4 g03878(new_n4264, new_n4263, new_n1703);
nand_4 g03879(new_n4265, new_n4264, new_n1860);
nand_4 g03880(new_n4266, new_n4265, new_n1864);
nand_4 g03881(new_n4267, new_n4266, new_n1699);
nand_4 g03882(new_n4268, new_n4267, new_n1697);
nand_4 g03883(new_n4269, new_n4268, new_n1871);
nand_4 g03884(new_n4270, new_n4269, new_n1694);
nand_4 g03885(new_n4271, new_n4270, new_n1690);
nand_4 g03886(new_n4272, new_n4271, new_n1878);
nand_4 g03887(new_n4273, new_n4272, new_n1882);
nand_4 g03888(new_n4274, new_n4273, new_n1686);
nand_4 g03889(new_n4275, new_n4274, new_n1682);
nand_4 g03890(new_n4276, new_n4275, new_n1678);
nand_4 g03891(new_n4277, new_n4276, new_n1674);
nand_4 g03892(new_n4278, new_n4277, new_n1890);
nand_4 g03893(new_n4279_1, new_n4278, new_n1669);
nand_4 g03894(new_n4280, new_n4279_1, new_n1665);
nand_4 g03895(new_n4281, new_n4280, new_n1661);
nand_4 g03896(new_n4282_1, new_n4281, new_n1657);
nand_4 g03897(new_n4283, new_n4282_1, new_n1652);
nand_4 g03898(new_n4284, new_n4283, new_n1648);
nand_4 g03899(new_n4285, new_n4284, new_n1644);
nand_4 g03900(new_n4286, new_n4285, new_n1640);
nand_4 g03901(new_n4287, new_n4286, new_n1636);
nand_4 g03902(new_n4288, new_n4287, new_n1632);
nand_4 g03903(new_n4289, new_n4288, new_n1378);
nand_4 g03904(new_n4290, new_n4289, new_n1372);
nand_4 g03905(new_n4291, new_n4290, new_n1367);
nand_4 g03906(new_n4292_1, new_n4291, new_n1363);
nand_4 g03907(new_n4293, new_n4292_1, new_n1360);
nand_4 g03908(new_n4294, new_n4293, new_n1357);
nand_4 g03909(new_n4295, new_n4294, new_n1354);
nand_4 g03910(new_n4296, new_n4295, new_n1352);
nand_4 g03911(new_n4297, new_n4296, new_n1350);
nand_4 g03912(new_n4298, new_n4297, new_n1347_1);
nand_4 g03913(new_n4299, new_n4298, new_n1344);
nand_4 g03914(new_n4300, new_n4299, new_n1341);
nand_4 g03915(new_n4301, new_n4300, new_n1338);
nand_4 g03916(new_n4302, new_n4301, new_n1395);
nand_4 g03917(new_n4303, new_n4302, new_n1335);
nand_4 g03918(new_n4304, new_n4303, new_n1332);
nand_4 g03919(new_n4305_1, new_n4304, new_n1328);
not_3  g03920(new_n4306, new_n4305_1);
nor_4  g03921(new_n4307, new_n4306, new_n2412);
nor_4  g03922(new_n4308, new_n4307, new_n2411);
nor_4  g03923(new_n4309, new_n4308, new_n2410);
nor_4  g03924(new_n4310, new_n4309, new_n2409);
nor_4  g03925(new_n4311, new_n4310, new_n2408);
nor_4  g03926(new_n4312, new_n4311, new_n2407_1);
nor_4  g03927(new_n4313, new_n4312, new_n2406);
nor_4  g03928(new_n4314, new_n4313, new_n2405);
nor_4  g03929(new_n4315, new_n4314, new_n2404);
nor_4  g03930(new_n4316, new_n4315, new_n2403);
nor_4  g03931(new_n4317, new_n4316, new_n2402);
nor_4  g03932(new_n4318, new_n4317, new_n2401);
nor_4  g03933(new_n4319, new_n4318, new_n2400);
nor_4  g03934(new_n4320, new_n4319, new_n2399);
nor_4  g03935(new_n4321, new_n4320, new_n2398);
nor_4  g03936(new_n4322, new_n4321, new_n2397);
nor_4  g03937(new_n4323, new_n4322, new_n2396);
nor_4  g03938(new_n4324, new_n4323, new_n2395);
nor_4  g03939(new_n4325, new_n4324, new_n1281);
nor_4  g03940(new_n4326, new_n4325, new_n1276);
nor_4  g03941(new_n4327, new_n4326, new_n1446);
nor_4  g03942(new_n4328, new_n4327, new_n1271);
nor_4  g03943(new_n4329, new_n4328, new_n1266);
nor_4  g03944(new_n4330, new_n4329, new_n1261);
nor_4  g03945(new_n4331, new_n4330, new_n1257);
nor_4  g03946(new_n4332, new_n4331, new_n1252);
nor_4  g03947(new_n4333, new_n4332, new_n1458);
not_3  g03948(new_n4334, new_n4333);
nand_4 g03949(new_n4335, new_n4334, new_n1462);
nand_4 g03950(new_n4336, new_n4335, new_n1468);
nand_4 g03951(new_n4337, new_n4336, new_n1247);
nand_4 g03952(new_n4338, new_n4337, new_n1474);
nand_4 g03953(new_n4339, new_n4338, new_n592);
nand_4 g03954(new_n4340, new_n4339, new_n585);
nand_4 g03955(new_n4341, new_n4340, n7832);
nor_4  g03956(n2559, new_n4341, new_n577);
not_3  g03957(new_n4343, new_n450);
nand_4 g03958(new_n4344, new_n1413, new_n4343);
nand_4 g03959(new_n4345_1, new_n4344, new_n1322);
nand_4 g03960(new_n4346, new_n4345_1, new_n1317);
nand_4 g03961(new_n4347, new_n4346, new_n1315);
nand_4 g03962(new_n4348, new_n4347, new_n1419);
nand_4 g03963(new_n4349, new_n4348, new_n1310);
nand_4 g03964(new_n4350, new_n4349, new_n1305);
nand_4 g03965(new_n4351, new_n4350, new_n1427);
nand_4 g03966(new_n4352, new_n4351, new_n1431);
nand_4 g03967(new_n4353, new_n4352, new_n1302);
nand_4 g03968(new_n4354, new_n4353, new_n1298);
nand_4 g03969(new_n4355, new_n4354, new_n1295);
nand_4 g03970(new_n4356, new_n4355, new_n1291);
nand_4 g03971(new_n4357, new_n4356, new_n1288);
nand_4 g03972(new_n4358, new_n4357, new_n1284);
nand_4 g03973(new_n4359, new_n4358, new_n1280);
nand_4 g03974(new_n4360, new_n4359, new_n1275);
nand_4 g03975(new_n4361, new_n4360, new_n1445);
nand_4 g03976(new_n4362, new_n4361, new_n1270);
nand_4 g03977(new_n4363, new_n4362, new_n1265_1);
nand_4 g03978(new_n4364, new_n4363, new_n1260);
nand_4 g03979(new_n4365, new_n4364, new_n1256);
nand_4 g03980(new_n4366, new_n4365, new_n1251);
nand_4 g03981(new_n4367, new_n4366, new_n1457);
nand_4 g03982(new_n4368, new_n4367, new_n1462);
nand_4 g03983(new_n4369, new_n4368, new_n1468);
nand_4 g03984(new_n4370, new_n4369, new_n1247);
nand_4 g03985(new_n4371, new_n4370, new_n1474);
nand_4 g03986(new_n4372, new_n4371, new_n592);
nand_4 g03987(new_n4373, new_n4372, new_n585);
nand_4 g03988(new_n4374, new_n4373, new_n580);
nand_4 g03989(new_n4375, new_n4374, new_n600);
nand_4 g03990(new_n4376, new_n4375, new_n606);
nand_4 g03991(new_n4377, new_n4376, new_n612);
nand_4 g03992(new_n4378, new_n4377, new_n575);
not_3  g03993(new_n4379, new_n4378);
nor_4  g03994(new_n4380, new_n4379, new_n3081);
nor_4  g03995(new_n4381, new_n4380, new_n3080);
nor_4  g03996(new_n4382, new_n4381, new_n3079);
nor_4  g03997(new_n4383, new_n4382, new_n3078);
nor_4  g03998(new_n4384, new_n4383, new_n3077);
nor_4  g03999(new_n4385, new_n4384, new_n3076);
nor_4  g04000(new_n4386, new_n4385, new_n3075);
nor_4  g04001(new_n4387, new_n4386, new_n3074);
nor_4  g04002(new_n4388, new_n4387, new_n3073);
nor_4  g04003(new_n4389, new_n4388, new_n3072);
nor_4  g04004(new_n4390, new_n4389, new_n3071);
nor_4  g04005(new_n4391, new_n4390, new_n3070);
nor_4  g04006(new_n4392, new_n4391, new_n3069);
nor_4  g04007(new_n4393, new_n4392, new_n3068);
nor_4  g04008(new_n4394, new_n4393, new_n3067);
nor_4  g04009(new_n4395, new_n4394, new_n3066);
nor_4  g04010(new_n4396, new_n4395, new_n3065);
nor_4  g04011(new_n4397, new_n4396, new_n3064);
nor_4  g04012(new_n4398, new_n4397, new_n3063);
not_3  g04013(new_n4399, new_n4398);
nand_4 g04014(new_n4400, new_n4399, new_n523);
nand_4 g04015(new_n4401, new_n4400, new_n687);
nand_4 g04016(new_n4402, new_n4401, new_n693);
nand_4 g04017(new_n4403, new_n4402, new_n699);
nand_4 g04018(new_n4404, new_n4403, new_n517);
nand_4 g04019(new_n4405, new_n4404, new_n705);
nand_4 g04020(new_n4406, new_n4405, new_n511);
nand_4 g04021(new_n4407, new_n4406, new_n711);
nand_4 g04022(new_n4408, new_n4407, new_n506);
nand_4 g04023(new_n4409, new_n4408, new_n719);
nand_4 g04024(new_n4410, new_n4409, new_n500);
nand_4 g04025(new_n4411, new_n4410, new_n727);
nand_4 g04026(new_n4412, new_n4411, new_n494);
nand_4 g04027(new_n4413, new_n4412, new_n735);
nand_4 g04028(new_n4414, new_n4413, new_n488);
nand_4 g04029(new_n4415, new_n4414, new_n743);
nand_4 g04030(new_n4416, new_n4415, new_n482);
nand_4 g04031(new_n4417, new_n4416, new_n751);
nand_4 g04032(new_n4418, new_n4417, new_n758);
nand_4 g04033(new_n4419, new_n4418, new_n765);
nand_4 g04034(new_n4420, new_n4419, new_n476);
nand_4 g04035(new_n4421, new_n4420, new_n773);
nand_4 g04036(new_n4422, new_n4421, new_n780);
nand_4 g04037(new_n4423, new_n4422, new_n787);
nand_4 g04038(new_n4424, new_n4423, new_n470);
nand_4 g04039(new_n4425, new_n4424, new_n795);
nand_4 g04040(new_n4426, new_n4425, new_n803);
nand_4 g04041(new_n4427, new_n4426, new_n809);
nand_4 g04042(new_n4428, new_n4427, new_n465);
nand_4 g04043(new_n4429, new_n4428, new_n818);
nand_4 g04044(new_n4430, new_n4429, n3263);
nor_4  g04045(n2572, new_n4430, new_n457);
not_3  g04046(new_n4432, new_n1093_1);
not_3  g04047(new_n4433, new_n1089);
nand_4 g04048(new_n4434, new_n4433, new_n638);
nand_4 g04049(new_n4435, new_n4434, new_n559);
nand_4 g04050(new_n4436, new_n4435, new_n554);
nand_4 g04051(new_n4437_1, new_n4436, new_n646);
nand_4 g04052(new_n4438, new_n4437_1, new_n652);
nand_4 g04053(new_n4439, new_n4438, new_n549);
nand_4 g04054(new_n4440, new_n4439, new_n544);
nand_4 g04055(new_n4441, new_n4440, new_n660);
nand_4 g04056(new_n4442, new_n4441, new_n539);
nand_4 g04057(new_n4443, new_n4442, new_n534);
nand_4 g04058(new_n4444, new_n4443, new_n529);
nand_4 g04059(new_n4445, new_n4444, new_n668);
nand_4 g04060(new_n4446, new_n4445, new_n674_1);
nand_4 g04061(new_n4447, new_n4446, new_n681);
nand_4 g04062(new_n4448, new_n4447, new_n523);
nand_4 g04063(new_n4449, new_n4448, new_n687);
nand_4 g04064(new_n4450, new_n4449, new_n693);
nand_4 g04065(new_n4451, new_n4450, new_n699);
nand_4 g04066(new_n4452, new_n4451, new_n517);
nand_4 g04067(new_n4453, new_n4452, new_n705);
nand_4 g04068(new_n4454, new_n4453, new_n511);
nand_4 g04069(new_n4455, new_n4454, new_n711);
nand_4 g04070(new_n4456, new_n4455, new_n506);
nand_4 g04071(new_n4457, new_n4456, new_n719);
nand_4 g04072(new_n4458, new_n4457, new_n500);
nand_4 g04073(new_n4459, new_n4458, new_n727);
nand_4 g04074(new_n4460, new_n4459, new_n494);
nand_4 g04075(new_n4461, new_n4460, new_n735);
nand_4 g04076(new_n4462, new_n4461, new_n488);
nand_4 g04077(new_n4463, new_n4462, new_n743);
nand_4 g04078(new_n4464, new_n4463, new_n482);
nand_4 g04079(new_n4465, new_n4464, new_n751);
nand_4 g04080(new_n4466, new_n4465, new_n758);
nand_4 g04081(new_n4467, new_n4466, new_n765);
nand_4 g04082(new_n4468, new_n4467, new_n476);
nand_4 g04083(new_n4469, new_n4468, new_n773);
nand_4 g04084(new_n4470, new_n4469, new_n780);
nand_4 g04085(new_n4471, new_n4470, new_n787);
nand_4 g04086(new_n4472, new_n4471, new_n470);
nand_4 g04087(new_n4473, new_n4472, new_n795);
nand_4 g04088(new_n4474, new_n4473, new_n803);
nand_4 g04089(new_n4475, new_n4474, new_n809);
nand_4 g04090(new_n4476, new_n4475, new_n465);
nand_4 g04091(new_n4477, new_n4476, new_n818);
nand_4 g04092(new_n4478, new_n4477, new_n460);
nand_4 g04093(new_n4479, new_n4478, new_n455);
nand_4 g04094(new_n4480, new_n4479, new_n449);
nand_4 g04095(new_n4481, new_n4480, new_n827);
nand_4 g04096(new_n4482, new_n4481, new_n833);
nand_4 g04097(new_n4483, new_n4482, new_n444);
nand_4 g04098(new_n4484, new_n4483, new_n439);
not_3  g04099(new_n4485, new_n4484);
nor_4  g04100(new_n4486, new_n4485, new_n2034);
nor_4  g04101(new_n4487, new_n4486, new_n2033);
nor_4  g04102(new_n4488, new_n4487, new_n2032);
nor_4  g04103(new_n4489, new_n4488, new_n2031);
nor_4  g04104(new_n4490, new_n4489, new_n2030);
nor_4  g04105(new_n4491, new_n4490, new_n2029);
nor_4  g04106(new_n4492, new_n4491, new_n2028);
nor_4  g04107(new_n4493, new_n4492, new_n2027_1);
nor_4  g04108(new_n4494, new_n4493, new_n2026);
nor_4  g04109(new_n4495, new_n4494, new_n2025);
nor_4  g04110(new_n4496, new_n4495, new_n2024);
nor_4  g04111(new_n4497, new_n4496, new_n2023);
nor_4  g04112(new_n4498, new_n4497, new_n2022);
nor_4  g04113(new_n4499, new_n4498, new_n2021);
nor_4  g04114(new_n4500, new_n4499, new_n2020);
nor_4  g04115(new_n4501, new_n4500, new_n2019);
nor_4  g04116(new_n4502, new_n4501, new_n1537);
nor_4  g04117(new_n4503, new_n4502, new_n1536);
nor_4  g04118(new_n4504, new_n4503, new_n1535);
nor_4  g04119(new_n4505, new_n4504, new_n1534);
nor_4  g04120(new_n4506, new_n4505, new_n1533);
nor_4  g04121(new_n4507, new_n4506, new_n1532);
nor_4  g04122(new_n4508, new_n4507, new_n1531);
nor_4  g04123(new_n4509, new_n4508, new_n1530);
nor_4  g04124(new_n4510, new_n4509, new_n1529);
nor_4  g04125(new_n4511, new_n4510, new_n1528);
nor_4  g04126(new_n4512, new_n4511, new_n1527);
not_3  g04127(new_n4513, new_n4512);
nand_4 g04128(new_n4514, new_n4513, new_n1106);
nand_4 g04129(new_n4515, new_n4514, new_n1178);
nand_4 g04130(new_n4516, new_n4515, new_n1183);
nand_4 g04131(new_n4517, new_n4516, new_n1102);
nand_4 g04132(new_n4518, new_n4517, new_n1099);
nand_4 g04133(new_n4519, new_n4518, new_n1191);
nand_4 g04134(new_n4520, new_n4519, n9977);
nor_4  g04135(n2672, new_n4520, new_n4432);
nand_4 g04136(new_n4522, new_n1014, new_n691);
nand_4 g04137(new_n4523, new_n4522, new_n699);
nand_4 g04138(new_n4524, new_n4523, new_n517);
nand_4 g04139(new_n4525, new_n4524, new_n705);
nand_4 g04140(new_n4526, new_n4525, new_n511);
nand_4 g04141(new_n4527, new_n4526, new_n711);
nand_4 g04142(new_n4528, new_n4527, new_n506);
nand_4 g04143(new_n4529, new_n4528, new_n719);
nand_4 g04144(new_n4530, new_n4529, new_n500);
nand_4 g04145(new_n4531, new_n4530, new_n727);
nand_4 g04146(new_n4532, new_n4531, new_n494);
nand_4 g04147(new_n4533, new_n4532, new_n735);
nand_4 g04148(new_n4534, new_n4533, new_n488);
nand_4 g04149(new_n4535, new_n4534, new_n743);
nand_4 g04150(new_n4536, new_n4535, new_n482);
nand_4 g04151(new_n4537, new_n4536, new_n751);
nand_4 g04152(new_n4538, new_n4537, new_n758);
nand_4 g04153(new_n4539, new_n4538, new_n765);
nand_4 g04154(new_n4540, new_n4539, new_n476);
nand_4 g04155(new_n4541_1, new_n4540, new_n773);
nand_4 g04156(new_n4542, new_n4541_1, new_n780);
nand_4 g04157(new_n4543, new_n4542, new_n787);
nand_4 g04158(new_n4544, new_n4543, new_n470);
nand_4 g04159(new_n4545, new_n4544, new_n795);
nand_4 g04160(new_n4546, new_n4545, new_n803);
nand_4 g04161(new_n4547, new_n4546, new_n809);
nand_4 g04162(new_n4548, new_n4547, new_n465);
nand_4 g04163(new_n4549, new_n4548, new_n818);
nand_4 g04164(new_n4550, new_n4549, new_n460);
nand_4 g04165(new_n4551, new_n4550, new_n455);
nand_4 g04166(new_n4552, new_n4551, new_n449);
nand_4 g04167(new_n4553, new_n4552, new_n827);
nand_4 g04168(new_n4554, new_n4553, new_n833);
nand_4 g04169(new_n4555, new_n4554, new_n444);
nand_4 g04170(new_n4556, new_n4555, new_n439);
nand_4 g04171(new_n4557, new_n4556, new_n841);
nand_4 g04172(new_n4558, new_n4557, new_n434);
nand_4 g04173(new_n4559, new_n4558, new_n429);
nand_4 g04174(new_n4560, new_n4559, new_n424);
nand_4 g04175(new_n4561, new_n4560, new_n850);
nand_4 g04176(new_n4562, new_n4561, new_n856);
nand_4 g04177(new_n4563, new_n4562, new_n863);
nand_4 g04178(new_n4564, new_n4563, new_n419);
nand_4 g04179(new_n4565, new_n4564, new_n869);
nand_4 g04180(new_n4566, new_n4565, new_n875);
not_3  g04181(new_n4567, new_n4566);
nor_4  g04182(new_n4568, new_n4567, new_n2024);
nor_4  g04183(new_n4569, new_n4568, new_n2023);
nor_4  g04184(new_n4570, new_n4569, new_n2022);
nor_4  g04185(new_n4571, new_n4570, new_n2021);
nor_4  g04186(new_n4572, new_n4571, new_n2020);
nor_4  g04187(new_n4573, new_n4572, new_n2019);
nor_4  g04188(new_n4574, new_n4573, new_n1537);
nor_4  g04189(new_n4575, new_n4574, new_n1536);
nor_4  g04190(new_n4576, new_n4575, new_n1535);
nor_4  g04191(new_n4577, new_n4576, new_n1534);
nor_4  g04192(new_n4578, new_n4577, new_n1533);
nor_4  g04193(new_n4579, new_n4578, new_n1532);
nor_4  g04194(new_n4580, new_n4579, new_n1531);
nor_4  g04195(new_n4581, new_n4580, new_n1530);
nor_4  g04196(new_n4582, new_n4581, new_n1529);
nor_4  g04197(new_n4583, new_n4582, new_n1528);
nor_4  g04198(new_n4584, new_n4583, new_n1527);
nor_4  g04199(new_n4585, new_n4584, new_n1526);
nor_4  g04200(new_n4586, new_n4585, new_n1525);
nor_4  g04201(new_n4587, new_n4586, new_n1524);
nor_4  g04202(new_n4588, new_n4587, new_n1523);
nor_4  g04203(new_n4589, new_n4588, new_n1522);
nor_4  g04204(new_n4590, new_n4589, new_n1521);
nor_4  g04205(new_n4591, new_n4590, new_n1520);
not_3  g04206(new_n4592, new_n4591);
nand_4 g04207(new_n4593, new_n4592, new_n1091);
nand_4 g04208(new_n4594, new_n4593, new_n1088);
nand_4 g04209(new_n4595, new_n4594, new_n1084);
nand_4 g04210(new_n4596, new_n4595, new_n1079);
nand_4 g04211(new_n4597, new_n4596, new_n1074);
nand_4 g04212(new_n4598, new_n4597, new_n1070);
nand_4 g04213(new_n4599, new_n4598, new_n1064);
nand_4 g04214(new_n4600, new_n4599, new_n1061);
nand_4 g04215(new_n4601, new_n4600, new_n1055);
nand_4 g04216(new_n4602, new_n4601, new_n1050);
nand_4 g04217(new_n4603, new_n4602, new_n1045);
nand_4 g04218(new_n4604_1, new_n4603, new_n1041);
nand_4 g04219(new_n4605, new_n4604_1, new_n1036);
nand_4 g04220(new_n4606, new_n4605, new_n1031);
nand_4 g04221(new_n4607, new_n4606, new_n1025);
nand_4 g04222(new_n4608, new_n4607, n6703);
nor_4  g04223(n2734, new_n4608, new_n1017);
nand_4 g04224(new_n4610, new_n1035, new_n672);
nand_4 g04225(new_n4611, new_n4610, new_n681);
nand_4 g04226(new_n4612, new_n4611, new_n523);
nand_4 g04227(new_n4613, new_n4612, new_n687);
nand_4 g04228(new_n4614, new_n4613, new_n693);
nand_4 g04229(new_n4615_1, new_n4614, new_n699);
nand_4 g04230(new_n4616, new_n4615_1, new_n517);
nand_4 g04231(new_n4617, new_n4616, new_n705);
nand_4 g04232(new_n4618, new_n4617, new_n511);
nand_4 g04233(new_n4619, new_n4618, new_n711);
nand_4 g04234(new_n4620, new_n4619, new_n506);
nand_4 g04235(new_n4621, new_n4620, new_n719);
nand_4 g04236(new_n4622, new_n4621, new_n500);
nand_4 g04237(new_n4623, new_n4622, new_n727);
nand_4 g04238(new_n4624, new_n4623, new_n494);
nand_4 g04239(new_n4625, new_n4624, new_n735);
nand_4 g04240(new_n4626, new_n4625, new_n488);
nand_4 g04241(new_n4627, new_n4626, new_n743);
nand_4 g04242(new_n4628, new_n4627, new_n482);
nand_4 g04243(new_n4629, new_n4628, new_n751);
nand_4 g04244(new_n4630, new_n4629, new_n758);
nand_4 g04245(new_n4631, new_n4630, new_n765);
nand_4 g04246(new_n4632, new_n4631, new_n476);
nand_4 g04247(new_n4633, new_n4632, new_n773);
nand_4 g04248(new_n4634, new_n4633, new_n780);
nand_4 g04249(new_n4635, new_n4634, new_n787);
nand_4 g04250(new_n4636, new_n4635, new_n470);
nand_4 g04251(new_n4637, new_n4636, new_n795);
nand_4 g04252(new_n4638, new_n4637, new_n803);
nand_4 g04253(new_n4639, new_n4638, new_n809);
nand_4 g04254(new_n4640, new_n4639, new_n465);
nand_4 g04255(new_n4641, new_n4640, new_n818);
nand_4 g04256(new_n4642, new_n4641, new_n460);
nand_4 g04257(new_n4643, new_n4642, new_n455);
nand_4 g04258(new_n4644, new_n4643, new_n449);
nand_4 g04259(new_n4645, new_n4644, new_n827);
nand_4 g04260(new_n4646, new_n4645, new_n833);
nand_4 g04261(new_n4647, new_n4646, new_n444);
nand_4 g04262(new_n4648, new_n4647, new_n439);
nand_4 g04263(new_n4649, new_n4648, new_n841);
nand_4 g04264(new_n4650, new_n4649, new_n434);
nand_4 g04265(new_n4651, new_n4650, new_n429);
nand_4 g04266(new_n4652, new_n4651, new_n424);
nand_4 g04267(new_n4653, new_n4652, new_n850);
nand_4 g04268(new_n4654, new_n4653, new_n856);
nand_4 g04269(new_n4655, new_n4654, new_n863);
nand_4 g04270(new_n4656, new_n4655, new_n419);
nand_4 g04271(new_n4657, new_n4656, new_n869);
nand_4 g04272(new_n4658, new_n4657, new_n875);
nand_4 g04273(new_n4659_1, new_n4658, new_n881);
not_3  g04274(new_n4660, new_n4659_1);
nor_4  g04275(new_n4661, new_n4660, new_n2023);
nor_4  g04276(new_n4662, new_n4661, new_n2022);
nor_4  g04277(new_n4663, new_n4662, new_n2021);
nor_4  g04278(new_n4664, new_n4663, new_n2020);
nor_4  g04279(new_n4665, new_n4664, new_n2019);
nor_4  g04280(new_n4666, new_n4665, new_n1537);
nor_4  g04281(new_n4667, new_n4666, new_n1536);
nor_4  g04282(new_n4668, new_n4667, new_n1535);
nor_4  g04283(new_n4669, new_n4668, new_n1534);
nor_4  g04284(new_n4670, new_n4669, new_n1533);
nor_4  g04285(new_n4671, new_n4670, new_n1532);
nor_4  g04286(new_n4672_1, new_n4671, new_n1531);
nor_4  g04287(new_n4673, new_n4672_1, new_n1530);
nor_4  g04288(new_n4674, new_n4673, new_n1529);
nor_4  g04289(new_n4675, new_n4674, new_n1528);
nor_4  g04290(new_n4676, new_n4675, new_n1527);
nor_4  g04291(new_n4677, new_n4676, new_n1526);
nor_4  g04292(new_n4678, new_n4677, new_n1525);
nor_4  g04293(new_n4679, new_n4678, new_n1524);
nor_4  g04294(new_n4680, new_n4679, new_n1523);
nor_4  g04295(new_n4681, new_n4680, new_n1522);
nor_4  g04296(new_n4682, new_n4681, new_n1521);
nor_4  g04297(new_n4683, new_n4682, new_n1520);
nor_4  g04298(new_n4684, new_n4683, new_n1519);
nor_4  g04299(new_n4685, new_n4684, new_n1518);
not_3  g04300(new_n4686, new_n4685);
nand_4 g04301(new_n4687, new_n4686, new_n1084);
nand_4 g04302(new_n4688, new_n4687, new_n1079);
nand_4 g04303(new_n4689, new_n4688, new_n1074);
nand_4 g04304(new_n4690, new_n4689, new_n1070);
nand_4 g04305(new_n4691, new_n4690, new_n1064);
nand_4 g04306(new_n4692, new_n4691, new_n1061);
nand_4 g04307(new_n4693, new_n4692, new_n1055);
nand_4 g04308(new_n4694, new_n4693, new_n1050);
nand_4 g04309(new_n4695, new_n4694, new_n1045);
nand_4 g04310(new_n4696, new_n4695, n650);
nor_4  g04311(n3090, new_n4696, new_n1038);
not_3  g04312(new_n4698, new_n590);
not_3  g04313(new_n4699, new_n1357);
not_3  g04314(new_n4700, new_n1360);
not_3  g04315(new_n4701, new_n583);
nand_4 g04316(new_n4702, new_n1736, new_n4701);
nand_4 g04317(new_n4703, new_n4702, new_n1732);
nand_4 g04318(new_n4704, new_n4703, new_n1729);
nand_4 g04319(new_n4705, new_n4704, new_n1726);
nand_4 g04320(new_n4706, new_n4705, new_n1724);
nand_4 g04321(new_n4707, new_n4706, new_n1721);
nand_4 g04322(new_n4708, new_n4707, new_n1718);
nand_4 g04323(new_n4709, new_n4708, new_n1715);
nand_4 g04324(new_n4710, new_n4709, new_n1711);
nand_4 g04325(new_n4711, new_n4710, new_n1708);
nand_4 g04326(new_n4712, new_n4711, new_n1705);
nand_4 g04327(new_n4713, new_n4712, new_n1703);
nand_4 g04328(new_n4714, new_n4713, new_n1860);
nand_4 g04329(new_n4715, new_n4714, new_n1864);
nand_4 g04330(new_n4716, new_n4715, new_n1699);
nand_4 g04331(new_n4717, new_n4716, new_n1697);
nand_4 g04332(new_n4718, new_n4717, new_n1871);
nand_4 g04333(new_n4719, new_n4718, new_n1694);
nand_4 g04334(new_n4720, new_n4719, new_n1690);
nand_4 g04335(new_n4721, new_n4720, new_n1878);
nand_4 g04336(new_n4722, new_n4721, new_n1882);
nand_4 g04337(new_n4723, new_n4722, new_n1686);
nand_4 g04338(new_n4724, new_n4723, new_n1682);
nand_4 g04339(new_n4725, new_n4724, new_n1678);
nand_4 g04340(new_n4726, new_n4725, new_n1674);
nand_4 g04341(new_n4727, new_n4726, new_n1890);
nand_4 g04342(new_n4728, new_n4727, new_n1669);
nand_4 g04343(new_n4729, new_n4728, new_n1665);
nand_4 g04344(new_n4730, new_n4729, new_n1661);
nand_4 g04345(new_n4731, new_n4730, new_n1657);
nand_4 g04346(new_n4732, new_n4731, new_n1652);
nand_4 g04347(new_n4733, new_n4732, new_n1648);
nand_4 g04348(new_n4734, new_n4733, new_n1644);
nand_4 g04349(new_n4735, new_n4734, new_n1640);
nand_4 g04350(new_n4736, new_n4735, new_n1636);
not_3  g04351(new_n4737, new_n4736);
nor_4  g04352(new_n4738, new_n4737, new_n1633);
nor_4  g04353(new_n4739, new_n4738, new_n1629);
nor_4  g04354(new_n4740, new_n4739, new_n1628);
nor_4  g04355(new_n4741, new_n4740, new_n1627);
nor_4  g04356(new_n4742, new_n4741, new_n1626);
nor_4  g04357(new_n4743, new_n4742, new_n4700);
nor_4  g04358(new_n4744, new_n4743, new_n4699);
nor_4  g04359(new_n4745, new_n4744, new_n3722);
nor_4  g04360(new_n4746, new_n4745, new_n3721);
nor_4  g04361(new_n4747, new_n4746, new_n3720);
nor_4  g04362(new_n4748, new_n4747, new_n3719);
nor_4  g04363(new_n4749, new_n4748, new_n3718);
nor_4  g04364(new_n4750, new_n4749, new_n3717);
nor_4  g04365(new_n4751, new_n4750, new_n3716);
nor_4  g04366(new_n4752, new_n4751, new_n2611);
nor_4  g04367(new_n4753, new_n4752, new_n2610);
nor_4  g04368(new_n4754, new_n4753, new_n2609);
nor_4  g04369(new_n4755_1, new_n4754, new_n2413);
nor_4  g04370(new_n4756, new_n4755_1, new_n2412);
not_3  g04371(new_n4757, new_n4756);
nand_4 g04372(new_n4758, new_n4757, new_n1325);
nand_4 g04373(new_n4759, new_n4758, new_n1410);
nand_4 g04374(new_n4760, new_n4759, new_n1413);
nand_4 g04375(new_n4761, new_n4760, new_n1322);
nand_4 g04376(new_n4762, new_n4761, new_n1317);
nand_4 g04377(new_n4763, new_n4762, new_n1315);
nand_4 g04378(new_n4764, new_n4763, new_n1419);
nand_4 g04379(new_n4765, new_n4764, new_n1310);
nand_4 g04380(new_n4766, new_n4765, new_n1305);
nand_4 g04381(new_n4767, new_n4766, new_n1427);
nand_4 g04382(new_n4768, new_n4767, new_n1431);
nand_4 g04383(new_n4769, new_n4768, new_n1302);
nand_4 g04384(new_n4770, new_n4769, new_n1298);
nand_4 g04385(new_n4771, new_n4770, new_n1295);
nand_4 g04386(new_n4772, new_n4771, new_n1291);
nand_4 g04387(new_n4773, new_n4772, new_n1288);
nand_4 g04388(new_n4774_1, new_n4773, new_n1284);
nand_4 g04389(new_n4775, new_n4774_1, new_n1280);
nand_4 g04390(new_n4776, new_n4775, new_n1275);
nand_4 g04391(new_n4777, new_n4776, new_n1445);
nand_4 g04392(new_n4778, new_n4777, new_n1270);
nand_4 g04393(new_n4779, new_n4778, new_n1265_1);
nand_4 g04394(new_n4780, new_n4779, new_n1260);
nand_4 g04395(new_n4781, new_n4780, new_n1256);
nand_4 g04396(new_n4782, new_n4781, new_n1251);
nand_4 g04397(new_n4783, new_n4782, new_n1457);
nand_4 g04398(new_n4784, new_n4783, new_n1462);
nand_4 g04399(new_n4785_1, new_n4784, new_n1468);
nand_4 g04400(new_n4786, new_n4785_1, new_n1247);
nand_4 g04401(new_n4787, new_n4786, new_n1474);
nand_4 g04402(new_n4788, new_n4787, n6147);
nor_4  g04403(n3242, new_n4788, new_n4698);
nor_4  g04404(new_n4790, new_n505, new_n418);
nor_4  g04405(new_n4791, new_n448, new_n438);
nor_4  g04406(new_n4792, new_n528, new_n392);
nand_4 g04407(new_n4793, new_n4792, new_n4791);
nor_4  g04408(new_n4794, new_n2193, new_n1793);
nand_4 g04409(new_n4795, new_n4794, new_n1778);
nor_4  g04410(new_n4796, new_n4795, new_n4793);
and_4  g04411(new_n4797, new_n4796, new_n4790);
nor_4  g04412(new_n4798, new_n1728, new_n1353);
nor_4  g04413(new_n4799, new_n481, new_n475);
nor_4  g04414(new_n4800, new_n1741, new_n1324);
and_4  g04415(new_n4801, new_n4800, new_n4799);
nand_4 g04416(new_n4802, new_n4801, new_n4798);
nor_4  g04417(new_n4803, new_n4802, new_n1030);
nand_4 g04418(new_n4804, new_n4803, new_n4797);
nor_4  g04419(new_n4805, new_n1304, new_n1297);
nor_4  g04420(new_n4806, new_n2182, new_n1805);
and_4  g04421(new_n4807, new_n4806, new_n1767);
nand_4 g04422(new_n4808, new_n4807, new_n4805);
nor_4  g04423(new_n4809, new_n464, new_n423);
nor_4  g04424(new_n4810, new_n516, new_n412);
nor_4  g04425(new_n4811, new_n522, new_n407);
and_4  g04426(new_n4812, new_n4811, new_n4810);
nand_4 g04427(new_n4813, new_n4812, new_n4809);
nor_4  g04428(new_n4814, new_n4813, new_n4808);
nor_4  g04429(new_n4815, new_n1366, new_n1269);
nor_4  g04430(new_n4816, new_n956, new_n937);
nor_4  g04431(new_n4817, new_n1668, new_n1119);
and_4  g04432(new_n4818, new_n4817, new_n4816);
nand_4 g04433(new_n4819, new_n4818, new_n4815);
nor_4  g04434(new_n4820, new_n1087, new_n553);
and_4  g04435(new_n4821, new_n4820, new_n562);
nor_4  g04436(new_n4822, new_n2154, new_n1704);
and_4  g04437(new_n4823, new_n4822, new_n1680);
nand_4 g04438(new_n4824, new_n4823, new_n4821);
nor_4  g04439(new_n4825, new_n4824, new_n4819);
nand_4 g04440(new_n4826, new_n4825, new_n4814);
nor_4  g04441(new_n4827, new_n4826, new_n4804);
not_3  g04442(new_n4828, new_n1049);
nor_4  g04443(new_n4829, new_n1098, new_n993);
nand_4 g04444(new_n4830, new_n4829, new_n4828);
nor_4  g04445(new_n4831, new_n1717, new_n1343);
nor_4  g04446(new_n4832, new_n493, new_n469);
nor_4  g04447(new_n4833, new_n1753, new_n1334);
and_4  g04448(new_n4834, new_n4833, new_n4832);
nand_4 g04449(new_n4835, new_n4834, new_n4831);
nor_4  g04450(new_n4836, new_n972, new_n579);
nor_4  g04451(new_n4837, new_n1651, new_n1246);
and_4  g04452(new_n4838, new_n4837, new_n4836);
nor_4  g04453(new_n4839, new_n1316, new_n1283);
nor_4  g04454(new_n4840, new_n1635, new_n1250);
and_4  g04455(new_n4841, new_n4840, new_n4839);
nand_4 g04456(new_n4842, new_n4841, new_n4838);
nor_4  g04457(new_n4843, new_n4842, new_n4835);
nor_4  g04458(new_n4844, new_n1105, new_n1009);
nor_4  g04459(new_n4845, new_n1069, new_n543_1);
nand_4 g04460(new_n4846, new_n4845, new_n573);
nor_4  g04461(new_n4847, new_n2167, new_n1698);
nand_4 g04462(new_n4848, new_n4847, new_n1688);
nor_4  g04463(new_n4849, new_n4848, new_n4846);
and_4  g04464(new_n4850, new_n4849, new_n4844);
nand_4 g04465(new_n4851, new_n4850, new_n4843);
nor_4  g04466(new_n4852, new_n4851, new_n4830);
nand_4 g04467(n3340, new_n4852, new_n4827);
not_3  g04468(new_n4854, n6460);
not_3  g04469(new_n4855, new_n2150);
nand_4 g04470(new_n4856, new_n4855, new_n4854);
nand_4 g04471(new_n4857, new_n4856, new_n437);
nand_4 g04472(new_n4858_1, new_n4857, new_n841);
nand_4 g04473(new_n4859, new_n4858_1, new_n434);
nand_4 g04474(new_n4860, new_n4859, new_n429);
nand_4 g04475(new_n4861, new_n4860, new_n424);
nand_4 g04476(new_n4862, new_n4861, new_n850);
nand_4 g04477(new_n4863, new_n4862, new_n856);
nand_4 g04478(new_n4864, new_n4863, new_n863);
nand_4 g04479(new_n4865, new_n4864, new_n419);
nand_4 g04480(new_n4866, new_n4865, new_n869);
nand_4 g04481(new_n4867, new_n4866, new_n875);
nand_4 g04482(new_n4868, new_n4867, new_n881);
nand_4 g04483(new_n4869, new_n4868, new_n413);
nand_4 g04484(new_n4870, new_n4869, new_n889);
nand_4 g04485(new_n4871, new_n4870, new_n896);
nand_4 g04486(new_n4872, new_n4871, new_n901);
nand_4 g04487(new_n4873, new_n4872, new_n408);
nand_4 g04488(new_n4874, new_n4873, new_n908);
nand_4 g04489(new_n4875, new_n4874, new_n403);
nand_4 g04490(new_n4876, new_n4875, new_n398);
nand_4 g04491(new_n4877, new_n4876, new_n393);
nand_4 g04492(new_n4878, new_n4877, new_n916);
nand_4 g04493(new_n4879, new_n4878, new_n1123);
nand_4 g04494(new_n4880, new_n4879, new_n1164);
nand_4 g04495(new_n4881, new_n4880, new_n1120);
nand_4 g04496(new_n4882, new_n4881, new_n1169);
nand_4 g04497(new_n4883, new_n4882, new_n1116);
nand_4 g04498(new_n4884, new_n4883, new_n1111);
nand_4 g04499(new_n4885, new_n4884, new_n1106);
nand_4 g04500(new_n4886, new_n4885, new_n1178);
nand_4 g04501(new_n4887, new_n4886, new_n1183);
nand_4 g04502(new_n4888, new_n4887, new_n1102);
nand_4 g04503(new_n4889, new_n4888, new_n1099);
nand_4 g04504(new_n4890, new_n4889, new_n1191);
nand_4 g04505(new_n4891, new_n4890, new_n1095);
nand_4 g04506(new_n4892, new_n4891, new_n1091);
nand_4 g04507(new_n4893, new_n4892, new_n1088);
nand_4 g04508(new_n4894, new_n4893, new_n1084);
nand_4 g04509(new_n4895_1, new_n4894, new_n1079);
nand_4 g04510(new_n4896, new_n4895_1, new_n1074);
nand_4 g04511(new_n4897, new_n4896, new_n1070);
nand_4 g04512(new_n4898, new_n4897, new_n1064);
nand_4 g04513(new_n4899, new_n4898, new_n1061);
nand_4 g04514(new_n4900, new_n4899, new_n1055);
nand_4 g04515(new_n4901, new_n4900, new_n1050);
not_3  g04516(new_n4902, new_n4901);
nor_4  g04517(new_n4903, new_n4902, new_n1046);
nor_4  g04518(new_n4904, new_n4903, new_n1042);
nor_4  g04519(new_n4905, new_n4904, new_n1037);
nor_4  g04520(new_n4906, new_n4905, new_n1032);
nor_4  g04521(new_n4907_1, new_n4906, new_n1026);
nor_4  g04522(new_n4908, new_n4907_1, new_n1021);
nor_4  g04523(new_n4909, new_n4908, new_n1016);
nor_4  g04524(new_n4910, new_n4909, new_n1011);
nor_4  g04525(new_n4911, new_n4910, new_n1216);
nor_4  g04526(new_n4912, new_n4911, new_n1006);
nor_4  g04527(new_n4913, new_n4912, new_n1001);
nor_4  g04528(new_n4914, new_n4913, new_n995);
nor_4  g04529(new_n4915, new_n4914, new_n990);
nor_4  g04530(new_n4916, new_n4915, new_n985);
nor_4  g04531(new_n4917, new_n4916, new_n979);
nor_4  g04532(new_n4918, new_n4917, new_n974);
nor_4  g04533(new_n4919, new_n4918, new_n968);
nor_4  g04534(new_n4920, new_n4919, new_n965);
nor_4  g04535(new_n4921, new_n4920, new_n961);
nor_4  g04536(new_n4922, new_n4921, new_n958);
nor_4  g04537(new_n4923, new_n4922, new_n953);
nor_4  g04538(new_n4924, new_n4923, new_n3536);
nor_4  g04539(new_n4925, new_n4924, new_n3535);
nor_4  g04540(new_n4926, new_n4925, new_n3534);
not_3  g04541(new_n4927, new_n4926);
nand_4 g04542(new_n4928, new_n4927, new_n934);
nand_4 g04543(new_n4929, new_n4928, new_n929);
nand_4 g04544(new_n4930, new_n4929, new_n925);
nand_4 g04545(new_n4931, new_n4930, new_n2194);
nand_4 g04546(new_n4932, new_n4931, new_n2191);
nand_4 g04547(new_n4933, new_n4932, new_n2190);
nand_4 g04548(new_n4934, new_n4933, new_n2186);
nand_4 g04549(new_n4935, new_n4934, new_n2183);
nand_4 g04550(new_n4936, new_n4935, new_n2179);
nand_4 g04551(new_n4937, new_n4936, new_n2175_1);
nand_4 g04552(new_n4938, new_n4937, new_n2171);
nand_4 g04553(new_n4939, new_n4938, new_n2168);
nand_4 g04554(new_n4940, new_n4939, new_n2165);
nand_4 g04555(new_n4941, new_n4940, new_n2162);
nand_4 g04556(new_n4942, new_n4941, new_n2158);
nand_4 g04557(new_n4943, new_n4942, n3130);
nor_4  g04558(n3603, new_n4943, new_n2152);
nand_4 g04559(new_n4945, new_n1063, new_n542);
nand_4 g04560(new_n4946, new_n4945, new_n660);
nand_4 g04561(new_n4947, new_n4946, new_n539);
nand_4 g04562(new_n4948, new_n4947, new_n534);
nand_4 g04563(new_n4949, new_n4948, new_n529);
nand_4 g04564(new_n4950, new_n4949, new_n668);
nand_4 g04565(new_n4951, new_n4950, new_n674_1);
nand_4 g04566(new_n4952, new_n4951, new_n681);
nand_4 g04567(new_n4953, new_n4952, new_n523);
nand_4 g04568(new_n4954, new_n4953, new_n687);
nand_4 g04569(new_n4955, new_n4954, new_n693);
nand_4 g04570(new_n4956, new_n4955, new_n699);
nand_4 g04571(new_n4957, new_n4956, new_n517);
nand_4 g04572(new_n4958, new_n4957, new_n705);
nand_4 g04573(new_n4959, new_n4958, new_n511);
nand_4 g04574(new_n4960, new_n4959, new_n711);
nand_4 g04575(new_n4961, new_n4960, new_n506);
nand_4 g04576(new_n4962, new_n4961, new_n719);
nand_4 g04577(new_n4963, new_n4962, new_n500);
nand_4 g04578(new_n4964, new_n4963, new_n727);
nand_4 g04579(new_n4965, new_n4964, new_n494);
nand_4 g04580(new_n4966, new_n4965, new_n735);
nand_4 g04581(new_n4967, new_n4966, new_n488);
nand_4 g04582(new_n4968, new_n4967, new_n743);
nand_4 g04583(new_n4969, new_n4968, new_n482);
nand_4 g04584(new_n4970, new_n4969, new_n751);
nand_4 g04585(new_n4971_1, new_n4970, new_n758);
nand_4 g04586(new_n4972, new_n4971_1, new_n765);
nand_4 g04587(new_n4973, new_n4972, new_n476);
nand_4 g04588(new_n4974, new_n4973, new_n773);
nand_4 g04589(new_n4975, new_n4974, new_n780);
nand_4 g04590(new_n4976, new_n4975, new_n787);
nand_4 g04591(new_n4977, new_n4976, new_n470);
nand_4 g04592(new_n4978, new_n4977, new_n795);
nand_4 g04593(new_n4979, new_n4978, new_n803);
nand_4 g04594(new_n4980, new_n4979, new_n809);
nand_4 g04595(new_n4981, new_n4980, new_n465);
nand_4 g04596(new_n4982, new_n4981, new_n818);
nand_4 g04597(new_n4983, new_n4982, new_n460);
nand_4 g04598(new_n4984, new_n4983, new_n455);
nand_4 g04599(new_n4985, new_n4984, new_n449);
nand_4 g04600(new_n4986, new_n4985, new_n827);
nand_4 g04601(new_n4987, new_n4986, new_n833);
nand_4 g04602(new_n4988, new_n4987, new_n444);
nand_4 g04603(new_n4989, new_n4988, new_n439);
nand_4 g04604(new_n4990, new_n4989, new_n841);
nand_4 g04605(new_n4991, new_n4990, new_n434);
nand_4 g04606(new_n4992, new_n4991, new_n429);
nand_4 g04607(new_n4993, new_n4992, new_n424);
nand_4 g04608(new_n4994, new_n4993, new_n850);
nand_4 g04609(new_n4995, new_n4994, new_n856);
not_3  g04610(new_n4996, new_n4995);
nor_4  g04611(new_n4997, new_n4996, new_n2028);
nor_4  g04612(new_n4998, new_n4997, new_n2027_1);
nor_4  g04613(new_n4999, new_n4998, new_n2026);
nor_4  g04614(new_n5000, new_n4999, new_n2025);
nor_4  g04615(new_n5001, new_n5000, new_n2024);
nor_4  g04616(new_n5002, new_n5001, new_n2023);
nor_4  g04617(new_n5003, new_n5002, new_n2022);
nor_4  g04618(new_n5004, new_n5003, new_n2021);
nor_4  g04619(new_n5005, new_n5004, new_n2020);
nor_4  g04620(new_n5006, new_n5005, new_n2019);
nor_4  g04621(new_n5007, new_n5006, new_n1537);
nor_4  g04622(new_n5008, new_n5007, new_n1536);
nor_4  g04623(new_n5009_1, new_n5008, new_n1535);
nor_4  g04624(new_n5010, new_n5009_1, new_n1534);
nor_4  g04625(new_n5011, new_n5010, new_n1533);
nor_4  g04626(new_n5012, new_n5011, new_n1532);
nor_4  g04627(new_n5013, new_n5012, new_n1531);
nor_4  g04628(new_n5014_1, new_n5013, new_n1530);
nor_4  g04629(new_n5015, new_n5014_1, new_n1529);
nor_4  g04630(new_n5016, new_n5015, new_n1528);
nor_4  g04631(new_n5017, new_n5016, new_n1527);
nor_4  g04632(new_n5018, new_n5017, new_n1526);
nor_4  g04633(new_n5019, new_n5018, new_n1525);
nor_4  g04634(new_n5020, new_n5019, new_n1524);
nor_4  g04635(new_n5021, new_n5020, new_n1523);
nor_4  g04636(new_n5022, new_n5021, new_n1522);
nor_4  g04637(new_n5023_1, new_n5022, new_n1521);
not_3  g04638(new_n5024, new_n5023_1);
nand_4 g04639(new_n5025, new_n5024, new_n1095);
nand_4 g04640(new_n5026, new_n5025, new_n1091);
nand_4 g04641(new_n5027, new_n5026, new_n1088);
nand_4 g04642(new_n5028, new_n5027, new_n1084);
nand_4 g04643(new_n5029, new_n5028, new_n1079);
nand_4 g04644(new_n5030, new_n5029, new_n1074);
nand_4 g04645(new_n5031, new_n5030, n3799);
nor_4  g04646(n3854, new_n5031, new_n1067);
nand_4 g04647(new_n5033_1, new_n1358, new_n742);
nand_4 g04648(new_n5034, new_n5033_1, new_n1357);
nand_4 g04649(new_n5035, new_n5034, new_n1354);
nand_4 g04650(new_n5036, new_n5035, new_n1352);
nand_4 g04651(new_n5037, new_n5036, new_n1350);
nand_4 g04652(new_n5038, new_n5037, new_n1347_1);
nand_4 g04653(new_n5039, new_n5038, new_n1344);
nand_4 g04654(new_n5040, new_n5039, new_n1341);
nand_4 g04655(new_n5041, new_n5040, new_n1338);
nand_4 g04656(new_n5042, new_n5041, new_n1395);
nand_4 g04657(new_n5043, new_n5042, new_n1335);
nand_4 g04658(new_n5044, new_n5043, new_n1332);
nand_4 g04659(new_n5045, new_n5044, new_n1328);
nand_4 g04660(new_n5046_1, new_n5045, new_n1403);
nand_4 g04661(new_n5047, new_n5046_1, new_n1325);
nand_4 g04662(new_n5048, new_n5047, new_n1410);
nand_4 g04663(new_n5049, new_n5048, new_n1413);
nand_4 g04664(new_n5050, new_n5049, new_n1322);
nand_4 g04665(new_n5051, new_n5050, new_n1317);
nand_4 g04666(new_n5052, new_n5051, new_n1315);
nand_4 g04667(new_n5053, new_n5052, new_n1419);
nand_4 g04668(new_n5054, new_n5053, new_n1310);
nand_4 g04669(new_n5055, new_n5054, new_n1305);
nand_4 g04670(new_n5056, new_n5055, new_n1427);
nand_4 g04671(new_n5057, new_n5056, new_n1431);
nand_4 g04672(new_n5058, new_n5057, new_n1302);
nand_4 g04673(new_n5059, new_n5058, new_n1298);
nand_4 g04674(new_n5060, new_n5059, new_n1295);
nand_4 g04675(new_n5061, new_n5060, new_n1291);
nand_4 g04676(new_n5062, new_n5061, new_n1288);
nand_4 g04677(new_n5063, new_n5062, new_n1284);
nand_4 g04678(new_n5064, new_n5063, new_n1280);
nand_4 g04679(new_n5065, new_n5064, new_n1275);
nand_4 g04680(new_n5066, new_n5065, new_n1445);
nand_4 g04681(new_n5067, new_n5066, new_n1270);
nand_4 g04682(new_n5068, new_n5067, new_n1265_1);
nand_4 g04683(new_n5069, new_n5068, new_n1260);
nand_4 g04684(new_n5070, new_n5069, new_n1256);
nand_4 g04685(new_n5071, new_n5070, new_n1251);
nand_4 g04686(new_n5072, new_n5071, new_n1457);
nand_4 g04687(new_n5073, new_n5072, new_n1462);
nand_4 g04688(new_n5074, new_n5073, new_n1468);
nand_4 g04689(new_n5075, new_n5074, new_n1247);
nand_4 g04690(new_n5076, new_n5075, new_n1474);
nand_4 g04691(new_n5077_1, new_n5076, new_n592);
nand_4 g04692(new_n5078, new_n5077_1, new_n585);
nand_4 g04693(new_n5079, new_n5078, new_n580);
nand_4 g04694(new_n5080, new_n5079, new_n600);
nand_4 g04695(new_n5081, new_n5080, new_n606);
nand_4 g04696(new_n5082, new_n5081, new_n612);
nand_4 g04697(new_n5083, new_n5082, new_n575);
not_3  g04698(new_n5084, new_n5083);
nor_4  g04699(new_n5085, new_n5084, new_n3081);
nor_4  g04700(new_n5086, new_n5085, new_n3080);
nor_4  g04701(new_n5087, new_n5086, new_n3079);
nor_4  g04702(new_n5088, new_n5087, new_n3078);
nor_4  g04703(new_n5089, new_n5088, new_n3077);
nor_4  g04704(new_n5090, new_n5089, new_n3076);
nor_4  g04705(new_n5091, new_n5090, new_n3075);
nor_4  g04706(new_n5092, new_n5091, new_n3074);
nor_4  g04707(new_n5093, new_n5092, new_n3073);
nor_4  g04708(new_n5094, new_n5093, new_n3072);
nor_4  g04709(new_n5095, new_n5094, new_n3071);
nor_4  g04710(new_n5096, new_n5095, new_n3070);
nor_4  g04711(new_n5097, new_n5096, new_n3069);
nor_4  g04712(new_n5098, new_n5097, new_n3068);
nor_4  g04713(new_n5099, new_n5098, new_n3067);
nor_4  g04714(new_n5100, new_n5099, new_n3066);
nor_4  g04715(new_n5101, new_n5100, new_n3065);
nor_4  g04716(new_n5102, new_n5101, new_n3064);
nor_4  g04717(new_n5103, new_n5102, new_n3063);
nor_4  g04718(new_n5104, new_n5103, new_n3062);
nor_4  g04719(new_n5105, new_n5104, new_n3061);
nor_4  g04720(new_n5106, new_n5105, new_n3354);
nor_4  g04721(new_n5107, new_n5106, new_n3353);
nor_4  g04722(new_n5108, new_n5107, new_n3352);
nor_4  g04723(new_n5109, new_n5108, new_n3351);
nor_4  g04724(new_n5110, new_n5109, new_n3350);
nor_4  g04725(new_n5111, new_n5110, new_n3349);
not_3  g04726(new_n5112, new_n5111);
nand_4 g04727(new_n5113, new_n5112, new_n506);
nand_4 g04728(new_n5114, new_n5113, new_n719);
nand_4 g04729(new_n5115, new_n5114, new_n500);
nand_4 g04730(new_n5116, new_n5115, new_n727);
nand_4 g04731(new_n5117, new_n5116, new_n494);
nand_4 g04732(new_n5118, new_n5117, new_n735);
nand_4 g04733(new_n5119, new_n5118, n12573);
nor_4  g04734(n3901, new_n5119, new_n485);
nand_4 g04735(new_n5121, new_n2187, new_n1393);
nand_4 g04736(new_n5122, new_n5121, new_n2190);
nand_4 g04737(new_n5123, new_n5122, new_n2186);
nand_4 g04738(new_n5124, new_n5123, new_n2183);
nand_4 g04739(new_n5125, new_n5124, new_n2179);
nand_4 g04740(new_n5126, new_n5125, new_n2175_1);
nand_4 g04741(new_n5127, new_n5126, new_n2171);
nand_4 g04742(new_n5128, new_n5127, new_n2168);
nand_4 g04743(new_n5129, new_n5128, new_n2165);
nand_4 g04744(new_n5130, new_n5129, new_n2162);
nand_4 g04745(new_n5131, new_n5130, new_n2158);
nand_4 g04746(new_n5132, new_n5131, new_n2155);
nand_4 g04747(new_n5133, new_n5132, new_n2151);
nand_4 g04748(new_n5134, new_n5133, new_n2147);
nand_4 g04749(new_n5135, new_n5134, new_n1810);
nand_4 g04750(new_n5136, new_n5135, new_n1806);
nand_4 g04751(new_n5137, new_n5136, new_n1802);
nand_4 g04752(new_n5138, new_n5137, new_n1798);
nand_4 g04753(new_n5139, new_n5138, new_n1820);
nand_4 g04754(new_n5140, new_n5139, new_n1794);
nand_4 g04755(new_n5141, new_n5140, new_n1825);
nand_4 g04756(new_n5142, new_n5141, new_n1789);
nand_4 g04757(new_n5143, new_n5142, new_n1785);
nand_4 g04758(new_n5144, new_n5143, new_n1780);
nand_4 g04759(new_n5145, new_n5144, new_n1777);
nand_4 g04760(new_n5146, new_n5145, new_n1774);
nand_4 g04761(new_n5147, new_n5146, new_n1834);
nand_4 g04762(new_n5148, new_n5147, new_n1769);
nand_4 g04763(new_n5149, new_n5148, new_n1766);
nand_4 g04764(new_n5150, new_n5149, new_n1762);
nand_4 g04765(new_n5151, new_n5150, new_n1758);
nand_4 g04766(new_n5152, new_n5151, new_n1754);
nand_4 g04767(new_n5153, new_n5152, new_n1751);
nand_4 g04768(new_n5154, new_n5153, new_n1748);
nand_4 g04769(new_n5155, new_n5154, new_n1746);
nand_4 g04770(new_n5156, new_n5155, new_n1742);
not_3  g04771(new_n5157, new_n5156);
nor_4  g04772(new_n5158, new_n5157, new_n2287);
nor_4  g04773(new_n5159, new_n5158, new_n2286);
nor_4  g04774(new_n5160, new_n5159, new_n2285);
nor_4  g04775(new_n5161, new_n5160, new_n2284);
nor_4  g04776(new_n5162, new_n5161, new_n2283);
nor_4  g04777(new_n5163, new_n5162, new_n2145);
nor_4  g04778(new_n5164, new_n5163, new_n2144);
nor_4  g04779(new_n5165, new_n5164, new_n2143);
nor_4  g04780(new_n5166, new_n5165, new_n2142);
nor_4  g04781(new_n5167, new_n5166, new_n2141);
nor_4  g04782(new_n5168, new_n5167, new_n2140);
nor_4  g04783(new_n5169, new_n5168, new_n2139);
nor_4  g04784(new_n5170, new_n5169, new_n2138);
nor_4  g04785(new_n5171, new_n5170, new_n2137);
nor_4  g04786(new_n5172, new_n5171, new_n2136);
nor_4  g04787(new_n5173, new_n5172, new_n2135);
nor_4  g04788(new_n5174, new_n5173, new_n2134);
nor_4  g04789(new_n5175, new_n5174, new_n2133);
nor_4  g04790(new_n5176, new_n5175, new_n2132);
not_3  g04791(new_n5177, new_n5176);
nand_4 g04792(new_n5178, new_n5177, new_n1690);
nand_4 g04793(new_n5179, new_n5178, new_n1878);
nand_4 g04794(new_n5180, new_n5179, new_n1882);
nand_4 g04795(new_n5181, new_n5180, new_n1686);
nand_4 g04796(new_n5182, new_n5181, new_n1682);
nand_4 g04797(new_n5183, new_n5182, new_n1678);
nand_4 g04798(new_n5184_1, new_n5183, new_n1674);
nand_4 g04799(new_n5185_1, new_n5184_1, new_n1890);
nand_4 g04800(new_n5186, new_n5185_1, new_n1669);
nand_4 g04801(new_n5187, new_n5186, new_n1665);
nand_4 g04802(new_n5188, new_n5187, new_n1661);
nand_4 g04803(new_n5189, new_n5188, new_n1657);
nand_4 g04804(new_n5190, new_n5189, new_n1652);
nand_4 g04805(new_n5191, new_n5190, new_n1648);
nand_4 g04806(new_n5192, new_n5191, new_n1644);
nand_4 g04807(new_n5193, new_n5192, new_n1640);
nand_4 g04808(new_n5194, new_n5193, new_n1636);
nand_4 g04809(new_n5195, new_n5194, new_n1632);
nand_4 g04810(new_n5196, new_n5195, new_n1378);
nand_4 g04811(new_n5197, new_n5196, new_n1372);
nand_4 g04812(new_n5198, new_n5197, new_n1367);
nand_4 g04813(new_n5199, new_n5198, new_n1363);
nand_4 g04814(new_n5200, new_n5199, new_n1360);
nand_4 g04815(new_n5201, new_n5200, new_n1357);
nand_4 g04816(new_n5202, new_n5201, new_n1354);
nand_4 g04817(new_n5203, new_n5202, new_n1352);
nand_4 g04818(new_n5204, new_n5203, new_n1350);
nand_4 g04819(new_n5205, new_n5204, new_n1347_1);
nand_4 g04820(new_n5206, new_n5205, new_n1344);
nand_4 g04821(new_n5207, new_n5206, new_n1341);
nand_4 g04822(new_n5208, new_n5207, n427);
nor_4  g04823(n4125, new_n5208, new_n784);
not_3  g04824(new_n5210, new_n749);
nand_4 g04825(new_n5211, new_n1354, new_n5210);
nand_4 g04826(new_n5212, new_n5211, new_n1352);
nand_4 g04827(new_n5213, new_n5212, new_n1350);
nand_4 g04828(new_n5214, new_n5213, new_n1347_1);
nand_4 g04829(new_n5215, new_n5214, new_n1344);
nand_4 g04830(new_n5216, new_n5215, new_n1341);
nand_4 g04831(new_n5217, new_n5216, new_n1338);
nand_4 g04832(new_n5218, new_n5217, new_n1395);
nand_4 g04833(new_n5219, new_n5218, new_n1335);
nand_4 g04834(new_n5220, new_n5219, new_n1332);
nand_4 g04835(new_n5221, new_n5220, new_n1328);
nand_4 g04836(new_n5222, new_n5221, new_n1403);
nand_4 g04837(new_n5223, new_n5222, new_n1325);
nand_4 g04838(new_n5224, new_n5223, new_n1410);
nand_4 g04839(new_n5225_1, new_n5224, new_n1413);
nand_4 g04840(new_n5226, new_n5225_1, new_n1322);
nand_4 g04841(new_n5227, new_n5226, new_n1317);
nand_4 g04842(new_n5228, new_n5227, new_n1315);
nand_4 g04843(new_n5229, new_n5228, new_n1419);
nand_4 g04844(new_n5230, new_n5229, new_n1310);
nand_4 g04845(new_n5231, new_n5230, new_n1305);
nand_4 g04846(new_n5232, new_n5231, new_n1427);
nand_4 g04847(new_n5233, new_n5232, new_n1431);
nand_4 g04848(new_n5234, new_n5233, new_n1302);
nand_4 g04849(new_n5235, new_n5234, new_n1298);
nand_4 g04850(new_n5236, new_n5235, new_n1295);
nand_4 g04851(new_n5237, new_n5236, new_n1291);
nand_4 g04852(new_n5238, new_n5237, new_n1288);
nand_4 g04853(new_n5239, new_n5238, new_n1284);
nand_4 g04854(new_n5240, new_n5239, new_n1280);
nand_4 g04855(new_n5241, new_n5240, new_n1275);
nand_4 g04856(new_n5242, new_n5241, new_n1445);
nand_4 g04857(new_n5243, new_n5242, new_n1270);
nand_4 g04858(new_n5244, new_n5243, new_n1265_1);
nand_4 g04859(new_n5245, new_n5244, new_n1260);
nand_4 g04860(new_n5246, new_n5245, new_n1256);
nand_4 g04861(new_n5247, new_n5246, new_n1251);
nand_4 g04862(new_n5248, new_n5247, new_n1457);
nand_4 g04863(new_n5249, new_n5248, new_n1462);
nand_4 g04864(new_n5250, new_n5249, new_n1468);
nand_4 g04865(new_n5251, new_n5250, new_n1247);
nand_4 g04866(new_n5252, new_n5251, new_n1474);
nand_4 g04867(new_n5253, new_n5252, new_n592);
nand_4 g04868(new_n5254, new_n5253, new_n585);
nand_4 g04869(new_n5255, new_n5254, new_n580);
nand_4 g04870(new_n5256, new_n5255, new_n600);
nand_4 g04871(new_n5257, new_n5256, new_n606);
nand_4 g04872(new_n5258, new_n5257, new_n612);
nand_4 g04873(new_n5259, new_n5258, new_n575);
nand_4 g04874(new_n5260, new_n5259, new_n619);
nand_4 g04875(new_n5261, new_n5260, new_n570);
not_3  g04876(new_n5262, new_n5261);
nor_4  g04877(new_n5263, new_n5262, new_n3079);
nor_4  g04878(new_n5264, new_n5263, new_n3078);
nor_4  g04879(new_n5265, new_n5264, new_n3077);
nor_4  g04880(new_n5266, new_n5265, new_n3076);
nor_4  g04881(new_n5267, new_n5266, new_n3075);
nor_4  g04882(new_n5268, new_n5267, new_n3074);
nor_4  g04883(new_n5269, new_n5268, new_n3073);
nor_4  g04884(new_n5270, new_n5269, new_n3072);
nor_4  g04885(new_n5271, new_n5270, new_n3071);
nor_4  g04886(new_n5272, new_n5271, new_n3070);
nor_4  g04887(new_n5273, new_n5272, new_n3069);
nor_4  g04888(new_n5274, new_n5273, new_n3068);
nor_4  g04889(new_n5275, new_n5274, new_n3067);
nor_4  g04890(new_n5276, new_n5275, new_n3066);
nor_4  g04891(new_n5277, new_n5276, new_n3065);
nor_4  g04892(new_n5278, new_n5277, new_n3064);
nor_4  g04893(new_n5279, new_n5278, new_n3063);
nor_4  g04894(new_n5280, new_n5279, new_n3062);
nor_4  g04895(new_n5281, new_n5280, new_n3061);
nor_4  g04896(new_n5282, new_n5281, new_n3354);
nor_4  g04897(new_n5283, new_n5282, new_n3353);
nor_4  g04898(new_n5284, new_n5283, new_n3352);
nor_4  g04899(new_n5285, new_n5284, new_n3351);
nor_4  g04900(new_n5286, new_n5285, new_n3350);
nor_4  g04901(new_n5287, new_n5286, new_n3349);
nor_4  g04902(new_n5288, new_n5287, new_n3348);
nor_4  g04903(new_n5289, new_n5288, new_n720);
not_3  g04904(new_n5290, new_n5289);
nand_4 g04905(new_n5291, new_n5290, new_n500);
nand_4 g04906(new_n5292, new_n5291, new_n727);
nand_4 g04907(new_n5293, new_n5292, new_n494);
nand_4 g04908(new_n5294, new_n5293, new_n735);
nand_4 g04909(new_n5295, new_n5294, new_n488);
nand_4 g04910(new_n5296, new_n5295, new_n743);
nand_4 g04911(new_n5297, new_n5296, n10736);
nor_4  g04912(n4279, new_n5297, new_n479);
nand_4 g04913(new_n5299, new_n1659, new_n698);
nand_4 g04914(new_n5300, new_n5299, new_n1657);
nand_4 g04915(new_n5301, new_n5300, new_n1652);
nand_4 g04916(new_n5302, new_n5301, new_n1648);
nand_4 g04917(new_n5303, new_n5302, new_n1644);
nand_4 g04918(new_n5304, new_n5303, new_n1640);
nand_4 g04919(new_n5305, new_n5304, new_n1636);
nand_4 g04920(new_n5306, new_n5305, new_n1632);
nand_4 g04921(new_n5307, new_n5306, new_n1378);
nand_4 g04922(new_n5308, new_n5307, new_n1372);
nand_4 g04923(new_n5309, new_n5308, new_n1367);
nand_4 g04924(new_n5310, new_n5309, new_n1363);
nand_4 g04925(new_n5311, new_n5310, new_n1360);
nand_4 g04926(new_n5312, new_n5311, new_n1357);
nand_4 g04927(new_n5313, new_n5312, new_n1354);
nand_4 g04928(new_n5314, new_n5313, new_n1352);
nand_4 g04929(new_n5315, new_n5314, new_n1350);
nand_4 g04930(new_n5316, new_n5315, new_n1347_1);
nand_4 g04931(new_n5317, new_n5316, new_n1344);
nand_4 g04932(new_n5318, new_n5317, new_n1341);
nand_4 g04933(new_n5319, new_n5318, new_n1338);
nand_4 g04934(new_n5320, new_n5319, new_n1395);
nand_4 g04935(new_n5321, new_n5320, new_n1335);
nand_4 g04936(new_n5322, new_n5321, new_n1332);
nand_4 g04937(new_n5323, new_n5322, new_n1328);
nand_4 g04938(new_n5324, new_n5323, new_n1403);
nand_4 g04939(new_n5325, new_n5324, new_n1325);
nand_4 g04940(new_n5326, new_n5325, new_n1410);
nand_4 g04941(new_n5327, new_n5326, new_n1413);
nand_4 g04942(new_n5328, new_n5327, new_n1322);
nand_4 g04943(new_n5329, new_n5328, new_n1317);
nand_4 g04944(new_n5330, new_n5329, new_n1315);
nand_4 g04945(new_n5331, new_n5330, new_n1419);
nand_4 g04946(new_n5332, new_n5331, new_n1310);
nand_4 g04947(new_n5333, new_n5332, new_n1305);
nand_4 g04948(new_n5334, new_n5333, new_n1427);
nand_4 g04949(new_n5335, new_n5334, new_n1431);
nand_4 g04950(new_n5336, new_n5335, new_n1302);
nand_4 g04951(new_n5337, new_n5336, new_n1298);
nand_4 g04952(new_n5338, new_n5337, new_n1295);
nand_4 g04953(new_n5339, new_n5338, new_n1291);
nand_4 g04954(new_n5340, new_n5339, new_n1288);
not_3  g04955(new_n5341, new_n5340);
nor_4  g04956(new_n5342, new_n5341, new_n2395);
nor_4  g04957(new_n5343, new_n5342, new_n1281);
nor_4  g04958(new_n5344, new_n5343, new_n1276);
nor_4  g04959(new_n5345, new_n5344, new_n1446);
nor_4  g04960(new_n5346, new_n5345, new_n1271);
nor_4  g04961(new_n5347, new_n5346, new_n1266);
nor_4  g04962(new_n5348, new_n5347, new_n1261);
nor_4  g04963(new_n5349, new_n5348, new_n1257);
nor_4  g04964(new_n5350, new_n5349, new_n1252);
nor_4  g04965(new_n5351, new_n5350, new_n1458);
nor_4  g04966(new_n5352, new_n5351, new_n1463);
nor_4  g04967(new_n5353, new_n5352, new_n1469);
nor_4  g04968(new_n5354, new_n5353, new_n1248);
nor_4  g04969(new_n5355, new_n5354, new_n1475);
nor_4  g04970(new_n5356, new_n5355, new_n1244);
nor_4  g04971(new_n5357, new_n5356, new_n1243);
nor_4  g04972(new_n5358, new_n5357, new_n1242);
nor_4  g04973(new_n5359, new_n5358, new_n1241);
nor_4  g04974(new_n5360, new_n5359, new_n1240);
nor_4  g04975(new_n5361, new_n5360, new_n1239);
nor_4  g04976(new_n5362, new_n5361, new_n3082);
nor_4  g04977(new_n5363, new_n5362, new_n3081);
not_3  g04978(new_n5364, new_n5363);
nand_4 g04979(new_n5365, new_n5364, new_n570);
nand_4 g04980(new_n5366, new_n5365, new_n625);
nand_4 g04981(new_n5367, new_n5366, new_n564);
nand_4 g04982(new_n5368, new_n5367, new_n632);
nand_4 g04983(new_n5369, new_n5368, new_n638);
nand_4 g04984(new_n5370, new_n5369, new_n559);
nand_4 g04985(new_n5371, new_n5370, new_n554);
nand_4 g04986(new_n5372, new_n5371, new_n646);
nand_4 g04987(new_n5373, new_n5372, new_n652);
nand_4 g04988(new_n5374, new_n5373, new_n549);
nand_4 g04989(new_n5375, new_n5374, new_n544);
nand_4 g04990(new_n5376, new_n5375, new_n660);
nand_4 g04991(new_n5377, new_n5376, new_n539);
nand_4 g04992(new_n5378, new_n5377, new_n534);
nand_4 g04993(new_n5379, new_n5378, new_n529);
nand_4 g04994(new_n5380, new_n5379, new_n668);
nand_4 g04995(new_n5381, new_n5380, new_n674_1);
nand_4 g04996(new_n5382, new_n5381, new_n681);
nand_4 g04997(new_n5383, new_n5382, new_n523);
nand_4 g04998(new_n5384, new_n5383, new_n687);
nand_4 g04999(new_n5385, new_n5384, n2454);
nor_4  g05000(n4305, new_n5385, new_n690);
nand_4 g05001(new_n5387, new_n1326, new_n808);
nand_4 g05002(new_n5388, new_n5387, new_n1403);
nand_4 g05003(new_n5389, new_n5388, new_n1325);
nand_4 g05004(new_n5390, new_n5389, new_n1410);
nand_4 g05005(new_n5391, new_n5390, new_n1413);
nand_4 g05006(new_n5392, new_n5391, new_n1322);
nand_4 g05007(new_n5393, new_n5392, new_n1317);
nand_4 g05008(new_n5394, new_n5393, new_n1315);
nand_4 g05009(new_n5395, new_n5394, new_n1419);
nand_4 g05010(new_n5396, new_n5395, new_n1310);
nand_4 g05011(new_n5397, new_n5396, new_n1305);
nand_4 g05012(new_n5398, new_n5397, new_n1427);
nand_4 g05013(new_n5399, new_n5398, new_n1431);
nand_4 g05014(new_n5400, new_n5399, new_n1302);
nand_4 g05015(new_n5401, new_n5400, new_n1298);
nand_4 g05016(new_n5402, new_n5401, new_n1295);
nand_4 g05017(new_n5403, new_n5402, new_n1291);
nand_4 g05018(new_n5404, new_n5403, new_n1288);
nand_4 g05019(new_n5405, new_n5404, new_n1284);
nand_4 g05020(new_n5406, new_n5405, new_n1280);
nand_4 g05021(new_n5407, new_n5406, new_n1275);
nand_4 g05022(new_n5408, new_n5407, new_n1445);
nand_4 g05023(new_n5409, new_n5408, new_n1270);
nand_4 g05024(new_n5410, new_n5409, new_n1265_1);
nand_4 g05025(new_n5411, new_n5410, new_n1260);
nand_4 g05026(new_n5412, new_n5411, new_n1256);
nand_4 g05027(new_n5413, new_n5412, new_n1251);
nand_4 g05028(new_n5414, new_n5413, new_n1457);
nand_4 g05029(new_n5415, new_n5414, new_n1462);
nand_4 g05030(new_n5416, new_n5415, new_n1468);
nand_4 g05031(new_n5417, new_n5416, new_n1247);
nand_4 g05032(new_n5418, new_n5417, new_n1474);
nand_4 g05033(new_n5419, new_n5418, new_n592);
nand_4 g05034(new_n5420, new_n5419, new_n585);
nand_4 g05035(new_n5421, new_n5420, new_n580);
nand_4 g05036(new_n5422, new_n5421, new_n600);
nand_4 g05037(new_n5423, new_n5422, new_n606);
nand_4 g05038(new_n5424, new_n5423, new_n612);
nand_4 g05039(new_n5425, new_n5424, new_n575);
nand_4 g05040(new_n5426, new_n5425, new_n619);
nand_4 g05041(new_n5427, new_n5426, new_n570);
nand_4 g05042(new_n5428, new_n5427, new_n625);
nand_4 g05043(new_n5429, new_n5428, new_n564);
nand_4 g05044(new_n5430_1, new_n5429, new_n632);
nand_4 g05045(new_n5431, new_n5430_1, new_n638);
nand_4 g05046(new_n5432, new_n5431, new_n559);
not_3  g05047(new_n5433, new_n5432);
nor_4  g05048(new_n5434, new_n5433, new_n3074);
nor_4  g05049(new_n5435, new_n5434, new_n3073);
nor_4  g05050(new_n5436, new_n5435, new_n3072);
nor_4  g05051(new_n5437, new_n5436, new_n3071);
nor_4  g05052(new_n5438, new_n5437, new_n3070);
nor_4  g05053(new_n5439, new_n5438, new_n3069);
nor_4  g05054(new_n5440, new_n5439, new_n3068);
nor_4  g05055(new_n5441, new_n5440, new_n3067);
nor_4  g05056(new_n5442, new_n5441, new_n3066);
nor_4  g05057(new_n5443, new_n5442, new_n3065);
nor_4  g05058(new_n5444, new_n5443, new_n3064);
nor_4  g05059(new_n5445, new_n5444, new_n3063);
nor_4  g05060(new_n5446, new_n5445, new_n3062);
nor_4  g05061(new_n5447, new_n5446, new_n3061);
nor_4  g05062(new_n5448, new_n5447, new_n3354);
nor_4  g05063(new_n5449_1, new_n5448, new_n3353);
nor_4  g05064(new_n5450, new_n5449_1, new_n3352);
nor_4  g05065(new_n5451, new_n5450, new_n3351);
nor_4  g05066(new_n5452, new_n5451, new_n3350);
nor_4  g05067(new_n5453, new_n5452, new_n3349);
nor_4  g05068(new_n5454, new_n5453, new_n3348);
nor_4  g05069(new_n5455, new_n5454, new_n720);
nor_4  g05070(new_n5456, new_n5455, new_n501);
nor_4  g05071(new_n5457, new_n5456, new_n728);
not_3  g05072(new_n5458, new_n5457);
nand_4 g05073(new_n5459, new_n5458, new_n494);
nand_4 g05074(new_n5460, new_n5459, new_n735);
nand_4 g05075(new_n5461, new_n5460, new_n488);
nand_4 g05076(new_n5462, new_n5461, new_n743);
nand_4 g05077(new_n5463, new_n5462, new_n482);
nand_4 g05078(new_n5464, new_n5463, new_n751);
nand_4 g05079(new_n5465, new_n5464, new_n758);
nand_4 g05080(new_n5466, new_n5465, new_n765);
nand_4 g05081(new_n5467_1, new_n5466, new_n476);
nand_4 g05082(new_n5468, new_n5467_1, new_n773);
nand_4 g05083(new_n5469, new_n5468, new_n780);
nand_4 g05084(new_n5470, new_n5469, new_n787);
nand_4 g05085(new_n5471, new_n5470, new_n470);
nand_4 g05086(new_n5472, new_n5471, new_n795);
nand_4 g05087(new_n5473, new_n5472, n2615);
nor_4  g05088(n4345, new_n5473, new_n799);
not_3  g05089(new_n5475, new_n1213);
nand_4 g05090(new_n5476, new_n5475, new_n517);
nand_4 g05091(new_n5477, new_n5476, new_n705);
nand_4 g05092(new_n5478, new_n5477, new_n511);
nand_4 g05093(new_n5479_1, new_n5478, new_n711);
nand_4 g05094(new_n5480, new_n5479_1, new_n506);
nand_4 g05095(new_n5481, new_n5480, new_n719);
nand_4 g05096(new_n5482, new_n5481, new_n500);
nand_4 g05097(new_n5483, new_n5482, new_n727);
nand_4 g05098(new_n5484, new_n5483, new_n494);
nand_4 g05099(new_n5485, new_n5484, new_n735);
nand_4 g05100(new_n5486, new_n5485, new_n488);
nand_4 g05101(new_n5487, new_n5486, new_n743);
nand_4 g05102(new_n5488, new_n5487, new_n482);
nand_4 g05103(new_n5489, new_n5488, new_n751);
nand_4 g05104(new_n5490, new_n5489, new_n758);
nand_4 g05105(new_n5491, new_n5490, new_n765);
nand_4 g05106(new_n5492, new_n5491, new_n476);
nand_4 g05107(new_n5493, new_n5492, new_n773);
nand_4 g05108(new_n5494, new_n5493, new_n780);
nand_4 g05109(new_n5495, new_n5494, new_n787);
nand_4 g05110(new_n5496, new_n5495, new_n470);
nand_4 g05111(new_n5497, new_n5496, new_n795);
nand_4 g05112(new_n5498, new_n5497, new_n803);
nand_4 g05113(new_n5499, new_n5498, new_n809);
nand_4 g05114(new_n5500, new_n5499, new_n465);
nand_4 g05115(new_n5501, new_n5500, new_n818);
nand_4 g05116(new_n5502_1, new_n5501, new_n460);
nand_4 g05117(new_n5503, new_n5502_1, new_n455);
nand_4 g05118(new_n5504, new_n5503, new_n449);
nand_4 g05119(new_n5505, new_n5504, new_n827);
nand_4 g05120(new_n5506, new_n5505, new_n833);
nand_4 g05121(new_n5507, new_n5506, new_n444);
nand_4 g05122(new_n5508, new_n5507, new_n439);
nand_4 g05123(new_n5509, new_n5508, new_n841);
nand_4 g05124(new_n5510, new_n5509, new_n434);
nand_4 g05125(new_n5511, new_n5510, new_n429);
nand_4 g05126(new_n5512, new_n5511, new_n424);
nand_4 g05127(new_n5513, new_n5512, new_n850);
nand_4 g05128(new_n5514, new_n5513, new_n856);
nand_4 g05129(new_n5515, new_n5514, new_n863);
nand_4 g05130(new_n5516, new_n5515, new_n419);
nand_4 g05131(new_n5517, new_n5516, new_n869);
nand_4 g05132(new_n5518, new_n5517, new_n875);
nand_4 g05133(new_n5519, new_n5518, new_n881);
nand_4 g05134(new_n5520, new_n5519, new_n413);
nand_4 g05135(new_n5521, new_n5520, new_n889);
nand_4 g05136(new_n5522, new_n5521, new_n896);
nand_4 g05137(new_n5523, new_n5522, new_n901);
nand_4 g05138(new_n5524, new_n5523, new_n408);
nand_4 g05139(new_n5525, new_n5524, new_n908);
nand_4 g05140(new_n5526, new_n5525, new_n403);
not_3  g05141(new_n5527, new_n5526);
nor_4  g05142(new_n5528, new_n5527, new_n1535);
nor_4  g05143(new_n5529, new_n5528, new_n1534);
nor_4  g05144(new_n5530, new_n5529, new_n1533);
nor_4  g05145(new_n5531, new_n5530, new_n1532);
nor_4  g05146(new_n5532, new_n5531, new_n1531);
nor_4  g05147(new_n5533, new_n5532, new_n1530);
nor_4  g05148(new_n5534, new_n5533, new_n1529);
nor_4  g05149(new_n5535, new_n5534, new_n1528);
nor_4  g05150(new_n5536, new_n5535, new_n1527);
nor_4  g05151(new_n5537, new_n5536, new_n1526);
nor_4  g05152(new_n5538, new_n5537, new_n1525);
nor_4  g05153(new_n5539, new_n5538, new_n1524);
nor_4  g05154(new_n5540, new_n5539, new_n1523);
nor_4  g05155(new_n5541, new_n5540, new_n1522);
nor_4  g05156(new_n5542, new_n5541, new_n1521);
nor_4  g05157(new_n5543, new_n5542, new_n1520);
nor_4  g05158(new_n5544, new_n5543, new_n1519);
nor_4  g05159(new_n5545, new_n5544, new_n1518);
nor_4  g05160(new_n5546, new_n5545, new_n1517);
nor_4  g05161(new_n5547, new_n5546, new_n1516);
nor_4  g05162(new_n5548, new_n5547, new_n1075);
nor_4  g05163(new_n5549, new_n5548, new_n1071);
nor_4  g05164(new_n5550_1, new_n5549, new_n1065);
nor_4  g05165(new_n5551, new_n5550_1, new_n1062);
nor_4  g05166(new_n5552, new_n5551, new_n1056);
nor_4  g05167(new_n5553, new_n5552, new_n1051);
nor_4  g05168(new_n5554, new_n5553, new_n1046);
not_3  g05169(new_n5555, new_n5554);
nand_4 g05170(new_n5556, new_n5555, new_n1041);
nand_4 g05171(new_n5557, new_n5556, new_n1036);
nand_4 g05172(new_n5558, new_n5557, new_n1031);
nand_4 g05173(new_n5559, new_n5558, new_n1025);
nand_4 g05174(new_n5560, new_n5559, new_n1020);
nand_4 g05175(new_n5561, new_n5560, new_n1015);
nand_4 g05176(new_n5562, new_n5561, n8044);
nor_4  g05177(n4437, new_n5562, new_n1008);
nand_4 g05178(new_n5564, new_n998, new_n508);
nand_4 g05179(new_n5565, new_n5564, new_n511);
nand_4 g05180(new_n5566, new_n5565, new_n711);
nand_4 g05181(new_n5567, new_n5566, new_n506);
nand_4 g05182(new_n5568, new_n5567, new_n719);
nand_4 g05183(new_n5569, new_n5568, new_n500);
nand_4 g05184(new_n5570, new_n5569, new_n727);
nand_4 g05185(new_n5571, new_n5570, new_n494);
nand_4 g05186(new_n5572, new_n5571, new_n735);
nand_4 g05187(new_n5573, new_n5572, new_n488);
nand_4 g05188(new_n5574, new_n5573, new_n743);
nand_4 g05189(new_n5575, new_n5574, new_n482);
nand_4 g05190(new_n5576, new_n5575, new_n751);
nand_4 g05191(new_n5577, new_n5576, new_n758);
nand_4 g05192(new_n5578, new_n5577, new_n765);
nand_4 g05193(new_n5579, new_n5578, new_n476);
nand_4 g05194(new_n5580, new_n5579, new_n773);
nand_4 g05195(new_n5581, new_n5580, new_n780);
nand_4 g05196(new_n5582, new_n5581, new_n787);
nand_4 g05197(new_n5583, new_n5582, new_n470);
nand_4 g05198(new_n5584, new_n5583, new_n795);
nand_4 g05199(new_n5585, new_n5584, new_n803);
nand_4 g05200(new_n5586_1, new_n5585, new_n809);
nand_4 g05201(new_n5587, new_n5586_1, new_n465);
nand_4 g05202(new_n5588, new_n5587, new_n818);
nand_4 g05203(new_n5589, new_n5588, new_n460);
nand_4 g05204(new_n5590, new_n5589, new_n455);
nand_4 g05205(new_n5591, new_n5590, new_n449);
nand_4 g05206(new_n5592, new_n5591, new_n827);
nand_4 g05207(new_n5593, new_n5592, new_n833);
nand_4 g05208(new_n5594, new_n5593, new_n444);
nand_4 g05209(new_n5595, new_n5594, new_n439);
nand_4 g05210(new_n5596, new_n5595, new_n841);
nand_4 g05211(new_n5597, new_n5596, new_n434);
nand_4 g05212(new_n5598, new_n5597, new_n429);
nand_4 g05213(new_n5599, new_n5598, new_n424);
not_3  g05214(new_n5600, new_n5599);
nor_4  g05215(new_n5601_1, new_n5600, new_n2030);
nor_4  g05216(new_n5602, new_n5601_1, new_n2029);
nor_4  g05217(new_n5603, new_n5602, new_n2028);
nor_4  g05218(new_n5604, new_n5603, new_n2027_1);
nor_4  g05219(new_n5605, new_n5604, new_n2026);
nor_4  g05220(new_n5606, new_n5605, new_n2025);
nor_4  g05221(new_n5607, new_n5606, new_n2024);
nor_4  g05222(new_n5608, new_n5607, new_n2023);
nor_4  g05223(new_n5609, new_n5608, new_n2022);
nor_4  g05224(new_n5610, new_n5609, new_n2021);
nor_4  g05225(new_n5611, new_n5610, new_n2020);
nor_4  g05226(new_n5612, new_n5611, new_n2019);
nor_4  g05227(new_n5613, new_n5612, new_n1537);
nor_4  g05228(new_n5614, new_n5613, new_n1536);
nor_4  g05229(new_n5615, new_n5614, new_n1535);
nor_4  g05230(new_n5616, new_n5615, new_n1534);
nor_4  g05231(new_n5617, new_n5616, new_n1533);
nor_4  g05232(new_n5618, new_n5617, new_n1532);
nor_4  g05233(new_n5619, new_n5618, new_n1531);
not_3  g05234(new_n5620, new_n5619);
nand_4 g05235(new_n5621, new_n5620, new_n1120);
nand_4 g05236(new_n5622, new_n5621, new_n1169);
nand_4 g05237(new_n5623, new_n5622, new_n1116);
nand_4 g05238(new_n5624, new_n5623, new_n1111);
nand_4 g05239(new_n5625, new_n5624, new_n1106);
nand_4 g05240(new_n5626, new_n5625, new_n1178);
nand_4 g05241(new_n5627, new_n5626, new_n1183);
nand_4 g05242(new_n5628, new_n5627, new_n1102);
nand_4 g05243(new_n5629, new_n5628, new_n1099);
nand_4 g05244(new_n5630, new_n5629, new_n1191);
nand_4 g05245(new_n5631, new_n5630, new_n1095);
nand_4 g05246(new_n5632, new_n5631, new_n1091);
nand_4 g05247(new_n5633, new_n5632, new_n1088);
nand_4 g05248(new_n5634, new_n5633, new_n1084);
nand_4 g05249(new_n5635, new_n5634, new_n1079);
nand_4 g05250(new_n5636, new_n5635, new_n1074);
nand_4 g05251(new_n5637, new_n5636, new_n1070);
nand_4 g05252(new_n5638, new_n5637, new_n1064);
nand_4 g05253(new_n5639, new_n5638, new_n1061);
nand_4 g05254(new_n5640, new_n5639, new_n1055);
nand_4 g05255(new_n5641, new_n5640, new_n1050);
nand_4 g05256(new_n5642, new_n5641, new_n1045);
nand_4 g05257(new_n5643, new_n5642, new_n1041);
nand_4 g05258(new_n5644, new_n5643, new_n1036);
nand_4 g05259(new_n5645, new_n5644, new_n1031);
nand_4 g05260(new_n5646, new_n5645, new_n1025);
nand_4 g05261(new_n5647, new_n5646, new_n1020);
nand_4 g05262(new_n5648, new_n5647, new_n1015);
nand_4 g05263(new_n5649, new_n5648, new_n1010);
nand_4 g05264(new_n5650, new_n5649, new_n1215);
nand_4 g05265(new_n5651, new_n5650, n5184);
nor_4  g05266(n4541, new_n5651, new_n1002);
not_3  g05267(new_n5653, new_n933);
nand_4 g05268(new_n5654, new_n5653, new_n930);
nand_4 g05269(new_n5655, new_n5654, new_n474);
nand_4 g05270(new_n5656, new_n5655, new_n773);
nand_4 g05271(new_n5657, new_n5656, new_n780);
nand_4 g05272(new_n5658, new_n5657, new_n787);
nand_4 g05273(new_n5659, new_n5658, new_n470);
nand_4 g05274(new_n5660, new_n5659, new_n795);
nand_4 g05275(new_n5661, new_n5660, new_n803);
nand_4 g05276(new_n5662, new_n5661, new_n809);
nand_4 g05277(new_n5663, new_n5662, new_n465);
nand_4 g05278(new_n5664, new_n5663, new_n818);
nand_4 g05279(new_n5665, new_n5664, new_n460);
nand_4 g05280(new_n5666, new_n5665, new_n455);
nand_4 g05281(new_n5667, new_n5666, new_n449);
nand_4 g05282(new_n5668, new_n5667, new_n827);
nand_4 g05283(new_n5669, new_n5668, new_n833);
nand_4 g05284(new_n5670, new_n5669, new_n444);
nand_4 g05285(new_n5671, new_n5670, new_n439);
nand_4 g05286(new_n5672, new_n5671, new_n841);
nand_4 g05287(new_n5673, new_n5672, new_n434);
nand_4 g05288(new_n5674, new_n5673, new_n429);
nand_4 g05289(new_n5675, new_n5674, new_n424);
nand_4 g05290(new_n5676, new_n5675, new_n850);
nand_4 g05291(new_n5677, new_n5676, new_n856);
nand_4 g05292(new_n5678, new_n5677, new_n863);
nand_4 g05293(new_n5679, new_n5678, new_n419);
nand_4 g05294(new_n5680, new_n5679, new_n869);
nand_4 g05295(new_n5681, new_n5680, new_n875);
nand_4 g05296(new_n5682, new_n5681, new_n881);
nand_4 g05297(new_n5683, new_n5682, new_n413);
nand_4 g05298(new_n5684, new_n5683, new_n889);
nand_4 g05299(new_n5685, new_n5684, new_n896);
nand_4 g05300(new_n5686, new_n5685, new_n901);
nand_4 g05301(new_n5687, new_n5686, new_n408);
nand_4 g05302(new_n5688, new_n5687, new_n908);
nand_4 g05303(new_n5689, new_n5688, new_n403);
nand_4 g05304(new_n5690, new_n5689, new_n398);
nand_4 g05305(new_n5691, new_n5690, new_n393);
nand_4 g05306(new_n5692, new_n5691, new_n916);
nand_4 g05307(new_n5693, new_n5692, new_n1123);
nand_4 g05308(new_n5694, new_n5693, new_n1164);
nand_4 g05309(new_n5695, new_n5694, new_n1120);
nand_4 g05310(new_n5696, new_n5695, new_n1169);
nand_4 g05311(new_n5697, new_n5696, new_n1116);
nand_4 g05312(new_n5698, new_n5697, new_n1111);
nand_4 g05313(new_n5699, new_n5698, new_n1106);
not_3  g05314(new_n5700, new_n5699);
nor_4  g05315(new_n5701, new_n5700, new_n1525);
nor_4  g05316(new_n5702, new_n5701, new_n1524);
nor_4  g05317(new_n5703, new_n5702, new_n1523);
nor_4  g05318(new_n5704, new_n5703, new_n1522);
nor_4  g05319(new_n5705, new_n5704, new_n1521);
nor_4  g05320(new_n5706, new_n5705, new_n1520);
nor_4  g05321(new_n5707, new_n5706, new_n1519);
nor_4  g05322(new_n5708, new_n5707, new_n1518);
nor_4  g05323(new_n5709, new_n5708, new_n1517);
nor_4  g05324(new_n5710, new_n5709, new_n1516);
nor_4  g05325(new_n5711, new_n5710, new_n1075);
nor_4  g05326(new_n5712, new_n5711, new_n1071);
nor_4  g05327(new_n5713, new_n5712, new_n1065);
nor_4  g05328(new_n5714, new_n5713, new_n1062);
nor_4  g05329(new_n5715, new_n5714, new_n1056);
nor_4  g05330(new_n5716, new_n5715, new_n1051);
nor_4  g05331(new_n5717, new_n5716, new_n1046);
nor_4  g05332(new_n5718, new_n5717, new_n1042);
nor_4  g05333(new_n5719, new_n5718, new_n1037);
nor_4  g05334(new_n5720, new_n5719, new_n1032);
nor_4  g05335(new_n5721, new_n5720, new_n1026);
nor_4  g05336(new_n5722, new_n5721, new_n1021);
nor_4  g05337(new_n5723, new_n5722, new_n1016);
nor_4  g05338(new_n5724, new_n5723, new_n1011);
not_3  g05339(new_n5725_1, new_n5724);
nand_4 g05340(new_n5726, new_n5725_1, new_n1215);
nand_4 g05341(new_n5727, new_n5726, new_n1005);
nand_4 g05342(new_n5728, new_n5727, new_n1000);
nand_4 g05343(new_n5729, new_n5728, new_n994);
nand_4 g05344(new_n5730, new_n5729, new_n989);
nand_4 g05345(new_n5731, new_n5730, new_n984);
nand_4 g05346(new_n5732, new_n5731, new_n978);
nand_4 g05347(new_n5733, new_n5732, new_n973);
nand_4 g05348(new_n5734, new_n5733, new_n967);
nand_4 g05349(new_n5735, new_n5734, new_n964);
nand_4 g05350(new_n5736, new_n5735, new_n960);
nand_4 g05351(new_n5737, new_n5736, new_n957);
nand_4 g05352(new_n5738, new_n5737, new_n952);
nand_4 g05353(new_n5739, new_n5738, new_n948_1);
nand_4 g05354(new_n5740, new_n5739, new_n943);
nand_4 g05355(new_n5741, new_n5740, n8302);
nor_4  g05356(n4604, new_n5741, new_n936);
not_3  g05357(new_n5743, new_n1796);
not_3  g05358(new_n5744, new_n1819);
nand_4 g05359(new_n5745, new_n5744, new_n1293);
nand_4 g05360(new_n5746, new_n5745, new_n854);
nand_4 g05361(new_n5747, new_n5746, new_n863);
nand_4 g05362(new_n5748, new_n5747, new_n419);
nand_4 g05363(new_n5749, new_n5748, new_n869);
nand_4 g05364(new_n5750, new_n5749, new_n875);
nand_4 g05365(new_n5751, new_n5750, new_n881);
nand_4 g05366(new_n5752, new_n5751, new_n413);
nand_4 g05367(new_n5753, new_n5752, new_n889);
nand_4 g05368(new_n5754, new_n5753, new_n896);
nand_4 g05369(new_n5755, new_n5754, new_n901);
nand_4 g05370(new_n5756, new_n5755, new_n408);
nand_4 g05371(new_n5757, new_n5756, new_n908);
nand_4 g05372(new_n5758, new_n5757, new_n403);
nand_4 g05373(new_n5759, new_n5758, new_n398);
nand_4 g05374(new_n5760, new_n5759, new_n393);
nand_4 g05375(new_n5761, new_n5760, new_n916);
nand_4 g05376(new_n5762, new_n5761, new_n1123);
nand_4 g05377(new_n5763, new_n5762, new_n1164);
nand_4 g05378(new_n5764, new_n5763, new_n1120);
nand_4 g05379(new_n5765, new_n5764, new_n1169);
nand_4 g05380(new_n5766, new_n5765, new_n1116);
nand_4 g05381(new_n5767, new_n5766, new_n1111);
nand_4 g05382(new_n5768, new_n5767, new_n1106);
nand_4 g05383(new_n5769, new_n5768, new_n1178);
nand_4 g05384(new_n5770, new_n5769, new_n1183);
nand_4 g05385(new_n5771, new_n5770, new_n1102);
nand_4 g05386(new_n5772, new_n5771, new_n1099);
nand_4 g05387(new_n5773, new_n5772, new_n1191);
nand_4 g05388(new_n5774, new_n5773, new_n1095);
nand_4 g05389(new_n5775, new_n5774, new_n1091);
nand_4 g05390(new_n5776, new_n5775, new_n1088);
nand_4 g05391(new_n5777, new_n5776, new_n1084);
nand_4 g05392(new_n5778, new_n5777, new_n1079);
nand_4 g05393(new_n5779, new_n5778, new_n1074);
nand_4 g05394(new_n5780, new_n5779, new_n1070);
nand_4 g05395(new_n5781, new_n5780, new_n1064);
nand_4 g05396(new_n5782, new_n5781, new_n1061);
nand_4 g05397(new_n5783, new_n5782, new_n1055);
nand_4 g05398(new_n5784, new_n5783, new_n1050);
nand_4 g05399(new_n5785, new_n5784, new_n1045);
nand_4 g05400(new_n5786_1, new_n5785, new_n1041);
nand_4 g05401(new_n5787, new_n5786_1, new_n1036);
nand_4 g05402(new_n5788, new_n5787, new_n1031);
nand_4 g05403(new_n5789, new_n5788, new_n1025);
nand_4 g05404(new_n5790, new_n5789, new_n1020);
nand_4 g05405(new_n5791, new_n5790, new_n1015);
nand_4 g05406(new_n5792, new_n5791, new_n1010);
nand_4 g05407(new_n5793, new_n5792, new_n1215);
nand_4 g05408(new_n5794, new_n5793, new_n1005);
nand_4 g05409(new_n5795, new_n5794, new_n1000);
not_3  g05410(new_n5796, new_n5795);
nor_4  g05411(new_n5797, new_n5796, new_n995);
nor_4  g05412(new_n5798, new_n5797, new_n990);
nor_4  g05413(new_n5799, new_n5798, new_n985);
nor_4  g05414(new_n5800, new_n5799, new_n979);
nor_4  g05415(new_n5801, new_n5800, new_n974);
nor_4  g05416(new_n5802, new_n5801, new_n968);
nor_4  g05417(new_n5803, new_n5802, new_n965);
nor_4  g05418(new_n5804, new_n5803, new_n961);
nor_4  g05419(new_n5805, new_n5804, new_n958);
nor_4  g05420(new_n5806_1, new_n5805, new_n953);
nor_4  g05421(new_n5807, new_n5806_1, new_n3536);
nor_4  g05422(new_n5808, new_n5807, new_n3535);
nor_4  g05423(new_n5809, new_n5808, new_n3534);
nor_4  g05424(new_n5810, new_n5809, new_n2520);
nor_4  g05425(new_n5811, new_n5810, new_n2519);
nor_4  g05426(new_n5812, new_n5811, new_n2518);
nor_4  g05427(new_n5813, new_n5812, new_n2517);
nor_4  g05428(new_n5814, new_n5813, new_n2516);
nor_4  g05429(new_n5815, new_n5814, new_n2515);
nor_4  g05430(new_n5816, new_n5815, new_n2514);
nor_4  g05431(new_n5817, new_n5816, new_n2513);
nor_4  g05432(new_n5818, new_n5817, new_n2512);
nor_4  g05433(new_n5819, new_n5818, new_n2511);
nor_4  g05434(new_n5820, new_n5819, new_n2510);
nor_4  g05435(new_n5821, new_n5820, new_n2509);
not_3  g05436(new_n5822, new_n5821);
nand_4 g05437(new_n5823, new_n5822, new_n2165);
nand_4 g05438(new_n5824, new_n5823, new_n2162);
nand_4 g05439(new_n5825, new_n5824, new_n2158);
nand_4 g05440(new_n5826, new_n5825, new_n2155);
nand_4 g05441(new_n5827, new_n5826, new_n2151);
nand_4 g05442(new_n5828, new_n5827, new_n2147);
nand_4 g05443(new_n5829, new_n5828, new_n1810);
nand_4 g05444(new_n5830, new_n5829, new_n1806);
nand_4 g05445(new_n5831, new_n5830, new_n1802);
nand_4 g05446(new_n5832, new_n5831, n12976);
nor_4  g05447(n4672, new_n5832, new_n5743);
nand_4 g05448(new_n5834, new_n547, new_n1868);
nand_4 g05449(new_n5835, new_n5834, new_n1871);
nand_4 g05450(new_n5836, new_n5835, new_n1694);
nand_4 g05451(new_n5837, new_n5836, new_n1690);
nand_4 g05452(new_n5838, new_n5837, new_n1878);
nand_4 g05453(new_n5839, new_n5838, new_n1882);
nand_4 g05454(new_n5840, new_n5839, new_n1686);
nand_4 g05455(new_n5841, new_n5840, new_n1682);
nand_4 g05456(new_n5842, new_n5841, new_n1678);
nand_4 g05457(new_n5843, new_n5842, new_n1674);
nand_4 g05458(new_n5844, new_n5843, new_n1890);
nand_4 g05459(new_n5845, new_n5844, new_n1669);
nand_4 g05460(new_n5846, new_n5845, new_n1665);
nand_4 g05461(new_n5847, new_n5846, new_n1661);
nand_4 g05462(new_n5848, new_n5847, new_n1657);
nand_4 g05463(new_n5849, new_n5848, new_n1652);
nand_4 g05464(new_n5850, new_n5849, new_n1648);
nand_4 g05465(new_n5851_1, new_n5850, new_n1644);
nand_4 g05466(new_n5852, new_n5851_1, new_n1640);
nand_4 g05467(new_n5853, new_n5852, new_n1636);
nand_4 g05468(new_n5854, new_n5853, new_n1632);
nand_4 g05469(new_n5855, new_n5854, new_n1378);
nand_4 g05470(new_n5856, new_n5855, new_n1372);
nand_4 g05471(new_n5857, new_n5856, new_n1367);
nand_4 g05472(new_n5858, new_n5857, new_n1363);
nand_4 g05473(new_n5859, new_n5858, new_n1360);
nand_4 g05474(new_n5860, new_n5859, new_n1357);
nand_4 g05475(new_n5861, new_n5860, new_n1354);
nand_4 g05476(new_n5862, new_n5861, new_n1352);
nand_4 g05477(new_n5863, new_n5862, new_n1350);
nand_4 g05478(new_n5864, new_n5863, new_n1347_1);
nand_4 g05479(new_n5865, new_n5864, new_n1344);
nand_4 g05480(new_n5866, new_n5865, new_n1341);
nand_4 g05481(new_n5867, new_n5866, new_n1338);
nand_4 g05482(new_n5868, new_n5867, new_n1395);
nand_4 g05483(new_n5869, new_n5868, new_n1335);
not_3  g05484(new_n5870, new_n5869);
nor_4  g05485(new_n5871, new_n5870, new_n2609);
nor_4  g05486(new_n5872, new_n5871, new_n2413);
nor_4  g05487(new_n5873, new_n5872, new_n2412);
nor_4  g05488(new_n5874, new_n5873, new_n2411);
nor_4  g05489(new_n5875, new_n5874, new_n2410);
nor_4  g05490(new_n5876, new_n5875, new_n2409);
nor_4  g05491(new_n5877, new_n5876, new_n2408);
nor_4  g05492(new_n5878, new_n5877, new_n2407_1);
nor_4  g05493(new_n5879, new_n5878, new_n2406);
nor_4  g05494(new_n5880, new_n5879, new_n2405);
nor_4  g05495(new_n5881, new_n5880, new_n2404);
nor_4  g05496(new_n5882, new_n5881, new_n2403);
nor_4  g05497(new_n5883, new_n5882, new_n2402);
nor_4  g05498(new_n5884, new_n5883, new_n2401);
nor_4  g05499(new_n5885, new_n5884, new_n2400);
nor_4  g05500(new_n5886, new_n5885, new_n2399);
nor_4  g05501(new_n5887, new_n5886, new_n2398);
nor_4  g05502(new_n5888, new_n5887, new_n2397);
nor_4  g05503(new_n5889, new_n5888, new_n2396);
not_3  g05504(new_n5890, new_n5889);
nand_4 g05505(new_n5891, new_n5890, new_n1284);
nand_4 g05506(new_n5892, new_n5891, new_n1280);
nand_4 g05507(new_n5893, new_n5892, new_n1275);
nand_4 g05508(new_n5894, new_n5893, new_n1445);
nand_4 g05509(new_n5895, new_n5894, new_n1270);
nand_4 g05510(new_n5896, new_n5895, new_n1265_1);
nand_4 g05511(new_n5897, new_n5896, new_n1260);
nand_4 g05512(new_n5898, new_n5897, new_n1256);
nand_4 g05513(new_n5899, new_n5898, new_n1251);
nand_4 g05514(new_n5900, new_n5899, new_n1457);
nand_4 g05515(new_n5901, new_n5900, new_n1462);
nand_4 g05516(new_n5902, new_n5901, new_n1468);
nand_4 g05517(new_n5903, new_n5902, new_n1247);
nand_4 g05518(new_n5904, new_n5903, new_n1474);
nand_4 g05519(new_n5905, new_n5904, new_n592);
nand_4 g05520(new_n5906, new_n5905, new_n585);
nand_4 g05521(new_n5907, new_n5906, new_n580);
nand_4 g05522(new_n5908, new_n5907, new_n600);
nand_4 g05523(new_n5909, new_n5908, new_n606);
nand_4 g05524(new_n5910, new_n5909, new_n612);
nand_4 g05525(new_n5911, new_n5910, new_n575);
nand_4 g05526(new_n5912, new_n5911, new_n619);
nand_4 g05527(new_n5913, new_n5912, new_n570);
nand_4 g05528(new_n5914, new_n5913, new_n625);
nand_4 g05529(new_n5915, new_n5914, new_n564);
nand_4 g05530(new_n5916, new_n5915, new_n632);
nand_4 g05531(new_n5917, new_n5916, new_n638);
nand_4 g05532(new_n5918, new_n5917, new_n559);
nand_4 g05533(new_n5919, new_n5918, new_n554);
nand_4 g05534(new_n5920, new_n5919, new_n646);
nand_4 g05535(new_n5921, new_n5920, n3652);
nor_4  g05536(n4858, new_n5921, new_n649);
nand_4 g05537(new_n5923, new_n1731, new_n1114);
nand_4 g05538(new_n5924, new_n5923, new_n1111);
nand_4 g05539(new_n5925, new_n5924, new_n1106);
nand_4 g05540(new_n5926, new_n5925, new_n1178);
nand_4 g05541(new_n5927, new_n5926, new_n1183);
nand_4 g05542(new_n5928, new_n5927, new_n1102);
nand_4 g05543(new_n5929, new_n5928, new_n1099);
nand_4 g05544(new_n5930, new_n5929, new_n1191);
nand_4 g05545(new_n5931, new_n5930, new_n1095);
nand_4 g05546(new_n5932, new_n5931, new_n1091);
nand_4 g05547(new_n5933, new_n5932, new_n1088);
nand_4 g05548(new_n5934, new_n5933, new_n1084);
nand_4 g05549(new_n5935, new_n5934, new_n1079);
nand_4 g05550(new_n5936, new_n5935, new_n1074);
nand_4 g05551(new_n5937, new_n5936, new_n1070);
nand_4 g05552(new_n5938, new_n5937, new_n1064);
nand_4 g05553(new_n5939, new_n5938, new_n1061);
nand_4 g05554(new_n5940, new_n5939, new_n1055);
nand_4 g05555(new_n5941, new_n5940, new_n1050);
nand_4 g05556(new_n5942, new_n5941, new_n1045);
nand_4 g05557(new_n5943_1, new_n5942, new_n1041);
nand_4 g05558(new_n5944, new_n5943_1, new_n1036);
nand_4 g05559(new_n5945, new_n5944, new_n1031);
nand_4 g05560(new_n5946, new_n5945, new_n1025);
nand_4 g05561(new_n5947, new_n5946, new_n1020);
nand_4 g05562(new_n5948, new_n5947, new_n1015);
nand_4 g05563(new_n5949, new_n5948, new_n1010);
nand_4 g05564(new_n5950_1, new_n5949, new_n1215);
nand_4 g05565(new_n5951, new_n5950_1, new_n1005);
nand_4 g05566(new_n5952, new_n5951, new_n1000);
nand_4 g05567(new_n5953, new_n5952, new_n994);
nand_4 g05568(new_n5954, new_n5953, new_n989);
nand_4 g05569(new_n5955, new_n5954, new_n984);
nand_4 g05570(new_n5956, new_n5955, new_n978);
nand_4 g05571(new_n5957, new_n5956, new_n973);
nand_4 g05572(new_n5958, new_n5957, new_n967);
nand_4 g05573(new_n5959, new_n5958, new_n964);
nand_4 g05574(new_n5960_1, new_n5959, new_n960);
nand_4 g05575(new_n5961, new_n5960_1, new_n957);
nand_4 g05576(new_n5962, new_n5961, new_n952);
nand_4 g05577(new_n5963, new_n5962, new_n948_1);
nand_4 g05578(new_n5964, new_n5963, new_n943);
nand_4 g05579(new_n5965, new_n5964, new_n938);
nand_4 g05580(new_n5966, new_n5965, new_n934);
nand_4 g05581(new_n5967, new_n5966, new_n929);
nand_4 g05582(new_n5968, new_n5967, new_n925);
not_3  g05583(new_n5969, new_n5968);
nor_4  g05584(new_n5970, new_n5969, new_n2517);
nor_4  g05585(new_n5971, new_n5970, new_n2516);
nor_4  g05586(new_n5972, new_n5971, new_n2515);
nor_4  g05587(new_n5973, new_n5972, new_n2514);
nor_4  g05588(new_n5974, new_n5973, new_n2513);
nor_4  g05589(new_n5975, new_n5974, new_n2512);
nor_4  g05590(new_n5976, new_n5975, new_n2511);
nor_4  g05591(new_n5977, new_n5976, new_n2510);
nor_4  g05592(new_n5978, new_n5977, new_n2509);
nor_4  g05593(new_n5979, new_n5978, new_n2508);
nor_4  g05594(new_n5980, new_n5979, new_n2507);
nor_4  g05595(new_n5981, new_n5980, new_n2506);
nor_4  g05596(new_n5982, new_n5981, new_n2505);
nor_4  g05597(new_n5983, new_n5982, new_n2504);
nor_4  g05598(new_n5984, new_n5983, new_n2503);
nor_4  g05599(new_n5985, new_n5984, new_n2502);
nor_4  g05600(new_n5986, new_n5985, new_n2790);
nor_4  g05601(new_n5987_1, new_n5986, new_n2789);
nor_4  g05602(new_n5988, new_n5987_1, new_n2788);
nor_4  g05603(new_n5989, new_n5988, new_n2305);
nor_4  g05604(new_n5990, new_n5989, new_n2304);
nor_4  g05605(new_n5991, new_n5990, new_n2303);
nor_4  g05606(new_n5992, new_n5991, new_n2302);
nor_4  g05607(new_n5993, new_n5992, new_n2301);
not_3  g05608(new_n5994, new_n5993);
nand_4 g05609(new_n5995, new_n5994, new_n1780);
nand_4 g05610(new_n5996, new_n5995, new_n1777);
nand_4 g05611(new_n5997, new_n5996, new_n1774);
nand_4 g05612(new_n5998, new_n5997, new_n1834);
nand_4 g05613(new_n5999, new_n5998, new_n1769);
nand_4 g05614(new_n6000, new_n5999, new_n1766);
nand_4 g05615(new_n6001, new_n6000, new_n1762);
nand_4 g05616(new_n6002, new_n6001, new_n1758);
nand_4 g05617(new_n6003, new_n6002, new_n1754);
nand_4 g05618(new_n6004, new_n6003, new_n1751);
nand_4 g05619(new_n6005, new_n6004, new_n1748);
nand_4 g05620(new_n6006, new_n6005, new_n1746);
nand_4 g05621(new_n6007_1, new_n6006, new_n1742);
nand_4 g05622(new_n6008, new_n6007_1, new_n1738);
nand_4 g05623(new_n6009, new_n6008, n1222);
nor_4  g05624(n4971, new_n6009, new_n582);
not_3  g05625(new_n6011, new_n927);
nand_4 g05626(new_n6012_1, new_n924, new_n778);
nand_4 g05627(new_n6013, new_n6012_1, new_n787);
nand_4 g05628(new_n6014, new_n6013, new_n470);
nand_4 g05629(new_n6015, new_n6014, new_n795);
nand_4 g05630(new_n6016, new_n6015, new_n803);
nand_4 g05631(new_n6017, new_n6016, new_n809);
nand_4 g05632(new_n6018, new_n6017, new_n465);
nand_4 g05633(new_n6019, new_n6018, new_n818);
nand_4 g05634(new_n6020, new_n6019, new_n460);
nand_4 g05635(new_n6021, new_n6020, new_n455);
nand_4 g05636(new_n6022, new_n6021, new_n449);
nand_4 g05637(new_n6023, new_n6022, new_n827);
nand_4 g05638(new_n6024, new_n6023, new_n833);
nand_4 g05639(new_n6025, new_n6024, new_n444);
nand_4 g05640(new_n6026, new_n6025, new_n439);
nand_4 g05641(new_n6027, new_n6026, new_n841);
nand_4 g05642(new_n6028, new_n6027, new_n434);
nand_4 g05643(new_n6029, new_n6028, new_n429);
nand_4 g05644(new_n6030, new_n6029, new_n424);
nand_4 g05645(new_n6031, new_n6030, new_n850);
nand_4 g05646(new_n6032, new_n6031, new_n856);
nand_4 g05647(new_n6033, new_n6032, new_n863);
nand_4 g05648(new_n6034, new_n6033, new_n419);
nand_4 g05649(new_n6035, new_n6034, new_n869);
nand_4 g05650(new_n6036, new_n6035, new_n875);
nand_4 g05651(new_n6037, new_n6036, new_n881);
nand_4 g05652(new_n6038, new_n6037, new_n413);
nand_4 g05653(new_n6039, new_n6038, new_n889);
nand_4 g05654(new_n6040, new_n6039, new_n896);
nand_4 g05655(new_n6041, new_n6040, new_n901);
nand_4 g05656(new_n6042, new_n6041, new_n408);
nand_4 g05657(new_n6043, new_n6042, new_n908);
nand_4 g05658(new_n6044, new_n6043, new_n403);
nand_4 g05659(new_n6045, new_n6044, new_n398);
nand_4 g05660(new_n6046, new_n6045, new_n393);
nand_4 g05661(new_n6047, new_n6046, new_n916);
nand_4 g05662(new_n6048, new_n6047, new_n1123);
nand_4 g05663(new_n6049, new_n6048, new_n1164);
nand_4 g05664(new_n6050, new_n6049, new_n1120);
nand_4 g05665(new_n6051, new_n6050, new_n1169);
nand_4 g05666(new_n6052, new_n6051, new_n1116);
nand_4 g05667(new_n6053, new_n6052, new_n1111);
nand_4 g05668(new_n6054_1, new_n6053, new_n1106);
nand_4 g05669(new_n6055, new_n6054_1, new_n1178);
nand_4 g05670(new_n6056, new_n6055, new_n1183);
not_3  g05671(new_n6057, new_n6056);
nor_4  g05672(new_n6058, new_n6057, new_n1523);
nor_4  g05673(new_n6059, new_n6058, new_n1522);
nor_4  g05674(new_n6060, new_n6059, new_n1521);
nor_4  g05675(new_n6061, new_n6060, new_n1520);
nor_4  g05676(new_n6062, new_n6061, new_n1519);
nor_4  g05677(new_n6063, new_n6062, new_n1518);
nor_4  g05678(new_n6064, new_n6063, new_n1517);
nor_4  g05679(new_n6065, new_n6064, new_n1516);
nor_4  g05680(new_n6066, new_n6065, new_n1075);
nor_4  g05681(new_n6067, new_n6066, new_n1071);
nor_4  g05682(new_n6068, new_n6067, new_n1065);
nor_4  g05683(new_n6069, new_n6068, new_n1062);
nor_4  g05684(new_n6070, new_n6069, new_n1056);
nor_4  g05685(new_n6071, new_n6070, new_n1051);
nor_4  g05686(new_n6072, new_n6071, new_n1046);
nor_4  g05687(new_n6073, new_n6072, new_n1042);
nor_4  g05688(new_n6074, new_n6073, new_n1037);
nor_4  g05689(new_n6075, new_n6074, new_n1032);
nor_4  g05690(new_n6076, new_n6075, new_n1026);
nor_4  g05691(new_n6077, new_n6076, new_n1021);
nor_4  g05692(new_n6078, new_n6077, new_n1016);
nor_4  g05693(new_n6079, new_n6078, new_n1011);
nor_4  g05694(new_n6080, new_n6079, new_n1216);
nor_4  g05695(new_n6081, new_n6080, new_n1006);
not_3  g05696(new_n6082, new_n6081);
nand_4 g05697(new_n6083, new_n6082, new_n1000);
nand_4 g05698(new_n6084, new_n6083, new_n994);
nand_4 g05699(new_n6085, new_n6084, new_n989);
nand_4 g05700(new_n6086, new_n6085, new_n984);
nand_4 g05701(new_n6087, new_n6086, new_n978);
nand_4 g05702(new_n6088, new_n6087, new_n973);
nand_4 g05703(new_n6089, new_n6088, new_n967);
nand_4 g05704(new_n6090, new_n6089, new_n964);
nand_4 g05705(new_n6091, new_n6090, new_n960);
nand_4 g05706(new_n6092, new_n6091, new_n957);
nand_4 g05707(new_n6093, new_n6092, new_n952);
nand_4 g05708(new_n6094, new_n6093, new_n948_1);
nand_4 g05709(new_n6095, new_n6094, new_n943);
nand_4 g05710(new_n6096, new_n6095, new_n938);
nand_4 g05711(new_n6097, new_n6096, new_n934);
nand_4 g05712(new_n6098, new_n6097, n14072);
nor_4  g05713(n5479, new_n6098, new_n6011);
nand_4 g05714(new_n6100, new_n1752, new_n1456);
nand_4 g05715(new_n6101, new_n6100, new_n1751);
nand_4 g05716(new_n6102, new_n6101, new_n1748);
nand_4 g05717(new_n6103, new_n6102, new_n1746);
nand_4 g05718(new_n6104, new_n6103, new_n1742);
nand_4 g05719(new_n6105, new_n6104, new_n1738);
nand_4 g05720(new_n6106, new_n6105, new_n1736);
nand_4 g05721(new_n6107, new_n6106, new_n1732);
nand_4 g05722(new_n6108, new_n6107, new_n1729);
nand_4 g05723(new_n6109, new_n6108, new_n1726);
nand_4 g05724(new_n6110, new_n6109, new_n1724);
nand_4 g05725(new_n6111, new_n6110, new_n1721);
nand_4 g05726(new_n6112, new_n6111, new_n1718);
nand_4 g05727(new_n6113, new_n6112, new_n1715);
nand_4 g05728(new_n6114_1, new_n6113, new_n1711);
nand_4 g05729(new_n6115, new_n6114_1, new_n1708);
nand_4 g05730(new_n6116, new_n6115, new_n1705);
nand_4 g05731(new_n6117, new_n6116, new_n1703);
nand_4 g05732(new_n6118, new_n6117, new_n1860);
nand_4 g05733(new_n6119, new_n6118, new_n1864);
nand_4 g05734(new_n6120, new_n6119, new_n1699);
nand_4 g05735(new_n6121, new_n6120, new_n1697);
nand_4 g05736(new_n6122, new_n6121, new_n1871);
nand_4 g05737(new_n6123, new_n6122, new_n1694);
nand_4 g05738(new_n6124, new_n6123, new_n1690);
nand_4 g05739(new_n6125, new_n6124, new_n1878);
nand_4 g05740(new_n6126, new_n6125, new_n1882);
nand_4 g05741(new_n6127, new_n6126, new_n1686);
nand_4 g05742(new_n6128, new_n6127, new_n1682);
nand_4 g05743(new_n6129, new_n6128, new_n1678);
nand_4 g05744(new_n6130, new_n6129, new_n1674);
nand_4 g05745(new_n6131, new_n6130, new_n1890);
nand_4 g05746(new_n6132, new_n6131, new_n1669);
nand_4 g05747(new_n6133, new_n6132, new_n1665);
nand_4 g05748(new_n6134, new_n6133, new_n1661);
nand_4 g05749(new_n6135, new_n6134, new_n1657);
nand_4 g05750(new_n6136, new_n6135, new_n1652);
nand_4 g05751(new_n6137, new_n6136, new_n1648);
nand_4 g05752(new_n6138, new_n6137, new_n1644);
nand_4 g05753(new_n6139, new_n6138, new_n1640);
nand_4 g05754(new_n6140, new_n6139, new_n1636);
nand_4 g05755(new_n6141, new_n6140, new_n1632);
nand_4 g05756(new_n6142, new_n6141, new_n1378);
nand_4 g05757(new_n6143, new_n6142, new_n1372);
nand_4 g05758(new_n6144, new_n6143, new_n1367);
nand_4 g05759(new_n6145, new_n6144, new_n1363);
nand_4 g05760(new_n6146, new_n6145, new_n1360);
nand_4 g05761(new_n6147_1, new_n6146, new_n1357);
nand_4 g05762(new_n6148, new_n6147_1, new_n1354);
nand_4 g05763(new_n6149, new_n6148, new_n1352);
nand_4 g05764(new_n6150, new_n6149, new_n1350);
not_3  g05765(new_n6151, new_n6150);
nor_4  g05766(new_n6152, new_n6151, new_n3719);
nor_4  g05767(new_n6153, new_n6152, new_n3718);
nor_4  g05768(new_n6154, new_n6153, new_n3717);
nor_4  g05769(new_n6155, new_n6154, new_n3716);
nor_4  g05770(new_n6156, new_n6155, new_n2611);
nor_4  g05771(new_n6157, new_n6156, new_n2610);
nor_4  g05772(new_n6158, new_n6157, new_n2609);
nor_4  g05773(new_n6159, new_n6158, new_n2413);
nor_4  g05774(new_n6160, new_n6159, new_n2412);
nor_4  g05775(new_n6161, new_n6160, new_n2411);
nor_4  g05776(new_n6162, new_n6161, new_n2410);
nor_4  g05777(new_n6163, new_n6162, new_n2409);
nor_4  g05778(new_n6164, new_n6163, new_n2408);
nor_4  g05779(new_n6165, new_n6164, new_n2407_1);
nor_4  g05780(new_n6166, new_n6165, new_n2406);
nor_4  g05781(new_n6167, new_n6166, new_n2405);
nor_4  g05782(new_n6168, new_n6167, new_n2404);
nor_4  g05783(new_n6169, new_n6168, new_n2403);
nor_4  g05784(new_n6170, new_n6169, new_n2402);
nor_4  g05785(new_n6171, new_n6170, new_n2401);
nor_4  g05786(new_n6172, new_n6171, new_n2400);
nor_4  g05787(new_n6173, new_n6172, new_n2399);
nor_4  g05788(new_n6174, new_n6173, new_n2398);
nor_4  g05789(new_n6175, new_n6174, new_n2397);
nor_4  g05790(new_n6176, new_n6175, new_n2396);
nor_4  g05791(new_n6177, new_n6176, new_n2395);
nor_4  g05792(new_n6178, new_n6177, new_n1281);
not_3  g05793(new_n6179, new_n6178);
nand_4 g05794(new_n6180, new_n6179, new_n1275);
nand_4 g05795(new_n6181, new_n6180, new_n1445);
nand_4 g05796(new_n6182, new_n6181, new_n1270);
nand_4 g05797(new_n6183, new_n6182, new_n1265_1);
nand_4 g05798(new_n6184, new_n6183, new_n1260);
nand_4 g05799(new_n6185, new_n6184, new_n1256);
nand_4 g05800(new_n6186, new_n6185, n5046);
nor_4  g05801(n5550, new_n6186, new_n905);
not_3  g05802(new_n6188, new_n825);
nand_4 g05803(new_n6189, new_n1317, new_n6188);
nand_4 g05804(new_n6190, new_n6189, new_n1315);
nand_4 g05805(new_n6191, new_n6190, new_n1419);
nand_4 g05806(new_n6192, new_n6191, new_n1310);
nand_4 g05807(new_n6193, new_n6192, new_n1305);
nand_4 g05808(new_n6194, new_n6193, new_n1427);
nand_4 g05809(new_n6195, new_n6194, new_n1431);
nand_4 g05810(new_n6196, new_n6195, new_n1302);
nand_4 g05811(new_n6197, new_n6196, new_n1298);
nand_4 g05812(new_n6198_1, new_n6197, new_n1295);
nand_4 g05813(new_n6199, new_n6198_1, new_n1291);
nand_4 g05814(new_n6200, new_n6199, new_n1288);
nand_4 g05815(new_n6201, new_n6200, new_n1284);
nand_4 g05816(new_n6202, new_n6201, new_n1280);
nand_4 g05817(new_n6203, new_n6202, new_n1275);
nand_4 g05818(new_n6204, new_n6203, new_n1445);
nand_4 g05819(new_n6205, new_n6204, new_n1270);
nand_4 g05820(new_n6206, new_n6205, new_n1265_1);
nand_4 g05821(new_n6207, new_n6206, new_n1260);
nand_4 g05822(new_n6208, new_n6207, new_n1256);
nand_4 g05823(new_n6209, new_n6208, new_n1251);
nand_4 g05824(new_n6210, new_n6209, new_n1457);
nand_4 g05825(new_n6211, new_n6210, new_n1462);
nand_4 g05826(new_n6212, new_n6211, new_n1468);
nand_4 g05827(new_n6213, new_n6212, new_n1247);
nand_4 g05828(new_n6214, new_n6213, new_n1474);
nand_4 g05829(new_n6215, new_n6214, new_n592);
nand_4 g05830(new_n6216, new_n6215, new_n585);
nand_4 g05831(new_n6217, new_n6216, new_n580);
nand_4 g05832(new_n6218, new_n6217, new_n600);
nand_4 g05833(new_n6219, new_n6218, new_n606);
nand_4 g05834(new_n6220, new_n6219, new_n612);
nand_4 g05835(new_n6221, new_n6220, new_n575);
nand_4 g05836(new_n6222, new_n6221, new_n619);
nand_4 g05837(new_n6223, new_n6222, new_n570);
nand_4 g05838(new_n6224, new_n6223, new_n625);
nand_4 g05839(new_n6225, new_n6224, new_n564);
nand_4 g05840(new_n6226, new_n6225, new_n632);
nand_4 g05841(new_n6227, new_n6226, new_n638);
nand_4 g05842(new_n6228, new_n6227, new_n559);
nand_4 g05843(new_n6229, new_n6228, new_n554);
nand_4 g05844(new_n6230, new_n6229, new_n646);
not_3  g05845(new_n6231, new_n6230);
nor_4  g05846(new_n6232, new_n6231, new_n3072);
nor_4  g05847(new_n6233, new_n6232, new_n3071);
nor_4  g05848(new_n6234, new_n6233, new_n3070);
nor_4  g05849(new_n6235, new_n6234, new_n3069);
nor_4  g05850(new_n6236, new_n6235, new_n3068);
nor_4  g05851(new_n6237, new_n6236, new_n3067);
nor_4  g05852(new_n6238, new_n6237, new_n3066);
nor_4  g05853(new_n6239, new_n6238, new_n3065);
nor_4  g05854(new_n6240, new_n6239, new_n3064);
nor_4  g05855(new_n6241, new_n6240, new_n3063);
nor_4  g05856(new_n6242, new_n6241, new_n3062);
nor_4  g05857(new_n6243, new_n6242, new_n3061);
nor_4  g05858(new_n6244, new_n6243, new_n3354);
nor_4  g05859(new_n6245, new_n6244, new_n3353);
nor_4  g05860(new_n6246, new_n6245, new_n3352);
nor_4  g05861(new_n6247, new_n6246, new_n3351);
nor_4  g05862(new_n6248, new_n6247, new_n3350);
nor_4  g05863(new_n6249, new_n6248, new_n3349);
nor_4  g05864(new_n6250, new_n6249, new_n3348);
nor_4  g05865(new_n6251_1, new_n6250, new_n720);
nor_4  g05866(new_n6252, new_n6251_1, new_n501);
nor_4  g05867(new_n6253, new_n6252, new_n728);
not_3  g05868(new_n6254, new_n6253);
nand_4 g05869(new_n6255, new_n6254, new_n494);
nand_4 g05870(new_n6256, new_n6255, new_n735);
nand_4 g05871(new_n6257, new_n6256, new_n488);
nand_4 g05872(new_n6258_1, new_n6257, new_n743);
nand_4 g05873(new_n6259, new_n6258_1, new_n482);
nand_4 g05874(new_n6260, new_n6259, new_n751);
nand_4 g05875(new_n6261, new_n6260, new_n758);
nand_4 g05876(new_n6262, new_n6261, new_n765);
nand_4 g05877(new_n6263, new_n6262, new_n476);
nand_4 g05878(new_n6264, new_n6263, new_n773);
nand_4 g05879(new_n6265, new_n6264, new_n780);
nand_4 g05880(new_n6266, new_n6265, new_n787);
nand_4 g05881(new_n6267, new_n6266, new_n470);
nand_4 g05882(new_n6268, new_n6267, new_n795);
nand_4 g05883(new_n6269, new_n6268, new_n803);
nand_4 g05884(new_n6270_1, new_n6269, new_n809);
nand_4 g05885(new_n6271, new_n6270_1, new_n465);
nand_4 g05886(new_n6272, new_n6271, new_n818);
nand_4 g05887(new_n6273, new_n6272, new_n460);
nand_4 g05888(new_n6274, new_n6273, new_n455);
nand_4 g05889(new_n6275_1, new_n6274, n8552);
nor_4  g05890(n5586, new_n6275_1, new_n446);
nand_4 g05891(new_n6277, new_n1685, new_n1039);
nand_4 g05892(new_n6278, new_n6277, new_n1036);
nand_4 g05893(new_n6279, new_n6278, new_n1031);
nand_4 g05894(new_n6280, new_n6279, new_n1025);
nand_4 g05895(new_n6281, new_n6280, new_n1020);
nand_4 g05896(new_n6282, new_n6281, new_n1015);
nand_4 g05897(new_n6283, new_n6282, new_n1010);
nand_4 g05898(new_n6284, new_n6283, new_n1215);
nand_4 g05899(new_n6285, new_n6284, new_n1005);
nand_4 g05900(new_n6286, new_n6285, new_n1000);
nand_4 g05901(new_n6287, new_n6286, new_n994);
nand_4 g05902(new_n6288, new_n6287, new_n989);
nand_4 g05903(new_n6289, new_n6288, new_n984);
nand_4 g05904(new_n6290, new_n6289, new_n978);
nand_4 g05905(new_n6291, new_n6290, new_n973);
nand_4 g05906(new_n6292, new_n6291, new_n967);
nand_4 g05907(new_n6293, new_n6292, new_n964);
nand_4 g05908(new_n6294, new_n6293, new_n960);
nand_4 g05909(new_n6295, new_n6294, new_n957);
nand_4 g05910(new_n6296, new_n6295, new_n952);
nand_4 g05911(new_n6297, new_n6296, new_n948_1);
nand_4 g05912(new_n6298, new_n6297, new_n943);
nand_4 g05913(new_n6299, new_n6298, new_n938);
nand_4 g05914(new_n6300, new_n6299, new_n934);
nand_4 g05915(new_n6301, new_n6300, new_n929);
nand_4 g05916(new_n6302, new_n6301, new_n925);
nand_4 g05917(new_n6303, new_n6302, new_n2194);
nand_4 g05918(new_n6304, new_n6303, new_n2191);
nand_4 g05919(new_n6305, new_n6304, new_n2190);
nand_4 g05920(new_n6306, new_n6305, new_n2186);
nand_4 g05921(new_n6307, new_n6306, new_n2183);
nand_4 g05922(new_n6308, new_n6307, new_n2179);
nand_4 g05923(new_n6309, new_n6308, new_n2175_1);
nand_4 g05924(new_n6310, new_n6309, new_n2171);
nand_4 g05925(new_n6311, new_n6310, new_n2168);
nand_4 g05926(new_n6312, new_n6311, new_n2165);
nand_4 g05927(new_n6313, new_n6312, new_n2162);
nand_4 g05928(new_n6314_1, new_n6313, new_n2158);
nand_4 g05929(new_n6315, new_n6314_1, new_n2155);
nand_4 g05930(new_n6316, new_n6315, new_n2151);
nand_4 g05931(new_n6317, new_n6316, new_n2147);
nand_4 g05932(new_n6318, new_n6317, new_n1810);
not_3  g05933(new_n6319, new_n6318);
nor_4  g05934(new_n6320, new_n6319, new_n2790);
nor_4  g05935(new_n6321, new_n6320, new_n2789);
nor_4  g05936(new_n6322, new_n6321, new_n2788);
nor_4  g05937(new_n6323, new_n6322, new_n2305);
nor_4  g05938(new_n6324, new_n6323, new_n2304);
nor_4  g05939(new_n6325, new_n6324, new_n2303);
nor_4  g05940(new_n6326, new_n6325, new_n2302);
nor_4  g05941(new_n6327, new_n6326, new_n2301);
nor_4  g05942(new_n6328, new_n6327, new_n2300);
nor_4  g05943(new_n6329, new_n6328, new_n2299);
nor_4  g05944(new_n6330, new_n6329, new_n2298);
nor_4  g05945(new_n6331, new_n6330, new_n2297);
nor_4  g05946(new_n6332, new_n6331, new_n2296);
nor_4  g05947(new_n6333, new_n6332, new_n2295);
nor_4  g05948(new_n6334, new_n6333, new_n2294);
nor_4  g05949(new_n6335, new_n6334, new_n2293);
nor_4  g05950(new_n6336, new_n6335, new_n2292);
nor_4  g05951(new_n6337, new_n6336, new_n2291);
nor_4  g05952(new_n6338, new_n6337, new_n2290);
nor_4  g05953(new_n6339, new_n6338, new_n2289);
nor_4  g05954(new_n6340, new_n6339, new_n2288);
nor_4  g05955(new_n6341, new_n6340, new_n2287);
not_3  g05956(new_n6342, new_n6341);
nand_4 g05957(new_n6343, new_n6342, new_n1736);
nand_4 g05958(new_n6344, new_n6343, new_n1732);
nand_4 g05959(new_n6345, new_n6344, new_n1729);
nand_4 g05960(new_n6346, new_n6345, new_n1726);
nand_4 g05961(new_n6347, new_n6346, new_n1724);
nand_4 g05962(new_n6348, new_n6347, new_n1721);
nand_4 g05963(new_n6349, new_n6348, new_n1718);
nand_4 g05964(new_n6350, new_n6349, new_n1715);
nand_4 g05965(new_n6351, new_n6350, new_n1711);
nand_4 g05966(new_n6352, new_n6351, new_n1708);
nand_4 g05967(new_n6353, new_n6352, new_n1705);
nand_4 g05968(new_n6354, new_n6353, new_n1703);
nand_4 g05969(new_n6355, new_n6354, new_n1860);
nand_4 g05970(new_n6356, new_n6355, new_n1864);
nand_4 g05971(new_n6357, new_n6356, new_n1699);
nand_4 g05972(new_n6358, new_n6357, new_n1697);
nand_4 g05973(new_n6359, new_n6358, new_n1871);
nand_4 g05974(new_n6360, new_n6359, new_n1694);
nand_4 g05975(new_n6361, new_n6360, new_n1690);
nand_4 g05976(new_n6362_1, new_n6361, new_n1878);
nand_4 g05977(new_n6363, new_n6362_1, n7652);
nor_4  g05978(n5806, new_n6363, new_n531);
not_3  g05979(new_n6365, new_n1765);
nand_4 g05980(new_n6366, new_n6365, new_n1254);
nand_4 g05981(new_n6367, new_n6366, new_n406);
nand_4 g05982(new_n6368, new_n6367, new_n908);
nand_4 g05983(new_n6369, new_n6368, new_n403);
nand_4 g05984(new_n6370, new_n6369, new_n398);
nand_4 g05985(new_n6371, new_n6370, new_n393);
nand_4 g05986(new_n6372, new_n6371, new_n916);
nand_4 g05987(new_n6373, new_n6372, new_n1123);
nand_4 g05988(new_n6374, new_n6373, new_n1164);
nand_4 g05989(new_n6375, new_n6374, new_n1120);
nand_4 g05990(new_n6376, new_n6375, new_n1169);
nand_4 g05991(new_n6377, new_n6376, new_n1116);
nand_4 g05992(new_n6378, new_n6377, new_n1111);
nand_4 g05993(new_n6379, new_n6378, new_n1106);
nand_4 g05994(new_n6380, new_n6379, new_n1178);
nand_4 g05995(new_n6381, new_n6380, new_n1183);
nand_4 g05996(new_n6382, new_n6381, new_n1102);
nand_4 g05997(new_n6383, new_n6382, new_n1099);
nand_4 g05998(new_n6384, new_n6383, new_n1191);
nand_4 g05999(new_n6385, new_n6384, new_n1095);
nand_4 g06000(new_n6386, new_n6385, new_n1091);
nand_4 g06001(new_n6387, new_n6386, new_n1088);
nand_4 g06002(new_n6388, new_n6387, new_n1084);
nand_4 g06003(new_n6389, new_n6388, new_n1079);
nand_4 g06004(new_n6390, new_n6389, new_n1074);
nand_4 g06005(new_n6391, new_n6390, new_n1070);
nand_4 g06006(new_n6392, new_n6391, new_n1064);
nand_4 g06007(new_n6393, new_n6392, new_n1061);
nand_4 g06008(new_n6394, new_n6393, new_n1055);
nand_4 g06009(new_n6395, new_n6394, new_n1050);
nand_4 g06010(new_n6396, new_n6395, new_n1045);
nand_4 g06011(new_n6397, new_n6396, new_n1041);
nand_4 g06012(new_n6398, new_n6397, new_n1036);
nand_4 g06013(new_n6399, new_n6398, new_n1031);
nand_4 g06014(new_n6400, new_n6399, new_n1025);
nand_4 g06015(new_n6401, new_n6400, new_n1020);
nand_4 g06016(new_n6402, new_n6401, new_n1015);
nand_4 g06017(new_n6403, new_n6402, new_n1010);
nand_4 g06018(new_n6404, new_n6403, new_n1215);
nand_4 g06019(new_n6405, new_n6404, new_n1005);
nand_4 g06020(new_n6406, new_n6405, new_n1000);
nand_4 g06021(new_n6407, new_n6406, new_n994);
nand_4 g06022(new_n6408, new_n6407, new_n989);
nand_4 g06023(new_n6409, new_n6408, new_n984);
nand_4 g06024(new_n6410, new_n6409, new_n978);
nand_4 g06025(new_n6411, new_n6410, new_n973);
not_3  g06026(new_n6412, new_n6411);
nor_4  g06027(new_n6413, new_n6412, new_n968);
nor_4  g06028(new_n6414, new_n6413, new_n965);
nor_4  g06029(new_n6415, new_n6414, new_n961);
nor_4  g06030(new_n6416, new_n6415, new_n958);
nor_4  g06031(new_n6417, new_n6416, new_n953);
nor_4  g06032(new_n6418, new_n6417, new_n3536);
nor_4  g06033(new_n6419, new_n6418, new_n3535);
nor_4  g06034(new_n6420, new_n6419, new_n3534);
nor_4  g06035(new_n6421, new_n6420, new_n2520);
nor_4  g06036(new_n6422, new_n6421, new_n2519);
nor_4  g06037(new_n6423, new_n6422, new_n2518);
nor_4  g06038(new_n6424, new_n6423, new_n2517);
nor_4  g06039(new_n6425, new_n6424, new_n2516);
nor_4  g06040(new_n6426, new_n6425, new_n2515);
nor_4  g06041(new_n6427, new_n6426, new_n2514);
nor_4  g06042(new_n6428, new_n6427, new_n2513);
nor_4  g06043(new_n6429, new_n6428, new_n2512);
nor_4  g06044(new_n6430, new_n6429, new_n2511);
nor_4  g06045(new_n6431, new_n6430, new_n2510);
nor_4  g06046(new_n6432, new_n6431, new_n2509);
nor_4  g06047(new_n6433, new_n6432, new_n2508);
nor_4  g06048(new_n6434, new_n6433, new_n2507);
nor_4  g06049(new_n6435, new_n6434, new_n2506);
nor_4  g06050(new_n6436_1, new_n6435, new_n2505);
not_3  g06051(new_n6437, new_n6436_1);
nand_4 g06052(new_n6438, new_n6437, new_n2151);
nand_4 g06053(new_n6439, new_n6438, new_n2147);
nand_4 g06054(new_n6440, new_n6439, new_n1810);
nand_4 g06055(new_n6441, new_n6440, new_n1806);
nand_4 g06056(new_n6442, new_n6441, new_n1802);
nand_4 g06057(new_n6443, new_n6442, new_n1798);
nand_4 g06058(new_n6444, new_n6443, new_n1820);
nand_4 g06059(new_n6445, new_n6444, new_n1794);
nand_4 g06060(new_n6446, new_n6445, new_n1825);
nand_4 g06061(new_n6447, new_n6446, new_n1789);
nand_4 g06062(new_n6448, new_n6447, new_n1785);
nand_4 g06063(new_n6449, new_n6448, new_n1780);
nand_4 g06064(new_n6450, new_n6449, new_n1777);
nand_4 g06065(new_n6451, new_n6450, new_n1774);
nand_4 g06066(new_n6452, new_n6451, new_n1834);
nand_4 g06067(new_n6453, new_n6452, n13944);
nor_4  g06068(n5851, new_n6453, new_n1262);
not_3  g06069(new_n6455, new_n1361);
nand_4 g06070(new_n6456, new_n6455, new_n957);
nand_4 g06071(new_n6457, new_n6456, new_n952);
nand_4 g06072(new_n6458, new_n6457, new_n948_1);
nand_4 g06073(new_n6459, new_n6458, new_n943);
nand_4 g06074(new_n6460_1, new_n6459, new_n938);
nand_4 g06075(new_n6461, new_n6460_1, new_n934);
nand_4 g06076(new_n6462, new_n6461, new_n929);
nand_4 g06077(new_n6463, new_n6462, new_n925);
nand_4 g06078(new_n6464, new_n6463, new_n2194);
nand_4 g06079(new_n6465, new_n6464, new_n2191);
nand_4 g06080(new_n6466, new_n6465, new_n2190);
nand_4 g06081(new_n6467, new_n6466, new_n2186);
nand_4 g06082(new_n6468, new_n6467, new_n2183);
nand_4 g06083(new_n6469, new_n6468, new_n2179);
nand_4 g06084(new_n6470, new_n6469, new_n2175_1);
nand_4 g06085(new_n6471, new_n6470, new_n2171);
nand_4 g06086(new_n6472, new_n6471, new_n2168);
nand_4 g06087(new_n6473, new_n6472, new_n2165);
nand_4 g06088(new_n6474, new_n6473, new_n2162);
nand_4 g06089(new_n6475, new_n6474, new_n2158);
nand_4 g06090(new_n6476, new_n6475, new_n2155);
nand_4 g06091(new_n6477, new_n6476, new_n2151);
nand_4 g06092(new_n6478, new_n6477, new_n2147);
nand_4 g06093(new_n6479, new_n6478, new_n1810);
nand_4 g06094(new_n6480_1, new_n6479, new_n1806);
nand_4 g06095(new_n6481, new_n6480_1, new_n1802);
nand_4 g06096(new_n6482, new_n6481, new_n1798);
nand_4 g06097(new_n6483, new_n6482, new_n1820);
nand_4 g06098(new_n6484, new_n6483, new_n1794);
nand_4 g06099(new_n6485, new_n6484, new_n1825);
nand_4 g06100(new_n6486, new_n6485, new_n1789);
nand_4 g06101(new_n6487, new_n6486, new_n1785);
nand_4 g06102(new_n6488, new_n6487, new_n1780);
nand_4 g06103(new_n6489, new_n6488, new_n1777);
nand_4 g06104(new_n6490, new_n6489, new_n1774);
nand_4 g06105(new_n6491, new_n6490, new_n1834);
nand_4 g06106(new_n6492, new_n6491, new_n1769);
nand_4 g06107(new_n6493, new_n6492, new_n1766);
nand_4 g06108(new_n6494, new_n6493, new_n1762);
nand_4 g06109(new_n6495, new_n6494, new_n1758);
nand_4 g06110(new_n6496, new_n6495, new_n1754);
nand_4 g06111(new_n6497, new_n6496, new_n1751);
not_3  g06112(new_n6498, new_n6497);
nor_4  g06113(new_n6499, new_n6498, new_n2290);
nor_4  g06114(new_n6500, new_n6499, new_n2289);
nor_4  g06115(new_n6501, new_n6500, new_n2288);
nor_4  g06116(new_n6502, new_n6501, new_n2287);
nor_4  g06117(new_n6503, new_n6502, new_n2286);
nor_4  g06118(new_n6504, new_n6503, new_n2285);
nor_4  g06119(new_n6505, new_n6504, new_n2284);
nor_4  g06120(new_n6506, new_n6505, new_n2283);
nor_4  g06121(new_n6507, new_n6506, new_n2145);
nor_4  g06122(new_n6508, new_n6507, new_n2144);
nor_4  g06123(new_n6509, new_n6508, new_n2143);
nor_4  g06124(new_n6510, new_n6509, new_n2142);
nor_4  g06125(new_n6511, new_n6510, new_n2141);
nor_4  g06126(new_n6512, new_n6511, new_n2140);
nor_4  g06127(new_n6513, new_n6512, new_n2139);
nor_4  g06128(new_n6514, new_n6513, new_n2138);
nor_4  g06129(new_n6515, new_n6514, new_n2137);
nor_4  g06130(new_n6516, new_n6515, new_n2136);
nor_4  g06131(new_n6517_1, new_n6516, new_n2135);
nor_4  g06132(new_n6518, new_n6517_1, new_n2134);
nor_4  g06133(new_n6519, new_n6518, new_n2133);
nor_4  g06134(new_n6520, new_n6519, new_n2132);
not_3  g06135(new_n6521, new_n6520);
nand_4 g06136(new_n6522, new_n6521, new_n1690);
nand_4 g06137(new_n6523, new_n6522, new_n1878);
nand_4 g06138(new_n6524, new_n6523, new_n1882);
nand_4 g06139(new_n6525, new_n6524, new_n1686);
nand_4 g06140(new_n6526, new_n6525, new_n1682);
nand_4 g06141(new_n6527, new_n6526, new_n1678);
nand_4 g06142(new_n6528, new_n6527, new_n1674);
nand_4 g06143(new_n6529, new_n6528, new_n1890);
nand_4 g06144(new_n6530, new_n6529, new_n1669);
nand_4 g06145(new_n6531, new_n6530, new_n1665);
nand_4 g06146(new_n6532, new_n6531, new_n1661);
nand_4 g06147(new_n6533, new_n6532, new_n1657);
nand_4 g06148(new_n6534, new_n6533, new_n1652);
nand_4 g06149(new_n6535, new_n6534, new_n1648);
nand_4 g06150(new_n6536, new_n6535, new_n1644);
nand_4 g06151(new_n6537, new_n6536, new_n1640);
nand_4 g06152(new_n6538, new_n6537, new_n1636);
nand_4 g06153(new_n6539, new_n6538, new_n1632);
nand_4 g06154(new_n6540, new_n6539, new_n1378);
nand_4 g06155(new_n6541, new_n6540, new_n1372);
nand_4 g06156(new_n6542, new_n6541, n4659);
nor_4  g06157(n5987, new_n6542, new_n1365);
nand_4 g06158(new_n6544, new_n1705, new_n1706);
nand_4 g06159(new_n6545, new_n6544, new_n1703);
nand_4 g06160(new_n6546, new_n6545, new_n1860);
nand_4 g06161(new_n6547, new_n6546, new_n1864);
nand_4 g06162(new_n6548, new_n6547, new_n1699);
nand_4 g06163(new_n6549, new_n6548, new_n1697);
nand_4 g06164(new_n6550, new_n6549, new_n1871);
nand_4 g06165(new_n6551, new_n6550, new_n1694);
nand_4 g06166(new_n6552, new_n6551, new_n1690);
nand_4 g06167(new_n6553, new_n6552, new_n1878);
nand_4 g06168(new_n6554, new_n6553, new_n1882);
nand_4 g06169(new_n6555_1, new_n6554, new_n1686);
nand_4 g06170(new_n6556, new_n6555_1, new_n1682);
nand_4 g06171(new_n6557, new_n6556, new_n1678);
nand_4 g06172(new_n6558, new_n6557, new_n1674);
nand_4 g06173(new_n6559, new_n6558, new_n1890);
nand_4 g06174(new_n6560, new_n6559, new_n1669);
nand_4 g06175(new_n6561, new_n6560, new_n1665);
nand_4 g06176(new_n6562, new_n6561, new_n1661);
nand_4 g06177(new_n6563, new_n6562, new_n1657);
nand_4 g06178(new_n6564, new_n6563, new_n1652);
nand_4 g06179(new_n6565, new_n6564, new_n1648);
nand_4 g06180(new_n6566, new_n6565, new_n1644);
nand_4 g06181(new_n6567, new_n6566, new_n1640);
nand_4 g06182(new_n6568, new_n6567, new_n1636);
nand_4 g06183(new_n6569, new_n6568, new_n1632);
nand_4 g06184(new_n6570, new_n6569, new_n1378);
nand_4 g06185(new_n6571, new_n6570, new_n1372);
nand_4 g06186(new_n6572, new_n6571, new_n1367);
nand_4 g06187(new_n6573, new_n6572, new_n1363);
nand_4 g06188(new_n6574, new_n6573, new_n1360);
nand_4 g06189(new_n6575, new_n6574, new_n1357);
nand_4 g06190(new_n6576, new_n6575, new_n1354);
nand_4 g06191(new_n6577, new_n6576, new_n1352);
nand_4 g06192(new_n6578, new_n6577, new_n1350);
nand_4 g06193(new_n6579, new_n6578, new_n1347_1);
nand_4 g06194(new_n6580, new_n6579, new_n1344);
nand_4 g06195(new_n6581, new_n6580, new_n1341);
nand_4 g06196(new_n6582, new_n6581, new_n1338);
nand_4 g06197(new_n6583, new_n6582, new_n1395);
nand_4 g06198(new_n6584, new_n6583, new_n1335);
nand_4 g06199(new_n6585, new_n6584, new_n1332);
not_3  g06200(new_n6586_1, new_n6585);
nor_4  g06201(new_n6587, new_n6586_1, new_n2413);
nor_4  g06202(new_n6588, new_n6587, new_n2412);
nor_4  g06203(new_n6589, new_n6588, new_n2411);
nor_4  g06204(new_n6590, new_n6589, new_n2410);
nor_4  g06205(new_n6591, new_n6590, new_n2409);
nor_4  g06206(new_n6592, new_n6591, new_n2408);
nor_4  g06207(new_n6593, new_n6592, new_n2407_1);
nor_4  g06208(new_n6594, new_n6593, new_n2406);
nor_4  g06209(new_n6595, new_n6594, new_n2405);
nor_4  g06210(new_n6596, new_n6595, new_n2404);
nor_4  g06211(new_n6597, new_n6596, new_n2403);
nor_4  g06212(new_n6598, new_n6597, new_n2402);
nor_4  g06213(new_n6599, new_n6598, new_n2401);
nor_4  g06214(new_n6600, new_n6599, new_n2400);
nor_4  g06215(new_n6601, new_n6600, new_n2399);
nor_4  g06216(new_n6602, new_n6601, new_n2398);
nor_4  g06217(new_n6603, new_n6602, new_n2397);
nor_4  g06218(new_n6604, new_n6603, new_n2396);
nor_4  g06219(new_n6605, new_n6604, new_n2395);
nor_4  g06220(new_n6606, new_n6605, new_n1281);
nor_4  g06221(new_n6607, new_n6606, new_n1276);
nor_4  g06222(new_n6608, new_n6607, new_n1446);
not_3  g06223(new_n6609, new_n6608);
nand_4 g06224(new_n6610, new_n6609, new_n1270);
nand_4 g06225(new_n6611, new_n6610, new_n1265_1);
nand_4 g06226(new_n6612, new_n6611, new_n1260);
nand_4 g06227(new_n6613, new_n6612, new_n1256);
nand_4 g06228(new_n6614, new_n6613, new_n1251);
nand_4 g06229(new_n6615, new_n6614, new_n1457);
nand_4 g06230(new_n6616, new_n6615, new_n1462);
nand_4 g06231(new_n6617, new_n6616, new_n1468);
nand_4 g06232(new_n6618, new_n6617, new_n1247);
nand_4 g06233(new_n6619, new_n6618, new_n1474);
nand_4 g06234(new_n6620, new_n6619, new_n592);
nand_4 g06235(new_n6621, new_n6620, new_n585);
nand_4 g06236(new_n6622, new_n6621, new_n580);
nand_4 g06237(new_n6623, new_n6622, new_n600);
nand_4 g06238(new_n6624, new_n6623, new_n606);
nand_4 g06239(new_n6625, new_n6624, new_n612);
nand_4 g06240(new_n6626, new_n6625, new_n575);
nand_4 g06241(new_n6627, new_n6626, new_n619);
nand_4 g06242(new_n6628, new_n6627, new_n570);
nand_4 g06243(new_n6629, new_n6628, new_n625);
nand_4 g06244(new_n6630, new_n6629, n5225);
nor_4  g06245(n6012, new_n6630, new_n561);
nand_4 g06246(new_n6632, new_n1303, new_n840);
nand_4 g06247(new_n6633, new_n6632, new_n1427);
nand_4 g06248(new_n6634, new_n6633, new_n1431);
nand_4 g06249(new_n6635, new_n6634, new_n1302);
nand_4 g06250(new_n6636, new_n6635, new_n1298);
nand_4 g06251(new_n6637, new_n6636, new_n1295);
nand_4 g06252(new_n6638, new_n6637, new_n1291);
nand_4 g06253(new_n6639, new_n6638, new_n1288);
nand_4 g06254(new_n6640, new_n6639, new_n1284);
nand_4 g06255(new_n6641, new_n6640, new_n1280);
nand_4 g06256(new_n6642, new_n6641, new_n1275);
nand_4 g06257(new_n6643, new_n6642, new_n1445);
nand_4 g06258(new_n6644, new_n6643, new_n1270);
nand_4 g06259(new_n6645, new_n6644, new_n1265_1);
nand_4 g06260(new_n6646, new_n6645, new_n1260);
nand_4 g06261(new_n6647, new_n6646, new_n1256);
nand_4 g06262(new_n6648, new_n6647, new_n1251);
nand_4 g06263(new_n6649, new_n6648, new_n1457);
nand_4 g06264(new_n6650, new_n6649, new_n1462);
nand_4 g06265(new_n6651, new_n6650, new_n1468);
nand_4 g06266(new_n6652, new_n6651, new_n1247);
nand_4 g06267(new_n6653, new_n6652, new_n1474);
nand_4 g06268(new_n6654, new_n6653, new_n592);
nand_4 g06269(new_n6655, new_n6654, new_n585);
nand_4 g06270(new_n6656, new_n6655, new_n580);
nand_4 g06271(new_n6657, new_n6656, new_n600);
nand_4 g06272(new_n6658, new_n6657, new_n606);
nand_4 g06273(new_n6659, new_n6658, new_n612);
nand_4 g06274(new_n6660, new_n6659, new_n575);
nand_4 g06275(new_n6661, new_n6660, new_n619);
nand_4 g06276(new_n6662, new_n6661, new_n570);
nand_4 g06277(new_n6663, new_n6662, new_n625);
nand_4 g06278(new_n6664, new_n6663, new_n564);
nand_4 g06279(new_n6665, new_n6664, new_n632);
nand_4 g06280(new_n6666, new_n6665, new_n638);
nand_4 g06281(new_n6667, new_n6666, new_n559);
nand_4 g06282(new_n6668, new_n6667, new_n554);
nand_4 g06283(new_n6669, new_n6668, new_n646);
nand_4 g06284(new_n6670, new_n6669, new_n652);
nand_4 g06285(new_n6671, new_n6670, new_n549);
nand_4 g06286(new_n6672, new_n6671, new_n544);
nand_4 g06287(new_n6673, new_n6672, new_n660);
not_3  g06288(new_n6674, new_n6673);
nor_4  g06289(new_n6675, new_n6674, new_n3068);
nor_4  g06290(new_n6676, new_n6675, new_n3067);
nor_4  g06291(new_n6677, new_n6676, new_n3066);
nor_4  g06292(new_n6678, new_n6677, new_n3065);
nor_4  g06293(new_n6679, new_n6678, new_n3064);
nor_4  g06294(new_n6680_1, new_n6679, new_n3063);
nor_4  g06295(new_n6681, new_n6680_1, new_n3062);
nor_4  g06296(new_n6682_1, new_n6681, new_n3061);
nor_4  g06297(new_n6683, new_n6682_1, new_n3354);
nor_4  g06298(new_n6684, new_n6683, new_n3353);
nor_4  g06299(new_n6685, new_n6684, new_n3352);
nor_4  g06300(new_n6686, new_n6685, new_n3351);
nor_4  g06301(new_n6687, new_n6686, new_n3350);
nor_4  g06302(new_n6688, new_n6687, new_n3349);
nor_4  g06303(new_n6689, new_n6688, new_n3348);
nor_4  g06304(new_n6690, new_n6689, new_n720);
nor_4  g06305(new_n6691, new_n6690, new_n501);
nor_4  g06306(new_n6692, new_n6691, new_n728);
nor_4  g06307(new_n6693_1, new_n6692, new_n495);
nor_4  g06308(new_n6694, new_n6693_1, new_n736);
nor_4  g06309(new_n6695, new_n6694, new_n489);
nor_4  g06310(new_n6696_1, new_n6695, new_n744);
not_3  g06311(new_n6697, new_n6696_1);
nand_4 g06312(new_n6698, new_n6697, new_n482);
nand_4 g06313(new_n6699, new_n6698, new_n751);
nand_4 g06314(new_n6700, new_n6699, new_n758);
nand_4 g06315(new_n6701, new_n6700, new_n765);
nand_4 g06316(new_n6702, new_n6701, new_n476);
nand_4 g06317(new_n6703_1, new_n6702, new_n773);
nand_4 g06318(new_n6704, new_n6703_1, new_n780);
nand_4 g06319(new_n6705, new_n6704, new_n787);
nand_4 g06320(new_n6706, new_n6705, new_n470);
nand_4 g06321(new_n6707, new_n6706, new_n795);
nand_4 g06322(new_n6708, new_n6707, new_n803);
nand_4 g06323(new_n6709, new_n6708, new_n809);
nand_4 g06324(new_n6710, new_n6709, new_n465);
nand_4 g06325(new_n6711, new_n6710, new_n818);
nand_4 g06326(new_n6712, new_n6711, new_n460);
nand_4 g06327(new_n6713, new_n6712, new_n455);
nand_4 g06328(new_n6714, new_n6713, new_n449);
nand_4 g06329(new_n6715, new_n6714, new_n827);
nand_4 g06330(new_n6716, new_n6715, new_n833);
nand_4 g06331(new_n6717, new_n6716, new_n444);
nand_4 g06332(new_n6718, new_n6717, n3673);
nor_4  g06333(n6198, new_n6718, new_n436);
nand_4 g06334(new_n6720, new_n1817, new_n1794);
nand_4 g06335(new_n6721, new_n6720, new_n1825);
nand_4 g06336(new_n6722, new_n6721, new_n1789);
nand_4 g06337(new_n6723, new_n6722, new_n1785);
nand_4 g06338(new_n6724, new_n6723, new_n1780);
nand_4 g06339(new_n6725, new_n6724, new_n1777);
nand_4 g06340(new_n6726, new_n6725, new_n1774);
nand_4 g06341(new_n6727, new_n6726, new_n1834);
nand_4 g06342(new_n6728, new_n6727, new_n1769);
nand_4 g06343(new_n6729, new_n6728, new_n1766);
nand_4 g06344(new_n6730, new_n6729, new_n1762);
nand_4 g06345(new_n6731, new_n6730, new_n1758);
nand_4 g06346(new_n6732, new_n6731, new_n1754);
nand_4 g06347(new_n6733, new_n6732, new_n1751);
nand_4 g06348(new_n6734, new_n6733, new_n1748);
nand_4 g06349(new_n6735, new_n6734, new_n1746);
nand_4 g06350(new_n6736, new_n6735, new_n1742);
nand_4 g06351(new_n6737, new_n6736, new_n1738);
nand_4 g06352(new_n6738, new_n6737, new_n1736);
nand_4 g06353(new_n6739, new_n6738, new_n1732);
nand_4 g06354(new_n6740, new_n6739, new_n1729);
nand_4 g06355(new_n6741, new_n6740, new_n1726);
nand_4 g06356(new_n6742, new_n6741, new_n1724);
nand_4 g06357(new_n6743, new_n6742, new_n1721);
nand_4 g06358(new_n6744, new_n6743, new_n1718);
nand_4 g06359(new_n6745, new_n6744, new_n1715);
nand_4 g06360(new_n6746, new_n6745, new_n1711);
nand_4 g06361(new_n6747, new_n6746, new_n1708);
nand_4 g06362(new_n6748, new_n6747, new_n1705);
nand_4 g06363(new_n6749, new_n6748, new_n1703);
nand_4 g06364(new_n6750, new_n6749, new_n1860);
nand_4 g06365(new_n6751, new_n6750, new_n1864);
nand_4 g06366(new_n6752, new_n6751, new_n1699);
nand_4 g06367(new_n6753, new_n6752, new_n1697);
nand_4 g06368(new_n6754, new_n6753, new_n1871);
nand_4 g06369(new_n6755, new_n6754, new_n1694);
nand_4 g06370(new_n6756, new_n6755, new_n1690);
nand_4 g06371(new_n6757, new_n6756, new_n1878);
nand_4 g06372(new_n6758_1, new_n6757, new_n1882);
nand_4 g06373(new_n6759, new_n6758_1, new_n1686);
nand_4 g06374(new_n6760, new_n6759, new_n1682);
nand_4 g06375(new_n6761, new_n6760, new_n1678);
nand_4 g06376(new_n6762, new_n6761, new_n1674);
nand_4 g06377(new_n6763, new_n6762, new_n1890);
nand_4 g06378(new_n6764, new_n6763, new_n1669);
nand_4 g06379(new_n6765, new_n6764, new_n1665);
not_3  g06380(new_n6766, new_n6765);
nor_4  g06381(new_n6767, new_n6766, new_n1662);
nor_4  g06382(new_n6768, new_n6767, new_n1658);
nor_4  g06383(new_n6769, new_n6768, new_n1653);
nor_4  g06384(new_n6770, new_n6769, new_n1649);
nor_4  g06385(new_n6771, new_n6770, new_n1645);
nor_4  g06386(new_n6772, new_n6771, new_n1641);
nor_4  g06387(new_n6773, new_n6772, new_n1637_1);
nor_4  g06388(new_n6774, new_n6773, new_n1633);
nor_4  g06389(new_n6775, new_n6774, new_n1629);
nor_4  g06390(new_n6776, new_n6775, new_n1628);
nor_4  g06391(new_n6777, new_n6776, new_n1627);
nor_4  g06392(new_n6778, new_n6777, new_n1626);
nor_4  g06393(new_n6779, new_n6778, new_n4700);
nor_4  g06394(new_n6780, new_n6779, new_n4699);
nor_4  g06395(new_n6781, new_n6780, new_n3722);
nor_4  g06396(new_n6782, new_n6781, new_n3721);
nor_4  g06397(new_n6783, new_n6782, new_n3720);
nor_4  g06398(new_n6784, new_n6783, new_n3719);
nor_4  g06399(new_n6785, new_n6784, new_n3718);
nor_4  g06400(new_n6786_1, new_n6785, new_n3717);
nor_4  g06401(new_n6787, new_n6786_1, new_n3716);
nor_4  g06402(new_n6788, new_n6787, new_n2611);
nor_4  g06403(new_n6789, new_n6788, new_n2610);
nor_4  g06404(new_n6790, new_n6789, new_n2609);
not_3  g06405(new_n6791_1, new_n6790);
nand_4 g06406(new_n6792, new_n6791_1, new_n1328);
nand_4 g06407(new_n6793, new_n6792, new_n1403);
nand_4 g06408(new_n6794, new_n6793, new_n1325);
nand_4 g06409(new_n6795, new_n6794, new_n1410);
nand_4 g06410(new_n6796, new_n6795, new_n1413);
nand_4 g06411(new_n6797, new_n6796, new_n1322);
nand_4 g06412(new_n6798, new_n6797, new_n1317);
nand_4 g06413(new_n6799, new_n6798, new_n1315);
nand_4 g06414(new_n6800, new_n6799, new_n1419);
nand_4 g06415(new_n6801, new_n6800, new_n1310);
nand_4 g06416(new_n6802, new_n6801, new_n1305);
nand_4 g06417(new_n6803, new_n6802, new_n1427);
nand_4 g06418(new_n6804, new_n6803, new_n1431);
nand_4 g06419(new_n6805, new_n6804, new_n1302);
nand_4 g06420(new_n6806, new_n6805, n666);
nor_4  g06421(n6275, new_n6806, new_n847);
not_3  g06422(new_n6808, new_n2188);
not_3  g06423(new_n6809, new_n2184);
nand_4 g06424(new_n6810_1, new_n6809, new_n803);
nand_4 g06425(new_n6811, new_n6810_1, new_n809);
nand_4 g06426(new_n6812, new_n6811, new_n465);
nand_4 g06427(new_n6813, new_n6812, new_n818);
nand_4 g06428(new_n6814, new_n6813, new_n460);
nand_4 g06429(new_n6815, new_n6814, new_n455);
nand_4 g06430(new_n6816, new_n6815, new_n449);
nand_4 g06431(new_n6817, new_n6816, new_n827);
nand_4 g06432(new_n6818, new_n6817, new_n833);
nand_4 g06433(new_n6819, new_n6818, new_n444);
nand_4 g06434(new_n6820, new_n6819, new_n439);
nand_4 g06435(new_n6821, new_n6820, new_n841);
nand_4 g06436(new_n6822, new_n6821, new_n434);
nand_4 g06437(new_n6823, new_n6822, new_n429);
nand_4 g06438(new_n6824, new_n6823, new_n424);
nand_4 g06439(new_n6825, new_n6824, new_n850);
nand_4 g06440(new_n6826, new_n6825, new_n856);
nand_4 g06441(new_n6827, new_n6826, new_n863);
nand_4 g06442(new_n6828, new_n6827, new_n419);
nand_4 g06443(new_n6829, new_n6828, new_n869);
nand_4 g06444(new_n6830, new_n6829, new_n875);
nand_4 g06445(new_n6831, new_n6830, new_n881);
nand_4 g06446(new_n6832, new_n6831, new_n413);
nand_4 g06447(new_n6833, new_n6832, new_n889);
nand_4 g06448(new_n6834, new_n6833, new_n896);
nand_4 g06449(new_n6835, new_n6834, new_n901);
nand_4 g06450(new_n6836, new_n6835, new_n408);
nand_4 g06451(new_n6837, new_n6836, new_n908);
nand_4 g06452(new_n6838, new_n6837, new_n403);
nand_4 g06453(new_n6839, new_n6838, new_n398);
nand_4 g06454(new_n6840, new_n6839, new_n393);
nand_4 g06455(new_n6841, new_n6840, new_n916);
nand_4 g06456(new_n6842, new_n6841, new_n1123);
nand_4 g06457(new_n6843, new_n6842, new_n1164);
nand_4 g06458(new_n6844, new_n6843, new_n1120);
nand_4 g06459(new_n6845, new_n6844, new_n1169);
nand_4 g06460(new_n6846, new_n6845, new_n1116);
nand_4 g06461(new_n6847, new_n6846, new_n1111);
nand_4 g06462(new_n6848, new_n6847, new_n1106);
nand_4 g06463(new_n6849, new_n6848, new_n1178);
nand_4 g06464(new_n6850, new_n6849, new_n1183);
nand_4 g06465(new_n6851, new_n6850, new_n1102);
nand_4 g06466(new_n6852, new_n6851, new_n1099);
nand_4 g06467(new_n6853_1, new_n6852, new_n1191);
nand_4 g06468(new_n6854, new_n6853_1, new_n1095);
nand_4 g06469(new_n6855, new_n6854, new_n1091);
nand_4 g06470(new_n6856, new_n6855, new_n1088);
nand_4 g06471(new_n6857, new_n6856, new_n1084);
nand_4 g06472(new_n6858, new_n6857, new_n1079);
nand_4 g06473(new_n6859, new_n6858, new_n1074);
nand_4 g06474(new_n6860, new_n6859, new_n1070);
not_3  g06475(new_n6861, new_n6860);
nor_4  g06476(new_n6862, new_n6861, new_n1065);
nor_4  g06477(new_n6863, new_n6862, new_n1062);
nor_4  g06478(new_n6864, new_n6863, new_n1056);
nor_4  g06479(new_n6865, new_n6864, new_n1051);
nor_4  g06480(new_n6866, new_n6865, new_n1046);
nor_4  g06481(new_n6867, new_n6866, new_n1042);
nor_4  g06482(new_n6868, new_n6867, new_n1037);
nor_4  g06483(new_n6869, new_n6868, new_n1032);
nor_4  g06484(new_n6870, new_n6869, new_n1026);
nor_4  g06485(new_n6871, new_n6870, new_n1021);
nor_4  g06486(new_n6872, new_n6871, new_n1016);
nor_4  g06487(new_n6873_1, new_n6872, new_n1011);
nor_4  g06488(new_n6874, new_n6873_1, new_n1216);
nor_4  g06489(new_n6875, new_n6874, new_n1006);
nor_4  g06490(new_n6876, new_n6875, new_n1001);
nor_4  g06491(new_n6877, new_n6876, new_n995);
nor_4  g06492(new_n6878, new_n6877, new_n990);
nor_4  g06493(new_n6879, new_n6878, new_n985);
nor_4  g06494(new_n6880, new_n6879, new_n979);
nor_4  g06495(new_n6881, new_n6880, new_n974);
nor_4  g06496(new_n6882, new_n6881, new_n968);
nor_4  g06497(new_n6883, new_n6882, new_n965);
nor_4  g06498(new_n6884, new_n6883, new_n961);
nor_4  g06499(new_n6885, new_n6884, new_n958);
nor_4  g06500(new_n6886, new_n6885, new_n953);
nor_4  g06501(new_n6887, new_n6886, new_n3536);
nor_4  g06502(new_n6888, new_n6887, new_n3535);
not_3  g06503(new_n6889, new_n6888);
nand_4 g06504(new_n6890, new_n6889, new_n938);
nand_4 g06505(new_n6891, new_n6890, new_n934);
nand_4 g06506(new_n6892, new_n6891, new_n929);
nand_4 g06507(new_n6893, new_n6892, new_n925);
nand_4 g06508(new_n6894, new_n6893, new_n2194);
nand_4 g06509(new_n6895, new_n6894, new_n2191);
nand_4 g06510(new_n6896, new_n6895, n6999);
nor_4  g06511(n6314, new_n6896, new_n6808);
nand_4 g06512(new_n6898, new_n1667, new_n686);
nand_4 g06513(new_n6899, new_n6898, new_n1665);
nand_4 g06514(new_n6900, new_n6899, new_n1661);
nand_4 g06515(new_n6901, new_n6900, new_n1657);
nand_4 g06516(new_n6902, new_n6901, new_n1652);
nand_4 g06517(new_n6903, new_n6902, new_n1648);
nand_4 g06518(new_n6904, new_n6903, new_n1644);
nand_4 g06519(new_n6905, new_n6904, new_n1640);
nand_4 g06520(new_n6906, new_n6905, new_n1636);
nand_4 g06521(new_n6907, new_n6906, new_n1632);
nand_4 g06522(new_n6908, new_n6907, new_n1378);
nand_4 g06523(new_n6909, new_n6908, new_n1372);
nand_4 g06524(new_n6910, new_n6909, new_n1367);
nand_4 g06525(new_n6911, new_n6910, new_n1363);
nand_4 g06526(new_n6912, new_n6911, new_n1360);
nand_4 g06527(new_n6913, new_n6912, new_n1357);
nand_4 g06528(new_n6914, new_n6913, new_n1354);
nand_4 g06529(new_n6915, new_n6914, new_n1352);
nand_4 g06530(new_n6916, new_n6915, new_n1350);
nand_4 g06531(new_n6917, new_n6916, new_n1347_1);
nand_4 g06532(new_n6918, new_n6917, new_n1344);
nand_4 g06533(new_n6919, new_n6918, new_n1341);
nand_4 g06534(new_n6920, new_n6919, new_n1338);
nand_4 g06535(new_n6921, new_n6920, new_n1395);
nand_4 g06536(new_n6922, new_n6921, new_n1335);
nand_4 g06537(new_n6923, new_n6922, new_n1332);
nand_4 g06538(new_n6924, new_n6923, new_n1328);
nand_4 g06539(new_n6925, new_n6924, new_n1403);
nand_4 g06540(new_n6926, new_n6925, new_n1325);
nand_4 g06541(new_n6927, new_n6926, new_n1410);
nand_4 g06542(new_n6928, new_n6927, new_n1413);
nand_4 g06543(new_n6929, new_n6928, new_n1322);
nand_4 g06544(new_n6930, new_n6929, new_n1317);
nand_4 g06545(new_n6931, new_n6930, new_n1315);
nand_4 g06546(new_n6932, new_n6931, new_n1419);
nand_4 g06547(new_n6933, new_n6932, new_n1310);
nand_4 g06548(new_n6934, new_n6933, new_n1305);
nand_4 g06549(new_n6935, new_n6934, new_n1427);
nand_4 g06550(new_n6936, new_n6935, new_n1431);
nand_4 g06551(new_n6937, new_n6936, new_n1302);
nand_4 g06552(new_n6938, new_n6937, new_n1298);
nand_4 g06553(new_n6939, new_n6938, new_n1295);
nand_4 g06554(new_n6940, new_n6939, new_n1291);
nand_4 g06555(new_n6941, new_n6940, new_n1288);
nand_4 g06556(new_n6942, new_n6941, new_n1284);
nand_4 g06557(new_n6943, new_n6942, new_n1280);
nand_4 g06558(new_n6944, new_n6943, new_n1275);
nand_4 g06559(new_n6945, new_n6944, new_n1445);
nand_4 g06560(new_n6946_1, new_n6945, new_n1270);
nand_4 g06561(new_n6947, new_n6946_1, new_n1265_1);
nand_4 g06562(new_n6948, new_n6947, new_n1260);
not_3  g06563(new_n6949, new_n6948);
nor_4  g06564(new_n6950, new_n6949, new_n1257);
nor_4  g06565(new_n6951, new_n6950, new_n1252);
nor_4  g06566(new_n6952_1, new_n6951, new_n1458);
nor_4  g06567(new_n6953, new_n6952_1, new_n1463);
nor_4  g06568(new_n6954, new_n6953, new_n1469);
nor_4  g06569(new_n6955, new_n6954, new_n1248);
nor_4  g06570(new_n6956, new_n6955, new_n1475);
nor_4  g06571(new_n6957, new_n6956, new_n1244);
nor_4  g06572(new_n6958, new_n6957, new_n1243);
nor_4  g06573(new_n6959, new_n6958, new_n1242);
nor_4  g06574(new_n6960, new_n6959, new_n1241);
nor_4  g06575(new_n6961, new_n6960, new_n1240);
nor_4  g06576(new_n6962, new_n6961, new_n1239);
nor_4  g06577(new_n6963, new_n6962, new_n3082);
nor_4  g06578(new_n6964, new_n6963, new_n3081);
nor_4  g06579(new_n6965, new_n6964, new_n3080);
nor_4  g06580(new_n6966, new_n6965, new_n3079);
nor_4  g06581(new_n6967, new_n6966, new_n3078);
nor_4  g06582(new_n6968, new_n6967, new_n3077);
nor_4  g06583(new_n6969, new_n6968, new_n3076);
nor_4  g06584(new_n6970, new_n6969, new_n3075);
nor_4  g06585(new_n6971, new_n6970, new_n3074);
nor_4  g06586(new_n6972, new_n6971, new_n3073);
nor_4  g06587(new_n6973, new_n6972, new_n3072);
nor_4  g06588(new_n6974, new_n6973, new_n3071);
nor_4  g06589(new_n6975, new_n6974, new_n3070);
nor_4  g06590(new_n6976, new_n6975, new_n3069);
not_3  g06591(new_n6977, new_n6976);
nand_4 g06592(new_n6978, new_n6977, new_n539);
nand_4 g06593(new_n6979_1, new_n6978, new_n534);
nand_4 g06594(new_n6980, new_n6979_1, new_n529);
nand_4 g06595(new_n6981, new_n6980, new_n668);
nand_4 g06596(new_n6982, new_n6981, new_n674_1);
nand_4 g06597(new_n6983, new_n6982, new_n681);
nand_4 g06598(new_n6984, new_n6983, n3506);
nor_4  g06599(n6682, new_n6984, new_n519);
nand_4 g06600(new_n6986, new_n1333, new_n794);
nand_4 g06601(new_n6987, new_n6986, new_n1332);
nand_4 g06602(new_n6988, new_n6987, new_n1328);
nand_4 g06603(new_n6989, new_n6988, new_n1403);
nand_4 g06604(new_n6990, new_n6989, new_n1325);
nand_4 g06605(new_n6991, new_n6990, new_n1410);
nand_4 g06606(new_n6992, new_n6991, new_n1413);
nand_4 g06607(new_n6993, new_n6992, new_n1322);
nand_4 g06608(new_n6994, new_n6993, new_n1317);
nand_4 g06609(new_n6995, new_n6994, new_n1315);
nand_4 g06610(new_n6996, new_n6995, new_n1419);
nand_4 g06611(new_n6997, new_n6996, new_n1310);
nand_4 g06612(new_n6998, new_n6997, new_n1305);
nand_4 g06613(new_n6999_1, new_n6998, new_n1427);
nand_4 g06614(new_n7000, new_n6999_1, new_n1431);
nand_4 g06615(new_n7001, new_n7000, new_n1302);
nand_4 g06616(new_n7002, new_n7001, new_n1298);
nand_4 g06617(new_n7003, new_n7002, new_n1295);
nand_4 g06618(new_n7004, new_n7003, new_n1291);
nand_4 g06619(new_n7005, new_n7004, new_n1288);
nand_4 g06620(new_n7006, new_n7005, new_n1284);
nand_4 g06621(new_n7007, new_n7006, new_n1280);
nand_4 g06622(new_n7008, new_n7007, new_n1275);
nand_4 g06623(new_n7009, new_n7008, new_n1445);
nand_4 g06624(new_n7010, new_n7009, new_n1270);
nand_4 g06625(new_n7011, new_n7010, new_n1265_1);
nand_4 g06626(new_n7012, new_n7011, new_n1260);
nand_4 g06627(new_n7013, new_n7012, new_n1256);
nand_4 g06628(new_n7014, new_n7013, new_n1251);
nand_4 g06629(new_n7015, new_n7014, new_n1457);
nand_4 g06630(new_n7016, new_n7015, new_n1462);
nand_4 g06631(new_n7017, new_n7016, new_n1468);
nand_4 g06632(new_n7018, new_n7017, new_n1247);
nand_4 g06633(new_n7019, new_n7018, new_n1474);
nand_4 g06634(new_n7020, new_n7019, new_n592);
nand_4 g06635(new_n7021, new_n7020, new_n585);
nand_4 g06636(new_n7022, new_n7021, new_n580);
nand_4 g06637(new_n7023, new_n7022, new_n600);
nand_4 g06638(new_n7024, new_n7023, new_n606);
nand_4 g06639(new_n7025, new_n7024, new_n612);
nand_4 g06640(new_n7026, new_n7025, new_n575);
nand_4 g06641(new_n7027, new_n7026, new_n619);
nand_4 g06642(new_n7028, new_n7027, new_n570);
nand_4 g06643(new_n7029, new_n7028, new_n625);
nand_4 g06644(new_n7030, new_n7029, new_n564);
nand_4 g06645(new_n7031, new_n7030, new_n632);
not_3  g06646(new_n7032, new_n7031);
nor_4  g06647(new_n7033, new_n7032, new_n3076);
nor_4  g06648(new_n7034, new_n7033, new_n3075);
nor_4  g06649(new_n7035, new_n7034, new_n3074);
nor_4  g06650(new_n7036, new_n7035, new_n3073);
nor_4  g06651(new_n7037, new_n7036, new_n3072);
nor_4  g06652(new_n7038, new_n7037, new_n3071);
nor_4  g06653(new_n7039, new_n7038, new_n3070);
nor_4  g06654(new_n7040, new_n7039, new_n3069);
nor_4  g06655(new_n7041, new_n7040, new_n3068);
nor_4  g06656(new_n7042, new_n7041, new_n3067);
nor_4  g06657(new_n7043, new_n7042, new_n3066);
nor_4  g06658(new_n7044, new_n7043, new_n3065);
nor_4  g06659(new_n7045, new_n7044, new_n3064);
nor_4  g06660(new_n7046, new_n7045, new_n3063);
nor_4  g06661(new_n7047, new_n7046, new_n3062);
nor_4  g06662(new_n7048, new_n7047, new_n3061);
nor_4  g06663(new_n7049, new_n7048, new_n3354);
nor_4  g06664(new_n7050, new_n7049, new_n3353);
nor_4  g06665(new_n7051, new_n7050, new_n3352);
nor_4  g06666(new_n7052, new_n7051, new_n3351);
nor_4  g06667(new_n7053, new_n7052, new_n3350);
nor_4  g06668(new_n7054, new_n7053, new_n3349);
nor_4  g06669(new_n7055, new_n7054, new_n3348);
nor_4  g06670(new_n7056, new_n7055, new_n720);
not_3  g06671(new_n7057, new_n7056);
nand_4 g06672(new_n7058, new_n7057, new_n500);
nand_4 g06673(new_n7059, new_n7058, new_n727);
nand_4 g06674(new_n7060, new_n7059, new_n494);
nand_4 g06675(new_n7061, new_n7060, new_n735);
nand_4 g06676(new_n7062, new_n7061, new_n488);
nand_4 g06677(new_n7063, new_n7062, new_n743);
nand_4 g06678(new_n7064, new_n7063, new_n482);
nand_4 g06679(new_n7065, new_n7064, new_n751);
nand_4 g06680(new_n7066, new_n7065, new_n758);
nand_4 g06681(new_n7067, new_n7066, new_n765);
nand_4 g06682(new_n7068, new_n7067, new_n476);
nand_4 g06683(new_n7069, new_n7068, new_n773);
nand_4 g06684(new_n7070, new_n7069, new_n780);
nand_4 g06685(new_n7071_1, new_n7070, new_n787);
nand_4 g06686(new_n7072, new_n7071_1, n6517);
nor_4  g06687(n6696, new_n7072, new_n467);
nand_4 g06688(new_n7074, new_n1639, new_n982);
nand_4 g06689(new_n7075, new_n7074, new_n978);
nand_4 g06690(new_n7076, new_n7075, new_n973);
nand_4 g06691(new_n7077, new_n7076, new_n967);
nand_4 g06692(new_n7078, new_n7077, new_n964);
nand_4 g06693(new_n7079, new_n7078, new_n960);
nand_4 g06694(new_n7080, new_n7079, new_n957);
nand_4 g06695(new_n7081, new_n7080, new_n952);
nand_4 g06696(new_n7082, new_n7081, new_n948_1);
nand_4 g06697(new_n7083, new_n7082, new_n943);
nand_4 g06698(new_n7084, new_n7083, new_n938);
nand_4 g06699(new_n7085, new_n7084, new_n934);
nand_4 g06700(new_n7086, new_n7085, new_n929);
nand_4 g06701(new_n7087, new_n7086, new_n925);
nand_4 g06702(new_n7088, new_n7087, new_n2194);
nand_4 g06703(new_n7089, new_n7088, new_n2191);
nand_4 g06704(new_n7090, new_n7089, new_n2190);
nand_4 g06705(new_n7091, new_n7090, new_n2186);
nand_4 g06706(new_n7092, new_n7091, new_n2183);
nand_4 g06707(new_n7093, new_n7092, new_n2179);
nand_4 g06708(new_n7094, new_n7093, new_n2175_1);
nand_4 g06709(new_n7095, new_n7094, new_n2171);
nand_4 g06710(new_n7096, new_n7095, new_n2168);
nand_4 g06711(new_n7097, new_n7096, new_n2165);
nand_4 g06712(new_n7098, new_n7097, new_n2162);
nand_4 g06713(new_n7099, new_n7098, new_n2158);
nand_4 g06714(new_n7100, new_n7099, new_n2155);
nand_4 g06715(new_n7101, new_n7100, new_n2151);
nand_4 g06716(new_n7102, new_n7101, new_n2147);
nand_4 g06717(new_n7103, new_n7102, new_n1810);
nand_4 g06718(new_n7104_1, new_n7103, new_n1806);
nand_4 g06719(new_n7105, new_n7104_1, new_n1802);
nand_4 g06720(new_n7106, new_n7105, new_n1798);
nand_4 g06721(new_n7107, new_n7106, new_n1820);
nand_4 g06722(new_n7108, new_n7107, new_n1794);
nand_4 g06723(new_n7109, new_n7108, new_n1825);
nand_4 g06724(new_n7110, new_n7109, new_n1789);
nand_4 g06725(new_n7111, new_n7110, new_n1785);
nand_4 g06726(new_n7112, new_n7111, new_n1780);
nand_4 g06727(new_n7113, new_n7112, new_n1777);
nand_4 g06728(new_n7114, new_n7113, new_n1774);
nand_4 g06729(new_n7115, new_n7114, new_n1834);
not_3  g06730(new_n7116, new_n7115);
nor_4  g06731(new_n7117, new_n7116, new_n2296);
nor_4  g06732(new_n7118, new_n7117, new_n2295);
nor_4  g06733(new_n7119, new_n7118, new_n2294);
nor_4  g06734(new_n7120, new_n7119, new_n2293);
nor_4  g06735(new_n7121, new_n7120, new_n2292);
nor_4  g06736(new_n7122, new_n7121, new_n2291);
nor_4  g06737(new_n7123, new_n7122, new_n2290);
nor_4  g06738(new_n7124, new_n7123, new_n2289);
nor_4  g06739(new_n7125, new_n7124, new_n2288);
nor_4  g06740(new_n7126, new_n7125, new_n2287);
nor_4  g06741(new_n7127, new_n7126, new_n2286);
nor_4  g06742(new_n7128, new_n7127, new_n2285);
nor_4  g06743(new_n7129, new_n7128, new_n2284);
nor_4  g06744(new_n7130, new_n7129, new_n2283);
nor_4  g06745(new_n7131, new_n7130, new_n2145);
nor_4  g06746(new_n7132_1, new_n7131, new_n2144);
nor_4  g06747(new_n7133, new_n7132_1, new_n2143);
nor_4  g06748(new_n7134, new_n7133, new_n2142);
nor_4  g06749(new_n7135, new_n7134, new_n2141);
nor_4  g06750(new_n7136, new_n7135, new_n2140);
nor_4  g06751(new_n7137, new_n7136, new_n2139);
nor_4  g06752(new_n7138, new_n7137, new_n2138);
not_3  g06753(new_n7139, new_n7138);
nand_4 g06754(new_n7140, new_n7139, new_n1860);
nand_4 g06755(new_n7141, new_n7140, new_n1864);
nand_4 g06756(new_n7142, new_n7141, new_n1699);
nand_4 g06757(new_n7143, new_n7142, new_n1697);
nand_4 g06758(new_n7144, new_n7143, new_n1871);
nand_4 g06759(new_n7145, new_n7144, new_n1694);
nand_4 g06760(new_n7146, new_n7145, new_n1690);
nand_4 g06761(new_n7147, new_n7146, new_n1878);
nand_4 g06762(new_n7148, new_n7147, new_n1882);
nand_4 g06763(new_n7149, new_n7148, new_n1686);
nand_4 g06764(new_n7150, new_n7149, new_n1682);
nand_4 g06765(new_n7151, new_n7150, new_n1678);
nand_4 g06766(new_n7152_1, new_n7151, new_n1674);
nand_4 g06767(new_n7153, new_n7152_1, new_n1890);
nand_4 g06768(new_n7154, new_n7153, new_n1669);
nand_4 g06769(new_n7155, new_n7154, new_n1665);
nand_4 g06770(new_n7156, new_n7155, new_n1661);
nand_4 g06771(new_n7157, new_n7156, new_n1657);
nand_4 g06772(new_n7158, new_n7157, new_n1652);
nand_4 g06773(new_n7159, new_n7158, new_n1648);
nand_4 g06774(new_n7160, new_n7159, n11875);
nor_4  g06775(n6786, new_n7160, new_n708);
nand_4 g06776(new_n7162, new_n2164_1, new_n447);
nand_4 g06777(new_n7163, new_n7162, new_n827);
nand_4 g06778(new_n7164, new_n7163, new_n833);
nand_4 g06779(new_n7165, new_n7164, new_n444);
nand_4 g06780(new_n7166, new_n7165, new_n439);
nand_4 g06781(new_n7167, new_n7166, new_n841);
nand_4 g06782(new_n7168, new_n7167, new_n434);
nand_4 g06783(new_n7169, new_n7168, new_n429);
nand_4 g06784(new_n7170, new_n7169, new_n424);
nand_4 g06785(new_n7171, new_n7170, new_n850);
nand_4 g06786(new_n7172, new_n7171, new_n856);
nand_4 g06787(new_n7173, new_n7172, new_n863);
nand_4 g06788(new_n7174, new_n7173, new_n419);
nand_4 g06789(new_n7175, new_n7174, new_n869);
nand_4 g06790(new_n7176, new_n7175, new_n875);
nand_4 g06791(new_n7177, new_n7176, new_n881);
nand_4 g06792(new_n7178, new_n7177, new_n413);
nand_4 g06793(new_n7179, new_n7178, new_n889);
nand_4 g06794(new_n7180, new_n7179, new_n896);
nand_4 g06795(new_n7181, new_n7180, new_n901);
nand_4 g06796(new_n7182, new_n7181, new_n408);
nand_4 g06797(new_n7183, new_n7182, new_n908);
nand_4 g06798(new_n7184, new_n7183, new_n403);
nand_4 g06799(new_n7185, new_n7184, new_n398);
nand_4 g06800(new_n7186, new_n7185, new_n393);
nand_4 g06801(new_n7187, new_n7186, new_n916);
nand_4 g06802(new_n7188, new_n7187, new_n1123);
nand_4 g06803(new_n7189, new_n7188, new_n1164);
nand_4 g06804(new_n7190, new_n7189, new_n1120);
nand_4 g06805(new_n7191, new_n7190, new_n1169);
nand_4 g06806(new_n7192, new_n7191, new_n1116);
nand_4 g06807(new_n7193, new_n7192, new_n1111);
nand_4 g06808(new_n7194, new_n7193, new_n1106);
nand_4 g06809(new_n7195, new_n7194, new_n1178);
nand_4 g06810(new_n7196, new_n7195, new_n1183);
nand_4 g06811(new_n7197, new_n7196, new_n1102);
nand_4 g06812(new_n7198, new_n7197, new_n1099);
nand_4 g06813(new_n7199, new_n7198, new_n1191);
nand_4 g06814(new_n7200, new_n7199, new_n1095);
nand_4 g06815(new_n7201, new_n7200, new_n1091);
nand_4 g06816(new_n7202, new_n7201, new_n1088);
nand_4 g06817(new_n7203, new_n7202, new_n1084);
nand_4 g06818(new_n7204, new_n7203, new_n1079);
nand_4 g06819(new_n7205, new_n7204, new_n1074);
nand_4 g06820(new_n7206, new_n7205, new_n1070);
nand_4 g06821(new_n7207, new_n7206, new_n1064);
nand_4 g06822(new_n7208, new_n7207, new_n1061);
nand_4 g06823(new_n7209, new_n7208, new_n1055);
nand_4 g06824(new_n7210, new_n7209, new_n1050);
nand_4 g06825(new_n7211, new_n7210, new_n1045);
nand_4 g06826(new_n7212, new_n7211, new_n1041);
not_3  g06827(new_n7213, new_n7212);
nor_4  g06828(new_n7214, new_n7213, new_n1037);
nor_4  g06829(new_n7215, new_n7214, new_n1032);
nor_4  g06830(new_n7216, new_n7215, new_n1026);
nor_4  g06831(new_n7217, new_n7216, new_n1021);
nor_4  g06832(new_n7218, new_n7217, new_n1016);
nor_4  g06833(new_n7219, new_n7218, new_n1011);
nor_4  g06834(new_n7220, new_n7219, new_n1216);
nor_4  g06835(new_n7221, new_n7220, new_n1006);
nor_4  g06836(new_n7222, new_n7221, new_n1001);
nor_4  g06837(new_n7223, new_n7222, new_n995);
nor_4  g06838(new_n7224, new_n7223, new_n990);
nor_4  g06839(new_n7225, new_n7224, new_n985);
nor_4  g06840(new_n7226, new_n7225, new_n979);
nor_4  g06841(new_n7227, new_n7226, new_n974);
nor_4  g06842(new_n7228, new_n7227, new_n968);
nor_4  g06843(new_n7229, new_n7228, new_n965);
nor_4  g06844(new_n7230, new_n7229, new_n961);
nor_4  g06845(new_n7231, new_n7230, new_n958);
nor_4  g06846(new_n7232, new_n7231, new_n953);
nor_4  g06847(new_n7233, new_n7232, new_n3536);
nor_4  g06848(new_n7234, new_n7233, new_n3535);
nor_4  g06849(new_n7235, new_n7234, new_n3534);
nor_4  g06850(new_n7236, new_n7235, new_n2520);
nor_4  g06851(new_n7237, new_n7236, new_n2519);
nor_4  g06852(new_n7238, new_n7237, new_n2518);
nor_4  g06853(new_n7239, new_n7238, new_n2517);
nor_4  g06854(new_n7240, new_n7239, new_n2516);
not_3  g06855(new_n7241, new_n7240);
nand_4 g06856(new_n7242, new_n7241, new_n2190);
nand_4 g06857(new_n7243, new_n7242, new_n2186);
nand_4 g06858(new_n7244, new_n7243, new_n2183);
nand_4 g06859(new_n7245, new_n7244, new_n2179);
nand_4 g06860(new_n7246_1, new_n7245, new_n2175_1);
nand_4 g06861(new_n7247, new_n7246_1, new_n2171);
nand_4 g06862(new_n7248, new_n7247, n11345);
nor_4  g06863(n6853, new_n7248, new_n1407);
nand_4 g06864(new_n7250, new_n1711, new_n1712);
nand_4 g06865(new_n7251, new_n7250, new_n1708);
nand_4 g06866(new_n7252, new_n7251, new_n1705);
nand_4 g06867(new_n7253, new_n7252, new_n1703);
nand_4 g06868(new_n7254, new_n7253, new_n1860);
nand_4 g06869(new_n7255, new_n7254, new_n1864);
nand_4 g06870(new_n7256, new_n7255, new_n1699);
nand_4 g06871(new_n7257, new_n7256, new_n1697);
nand_4 g06872(new_n7258, new_n7257, new_n1871);
nand_4 g06873(new_n7259, new_n7258, new_n1694);
nand_4 g06874(new_n7260, new_n7259, new_n1690);
nand_4 g06875(new_n7261, new_n7260, new_n1878);
nand_4 g06876(new_n7262, new_n7261, new_n1882);
nand_4 g06877(new_n7263, new_n7262, new_n1686);
nand_4 g06878(new_n7264, new_n7263, new_n1682);
nand_4 g06879(new_n7265_1, new_n7264, new_n1678);
nand_4 g06880(new_n7266, new_n7265_1, new_n1674);
nand_4 g06881(new_n7267, new_n7266, new_n1890);
nand_4 g06882(new_n7268, new_n7267, new_n1669);
nand_4 g06883(new_n7269, new_n7268, new_n1665);
nand_4 g06884(new_n7270, new_n7269, new_n1661);
nand_4 g06885(new_n7271, new_n7270, new_n1657);
nand_4 g06886(new_n7272_1, new_n7271, new_n1652);
nand_4 g06887(new_n7273, new_n7272_1, new_n1648);
nand_4 g06888(new_n7274, new_n7273, new_n1644);
nand_4 g06889(new_n7275, new_n7274, new_n1640);
nand_4 g06890(new_n7276, new_n7275, new_n1636);
nand_4 g06891(new_n7277, new_n7276, new_n1632);
nand_4 g06892(new_n7278, new_n7277, new_n1378);
nand_4 g06893(new_n7279, new_n7278, new_n1372);
nand_4 g06894(new_n7280, new_n7279, new_n1367);
nand_4 g06895(new_n7281, new_n7280, new_n1363);
nand_4 g06896(new_n7282_1, new_n7281, new_n1360);
nand_4 g06897(new_n7283, new_n7282_1, new_n1357);
nand_4 g06898(new_n7284, new_n7283, new_n1354);
nand_4 g06899(new_n7285, new_n7284, new_n1352);
nand_4 g06900(new_n7286, new_n7285, new_n1350);
nand_4 g06901(new_n7287, new_n7286, new_n1347_1);
nand_4 g06902(new_n7288, new_n7287, new_n1344);
nand_4 g06903(new_n7289, new_n7288, new_n1341);
nand_4 g06904(new_n7290, new_n7289, new_n1338);
nand_4 g06905(new_n7291, new_n7290, new_n1395);
nand_4 g06906(new_n7292, new_n7291, new_n1335);
nand_4 g06907(new_n7293, new_n7292, new_n1332);
nand_4 g06908(new_n7294, new_n7293, new_n1328);
nand_4 g06909(new_n7295, new_n7294, new_n1403);
not_3  g06910(new_n7296, new_n7295);
nor_4  g06911(new_n7297, new_n7296, new_n2411);
nor_4  g06912(new_n7298, new_n7297, new_n2410);
nor_4  g06913(new_n7299, new_n7298, new_n2409);
nor_4  g06914(new_n7300, new_n7299, new_n2408);
nor_4  g06915(new_n7301, new_n7300, new_n2407_1);
nor_4  g06916(new_n7302, new_n7301, new_n2406);
nor_4  g06917(new_n7303, new_n7302, new_n2405);
nor_4  g06918(new_n7304, new_n7303, new_n2404);
nor_4  g06919(new_n7305, new_n7304, new_n2403);
nor_4  g06920(new_n7306, new_n7305, new_n2402);
nor_4  g06921(new_n7307, new_n7306, new_n2401);
nor_4  g06922(new_n7308, new_n7307, new_n2400);
nor_4  g06923(new_n7309, new_n7308, new_n2399);
nor_4  g06924(new_n7310, new_n7309, new_n2398);
nor_4  g06925(new_n7311, new_n7310, new_n2397);
nor_4  g06926(new_n7312, new_n7311, new_n2396);
nor_4  g06927(new_n7313, new_n7312, new_n2395);
nor_4  g06928(new_n7314, new_n7313, new_n1281);
nor_4  g06929(new_n7315, new_n7314, new_n1276);
nor_4  g06930(new_n7316, new_n7315, new_n1446);
nor_4  g06931(new_n7317, new_n7316, new_n1271);
nor_4  g06932(new_n7318, new_n7317, new_n1266);
nor_4  g06933(new_n7319, new_n7318, new_n1261);
nor_4  g06934(new_n7320, new_n7319, new_n1257);
not_3  g06935(new_n7321, new_n7320);
nand_4 g06936(new_n7322, new_n7321, new_n1251);
nand_4 g06937(new_n7323, new_n7322, new_n1457);
nand_4 g06938(new_n7324, new_n7323, new_n1462);
nand_4 g06939(new_n7325, new_n7324, new_n1468);
nand_4 g06940(new_n7326, new_n7325, new_n1247);
nand_4 g06941(new_n7327, new_n7326, new_n1474);
nand_4 g06942(new_n7328, new_n7327, new_n592);
nand_4 g06943(new_n7329, new_n7328, new_n585);
nand_4 g06944(new_n7330, new_n7329, new_n580);
nand_4 g06945(new_n7331, new_n7330, new_n600);
nand_4 g06946(new_n7332, new_n7331, new_n606);
nand_4 g06947(new_n7333, new_n7332, new_n612);
nand_4 g06948(new_n7334, new_n7333, new_n575);
nand_4 g06949(new_n7335, new_n7334, new_n619);
nand_4 g06950(new_n7336, new_n7335, n13109);
nor_4  g06951(n6952, new_n7336, new_n566);
nand_4 g06952(new_n7338, new_n997, new_n994);
nand_4 g06953(new_n7339, new_n7338, new_n989);
nand_4 g06954(new_n7340, new_n7339, new_n984);
nand_4 g06955(new_n7341, new_n7340, new_n978);
nand_4 g06956(new_n7342, new_n7341, new_n973);
nand_4 g06957(new_n7343, new_n7342, new_n967);
nand_4 g06958(new_n7344, new_n7343, new_n964);
nand_4 g06959(new_n7345, new_n7344, new_n960);
nand_4 g06960(new_n7346, new_n7345, new_n957);
nand_4 g06961(new_n7347, new_n7346, new_n952);
nand_4 g06962(new_n7348, new_n7347, new_n948_1);
nand_4 g06963(new_n7349, new_n7348, new_n943);
nand_4 g06964(new_n7350, new_n7349, new_n938);
nand_4 g06965(new_n7351, new_n7350, new_n934);
nand_4 g06966(new_n7352, new_n7351, new_n929);
nand_4 g06967(new_n7353, new_n7352, new_n925);
nand_4 g06968(new_n7354_1, new_n7353, new_n2194);
nand_4 g06969(new_n7355, new_n7354_1, new_n2191);
nand_4 g06970(new_n7356, new_n7355, new_n2190);
nand_4 g06971(new_n7357, new_n7356, new_n2186);
nand_4 g06972(new_n7358, new_n7357, new_n2183);
nand_4 g06973(new_n7359, new_n7358, new_n2179);
nand_4 g06974(new_n7360, new_n7359, new_n2175_1);
nand_4 g06975(new_n7361, new_n7360, new_n2171);
nand_4 g06976(new_n7362, new_n7361, new_n2168);
nand_4 g06977(new_n7363, new_n7362, new_n2165);
nand_4 g06978(new_n7364, new_n7363, new_n2162);
nand_4 g06979(new_n7365, new_n7364, new_n2158);
nand_4 g06980(new_n7366, new_n7365, new_n2155);
nand_4 g06981(new_n7367, new_n7366, new_n2151);
nand_4 g06982(new_n7368, new_n7367, new_n2147);
nand_4 g06983(new_n7369, new_n7368, new_n1810);
nand_4 g06984(new_n7370, new_n7369, new_n1806);
nand_4 g06985(new_n7371, new_n7370, new_n1802);
nand_4 g06986(new_n7372, new_n7371, new_n1798);
nand_4 g06987(new_n7373, new_n7372, new_n1820);
nand_4 g06988(new_n7374, new_n7373, new_n1794);
nand_4 g06989(new_n7375, new_n7374, new_n1825);
nand_4 g06990(new_n7376, new_n7375, new_n1789);
nand_4 g06991(new_n7377, new_n7376, new_n1785);
nand_4 g06992(new_n7378, new_n7377, new_n1780);
nand_4 g06993(new_n7379, new_n7378, new_n1777);
not_3  g06994(new_n7380, new_n7379);
nor_4  g06995(new_n7381, new_n7380, new_n2298);
nor_4  g06996(new_n7382_1, new_n7381, new_n2297);
nor_4  g06997(new_n7383, new_n7382_1, new_n2296);
nor_4  g06998(new_n7384, new_n7383, new_n2295);
nor_4  g06999(new_n7385, new_n7384, new_n2294);
nor_4  g07000(new_n7386, new_n7385, new_n2293);
nor_4  g07001(new_n7387, new_n7386, new_n2292);
nor_4  g07002(new_n7388, new_n7387, new_n2291);
nor_4  g07003(new_n7389, new_n7388, new_n2290);
nor_4  g07004(new_n7390, new_n7389, new_n2289);
nor_4  g07005(new_n7391, new_n7390, new_n2288);
nor_4  g07006(new_n7392, new_n7391, new_n2287);
nor_4  g07007(new_n7393, new_n7392, new_n2286);
nor_4  g07008(new_n7394, new_n7393, new_n2285);
nor_4  g07009(new_n7395, new_n7394, new_n2284);
nor_4  g07010(new_n7396, new_n7395, new_n2283);
nor_4  g07011(new_n7397, new_n7396, new_n2145);
nor_4  g07012(new_n7398, new_n7397, new_n2144);
nor_4  g07013(new_n7399, new_n7398, new_n2143);
nor_4  g07014(new_n7400, new_n7399, new_n2142);
nor_4  g07015(new_n7401, new_n7400, new_n2141);
nor_4  g07016(new_n7402, new_n7401, new_n2140);
not_3  g07017(new_n7403, new_n7402);
nand_4 g07018(new_n7404, new_n7403, new_n1705);
nand_4 g07019(new_n7405, new_n7404, new_n1703);
nand_4 g07020(new_n7406, new_n7405, new_n1860);
nand_4 g07021(new_n7407, new_n7406, new_n1864);
nand_4 g07022(new_n7408, new_n7407, new_n1699);
nand_4 g07023(new_n7409, new_n7408, new_n1697);
nand_4 g07024(new_n7410, new_n7409, new_n1871);
nand_4 g07025(new_n7411, new_n7410, new_n1694);
nand_4 g07026(new_n7412, new_n7411, new_n1690);
nand_4 g07027(new_n7413, new_n7412, new_n1878);
nand_4 g07028(new_n7414, new_n7413, new_n1882);
nand_4 g07029(new_n7415, new_n7414, new_n1686);
nand_4 g07030(new_n7416, new_n7415, new_n1682);
nand_4 g07031(new_n7417, new_n7416, new_n1678);
nand_4 g07032(new_n7418, new_n7417, new_n1674);
nand_4 g07033(new_n7419, new_n7418, new_n1890);
nand_4 g07034(new_n7420, new_n7419, new_n1669);
nand_4 g07035(new_n7421, new_n7420, new_n1665);
nand_4 g07036(new_n7422, new_n7421, new_n1661);
nand_4 g07037(new_n7423, new_n7422, new_n1657);
nand_4 g07038(new_n7424, new_n7423, n8635);
nor_4  g07039(n6979, new_n7424, new_n702_1);
nand_4 g07040(new_n7426, new_n1804, new_n1426);
nand_4 g07041(new_n7427, new_n7426, new_n1802);
nand_4 g07042(new_n7428, new_n7427, new_n1798);
nand_4 g07043(new_n7429, new_n7428, new_n1820);
nand_4 g07044(new_n7430, new_n7429, new_n1794);
nand_4 g07045(new_n7431, new_n7430, new_n1825);
nand_4 g07046(new_n7432, new_n7431, new_n1789);
nand_4 g07047(new_n7433, new_n7432, new_n1785);
nand_4 g07048(new_n7434, new_n7433, new_n1780);
nand_4 g07049(new_n7435, new_n7434, new_n1777);
nand_4 g07050(new_n7436, new_n7435, new_n1774);
nand_4 g07051(new_n7437, new_n7436, new_n1834);
nand_4 g07052(new_n7438, new_n7437, new_n1769);
nand_4 g07053(new_n7439, new_n7438, new_n1766);
nand_4 g07054(new_n7440, new_n7439, new_n1762);
nand_4 g07055(new_n7441, new_n7440, new_n1758);
nand_4 g07056(new_n7442, new_n7441, new_n1754);
nand_4 g07057(new_n7443, new_n7442, new_n1751);
nand_4 g07058(new_n7444, new_n7443, new_n1748);
nand_4 g07059(new_n7445, new_n7444, new_n1746);
nand_4 g07060(new_n7446, new_n7445, new_n1742);
nand_4 g07061(new_n7447, new_n7446, new_n1738);
nand_4 g07062(new_n7448, new_n7447, new_n1736);
nand_4 g07063(new_n7449, new_n7448, new_n1732);
nand_4 g07064(new_n7450_1, new_n7449, new_n1729);
nand_4 g07065(new_n7451, new_n7450_1, new_n1726);
nand_4 g07066(new_n7452, new_n7451, new_n1724);
nand_4 g07067(new_n7453, new_n7452, new_n1721);
nand_4 g07068(new_n7454, new_n7453, new_n1718);
nand_4 g07069(new_n7455, new_n7454, new_n1715);
nand_4 g07070(new_n7456, new_n7455, new_n1711);
nand_4 g07071(new_n7457, new_n7456, new_n1708);
nand_4 g07072(new_n7458, new_n7457, new_n1705);
nand_4 g07073(new_n7459, new_n7458, new_n1703);
nand_4 g07074(new_n7460, new_n7459, new_n1860);
nand_4 g07075(new_n7461, new_n7460, new_n1864);
nand_4 g07076(new_n7462, new_n7461, new_n1699);
nand_4 g07077(new_n7463, new_n7462, new_n1697);
nand_4 g07078(new_n7464, new_n7463, new_n1871);
nand_4 g07079(new_n7465, new_n7464, new_n1694);
nand_4 g07080(new_n7466, new_n7465, new_n1690);
nand_4 g07081(new_n7467, new_n7466, new_n1878);
nand_4 g07082(new_n7468, new_n7467, new_n1882);
nand_4 g07083(new_n7469, new_n7468, new_n1686);
nand_4 g07084(new_n7470, new_n7469, new_n1682);
nand_4 g07085(new_n7471, new_n7470, new_n1678);
nand_4 g07086(new_n7472, new_n7471, new_n1674);
nand_4 g07087(new_n7473, new_n7472, new_n1890);
nand_4 g07088(new_n7474, new_n7473, new_n1669);
nand_4 g07089(new_n7475, new_n7474, new_n1665);
not_3  g07090(new_n7476, new_n7475);
nor_4  g07091(new_n7477, new_n7476, new_n1662);
nor_4  g07092(new_n7478, new_n7477, new_n1658);
nor_4  g07093(new_n7479, new_n7478, new_n1653);
nor_4  g07094(new_n7480, new_n7479, new_n1649);
nor_4  g07095(new_n7481, new_n7480, new_n1645);
nor_4  g07096(new_n7482, new_n7481, new_n1641);
nor_4  g07097(new_n7483, new_n7482, new_n1637_1);
nor_4  g07098(new_n7484, new_n7483, new_n1633);
nor_4  g07099(new_n7485, new_n7484, new_n1629);
nor_4  g07100(new_n7486, new_n7485, new_n1628);
nor_4  g07101(new_n7487, new_n7486, new_n1627);
nor_4  g07102(new_n7488, new_n7487, new_n1626);
nor_4  g07103(new_n7489, new_n7488, new_n4700);
nor_4  g07104(new_n7490, new_n7489, new_n4699);
nor_4  g07105(new_n7491, new_n7490, new_n3722);
nor_4  g07106(new_n7492, new_n7491, new_n3721);
nor_4  g07107(new_n7493, new_n7492, new_n3720);
nor_4  g07108(new_n7494, new_n7493, new_n3719);
nor_4  g07109(new_n7495, new_n7494, new_n3718);
nor_4  g07110(new_n7496, new_n7495, new_n3717);
nor_4  g07111(new_n7497, new_n7496, new_n3716);
nor_4  g07112(new_n7498, new_n7497, new_n2611);
nor_4  g07113(new_n7499, new_n7498, new_n2610);
nor_4  g07114(new_n7500, new_n7499, new_n2609);
nor_4  g07115(new_n7501, new_n7500, new_n2413);
not_3  g07116(new_n7502, new_n7501);
nand_4 g07117(new_n7503, new_n7502, new_n1403);
nand_4 g07118(new_n7504, new_n7503, new_n1325);
nand_4 g07119(new_n7505, new_n7504, new_n1410);
nand_4 g07120(new_n7506, new_n7505, new_n1413);
nand_4 g07121(new_n7507, new_n7506, new_n1322);
nand_4 g07122(new_n7508, new_n7507, new_n1317);
nand_4 g07123(new_n7509, new_n7508, new_n1315);
nand_4 g07124(new_n7510, new_n7509, new_n1419);
nand_4 g07125(new_n7511, new_n7510, new_n1310);
nand_4 g07126(new_n7512, new_n7511, n14408);
nor_4  g07127(n7071, new_n7512, new_n838);
nand_4 g07128(new_n7514, new_n1809, new_n432);
nand_4 g07129(new_n7515, new_n7514, new_n429);
nand_4 g07130(new_n7516, new_n7515, new_n424);
nand_4 g07131(new_n7517, new_n7516, new_n850);
nand_4 g07132(new_n7518, new_n7517, new_n856);
nand_4 g07133(new_n7519, new_n7518, new_n863);
nand_4 g07134(new_n7520, new_n7519, new_n419);
nand_4 g07135(new_n7521, new_n7520, new_n869);
nand_4 g07136(new_n7522, new_n7521, new_n875);
nand_4 g07137(new_n7523, new_n7522, new_n881);
nand_4 g07138(new_n7524, new_n7523, new_n413);
nand_4 g07139(new_n7525, new_n7524, new_n889);
nand_4 g07140(new_n7526, new_n7525, new_n896);
nand_4 g07141(new_n7527, new_n7526, new_n901);
nand_4 g07142(new_n7528, new_n7527, new_n408);
nand_4 g07143(new_n7529, new_n7528, new_n908);
nand_4 g07144(new_n7530, new_n7529, new_n403);
nand_4 g07145(new_n7531, new_n7530, new_n398);
nand_4 g07146(new_n7532, new_n7531, new_n393);
nand_4 g07147(new_n7533, new_n7532, new_n916);
nand_4 g07148(new_n7534, new_n7533, new_n1123);
nand_4 g07149(new_n7535, new_n7534, new_n1164);
nand_4 g07150(new_n7536, new_n7535, new_n1120);
nand_4 g07151(new_n7537, new_n7536, new_n1169);
nand_4 g07152(new_n7538, new_n7537, new_n1116);
nand_4 g07153(new_n7539, new_n7538, new_n1111);
nand_4 g07154(new_n7540, new_n7539, new_n1106);
nand_4 g07155(new_n7541, new_n7540, new_n1178);
nand_4 g07156(new_n7542, new_n7541, new_n1183);
nand_4 g07157(new_n7543, new_n7542, new_n1102);
nand_4 g07158(new_n7544, new_n7543, new_n1099);
nand_4 g07159(new_n7545, new_n7544, new_n1191);
nand_4 g07160(new_n7546, new_n7545, new_n1095);
nand_4 g07161(new_n7547, new_n7546, new_n1091);
nand_4 g07162(new_n7548, new_n7547, new_n1088);
nand_4 g07163(new_n7549, new_n7548, new_n1084);
nand_4 g07164(new_n7550, new_n7549, new_n1079);
nand_4 g07165(new_n7551, new_n7550, new_n1074);
nand_4 g07166(new_n7552, new_n7551, new_n1070);
nand_4 g07167(new_n7553, new_n7552, new_n1064);
nand_4 g07168(new_n7554, new_n7553, new_n1061);
nand_4 g07169(new_n7555, new_n7554, new_n1055);
nand_4 g07170(new_n7556, new_n7555, new_n1050);
nand_4 g07171(new_n7557, new_n7556, new_n1045);
nand_4 g07172(new_n7558, new_n7557, new_n1041);
not_3  g07173(new_n7559, new_n7558);
nor_4  g07174(new_n7560, new_n7559, new_n1037);
nor_4  g07175(new_n7561, new_n7560, new_n1032);
nor_4  g07176(new_n7562, new_n7561, new_n1026);
nor_4  g07177(new_n7563, new_n7562, new_n1021);
nor_4  g07178(new_n7564, new_n7563, new_n1016);
nor_4  g07179(new_n7565, new_n7564, new_n1011);
nor_4  g07180(new_n7566, new_n7565, new_n1216);
nor_4  g07181(new_n7567, new_n7566, new_n1006);
nor_4  g07182(new_n7568, new_n7567, new_n1001);
nor_4  g07183(new_n7569, new_n7568, new_n995);
nor_4  g07184(new_n7570, new_n7569, new_n990);
nor_4  g07185(new_n7571, new_n7570, new_n985);
nor_4  g07186(new_n7572, new_n7571, new_n979);
nor_4  g07187(new_n7573, new_n7572, new_n974);
nor_4  g07188(new_n7574, new_n7573, new_n968);
nor_4  g07189(new_n7575, new_n7574, new_n965);
nor_4  g07190(new_n7576, new_n7575, new_n961);
nor_4  g07191(new_n7577, new_n7576, new_n958);
nor_4  g07192(new_n7578, new_n7577, new_n953);
nor_4  g07193(new_n7579, new_n7578, new_n3536);
nor_4  g07194(new_n7580, new_n7579, new_n3535);
nor_4  g07195(new_n7581, new_n7580, new_n3534);
nor_4  g07196(new_n7582, new_n7581, new_n2520);
nor_4  g07197(new_n7583, new_n7582, new_n2519);
not_3  g07198(new_n7584, new_n7583);
nand_4 g07199(new_n7585, new_n7584, new_n925);
nand_4 g07200(new_n7586, new_n7585, new_n2194);
nand_4 g07201(new_n7587, new_n7586, new_n2191);
nand_4 g07202(new_n7588, new_n7587, new_n2190);
nand_4 g07203(new_n7589, new_n7588, new_n2186);
nand_4 g07204(new_n7590, new_n7589, new_n2183);
nand_4 g07205(new_n7591, new_n7590, new_n2179);
nand_4 g07206(new_n7592, new_n7591, new_n2175_1);
nand_4 g07207(new_n7593, new_n7592, new_n2171);
nand_4 g07208(new_n7594, new_n7593, new_n2168);
nand_4 g07209(new_n7595, new_n7594, new_n2165);
nand_4 g07210(new_n7596, new_n7595, new_n2162);
nand_4 g07211(new_n7597, new_n7596, new_n2158);
nand_4 g07212(new_n7598, new_n7597, new_n2155);
nand_4 g07213(new_n7599, new_n7598, new_n2151);
nand_4 g07214(new_n7600, new_n7599, n5023);
nor_4  g07215(n7073, new_n7600, new_n1307);
not_3  g07216(new_n7602, new_n1376);
nand_4 g07217(new_n7603, new_n733, new_n1370);
nand_4 g07218(new_n7604, new_n7603, new_n964);
nand_4 g07219(new_n7605, new_n7604, new_n960);
nand_4 g07220(new_n7606, new_n7605, new_n957);
nand_4 g07221(new_n7607, new_n7606, new_n952);
nand_4 g07222(new_n7608, new_n7607, new_n948_1);
nand_4 g07223(new_n7609, new_n7608, new_n943);
nand_4 g07224(new_n7610, new_n7609, new_n938);
nand_4 g07225(new_n7611, new_n7610, new_n934);
nand_4 g07226(new_n7612, new_n7611, new_n929);
nand_4 g07227(new_n7613, new_n7612, new_n925);
nand_4 g07228(new_n7614, new_n7613, new_n2194);
nand_4 g07229(new_n7615, new_n7614, new_n2191);
nand_4 g07230(new_n7616, new_n7615, new_n2190);
nand_4 g07231(new_n7617, new_n7616, new_n2186);
nand_4 g07232(new_n7618, new_n7617, new_n2183);
nand_4 g07233(new_n7619, new_n7618, new_n2179);
nand_4 g07234(new_n7620, new_n7619, new_n2175_1);
nand_4 g07235(new_n7621, new_n7620, new_n2171);
nand_4 g07236(new_n7622, new_n7621, new_n2168);
nand_4 g07237(new_n7623, new_n7622, new_n2165);
nand_4 g07238(new_n7624, new_n7623, new_n2162);
nand_4 g07239(new_n7625, new_n7624, new_n2158);
nand_4 g07240(new_n7626, new_n7625, new_n2155);
nand_4 g07241(new_n7627, new_n7626, new_n2151);
nand_4 g07242(new_n7628, new_n7627, new_n2147);
nand_4 g07243(new_n7629, new_n7628, new_n1810);
nand_4 g07244(new_n7630, new_n7629, new_n1806);
nand_4 g07245(new_n7631, new_n7630, new_n1802);
nand_4 g07246(new_n7632, new_n7631, new_n1798);
nand_4 g07247(new_n7633, new_n7632, new_n1820);
nand_4 g07248(new_n7634, new_n7633, new_n1794);
nand_4 g07249(new_n7635, new_n7634, new_n1825);
nand_4 g07250(new_n7636, new_n7635, new_n1789);
nand_4 g07251(new_n7637, new_n7636, new_n1785);
nand_4 g07252(new_n7638, new_n7637, new_n1780);
not_3  g07253(new_n7639, new_n7638);
nor_4  g07254(new_n7640, new_n7639, new_n2299);
nor_4  g07255(new_n7641, new_n7640, new_n2298);
nor_4  g07256(new_n7642, new_n7641, new_n2297);
nor_4  g07257(new_n7643, new_n7642, new_n2296);
nor_4  g07258(new_n7644, new_n7643, new_n2295);
nor_4  g07259(new_n7645, new_n7644, new_n2294);
nor_4  g07260(new_n7646, new_n7645, new_n2293);
nor_4  g07261(new_n7647, new_n7646, new_n2292);
nor_4  g07262(new_n7648, new_n7647, new_n2291);
nor_4  g07263(new_n7649, new_n7648, new_n2290);
nor_4  g07264(new_n7650, new_n7649, new_n2289);
nor_4  g07265(new_n7651, new_n7650, new_n2288);
nor_4  g07266(new_n7652_1, new_n7651, new_n2287);
nor_4  g07267(new_n7653, new_n7652_1, new_n2286);
nor_4  g07268(new_n7654, new_n7653, new_n2285);
nor_4  g07269(new_n7655_1, new_n7654, new_n2284);
nor_4  g07270(new_n7656, new_n7655_1, new_n2283);
nor_4  g07271(new_n7657, new_n7656, new_n2145);
nor_4  g07272(new_n7658, new_n7657, new_n2144);
not_3  g07273(new_n7659, new_n7658);
nand_4 g07274(new_n7660, new_n7659, new_n1718);
nand_4 g07275(new_n7661, new_n7660, new_n1715);
nand_4 g07276(new_n7662, new_n7661, new_n1711);
nand_4 g07277(new_n7663, new_n7662, new_n1708);
nand_4 g07278(new_n7664, new_n7663, new_n1705);
nand_4 g07279(new_n7665, new_n7664, new_n1703);
nand_4 g07280(new_n7666, new_n7665, new_n1860);
nand_4 g07281(new_n7667_1, new_n7666, new_n1864);
nand_4 g07282(new_n7668, new_n7667_1, new_n1699);
nand_4 g07283(new_n7669, new_n7668, new_n1697);
nand_4 g07284(new_n7670, new_n7669, new_n1871);
nand_4 g07285(new_n7671, new_n7670, new_n1694);
nand_4 g07286(new_n7672, new_n7671, new_n1690);
nand_4 g07287(new_n7673, new_n7672, new_n1878);
nand_4 g07288(new_n7674, new_n7673, new_n1882);
nand_4 g07289(new_n7675, new_n7674, new_n1686);
nand_4 g07290(new_n7676, new_n7675, new_n1682);
nand_4 g07291(new_n7677, new_n7676, new_n1678);
nand_4 g07292(new_n7678, new_n7677, new_n1674);
nand_4 g07293(new_n7679, new_n7678, new_n1890);
nand_4 g07294(new_n7680, new_n7679, new_n1669);
nand_4 g07295(new_n7681, new_n7680, new_n1665);
nand_4 g07296(new_n7682, new_n7681, new_n1661);
nand_4 g07297(new_n7683, new_n7682, new_n1657);
nand_4 g07298(new_n7684, new_n7683, new_n1652);
nand_4 g07299(new_n7685, new_n7684, new_n1648);
nand_4 g07300(new_n7686, new_n7685, new_n1644);
nand_4 g07301(new_n7687, new_n7686, new_n1640);
nand_4 g07302(new_n7688, new_n7687, new_n1636);
nand_4 g07303(new_n7689, new_n7688, new_n1632);
nand_4 g07304(new_n7690, new_n7689, n11590);
nor_4  g07305(n7132, new_n7690, new_n7602);
nand_4 g07306(new_n7692, new_n1348, new_n764);
nand_4 g07307(new_n7693, new_n7692, new_n1347_1);
nand_4 g07308(new_n7694, new_n7693, new_n1344);
nand_4 g07309(new_n7695, new_n7694, new_n1341);
nand_4 g07310(new_n7696, new_n7695, new_n1338);
nand_4 g07311(new_n7697, new_n7696, new_n1395);
nand_4 g07312(new_n7698, new_n7697, new_n1335);
nand_4 g07313(new_n7699, new_n7698, new_n1332);
nand_4 g07314(new_n7700, new_n7699, new_n1328);
nand_4 g07315(new_n7701, new_n7700, new_n1403);
nand_4 g07316(new_n7702, new_n7701, new_n1325);
nand_4 g07317(new_n7703, new_n7702, new_n1410);
nand_4 g07318(new_n7704, new_n7703, new_n1413);
nand_4 g07319(new_n7705, new_n7704, new_n1322);
nand_4 g07320(new_n7706, new_n7705, new_n1317);
nand_4 g07321(new_n7707, new_n7706, new_n1315);
nand_4 g07322(new_n7708, new_n7707, new_n1419);
nand_4 g07323(new_n7709, new_n7708, new_n1310);
nand_4 g07324(new_n7710, new_n7709, new_n1305);
nand_4 g07325(new_n7711, new_n7710, new_n1427);
nand_4 g07326(new_n7712, new_n7711, new_n1431);
nand_4 g07327(new_n7713, new_n7712, new_n1302);
nand_4 g07328(new_n7714, new_n7713, new_n1298);
nand_4 g07329(new_n7715, new_n7714, new_n1295);
nand_4 g07330(new_n7716, new_n7715, new_n1291);
nand_4 g07331(new_n7717, new_n7716, new_n1288);
nand_4 g07332(new_n7718, new_n7717, new_n1284);
nand_4 g07333(new_n7719, new_n7718, new_n1280);
nand_4 g07334(new_n7720, new_n7719, new_n1275);
nand_4 g07335(new_n7721, new_n7720, new_n1445);
nand_4 g07336(new_n7722, new_n7721, new_n1270);
nand_4 g07337(new_n7723, new_n7722, new_n1265_1);
nand_4 g07338(new_n7724, new_n7723, new_n1260);
nand_4 g07339(new_n7725, new_n7724, new_n1256);
nand_4 g07340(new_n7726, new_n7725, new_n1251);
nand_4 g07341(new_n7727, new_n7726, new_n1457);
nand_4 g07342(new_n7728, new_n7727, new_n1462);
nand_4 g07343(new_n7729, new_n7728, new_n1468);
nand_4 g07344(new_n7730, new_n7729, new_n1247);
nand_4 g07345(new_n7731, new_n7730, new_n1474);
nand_4 g07346(new_n7732, new_n7731, new_n592);
nand_4 g07347(new_n7733, new_n7732, new_n585);
nand_4 g07348(new_n7734, new_n7733, new_n580);
nand_4 g07349(new_n7735, new_n7734, new_n600);
nand_4 g07350(new_n7736, new_n7735, new_n606);
nand_4 g07351(new_n7737, new_n7736, new_n612);
not_3  g07352(new_n7738, new_n7737);
nor_4  g07353(new_n7739, new_n7738, new_n3082);
nor_4  g07354(new_n7740, new_n7739, new_n3081);
nor_4  g07355(new_n7741, new_n7740, new_n3080);
nor_4  g07356(new_n7742, new_n7741, new_n3079);
nor_4  g07357(new_n7743, new_n7742, new_n3078);
nor_4  g07358(new_n7744, new_n7743, new_n3077);
nor_4  g07359(new_n7745, new_n7744, new_n3076);
nor_4  g07360(new_n7746, new_n7745, new_n3075);
nor_4  g07361(new_n7747, new_n7746, new_n3074);
nor_4  g07362(new_n7748_1, new_n7747, new_n3073);
nor_4  g07363(new_n7749, new_n7748_1, new_n3072);
nor_4  g07364(new_n7750, new_n7749, new_n3071);
nor_4  g07365(new_n7751, new_n7750, new_n3070);
nor_4  g07366(new_n7752, new_n7751, new_n3069);
nor_4  g07367(new_n7753, new_n7752, new_n3068);
nor_4  g07368(new_n7754, new_n7753, new_n3067);
nor_4  g07369(new_n7755, new_n7754, new_n3066);
nor_4  g07370(new_n7756, new_n7755, new_n3065);
nor_4  g07371(new_n7757, new_n7756, new_n3064);
nor_4  g07372(new_n7758, new_n7757, new_n3063);
nor_4  g07373(new_n7759, new_n7758, new_n3062);
nor_4  g07374(new_n7760, new_n7759, new_n3061);
nor_4  g07375(new_n7761, new_n7760, new_n3354);
nor_4  g07376(new_n7762, new_n7761, new_n3353);
not_3  g07377(new_n7763, new_n7762);
nand_4 g07378(new_n7764, new_n7763, new_n517);
nand_4 g07379(new_n7765, new_n7764, new_n705);
nand_4 g07380(new_n7766, new_n7765, new_n511);
nand_4 g07381(new_n7767, new_n7766, new_n711);
nand_4 g07382(new_n7768, new_n7767, new_n506);
nand_4 g07383(new_n7769, new_n7768, new_n719);
nand_4 g07384(new_n7770, new_n7769, new_n500);
nand_4 g07385(new_n7771_1, new_n7770, new_n727);
nand_4 g07386(new_n7772, new_n7771_1, new_n494);
nand_4 g07387(new_n7773, new_n7772, new_n735);
nand_4 g07388(new_n7774, new_n7773, new_n488);
nand_4 g07389(new_n7775, new_n7774, new_n743);
nand_4 g07390(new_n7776, new_n7775, new_n482);
nand_4 g07391(new_n7777, new_n7776, new_n751);
nand_4 g07392(new_n7778, new_n7777, n9830);
nor_4  g07393(n7152, new_n7778, new_n755);
nand_4 g07394(new_n7780, new_n1680, new_n667);
nand_4 g07395(new_n7781, new_n7780, new_n1678);
nand_4 g07396(new_n7782, new_n7781, new_n1674);
nand_4 g07397(new_n7783, new_n7782, new_n1890);
nand_4 g07398(new_n7784, new_n7783, new_n1669);
nand_4 g07399(new_n7785, new_n7784, new_n1665);
nand_4 g07400(new_n7786, new_n7785, new_n1661);
nand_4 g07401(new_n7787, new_n7786, new_n1657);
nand_4 g07402(new_n7788, new_n7787, new_n1652);
nand_4 g07403(new_n7789, new_n7788, new_n1648);
nand_4 g07404(new_n7790, new_n7789, new_n1644);
nand_4 g07405(new_n7791, new_n7790, new_n1640);
nand_4 g07406(new_n7792, new_n7791, new_n1636);
nand_4 g07407(new_n7793, new_n7792, new_n1632);
nand_4 g07408(new_n7794, new_n7793, new_n1378);
nand_4 g07409(new_n7795, new_n7794, new_n1372);
nand_4 g07410(new_n7796, new_n7795, new_n1367);
nand_4 g07411(new_n7797, new_n7796, new_n1363);
nand_4 g07412(new_n7798, new_n7797, new_n1360);
nand_4 g07413(new_n7799, new_n7798, new_n1357);
nand_4 g07414(new_n7800, new_n7799, new_n1354);
nand_4 g07415(new_n7801, new_n7800, new_n1352);
nand_4 g07416(new_n7802, new_n7801, new_n1350);
nand_4 g07417(new_n7803, new_n7802, new_n1347_1);
nand_4 g07418(new_n7804, new_n7803, new_n1344);
nand_4 g07419(new_n7805, new_n7804, new_n1341);
nand_4 g07420(new_n7806, new_n7805, new_n1338);
nand_4 g07421(new_n7807, new_n7806, new_n1395);
nand_4 g07422(new_n7808, new_n7807, new_n1335);
nand_4 g07423(new_n7809, new_n7808, new_n1332);
nand_4 g07424(new_n7810, new_n7809, new_n1328);
nand_4 g07425(new_n7811, new_n7810, new_n1403);
nand_4 g07426(new_n7812, new_n7811, new_n1325);
nand_4 g07427(new_n7813, new_n7812, new_n1410);
nand_4 g07428(new_n7814, new_n7813, new_n1413);
nand_4 g07429(new_n7815, new_n7814, new_n1322);
nand_4 g07430(new_n7816, new_n7815, new_n1317);
nand_4 g07431(new_n7817, new_n7816, new_n1315);
nand_4 g07432(new_n7818, new_n7817, new_n1419);
nand_4 g07433(new_n7819, new_n7818, new_n1310);
nand_4 g07434(new_n7820, new_n7819, new_n1305);
nand_4 g07435(new_n7821, new_n7820, new_n1427);
nand_4 g07436(new_n7822, new_n7821, new_n1431);
nand_4 g07437(new_n7823, new_n7822, new_n1302);
nand_4 g07438(new_n7824, new_n7823, new_n1298);
nand_4 g07439(new_n7825_1, new_n7824, new_n1295);
nand_4 g07440(new_n7826, new_n7825_1, new_n1291);
nand_4 g07441(new_n7827, new_n7826, new_n1288);
nand_4 g07442(new_n7828, new_n7827, new_n1284);
nand_4 g07443(new_n7829, new_n7828, new_n1280);
nand_4 g07444(new_n7830, new_n7829, new_n1275);
not_3  g07445(new_n7831, new_n7830);
nor_4  g07446(new_n7832_1, new_n7831, new_n1446);
nor_4  g07447(new_n7833, new_n7832_1, new_n1271);
nor_4  g07448(new_n7834, new_n7833, new_n1266);
nor_4  g07449(new_n7835, new_n7834, new_n1261);
nor_4  g07450(new_n7836, new_n7835, new_n1257);
nor_4  g07451(new_n7837, new_n7836, new_n1252);
nor_4  g07452(new_n7838, new_n7837, new_n1458);
nor_4  g07453(new_n7839, new_n7838, new_n1463);
nor_4  g07454(new_n7840, new_n7839, new_n1469);
nor_4  g07455(new_n7841, new_n7840, new_n1248);
nor_4  g07456(new_n7842, new_n7841, new_n1475);
nor_4  g07457(new_n7843, new_n7842, new_n1244);
nor_4  g07458(new_n7844, new_n7843, new_n1243);
nor_4  g07459(new_n7845, new_n7844, new_n1242);
nor_4  g07460(new_n7846, new_n7845, new_n1241);
nor_4  g07461(new_n7847, new_n7846, new_n1240);
nor_4  g07462(new_n7848, new_n7847, new_n1239);
nor_4  g07463(new_n7849, new_n7848, new_n3082);
nor_4  g07464(new_n7850, new_n7849, new_n3081);
nor_4  g07465(new_n7851, new_n7850, new_n3080);
nor_4  g07466(new_n7852, new_n7851, new_n3079);
nor_4  g07467(new_n7853, new_n7852, new_n3078);
nor_4  g07468(new_n7854, new_n7853, new_n3077);
nor_4  g07469(new_n7855, new_n7854, new_n3076);
nor_4  g07470(new_n7856, new_n7855, new_n3075);
nor_4  g07471(new_n7857, new_n7856, new_n3074);
nor_4  g07472(new_n7858, new_n7857, new_n3073);
not_3  g07473(new_n7859, new_n7858);
nand_4 g07474(new_n7860, new_n7859, new_n652);
nand_4 g07475(new_n7861, new_n7860, new_n549);
nand_4 g07476(new_n7862, new_n7861, new_n544);
nand_4 g07477(new_n7863, new_n7862, new_n660);
nand_4 g07478(new_n7864, new_n7863, new_n539);
nand_4 g07479(new_n7865, new_n7864, new_n534);
nand_4 g07480(new_n7866, new_n7865, n13093);
nor_4  g07481(n7246, new_n7866, new_n525);
not_3  g07482(new_n7868, n10573);
not_3  g07483(new_n7869, new_n1110);
nand_4 g07484(new_n7870, new_n7869, new_n7868);
nand_4 g07485(new_n7871, new_n7870, new_n604);
nand_4 g07486(new_n7872, new_n7871, new_n612);
nand_4 g07487(new_n7873, new_n7872, new_n575);
nand_4 g07488(new_n7874, new_n7873, new_n619);
nand_4 g07489(new_n7875, new_n7874, new_n570);
nand_4 g07490(new_n7876, new_n7875, new_n625);
nand_4 g07491(new_n7877, new_n7876, new_n564);
nand_4 g07492(new_n7878, new_n7877, new_n632);
nand_4 g07493(new_n7879, new_n7878, new_n638);
nand_4 g07494(new_n7880, new_n7879, new_n559);
nand_4 g07495(new_n7881, new_n7880, new_n554);
nand_4 g07496(new_n7882, new_n7881, new_n646);
nand_4 g07497(new_n7883, new_n7882, new_n652);
nand_4 g07498(new_n7884, new_n7883, new_n549);
nand_4 g07499(new_n7885, new_n7884, new_n544);
nand_4 g07500(new_n7886, new_n7885, new_n660);
nand_4 g07501(new_n7887, new_n7886, new_n539);
nand_4 g07502(new_n7888, new_n7887, new_n534);
nand_4 g07503(new_n7889, new_n7888, new_n529);
nand_4 g07504(new_n7890, new_n7889, new_n668);
nand_4 g07505(new_n7891, new_n7890, new_n674_1);
nand_4 g07506(new_n7892, new_n7891, new_n681);
nand_4 g07507(new_n7893, new_n7892, new_n523);
nand_4 g07508(new_n7894, new_n7893, new_n687);
nand_4 g07509(new_n7895, new_n7894, new_n693);
nand_4 g07510(new_n7896, new_n7895, new_n699);
nand_4 g07511(new_n7897, new_n7896, new_n517);
nand_4 g07512(new_n7898, new_n7897, new_n705);
nand_4 g07513(new_n7899, new_n7898, new_n511);
nand_4 g07514(new_n7900, new_n7899, new_n711);
nand_4 g07515(new_n7901, new_n7900, new_n506);
nand_4 g07516(new_n7902, new_n7901, new_n719);
nand_4 g07517(new_n7903, new_n7902, new_n500);
nand_4 g07518(new_n7904, new_n7903, new_n727);
nand_4 g07519(new_n7905, new_n7904, new_n494);
nand_4 g07520(new_n7906, new_n7905, new_n735);
nand_4 g07521(new_n7907, new_n7906, new_n488);
nand_4 g07522(new_n7908, new_n7907, new_n743);
nand_4 g07523(new_n7909, new_n7908, new_n482);
nand_4 g07524(new_n7910, new_n7909, new_n751);
nand_4 g07525(new_n7911, new_n7910, new_n758);
nand_4 g07526(new_n7912, new_n7911, new_n765);
nand_4 g07527(new_n7913, new_n7912, new_n476);
nand_4 g07528(new_n7914, new_n7913, new_n773);
nand_4 g07529(new_n7915, new_n7914, new_n780);
not_3  g07530(new_n7916, new_n7915);
nor_4  g07531(new_n7917, new_n7916, new_n788);
nor_4  g07532(new_n7918, new_n7917, new_n471);
nor_4  g07533(new_n7919, new_n7918, new_n796);
nor_4  g07534(new_n7920, new_n7919, new_n804);
nor_4  g07535(new_n7921, new_n7920, new_n810);
nor_4  g07536(new_n7922, new_n7921, new_n2043);
nor_4  g07537(new_n7923, new_n7922, new_n2042);
nor_4  g07538(new_n7924, new_n7923, new_n2041);
nor_4  g07539(new_n7925, new_n7924, new_n2040);
nor_4  g07540(new_n7926, new_n7925, new_n2039);
nor_4  g07541(new_n7927, new_n7926, new_n2038);
nor_4  g07542(new_n7928, new_n7927, new_n2037);
nor_4  g07543(new_n7929, new_n7928, new_n2036);
nor_4  g07544(new_n7930, new_n7929, new_n2035);
nor_4  g07545(new_n7931, new_n7930, new_n2034);
nor_4  g07546(new_n7932, new_n7931, new_n2033);
nor_4  g07547(new_n7933, new_n7932, new_n2032);
nor_4  g07548(new_n7934, new_n7933, new_n2031);
nor_4  g07549(new_n7935, new_n7934, new_n2030);
nor_4  g07550(new_n7936, new_n7935, new_n2029);
nor_4  g07551(new_n7937, new_n7936, new_n2028);
nor_4  g07552(new_n7938, new_n7937, new_n2027_1);
nor_4  g07553(new_n7939, new_n7938, new_n2026);
nor_4  g07554(new_n7940, new_n7939, new_n2025);
not_3  g07555(new_n7941_1, new_n7940);
nand_4 g07556(new_n7942, new_n7941_1, new_n881);
nand_4 g07557(new_n7943, new_n7942, new_n413);
nand_4 g07558(new_n7944, new_n7943, new_n889);
nand_4 g07559(new_n7945, new_n7944, new_n896);
nand_4 g07560(new_n7946, new_n7945, new_n901);
nand_4 g07561(new_n7947, new_n7946, new_n408);
nand_4 g07562(new_n7948, new_n7947, new_n908);
nand_4 g07563(new_n7949, new_n7948, new_n403);
nand_4 g07564(new_n7950, new_n7949, new_n398);
nand_4 g07565(new_n7951, new_n7950, new_n393);
nand_4 g07566(new_n7952, new_n7951, new_n916);
nand_4 g07567(new_n7953, new_n7952, new_n1123);
nand_4 g07568(new_n7954, new_n7953, new_n1164);
nand_4 g07569(new_n7955, new_n7954, new_n1120);
nand_4 g07570(new_n7956, new_n7955, new_n1169);
nand_4 g07571(new_n7957, new_n7956, n1776);
nor_4  g07572(n7265, new_n7957, new_n1113);
nand_4 g07573(new_n7959, new_n1442, new_n1270);
nand_4 g07574(new_n7960, new_n7959, new_n1265_1);
nand_4 g07575(new_n7961, new_n7960, new_n1260);
nand_4 g07576(new_n7962, new_n7961, new_n1256);
nand_4 g07577(new_n7963, new_n7962, new_n1251);
nand_4 g07578(new_n7964, new_n7963, new_n1457);
nand_4 g07579(new_n7965, new_n7964, new_n1462);
nand_4 g07580(new_n7966, new_n7965, new_n1468);
nand_4 g07581(new_n7967, new_n7966, new_n1247);
nand_4 g07582(new_n7968, new_n7967, new_n1474);
nand_4 g07583(new_n7969, new_n7968, new_n592);
nand_4 g07584(new_n7970, new_n7969, new_n585);
nand_4 g07585(new_n7971, new_n7970, new_n580);
nand_4 g07586(new_n7972_1, new_n7971, new_n600);
nand_4 g07587(new_n7973, new_n7972_1, new_n606);
nand_4 g07588(new_n7974, new_n7973, new_n612);
nand_4 g07589(new_n7975, new_n7974, new_n575);
nand_4 g07590(new_n7976, new_n7975, new_n619);
nand_4 g07591(new_n7977, new_n7976, new_n570);
nand_4 g07592(new_n7978, new_n7977, new_n625);
nand_4 g07593(new_n7979, new_n7978, new_n564);
nand_4 g07594(new_n7980, new_n7979, new_n632);
nand_4 g07595(new_n7981, new_n7980, new_n638);
nand_4 g07596(new_n7982, new_n7981, new_n559);
nand_4 g07597(new_n7983, new_n7982, new_n554);
nand_4 g07598(new_n7984, new_n7983, new_n646);
nand_4 g07599(new_n7985, new_n7984, new_n652);
nand_4 g07600(new_n7986, new_n7985, new_n549);
nand_4 g07601(new_n7987, new_n7986, new_n544);
nand_4 g07602(new_n7988_1, new_n7987, new_n660);
nand_4 g07603(new_n7989, new_n7988_1, new_n539);
nand_4 g07604(new_n7990, new_n7989, new_n534);
nand_4 g07605(new_n7991, new_n7990, new_n529);
nand_4 g07606(new_n7992, new_n7991, new_n668);
nand_4 g07607(new_n7993, new_n7992, new_n674_1);
nand_4 g07608(new_n7994, new_n7993, new_n681);
nand_4 g07609(new_n7995, new_n7994, new_n523);
nand_4 g07610(new_n7996, new_n7995, new_n687);
nand_4 g07611(new_n7997, new_n7996, new_n693);
nand_4 g07612(new_n7998, new_n7997, new_n699);
nand_4 g07613(new_n7999, new_n7998, new_n517);
nand_4 g07614(new_n8000, new_n7999, new_n705);
nand_4 g07615(new_n8001, new_n8000, new_n511);
nand_4 g07616(new_n8002_1, new_n8001, new_n711);
nand_4 g07617(new_n8003, new_n8002_1, new_n506);
nand_4 g07618(new_n8004, new_n8003, new_n719);
nand_4 g07619(new_n8005, new_n8004, new_n500);
nand_4 g07620(new_n8006, new_n8005, new_n727);
nand_4 g07621(new_n8007, new_n8006, new_n494);
nand_4 g07622(new_n8008, new_n8007, new_n735);
nand_4 g07623(new_n8009, new_n8008, new_n488);
not_3  g07624(new_n8010, new_n8009);
nor_4  g07625(new_n8011, new_n8010, new_n744);
nor_4  g07626(new_n8012, new_n8011, new_n483);
nor_4  g07627(new_n8013, new_n8012, new_n752);
nor_4  g07628(new_n8014, new_n8013, new_n759);
nor_4  g07629(new_n8015, new_n8014, new_n766);
nor_4  g07630(new_n8016, new_n8015, new_n477);
nor_4  g07631(new_n8017, new_n8016, new_n774);
nor_4  g07632(new_n8018, new_n8017, new_n781);
nor_4  g07633(new_n8019, new_n8018, new_n788);
nor_4  g07634(new_n8020, new_n8019, new_n471);
nor_4  g07635(new_n8021, new_n8020, new_n796);
nor_4  g07636(new_n8022, new_n8021, new_n804);
nor_4  g07637(new_n8023, new_n8022, new_n810);
nor_4  g07638(new_n8024, new_n8023, new_n2043);
nor_4  g07639(new_n8025, new_n8024, new_n2042);
nor_4  g07640(new_n8026, new_n8025, new_n2041);
nor_4  g07641(new_n8027, new_n8026, new_n2040);
nor_4  g07642(new_n8028, new_n8027, new_n2039);
nor_4  g07643(new_n8029, new_n8028, new_n2038);
nor_4  g07644(new_n8030, new_n8029, new_n2037);
nor_4  g07645(new_n8031, new_n8030, new_n2036);
nor_4  g07646(new_n8032, new_n8031, new_n2035);
nor_4  g07647(new_n8033, new_n8032, new_n2034);
nor_4  g07648(new_n8034, new_n8033, new_n2033);
nor_4  g07649(new_n8035, new_n8034, new_n2032);
nor_4  g07650(new_n8036, new_n8035, new_n2031);
nor_4  g07651(new_n8037, new_n8036, new_n2030);
not_3  g07652(new_n8038, new_n8037);
nand_4 g07653(new_n8039, new_n8038, new_n856);
nand_4 g07654(new_n8040, new_n8039, new_n863);
nand_4 g07655(new_n8041, new_n8040, new_n419);
nand_4 g07656(new_n8042, new_n8041, new_n869);
nand_4 g07657(new_n8043, new_n8042, new_n875);
nand_4 g07658(new_n8044_1, new_n8043, new_n881);
nand_4 g07659(new_n8045, new_n8044_1, n844);
nor_4  g07660(n7382, new_n8045, new_n410);
not_3  g07661(new_n8047, new_n1876);
nand_4 g07662(new_n8048, new_n8047, new_n1050);
nand_4 g07663(new_n8049, new_n8048, new_n1045);
nand_4 g07664(new_n8050, new_n8049, new_n1041);
nand_4 g07665(new_n8051, new_n8050, new_n1036);
nand_4 g07666(new_n8052, new_n8051, new_n1031);
nand_4 g07667(new_n8053, new_n8052, new_n1025);
nand_4 g07668(new_n8054, new_n8053, new_n1020);
nand_4 g07669(new_n8055, new_n8054, new_n1015);
nand_4 g07670(new_n8056, new_n8055, new_n1010);
nand_4 g07671(new_n8057, new_n8056, new_n1215);
nand_4 g07672(new_n8058, new_n8057, new_n1005);
nand_4 g07673(new_n8059, new_n8058, new_n1000);
nand_4 g07674(new_n8060, new_n8059, new_n994);
nand_4 g07675(new_n8061, new_n8060, new_n989);
nand_4 g07676(new_n8062, new_n8061, new_n984);
nand_4 g07677(new_n8063, new_n8062, new_n978);
nand_4 g07678(new_n8064, new_n8063, new_n973);
nand_4 g07679(new_n8065, new_n8064, new_n967);
nand_4 g07680(new_n8066, new_n8065, new_n964);
nand_4 g07681(new_n8067, new_n8066, new_n960);
nand_4 g07682(new_n8068_1, new_n8067, new_n957);
nand_4 g07683(new_n8069, new_n8068_1, new_n952);
nand_4 g07684(new_n8070, new_n8069, new_n948_1);
nand_4 g07685(new_n8071, new_n8070, new_n943);
nand_4 g07686(new_n8072, new_n8071, new_n938);
nand_4 g07687(new_n8073_1, new_n8072, new_n934);
nand_4 g07688(new_n8074, new_n8073_1, new_n929);
nand_4 g07689(new_n8075, new_n8074, new_n925);
nand_4 g07690(new_n8076, new_n8075, new_n2194);
nand_4 g07691(new_n8077, new_n8076, new_n2191);
nand_4 g07692(new_n8078, new_n8077, new_n2190);
nand_4 g07693(new_n8079, new_n8078, new_n2186);
nand_4 g07694(new_n8080, new_n8079, new_n2183);
nand_4 g07695(new_n8081, new_n8080, new_n2179);
nand_4 g07696(new_n8082, new_n8081, new_n2175_1);
nand_4 g07697(new_n8083, new_n8082, new_n2171);
nand_4 g07698(new_n8084, new_n8083, new_n2168);
nand_4 g07699(new_n8085_1, new_n8084, new_n2165);
nand_4 g07700(new_n8086, new_n8085_1, new_n2162);
nand_4 g07701(new_n8087, new_n8086, new_n2158);
nand_4 g07702(new_n8088, new_n8087, new_n2155);
nand_4 g07703(new_n8089, new_n8088, new_n2151);
nand_4 g07704(new_n8090, new_n8089, new_n2147);
nand_4 g07705(new_n8091, new_n8090, new_n1810);
nand_4 g07706(new_n8092, new_n8091, new_n1806);
nand_4 g07707(new_n8093, new_n8092, new_n1802);
nand_4 g07708(new_n8094, new_n8093, new_n1798);
nand_4 g07709(new_n8095, new_n8094, new_n1820);
nand_4 g07710(new_n8096, new_n8095, new_n1794);
nand_4 g07711(new_n8097, new_n8096, new_n1825);
nand_4 g07712(new_n8098, new_n8097, new_n1789);
not_3  g07713(new_n8099, new_n8098);
nor_4  g07714(new_n8100, new_n8099, new_n2301);
nor_4  g07715(new_n8101, new_n8100, new_n2300);
nor_4  g07716(new_n8102, new_n8101, new_n2299);
nor_4  g07717(new_n8103, new_n8102, new_n2298);
nor_4  g07718(new_n8104, new_n8103, new_n2297);
nor_4  g07719(new_n8105, new_n8104, new_n2296);
nor_4  g07720(new_n8106, new_n8105, new_n2295);
nor_4  g07721(new_n8107, new_n8106, new_n2294);
nor_4  g07722(new_n8108, new_n8107, new_n2293);
nor_4  g07723(new_n8109, new_n8108, new_n2292);
nor_4  g07724(new_n8110, new_n8109, new_n2291);
nor_4  g07725(new_n8111, new_n8110, new_n2290);
nor_4  g07726(new_n8112, new_n8111, new_n2289);
nor_4  g07727(new_n8113, new_n8112, new_n2288);
nor_4  g07728(new_n8114, new_n8113, new_n2287);
nor_4  g07729(new_n8115, new_n8114, new_n2286);
nor_4  g07730(new_n8116, new_n8115, new_n2285);
nor_4  g07731(new_n8117, new_n8116, new_n2284);
nor_4  g07732(new_n8118, new_n8117, new_n2283);
nor_4  g07733(new_n8119, new_n8118, new_n2145);
nor_4  g07734(new_n8120, new_n8119, new_n2144);
nor_4  g07735(new_n8121, new_n8120, new_n2143);
nor_4  g07736(new_n8122, new_n8121, new_n2142);
nor_4  g07737(new_n8123, new_n8122, new_n2141);
nor_4  g07738(new_n8124_1, new_n8123, new_n2140);
nor_4  g07739(new_n8125, new_n8124_1, new_n2139);
nor_4  g07740(new_n8126, new_n8125, new_n2138);
not_3  g07741(new_n8127, new_n8126);
nand_4 g07742(new_n8128, new_n8127, new_n1860);
nand_4 g07743(new_n8129, new_n8128, new_n1864);
nand_4 g07744(new_n8130, new_n8129, new_n1699);
nand_4 g07745(new_n8131, new_n8130, new_n1697);
nand_4 g07746(new_n8132, new_n8131, new_n1871);
nand_4 g07747(new_n8133, new_n8132, new_n1694);
nand_4 g07748(new_n8134, new_n8133, n13882);
nor_4  g07749(n7655, new_n8134, new_n657);
nand_4 g07750(new_n8136, new_n1183, new_n1175);
nand_4 g07751(new_n8137, new_n8136, new_n1102);
nand_4 g07752(new_n8138, new_n8137, new_n1099);
nand_4 g07753(new_n8139, new_n8138, new_n1191);
nand_4 g07754(new_n8140, new_n8139, new_n1095);
nand_4 g07755(new_n8141, new_n8140, new_n1091);
nand_4 g07756(new_n8142, new_n8141, new_n1088);
nand_4 g07757(new_n8143, new_n8142, new_n1084);
nand_4 g07758(new_n8144_1, new_n8143, new_n1079);
nand_4 g07759(new_n8145, new_n8144_1, new_n1074);
nand_4 g07760(new_n8146, new_n8145, new_n1070);
nand_4 g07761(new_n8147, new_n8146, new_n1064);
nand_4 g07762(new_n8148, new_n8147, new_n1061);
nand_4 g07763(new_n8149, new_n8148, new_n1055);
nand_4 g07764(new_n8150, new_n8149, new_n1050);
nand_4 g07765(new_n8151, new_n8150, new_n1045);
nand_4 g07766(new_n8152, new_n8151, new_n1041);
nand_4 g07767(new_n8153, new_n8152, new_n1036);
nand_4 g07768(new_n8154, new_n8153, new_n1031);
nand_4 g07769(new_n8155, new_n8154, new_n1025);
nand_4 g07770(new_n8156, new_n8155, new_n1020);
nand_4 g07771(new_n8157, new_n8156, new_n1015);
nand_4 g07772(new_n8158, new_n8157, new_n1010);
nand_4 g07773(new_n8159, new_n8158, new_n1215);
nand_4 g07774(new_n8160, new_n8159, new_n1005);
nand_4 g07775(new_n8161, new_n8160, new_n1000);
nand_4 g07776(new_n8162, new_n8161, new_n994);
nand_4 g07777(new_n8163, new_n8162, new_n989);
nand_4 g07778(new_n8164, new_n8163, new_n984);
nand_4 g07779(new_n8165, new_n8164, new_n978);
nand_4 g07780(new_n8166, new_n8165, new_n973);
nand_4 g07781(new_n8167, new_n8166, new_n967);
nand_4 g07782(new_n8168, new_n8167, new_n964);
nand_4 g07783(new_n8169, new_n8168, new_n960);
nand_4 g07784(new_n8170, new_n8169, new_n957);
not_3  g07785(new_n8171, new_n8170);
nor_4  g07786(new_n8172, new_n8171, new_n953);
nor_4  g07787(new_n8173, new_n8172, new_n3536);
nor_4  g07788(new_n8174, new_n8173, new_n3535);
nor_4  g07789(new_n8175, new_n8174, new_n3534);
nor_4  g07790(new_n8176, new_n8175, new_n2520);
nor_4  g07791(new_n8177, new_n8176, new_n2519);
nor_4  g07792(new_n8178, new_n8177, new_n2518);
nor_4  g07793(new_n8179, new_n8178, new_n2517);
nor_4  g07794(new_n8180, new_n8179, new_n2516);
nor_4  g07795(new_n8181, new_n8180, new_n2515);
nor_4  g07796(new_n8182, new_n8181, new_n2514);
nor_4  g07797(new_n8183, new_n8182, new_n2513);
nor_4  g07798(new_n8184, new_n8183, new_n2512);
nor_4  g07799(new_n8185, new_n8184, new_n2511);
nor_4  g07800(new_n8186, new_n8185, new_n2510);
nor_4  g07801(new_n8187, new_n8186, new_n2509);
nor_4  g07802(new_n8188, new_n8187, new_n2508);
nor_4  g07803(new_n8189, new_n8188, new_n2507);
nor_4  g07804(new_n8190, new_n8189, new_n2506);
not_3  g07805(new_n8191, new_n8190);
nand_4 g07806(new_n8192, new_n8191, new_n2155);
nand_4 g07807(new_n8193, new_n8192, new_n2151);
nand_4 g07808(new_n8194, new_n8193, new_n2147);
nand_4 g07809(new_n8195, new_n8194, new_n1810);
nand_4 g07810(new_n8196, new_n8195, new_n1806);
nand_4 g07811(new_n8197, new_n8196, new_n1802);
nand_4 g07812(new_n8198, new_n8197, new_n1798);
nand_4 g07813(new_n8199, new_n8198, new_n1820);
nand_4 g07814(new_n8200, new_n8199, new_n1794);
nand_4 g07815(new_n8201, new_n8200, new_n1825);
nand_4 g07816(new_n8202, new_n8201, new_n1789);
nand_4 g07817(new_n8203, new_n8202, new_n1785);
nand_4 g07818(new_n8204_1, new_n8203, new_n1780);
nand_4 g07819(new_n8205, new_n8204_1, new_n1777);
nand_4 g07820(new_n8206, new_n8205, new_n1774);
nand_4 g07821(new_n8207, new_n8206, new_n1834);
nand_4 g07822(new_n8208, new_n8207, new_n1769);
nand_4 g07823(new_n8209, new_n8208, new_n1766);
nand_4 g07824(new_n8210, new_n8209, new_n1762);
nand_4 g07825(new_n8211, new_n8210, new_n1758);
nand_4 g07826(new_n8212, new_n8211, new_n1754);
nand_4 g07827(new_n8213, new_n8212, new_n1751);
nand_4 g07828(new_n8214, new_n8213, new_n1748);
nand_4 g07829(new_n8215_1, new_n8214, new_n1746);
nand_4 g07830(new_n8216, new_n8215_1, new_n1742);
nand_4 g07831(new_n8217, new_n8216, new_n1738);
nand_4 g07832(new_n8218, new_n8217, new_n1736);
nand_4 g07833(new_n8219, new_n8218, new_n1732);
nand_4 g07834(new_n8220, new_n8219, new_n1729);
nand_4 g07835(new_n8221, new_n8220, new_n1726);
nand_4 g07836(new_n8222, new_n8221, n1763);
nor_4  g07837(n7771, new_n8222, new_n609);
nand_4 g07838(new_n8224, new_n2153, new_n1314);
nand_4 g07839(new_n8225, new_n8224, new_n2151);
nand_4 g07840(new_n8226, new_n8225, new_n2147);
nand_4 g07841(new_n8227, new_n8226, new_n1810);
nand_4 g07842(new_n8228, new_n8227, new_n1806);
nand_4 g07843(new_n8229, new_n8228, new_n1802);
nand_4 g07844(new_n8230, new_n8229, new_n1798);
nand_4 g07845(new_n8231, new_n8230, new_n1820);
nand_4 g07846(new_n8232, new_n8231, new_n1794);
nand_4 g07847(new_n8233, new_n8232, new_n1825);
nand_4 g07848(new_n8234, new_n8233, new_n1789);
nand_4 g07849(new_n8235, new_n8234, new_n1785);
nand_4 g07850(new_n8236, new_n8235, new_n1780);
nand_4 g07851(new_n8237, new_n8236, new_n1777);
nand_4 g07852(new_n8238, new_n8237, new_n1774);
nand_4 g07853(new_n8239, new_n8238, new_n1834);
nand_4 g07854(new_n8240, new_n8239, new_n1769);
nand_4 g07855(new_n8241, new_n8240, new_n1766);
nand_4 g07856(new_n8242, new_n8241, new_n1762);
nand_4 g07857(new_n8243, new_n8242, new_n1758);
nand_4 g07858(new_n8244, new_n8243, new_n1754);
nand_4 g07859(new_n8245, new_n8244, new_n1751);
nand_4 g07860(new_n8246, new_n8245, new_n1748);
nand_4 g07861(new_n8247, new_n8246, new_n1746);
nand_4 g07862(new_n8248, new_n8247, new_n1742);
nand_4 g07863(new_n8249, new_n8248, new_n1738);
nand_4 g07864(new_n8250, new_n8249, new_n1736);
nand_4 g07865(new_n8251, new_n8250, new_n1732);
nand_4 g07866(new_n8252, new_n8251, new_n1729);
nand_4 g07867(new_n8253, new_n8252, new_n1726);
nand_4 g07868(new_n8254, new_n8253, new_n1724);
nand_4 g07869(new_n8255, new_n8254, new_n1721);
nand_4 g07870(new_n8256, new_n8255, new_n1718);
nand_4 g07871(new_n8257, new_n8256, new_n1715);
nand_4 g07872(new_n8258, new_n8257, new_n1711);
nand_4 g07873(new_n8259, new_n8258, new_n1708);
nand_4 g07874(new_n8260, new_n8259, new_n1705);
nand_4 g07875(new_n8261, new_n8260, new_n1703);
nand_4 g07876(new_n8262_1, new_n8261, new_n1860);
nand_4 g07877(new_n8263, new_n8262_1, new_n1864);
nand_4 g07878(new_n8264, new_n8263, new_n1699);
nand_4 g07879(new_n8265, new_n8264, new_n1697);
nand_4 g07880(new_n8266, new_n8265, new_n1871);
nand_4 g07881(new_n8267, new_n8266, new_n1694);
nand_4 g07882(new_n8268, new_n8267, new_n1690);
nand_4 g07883(new_n8269, new_n8268, new_n1878);
nand_4 g07884(new_n8270, new_n8269, new_n1882);
nand_4 g07885(new_n8271, new_n8270, new_n1686);
nand_4 g07886(new_n8272, new_n8271, new_n1682);
nand_4 g07887(new_n8273, new_n8272, new_n1678);
not_3  g07888(new_n8274, new_n8273);
nor_4  g07889(new_n8275, new_n8274, new_n1675);
nor_4  g07890(new_n8276, new_n8275, new_n1891);
nor_4  g07891(new_n8277, new_n8276, new_n1670);
nor_4  g07892(new_n8278, new_n8277, new_n1666);
nor_4  g07893(new_n8279, new_n8278, new_n1662);
nor_4  g07894(new_n8280, new_n8279, new_n1658);
nor_4  g07895(new_n8281, new_n8280, new_n1653);
nor_4  g07896(new_n8282, new_n8281, new_n1649);
nor_4  g07897(new_n8283, new_n8282, new_n1645);
nor_4  g07898(new_n8284, new_n8283, new_n1641);
nor_4  g07899(new_n8285, new_n8284, new_n1637_1);
nor_4  g07900(new_n8286, new_n8285, new_n1633);
nor_4  g07901(new_n8287, new_n8286, new_n1629);
nor_4  g07902(new_n8288, new_n8287, new_n1628);
nor_4  g07903(new_n8289, new_n8288, new_n1627);
nor_4  g07904(new_n8290, new_n8289, new_n1626);
nor_4  g07905(new_n8291, new_n8290, new_n4700);
nor_4  g07906(new_n8292, new_n8291, new_n4699);
nor_4  g07907(new_n8293, new_n8292, new_n3722);
nor_4  g07908(new_n8294, new_n8293, new_n3721);
nor_4  g07909(new_n8295, new_n8294, new_n3720);
nor_4  g07910(new_n8296, new_n8295, new_n3719);
nor_4  g07911(new_n8297, new_n8296, new_n3718);
nor_4  g07912(new_n8298, new_n8297, new_n3717);
nor_4  g07913(new_n8299, new_n8298, new_n3716);
not_3  g07914(new_n8300, new_n8299);
nand_4 g07915(new_n8301, new_n8300, new_n1395);
nand_4 g07916(new_n8302_1, new_n8301, new_n1335);
nand_4 g07917(new_n8303, new_n8302_1, new_n1332);
nand_4 g07918(new_n8304, new_n8303, new_n1328);
nand_4 g07919(new_n8305, new_n8304, new_n1403);
nand_4 g07920(new_n8306_1, new_n8305, new_n1325);
nand_4 g07921(new_n8307, new_n8306_1, new_n1410);
nand_4 g07922(new_n8308, new_n8307, new_n1413);
nand_4 g07923(new_n8309, new_n8308, new_n1322);
nand_4 g07924(new_n8310, new_n8309, n11404);
nor_4  g07925(n7825, new_n8310, new_n824);
not_3  g07926(new_n8312, n12009);
not_3  g07927(new_n8313, new_n1177);
nand_4 g07928(new_n8314, new_n8313, new_n8312);
nand_4 g07929(new_n8315_1, new_n8314, new_n573);
nand_4 g07930(new_n8316, new_n8315_1, new_n619);
nand_4 g07931(new_n8317, new_n8316, new_n570);
nand_4 g07932(new_n8318, new_n8317, new_n625);
nand_4 g07933(new_n8319, new_n8318, new_n564);
nand_4 g07934(new_n8320, new_n8319, new_n632);
nand_4 g07935(new_n8321, new_n8320, new_n638);
nand_4 g07936(new_n8322, new_n8321, new_n559);
nand_4 g07937(new_n8323, new_n8322, new_n554);
nand_4 g07938(new_n8324, new_n8323, new_n646);
nand_4 g07939(new_n8325, new_n8324, new_n652);
nand_4 g07940(new_n8326, new_n8325, new_n549);
nand_4 g07941(new_n8327, new_n8326, new_n544);
nand_4 g07942(new_n8328, new_n8327, new_n660);
nand_4 g07943(new_n8329, new_n8328, new_n539);
nand_4 g07944(new_n8330, new_n8329, new_n534);
nand_4 g07945(new_n8331, new_n8330, new_n529);
nand_4 g07946(new_n8332, new_n8331, new_n668);
nand_4 g07947(new_n8333, new_n8332, new_n674_1);
nand_4 g07948(new_n8334, new_n8333, new_n681);
nand_4 g07949(new_n8335, new_n8334, new_n523);
nand_4 g07950(new_n8336, new_n8335, new_n687);
nand_4 g07951(new_n8337, new_n8336, new_n693);
nand_4 g07952(new_n8338, new_n8337, new_n699);
nand_4 g07953(new_n8339, new_n8338, new_n517);
nand_4 g07954(new_n8340, new_n8339, new_n705);
nand_4 g07955(new_n8341, new_n8340, new_n511);
nand_4 g07956(new_n8342, new_n8341, new_n711);
nand_4 g07957(new_n8343, new_n8342, new_n506);
nand_4 g07958(new_n8344, new_n8343, new_n719);
nand_4 g07959(new_n8345, new_n8344, new_n500);
nand_4 g07960(new_n8346, new_n8345, new_n727);
nand_4 g07961(new_n8347, new_n8346, new_n494);
nand_4 g07962(new_n8348, new_n8347, new_n735);
nand_4 g07963(new_n8349, new_n8348, new_n488);
nand_4 g07964(new_n8350, new_n8349, new_n743);
nand_4 g07965(new_n8351, new_n8350, new_n482);
nand_4 g07966(new_n8352, new_n8351, new_n751);
nand_4 g07967(new_n8353, new_n8352, new_n758);
nand_4 g07968(new_n8354, new_n8353, new_n765);
nand_4 g07969(new_n8355, new_n8354, new_n476);
nand_4 g07970(new_n8356, new_n8355, new_n773);
nand_4 g07971(new_n8357, new_n8356, new_n780);
nand_4 g07972(new_n8358, new_n8357, new_n787);
nand_4 g07973(new_n8359, new_n8358, new_n470);
not_3  g07974(new_n8360, new_n8359);
nor_4  g07975(new_n8361, new_n8360, new_n796);
nor_4  g07976(new_n8362, new_n8361, new_n804);
nor_4  g07977(new_n8363, new_n8362, new_n810);
nor_4  g07978(new_n8364, new_n8363, new_n2043);
nor_4  g07979(new_n8365, new_n8364, new_n2042);
nor_4  g07980(new_n8366, new_n8365, new_n2041);
nor_4  g07981(new_n8367, new_n8366, new_n2040);
nor_4  g07982(new_n8368, new_n8367, new_n2039);
nor_4  g07983(new_n8369, new_n8368, new_n2038);
nor_4  g07984(new_n8370, new_n8369, new_n2037);
nor_4  g07985(new_n8371, new_n8370, new_n2036);
nor_4  g07986(new_n8372, new_n8371, new_n2035);
nor_4  g07987(new_n8373, new_n8372, new_n2034);
nor_4  g07988(new_n8374, new_n8373, new_n2033);
nor_4  g07989(new_n8375, new_n8374, new_n2032);
nor_4  g07990(new_n8376, new_n8375, new_n2031);
nor_4  g07991(new_n8377, new_n8376, new_n2030);
nor_4  g07992(new_n8378, new_n8377, new_n2029);
nor_4  g07993(new_n8379, new_n8378, new_n2028);
nor_4  g07994(new_n8380, new_n8379, new_n2027_1);
nor_4  g07995(new_n8381, new_n8380, new_n2026);
nor_4  g07996(new_n8382, new_n8381, new_n2025);
nor_4  g07997(new_n8383, new_n8382, new_n2024);
nor_4  g07998(new_n8384, new_n8383, new_n2023);
not_3  g07999(new_n8385, new_n8384);
nand_4 g08000(new_n8386, new_n8385, new_n889);
nand_4 g08001(new_n8387, new_n8386, new_n896);
nand_4 g08002(new_n8388, new_n8387, new_n901);
nand_4 g08003(new_n8389, new_n8388, new_n408);
nand_4 g08004(new_n8390, new_n8389, new_n908);
nand_4 g08005(new_n8391, new_n8390, new_n403);
nand_4 g08006(new_n8392, new_n8391, new_n398);
nand_4 g08007(new_n8393, new_n8392, new_n393);
nand_4 g08008(new_n8394, new_n8393, new_n916);
nand_4 g08009(new_n8395, new_n8394, new_n1123);
nand_4 g08010(new_n8396, new_n8395, new_n1164);
nand_4 g08011(new_n8397_1, new_n8396, new_n1120);
nand_4 g08012(new_n8398, new_n8397_1, new_n1169);
nand_4 g08013(new_n8399, new_n8398, new_n1116);
nand_4 g08014(new_n8400, new_n8399, new_n1111);
nand_4 g08015(new_n8401, new_n8400, n13363);
nor_4  g08016(n8068, new_n8401, new_n1104);
nand_4 g08017(new_n8403, new_n1656, new_n1003);
nand_4 g08018(new_n8404, new_n8403, new_n1000);
nand_4 g08019(new_n8405, new_n8404, new_n994);
nand_4 g08020(new_n8406, new_n8405, new_n989);
nand_4 g08021(new_n8407, new_n8406, new_n984);
nand_4 g08022(new_n8408, new_n8407, new_n978);
nand_4 g08023(new_n8409, new_n8408, new_n973);
nand_4 g08024(new_n8410, new_n8409, new_n967);
nand_4 g08025(new_n8411, new_n8410, new_n964);
nand_4 g08026(new_n8412, new_n8411, new_n960);
nand_4 g08027(new_n8413, new_n8412, new_n957);
nand_4 g08028(new_n8414, new_n8413, new_n952);
nand_4 g08029(new_n8415, new_n8414, new_n948_1);
nand_4 g08030(new_n8416, new_n8415, new_n943);
nand_4 g08031(new_n8417, new_n8416, new_n938);
nand_4 g08032(new_n8418, new_n8417, new_n934);
nand_4 g08033(new_n8419, new_n8418, new_n929);
nand_4 g08034(new_n8420, new_n8419, new_n925);
nand_4 g08035(new_n8421, new_n8420, new_n2194);
nand_4 g08036(new_n8422, new_n8421, new_n2191);
nand_4 g08037(new_n8423, new_n8422, new_n2190);
nand_4 g08038(new_n8424, new_n8423, new_n2186);
nand_4 g08039(new_n8425, new_n8424, new_n2183);
nand_4 g08040(new_n8426, new_n8425, new_n2179);
nand_4 g08041(new_n8427, new_n8426, new_n2175_1);
nand_4 g08042(new_n8428, new_n8427, new_n2171);
nand_4 g08043(new_n8429, new_n8428, new_n2168);
nand_4 g08044(new_n8430, new_n8429, new_n2165);
nand_4 g08045(new_n8431, new_n8430, new_n2162);
nand_4 g08046(new_n8432, new_n8431, new_n2158);
nand_4 g08047(new_n8433, new_n8432, new_n2155);
nand_4 g08048(new_n8434, new_n8433, new_n2151);
nand_4 g08049(new_n8435, new_n8434, new_n2147);
nand_4 g08050(new_n8436, new_n8435, new_n1810);
nand_4 g08051(new_n8437, new_n8436, new_n1806);
nand_4 g08052(new_n8438, new_n8437, new_n1802);
nand_4 g08053(new_n8439_1, new_n8438, new_n1798);
nand_4 g08054(new_n8440, new_n8439_1, new_n1820);
nand_4 g08055(new_n8441, new_n8440, new_n1794);
nand_4 g08056(new_n8442, new_n8441, new_n1825);
nand_4 g08057(new_n8443, new_n8442, new_n1789);
nand_4 g08058(new_n8444, new_n8443, new_n1785);
nand_4 g08059(new_n8445, new_n8444, new_n1780);
nand_4 g08060(new_n8446, new_n8445, new_n1777);
nand_4 g08061(new_n8447, new_n8446, new_n1774);
nand_4 g08062(new_n8448, new_n8447, new_n1834);
nand_4 g08063(new_n8449, new_n8448, new_n1769);
nand_4 g08064(new_n8450, new_n8449, new_n1766);
nand_4 g08065(new_n8451, new_n8450, new_n1762);
nand_4 g08066(new_n8452, new_n8451, new_n1758);
not_3  g08067(new_n8453, new_n8452);
nor_4  g08068(new_n8454, new_n8453, new_n2292);
nor_4  g08069(new_n8455, new_n8454, new_n2291);
nor_4  g08070(new_n8456, new_n8455, new_n2290);
nor_4  g08071(new_n8457, new_n8456, new_n2289);
nor_4  g08072(new_n8458, new_n8457, new_n2288);
nor_4  g08073(new_n8459, new_n8458, new_n2287);
nor_4  g08074(new_n8460, new_n8459, new_n2286);
nor_4  g08075(new_n8461, new_n8460, new_n2285);
nor_4  g08076(new_n8462, new_n8461, new_n2284);
nor_4  g08077(new_n8463_1, new_n8462, new_n2283);
nor_4  g08078(new_n8464, new_n8463_1, new_n2145);
nor_4  g08079(new_n8465, new_n8464, new_n2144);
nor_4  g08080(new_n8466, new_n8465, new_n2143);
nor_4  g08081(new_n8467, new_n8466, new_n2142);
nor_4  g08082(new_n8468, new_n8467, new_n2141);
nor_4  g08083(new_n8469, new_n8468, new_n2140);
nor_4  g08084(new_n8470, new_n8469, new_n2139);
nor_4  g08085(new_n8471_1, new_n8470, new_n2138);
nor_4  g08086(new_n8472, new_n8471_1, new_n2137);
nor_4  g08087(new_n8473, new_n8472, new_n2136);
nor_4  g08088(new_n8474, new_n8473, new_n2135);
nor_4  g08089(new_n8475, new_n8474, new_n2134);
nor_4  g08090(new_n8476, new_n8475, new_n2133);
nor_4  g08091(new_n8477, new_n8476, new_n2132);
nor_4  g08092(new_n8478, new_n8477, new_n1691);
not_3  g08093(new_n8479, new_n8478);
nand_4 g08094(new_n8480, new_n8479, new_n1878);
nand_4 g08095(new_n8481, new_n8480, new_n1882);
nand_4 g08096(new_n8482, new_n8481, new_n1686);
nand_4 g08097(new_n8483, new_n8482, new_n1682);
nand_4 g08098(new_n8484, new_n8483, new_n1678);
nand_4 g08099(new_n8485, new_n8484, new_n1674);
nand_4 g08100(new_n8486_1, new_n8485, new_n1890);
nand_4 g08101(new_n8487, new_n8486_1, new_n1669);
nand_4 g08102(new_n8488, new_n8487, new_n1665);
nand_4 g08103(new_n8489, new_n8488, n8800);
nor_4  g08104(n8085, new_n8489, new_n696);
nand_4 g08105(new_n8491, new_n1631, new_n971);
nand_4 g08106(new_n8492, new_n8491, new_n967);
nand_4 g08107(new_n8493, new_n8492, new_n964);
nand_4 g08108(new_n8494, new_n8493, new_n960);
nand_4 g08109(new_n8495, new_n8494, new_n957);
nand_4 g08110(new_n8496, new_n8495, new_n952);
nand_4 g08111(new_n8497, new_n8496, new_n948_1);
nand_4 g08112(new_n8498, new_n8497, new_n943);
nand_4 g08113(new_n8499, new_n8498, new_n938);
nand_4 g08114(new_n8500, new_n8499, new_n934);
nand_4 g08115(new_n8501, new_n8500, new_n929);
nand_4 g08116(new_n8502, new_n8501, new_n925);
nand_4 g08117(new_n8503, new_n8502, new_n2194);
nand_4 g08118(new_n8504, new_n8503, new_n2191);
nand_4 g08119(new_n8505, new_n8504, new_n2190);
nand_4 g08120(new_n8506, new_n8505, new_n2186);
nand_4 g08121(new_n8507, new_n8506, new_n2183);
nand_4 g08122(new_n8508, new_n8507, new_n2179);
nand_4 g08123(new_n8509, new_n8508, new_n2175_1);
nand_4 g08124(new_n8510, new_n8509, new_n2171);
nand_4 g08125(new_n8511, new_n8510, new_n2168);
nand_4 g08126(new_n8512, new_n8511, new_n2165);
nand_4 g08127(new_n8513, new_n8512, new_n2162);
nand_4 g08128(new_n8514, new_n8513, new_n2158);
nand_4 g08129(new_n8515, new_n8514, new_n2155);
nand_4 g08130(new_n8516, new_n8515, new_n2151);
nand_4 g08131(new_n8517, new_n8516, new_n2147);
nand_4 g08132(new_n8518, new_n8517, new_n1810);
nand_4 g08133(new_n8519, new_n8518, new_n1806);
nand_4 g08134(new_n8520, new_n8519, new_n1802);
nand_4 g08135(new_n8521, new_n8520, new_n1798);
nand_4 g08136(new_n8522, new_n8521, new_n1820);
nand_4 g08137(new_n8523, new_n8522, new_n1794);
nand_4 g08138(new_n8524, new_n8523, new_n1825);
nand_4 g08139(new_n8525, new_n8524, new_n1789);
nand_4 g08140(new_n8526, new_n8525, new_n1785);
nand_4 g08141(new_n8527, new_n8526, new_n1780);
nand_4 g08142(new_n8528, new_n8527, new_n1777);
nand_4 g08143(new_n8529, new_n8528, new_n1774);
nand_4 g08144(new_n8530, new_n8529, new_n1834);
nand_4 g08145(new_n8531, new_n8530, new_n1769);
nand_4 g08146(new_n8532, new_n8531, new_n1766);
nand_4 g08147(new_n8533, new_n8532, new_n1762);
nand_4 g08148(new_n8534, new_n8533, new_n1758);
nand_4 g08149(new_n8535, new_n8534, new_n1754);
nand_4 g08150(new_n8536, new_n8535, new_n1751);
nand_4 g08151(new_n8537, new_n8536, new_n1748);
nand_4 g08152(new_n8538, new_n8537, new_n1746);
nand_4 g08153(new_n8539, new_n8538, new_n1742);
nand_4 g08154(new_n8540, new_n8539, new_n1738);
nand_4 g08155(new_n8541, new_n8540, new_n1736);
not_3  g08156(new_n8542, new_n8541);
nor_4  g08157(new_n8543, new_n8542, new_n2285);
nor_4  g08158(new_n8544, new_n8543, new_n2284);
nor_4  g08159(new_n8545, new_n8544, new_n2283);
nor_4  g08160(new_n8546, new_n8545, new_n2145);
nor_4  g08161(new_n8547, new_n8546, new_n2144);
nor_4  g08162(new_n8548, new_n8547, new_n2143);
nor_4  g08163(new_n8549, new_n8548, new_n2142);
nor_4  g08164(new_n8550_1, new_n8549, new_n2141);
nor_4  g08165(new_n8551, new_n8550_1, new_n2140);
nor_4  g08166(new_n8552_1, new_n8551, new_n2139);
nor_4  g08167(new_n8553, new_n8552_1, new_n2138);
nor_4  g08168(new_n8554, new_n8553, new_n2137);
nor_4  g08169(new_n8555, new_n8554, new_n2136);
nor_4  g08170(new_n8556, new_n8555, new_n2135);
nor_4  g08171(new_n8557, new_n8556, new_n2134);
nor_4  g08172(new_n8558, new_n8557, new_n2133);
nor_4  g08173(new_n8559, new_n8558, new_n2132);
nor_4  g08174(new_n8560, new_n8559, new_n1691);
nor_4  g08175(new_n8561, new_n8560, new_n1879);
nor_4  g08176(new_n8562, new_n8561, new_n1883);
nor_4  g08177(new_n8563, new_n8562, new_n1687);
nor_4  g08178(new_n8564, new_n8563, new_n1683);
nor_4  g08179(new_n8565, new_n8564, new_n1679);
nor_4  g08180(new_n8566, new_n8565, new_n1675);
nor_4  g08181(new_n8567, new_n8566, new_n1891);
nor_4  g08182(new_n8568, new_n8567, new_n1670);
nor_4  g08183(new_n8569, new_n8568, new_n1666);
not_3  g08184(new_n8570, new_n8569);
nand_4 g08185(new_n8571, new_n8570, new_n1661);
nand_4 g08186(new_n8572, new_n8571, new_n1657);
nand_4 g08187(new_n8573, new_n8572, new_n1652);
nand_4 g08188(new_n8574, new_n8573, new_n1648);
nand_4 g08189(new_n8575, new_n8574, new_n1644);
nand_4 g08190(new_n8576, new_n8575, new_n1640);
nand_4 g08191(new_n8577, new_n8576, n9154);
nor_4  g08192(n8124, new_n8577, new_n716);
not_3  g08193(new_n8579, new_n914);
nand_4 g08194(new_n8580, new_n1247, new_n8579);
nand_4 g08195(new_n8581, new_n8580, new_n1474);
nand_4 g08196(new_n8582, new_n8581, new_n592);
nand_4 g08197(new_n8583, new_n8582, new_n585);
nand_4 g08198(new_n8584, new_n8583, new_n580);
nand_4 g08199(new_n8585, new_n8584, new_n600);
nand_4 g08200(new_n8586, new_n8585, new_n606);
nand_4 g08201(new_n8587, new_n8586, new_n612);
nand_4 g08202(new_n8588, new_n8587, new_n575);
nand_4 g08203(new_n8589, new_n8588, new_n619);
nand_4 g08204(new_n8590, new_n8589, new_n570);
nand_4 g08205(new_n8591, new_n8590, new_n625);
nand_4 g08206(new_n8592, new_n8591, new_n564);
nand_4 g08207(new_n8593, new_n8592, new_n632);
nand_4 g08208(new_n8594, new_n8593, new_n638);
nand_4 g08209(new_n8595, new_n8594, new_n559);
nand_4 g08210(new_n8596, new_n8595, new_n554);
nand_4 g08211(new_n8597, new_n8596, new_n646);
nand_4 g08212(new_n8598_1, new_n8597, new_n652);
nand_4 g08213(new_n8599, new_n8598_1, new_n549);
nand_4 g08214(new_n8600, new_n8599, new_n544);
nand_4 g08215(new_n8601, new_n8600, new_n660);
nand_4 g08216(new_n8602, new_n8601, new_n539);
nand_4 g08217(new_n8603, new_n8602, new_n534);
nand_4 g08218(new_n8604_1, new_n8603, new_n529);
nand_4 g08219(new_n8605, new_n8604_1, new_n668);
nand_4 g08220(new_n8606, new_n8605, new_n674_1);
nand_4 g08221(new_n8607, new_n8606, new_n681);
nand_4 g08222(new_n8608, new_n8607, new_n523);
nand_4 g08223(new_n8609, new_n8608, new_n687);
nand_4 g08224(new_n8610, new_n8609, new_n693);
nand_4 g08225(new_n8611, new_n8610, new_n699);
nand_4 g08226(new_n8612, new_n8611, new_n517);
nand_4 g08227(new_n8613, new_n8612, new_n705);
nand_4 g08228(new_n8614, new_n8613, new_n511);
nand_4 g08229(new_n8615, new_n8614, new_n711);
nand_4 g08230(new_n8616, new_n8615, new_n506);
nand_4 g08231(new_n8617, new_n8616, new_n719);
nand_4 g08232(new_n8618, new_n8617, new_n500);
nand_4 g08233(new_n8619, new_n8618, new_n727);
nand_4 g08234(new_n8620, new_n8619, new_n494);
nand_4 g08235(new_n8621, new_n8620, new_n735);
nand_4 g08236(new_n8622, new_n8621, new_n488);
nand_4 g08237(new_n8623, new_n8622, new_n743);
nand_4 g08238(new_n8624, new_n8623, new_n482);
nand_4 g08239(new_n8625, new_n8624, new_n751);
not_3  g08240(new_n8626, new_n8625);
nor_4  g08241(new_n8627, new_n8626, new_n759);
nor_4  g08242(new_n8628, new_n8627, new_n766);
nor_4  g08243(new_n8629, new_n8628, new_n477);
nor_4  g08244(new_n8630, new_n8629, new_n774);
nor_4  g08245(new_n8631, new_n8630, new_n781);
nor_4  g08246(new_n8632, new_n8631, new_n788);
nor_4  g08247(new_n8633, new_n8632, new_n471);
nor_4  g08248(new_n8634, new_n8633, new_n796);
nor_4  g08249(new_n8635_1, new_n8634, new_n804);
nor_4  g08250(new_n8636, new_n8635_1, new_n810);
nor_4  g08251(new_n8637, new_n8636, new_n2043);
nor_4  g08252(new_n8638, new_n8637, new_n2042);
nor_4  g08253(new_n8639, new_n8638, new_n2041);
nor_4  g08254(new_n8640, new_n8639, new_n2040);
nor_4  g08255(new_n8641, new_n8640, new_n2039);
nor_4  g08256(new_n8642, new_n8641, new_n2038);
nor_4  g08257(new_n8643, new_n8642, new_n2037);
nor_4  g08258(new_n8644, new_n8643, new_n2036);
nor_4  g08259(new_n8645, new_n8644, new_n2035);
nor_4  g08260(new_n8646, new_n8645, new_n2034);
nor_4  g08261(new_n8647, new_n8646, new_n2033);
nor_4  g08262(new_n8648, new_n8647, new_n2032);
nor_4  g08263(new_n8649_1, new_n8648, new_n2031);
nor_4  g08264(new_n8650, new_n8649_1, new_n2030);
not_3  g08265(new_n8651, new_n8650);
nand_4 g08266(new_n8652, new_n8651, new_n856);
nand_4 g08267(new_n8653, new_n8652, new_n863);
nand_4 g08268(new_n8654, new_n8653, new_n419);
nand_4 g08269(new_n8655, new_n8654, new_n869);
nand_4 g08270(new_n8656, new_n8655, new_n875);
nand_4 g08271(new_n8657, new_n8656, new_n881);
nand_4 g08272(new_n8658, new_n8657, new_n413);
nand_4 g08273(new_n8659, new_n8658, new_n889);
nand_4 g08274(new_n8660, new_n8659, new_n896);
nand_4 g08275(new_n8661, new_n8660, new_n901);
nand_4 g08276(new_n8662, new_n8661, new_n408);
nand_4 g08277(new_n8663, new_n8662, new_n908);
nand_4 g08278(new_n8664, new_n8663, new_n403);
nand_4 g08279(new_n8665, new_n8664, new_n398);
nand_4 g08280(new_n8666, new_n8665, n8780);
nor_4  g08281(n8144, new_n8666, new_n389_1);
not_3  g08282(new_n8668, new_n962);
nand_4 g08283(new_n8669, new_n959, new_n486);
nand_4 g08284(new_n8670, new_n8669, new_n743);
nand_4 g08285(new_n8671, new_n8670, new_n482);
nand_4 g08286(new_n8672, new_n8671, new_n751);
nand_4 g08287(new_n8673, new_n8672, new_n758);
nand_4 g08288(new_n8674, new_n8673, new_n765);
nand_4 g08289(new_n8675, new_n8674, new_n476);
nand_4 g08290(new_n8676, new_n8675, new_n773);
nand_4 g08291(new_n8677, new_n8676, new_n780);
nand_4 g08292(new_n8678, new_n8677, new_n787);
nand_4 g08293(new_n8679, new_n8678, new_n470);
nand_4 g08294(new_n8680, new_n8679, new_n795);
nand_4 g08295(new_n8681, new_n8680, new_n803);
nand_4 g08296(new_n8682, new_n8681, new_n809);
nand_4 g08297(new_n8683, new_n8682, new_n465);
nand_4 g08298(new_n8684, new_n8683, new_n818);
nand_4 g08299(new_n8685, new_n8684, new_n460);
nand_4 g08300(new_n8686, new_n8685, new_n455);
nand_4 g08301(new_n8687, new_n8686, new_n449);
nand_4 g08302(new_n8688, new_n8687, new_n827);
nand_4 g08303(new_n8689, new_n8688, new_n833);
nand_4 g08304(new_n8690, new_n8689, new_n444);
nand_4 g08305(new_n8691, new_n8690, new_n439);
nand_4 g08306(new_n8692, new_n8691, new_n841);
nand_4 g08307(new_n8693, new_n8692, new_n434);
nand_4 g08308(new_n8694, new_n8693, new_n429);
nand_4 g08309(new_n8695, new_n8694, new_n424);
nand_4 g08310(new_n8696, new_n8695, new_n850);
nand_4 g08311(new_n8697, new_n8696, new_n856);
nand_4 g08312(new_n8698, new_n8697, new_n863);
nand_4 g08313(new_n8699, new_n8698, new_n419);
nand_4 g08314(new_n8700, new_n8699, new_n869);
nand_4 g08315(new_n8701, new_n8700, new_n875);
nand_4 g08316(new_n8702, new_n8701, new_n881);
nand_4 g08317(new_n8703, new_n8702, new_n413);
nand_4 g08318(new_n8704, new_n8703, new_n889);
nand_4 g08319(new_n8705, new_n8704, new_n896);
nand_4 g08320(new_n8706, new_n8705, new_n901);
nand_4 g08321(new_n8707, new_n8706, new_n408);
nand_4 g08322(new_n8708, new_n8707, new_n908);
nand_4 g08323(new_n8709, new_n8708, new_n403);
nand_4 g08324(new_n8710, new_n8709, new_n398);
nand_4 g08325(new_n8711, new_n8710, new_n393);
nand_4 g08326(new_n8712, new_n8711, new_n916);
nand_4 g08327(new_n8713, new_n8712, new_n1123);
nand_4 g08328(new_n8714, new_n8713, new_n1164);
nand_4 g08329(new_n8715, new_n8714, new_n1120);
nand_4 g08330(new_n8716, new_n8715, new_n1169);
nand_4 g08331(new_n8717, new_n8716, new_n1116);
nand_4 g08332(new_n8718, new_n8717, new_n1111);
nand_4 g08333(new_n8719, new_n8718, new_n1106);
not_3  g08334(new_n8720, new_n8719);
nor_4  g08335(new_n8721, new_n8720, new_n1525);
nor_4  g08336(new_n8722, new_n8721, new_n1524);
nor_4  g08337(new_n8723, new_n8722, new_n1523);
nor_4  g08338(new_n8724, new_n8723, new_n1522);
nor_4  g08339(new_n8725, new_n8724, new_n1521);
nor_4  g08340(new_n8726, new_n8725, new_n1520);
nor_4  g08341(new_n8727, new_n8726, new_n1519);
nor_4  g08342(new_n8728, new_n8727, new_n1518);
nor_4  g08343(new_n8729, new_n8728, new_n1517);
nor_4  g08344(new_n8730, new_n8729, new_n1516);
nor_4  g08345(new_n8731, new_n8730, new_n1075);
nor_4  g08346(new_n8732, new_n8731, new_n1071);
nor_4  g08347(new_n8733, new_n8732, new_n1065);
nor_4  g08348(new_n8734, new_n8733, new_n1062);
nor_4  g08349(new_n8735, new_n8734, new_n1056);
nor_4  g08350(new_n8736, new_n8735, new_n1051);
nor_4  g08351(new_n8737_1, new_n8736, new_n1046);
nor_4  g08352(new_n8738, new_n8737_1, new_n1042);
nor_4  g08353(new_n8739, new_n8738, new_n1037);
nor_4  g08354(new_n8740, new_n8739, new_n1032);
nor_4  g08355(new_n8741, new_n8740, new_n1026);
nor_4  g08356(new_n8742, new_n8741, new_n1021);
nor_4  g08357(new_n8743, new_n8742, new_n1016);
nor_4  g08358(new_n8744, new_n8743, new_n1011);
nor_4  g08359(new_n8745, new_n8744, new_n1216);
nor_4  g08360(new_n8746_1, new_n8745, new_n1006);
nor_4  g08361(new_n8747, new_n8746_1, new_n1001);
not_3  g08362(new_n8748, new_n8747);
nand_4 g08363(new_n8749, new_n8748, new_n994);
nand_4 g08364(new_n8750, new_n8749, new_n989);
nand_4 g08365(new_n8751, new_n8750, new_n984);
nand_4 g08366(new_n8752, new_n8751, new_n978);
nand_4 g08367(new_n8753, new_n8752, new_n973);
nand_4 g08368(new_n8754, new_n8753, new_n967);
nand_4 g08369(new_n8755, new_n8754, n10407);
nor_4  g08370(n8215, new_n8755, new_n8668);
not_3  g08371(new_n8757, n656);
not_3  g08372(new_n8758, new_n1331);
nand_4 g08373(new_n8759, new_n8758, new_n8757);
nand_4 g08374(new_n8760, new_n8759, new_n2181);
nand_4 g08375(new_n8761, new_n8760, new_n2179);
nand_4 g08376(new_n8762, new_n8761, new_n2175_1);
nand_4 g08377(new_n8763, new_n8762, new_n2171);
nand_4 g08378(new_n8764, new_n8763, new_n2168);
nand_4 g08379(new_n8765, new_n8764, new_n2165);
nand_4 g08380(new_n8766, new_n8765, new_n2162);
nand_4 g08381(new_n8767, new_n8766, new_n2158);
nand_4 g08382(new_n8768, new_n8767, new_n2155);
nand_4 g08383(new_n8769, new_n8768, new_n2151);
nand_4 g08384(new_n8770, new_n8769, new_n2147);
nand_4 g08385(new_n8771, new_n8770, new_n1810);
nand_4 g08386(new_n8772, new_n8771, new_n1806);
nand_4 g08387(new_n8773, new_n8772, new_n1802);
nand_4 g08388(new_n8774, new_n8773, new_n1798);
nand_4 g08389(new_n8775, new_n8774, new_n1820);
nand_4 g08390(new_n8776, new_n8775, new_n1794);
nand_4 g08391(new_n8777, new_n8776, new_n1825);
nand_4 g08392(new_n8778, new_n8777, new_n1789);
nand_4 g08393(new_n8779, new_n8778, new_n1785);
nand_4 g08394(new_n8780_1, new_n8779, new_n1780);
nand_4 g08395(new_n8781, new_n8780_1, new_n1777);
nand_4 g08396(new_n8782, new_n8781, new_n1774);
nand_4 g08397(new_n8783, new_n8782, new_n1834);
nand_4 g08398(new_n8784, new_n8783, new_n1769);
nand_4 g08399(new_n8785, new_n8784, new_n1766);
nand_4 g08400(new_n8786, new_n8785, new_n1762);
nand_4 g08401(new_n8787, new_n8786, new_n1758);
nand_4 g08402(new_n8788, new_n8787, new_n1754);
nand_4 g08403(new_n8789, new_n8788, new_n1751);
nand_4 g08404(new_n8790, new_n8789, new_n1748);
nand_4 g08405(new_n8791, new_n8790, new_n1746);
nand_4 g08406(new_n8792, new_n8791, new_n1742);
nand_4 g08407(new_n8793, new_n8792, new_n1738);
nand_4 g08408(new_n8794, new_n8793, new_n1736);
nand_4 g08409(new_n8795, new_n8794, new_n1732);
nand_4 g08410(new_n8796, new_n8795, new_n1729);
nand_4 g08411(new_n8797, new_n8796, new_n1726);
nand_4 g08412(new_n8798, new_n8797, new_n1724);
nand_4 g08413(new_n8799_1, new_n8798, new_n1721);
nand_4 g08414(new_n8800_1, new_n8799_1, new_n1718);
nand_4 g08415(new_n8801, new_n8800_1, new_n1715);
nand_4 g08416(new_n8802, new_n8801, new_n1711);
nand_4 g08417(new_n8803, new_n8802, new_n1708);
nand_4 g08418(new_n8804, new_n8803, new_n1705);
nand_4 g08419(new_n8805, new_n8804, new_n1703);
nand_4 g08420(new_n8806, new_n8805, new_n1860);
nand_4 g08421(new_n8807, new_n8806, new_n1864);
nand_4 g08422(new_n8808, new_n8807, new_n1699);
nand_4 g08423(new_n8809, new_n8808, new_n1697);
not_3  g08424(new_n8810, new_n8809);
nor_4  g08425(new_n8811, new_n8810, new_n2133);
nor_4  g08426(new_n8812, new_n8811, new_n2132);
nor_4  g08427(new_n8813, new_n8812, new_n1691);
nor_4  g08428(new_n8814, new_n8813, new_n1879);
nor_4  g08429(new_n8815, new_n8814, new_n1883);
nor_4  g08430(new_n8816, new_n8815, new_n1687);
nor_4  g08431(new_n8817, new_n8816, new_n1683);
nor_4  g08432(new_n8818, new_n8817, new_n1679);
nor_4  g08433(new_n8819, new_n8818, new_n1675);
nor_4  g08434(new_n8820, new_n8819, new_n1891);
nor_4  g08435(new_n8821, new_n8820, new_n1670);
nor_4  g08436(new_n8822, new_n8821, new_n1666);
nor_4  g08437(new_n8823, new_n8822, new_n1662);
nor_4  g08438(new_n8824, new_n8823, new_n1658);
nor_4  g08439(new_n8825, new_n8824, new_n1653);
nor_4  g08440(new_n8826, new_n8825, new_n1649);
nor_4  g08441(new_n8827, new_n8826, new_n1645);
nor_4  g08442(new_n8828, new_n8827, new_n1641);
nor_4  g08443(new_n8829, new_n8828, new_n1637_1);
nor_4  g08444(new_n8830, new_n8829, new_n1633);
nor_4  g08445(new_n8831, new_n8830, new_n1629);
nor_4  g08446(new_n8832, new_n8831, new_n1628);
nor_4  g08447(new_n8833, new_n8832, new_n1627);
nor_4  g08448(new_n8834, new_n8833, new_n1626);
nor_4  g08449(new_n8835, new_n8834, new_n4700);
not_3  g08450(new_n8836, new_n8835);
nand_4 g08451(new_n8837, new_n8836, new_n1357);
nand_4 g08452(new_n8838, new_n8837, new_n1354);
nand_4 g08453(new_n8839, new_n8838, new_n1352);
nand_4 g08454(new_n8840, new_n8839, new_n1350);
nand_4 g08455(new_n8841, new_n8840, new_n1347_1);
nand_4 g08456(new_n8842, new_n8841, new_n1344);
nand_4 g08457(new_n8843, new_n8842, new_n1341);
nand_4 g08458(new_n8844, new_n8843, new_n1338);
nand_4 g08459(new_n8845, new_n8844, new_n1395);
nand_4 g08460(new_n8846, new_n8845, n1093);
nor_4  g08461(n8306, new_n8846, new_n792);
nand_4 g08462(new_n8848, new_n1342, new_n772);
nand_4 g08463(new_n8849, new_n8848, new_n1341);
nand_4 g08464(new_n8850, new_n8849, new_n1338);
nand_4 g08465(new_n8851, new_n8850, new_n1395);
nand_4 g08466(new_n8852, new_n8851, new_n1335);
nand_4 g08467(new_n8853, new_n8852, new_n1332);
nand_4 g08468(new_n8854, new_n8853, new_n1328);
nand_4 g08469(new_n8855, new_n8854, new_n1403);
nand_4 g08470(new_n8856, new_n8855, new_n1325);
nand_4 g08471(new_n8857, new_n8856, new_n1410);
nand_4 g08472(new_n8858, new_n8857, new_n1413);
nand_4 g08473(new_n8859, new_n8858, new_n1322);
nand_4 g08474(new_n8860, new_n8859, new_n1317);
nand_4 g08475(new_n8861, new_n8860, new_n1315);
nand_4 g08476(new_n8862, new_n8861, new_n1419);
nand_4 g08477(new_n8863, new_n8862, new_n1310);
nand_4 g08478(new_n8864, new_n8863, new_n1305);
nand_4 g08479(new_n8865, new_n8864, new_n1427);
nand_4 g08480(new_n8866, new_n8865, new_n1431);
nand_4 g08481(new_n8867, new_n8866, new_n1302);
nand_4 g08482(new_n8868, new_n8867, new_n1298);
nand_4 g08483(new_n8869, new_n8868, new_n1295);
nand_4 g08484(new_n8870, new_n8869, new_n1291);
nand_4 g08485(new_n8871, new_n8870, new_n1288);
nand_4 g08486(new_n8872, new_n8871, new_n1284);
nand_4 g08487(new_n8873_1, new_n8872, new_n1280);
nand_4 g08488(new_n8874, new_n8873_1, new_n1275);
nand_4 g08489(new_n8875, new_n8874, new_n1445);
nand_4 g08490(new_n8876, new_n8875, new_n1270);
nand_4 g08491(new_n8877, new_n8876, new_n1265_1);
nand_4 g08492(new_n8878, new_n8877, new_n1260);
nand_4 g08493(new_n8879, new_n8878, new_n1256);
nand_4 g08494(new_n8880, new_n8879, new_n1251);
nand_4 g08495(new_n8881, new_n8880, new_n1457);
nand_4 g08496(new_n8882, new_n8881, new_n1462);
nand_4 g08497(new_n8883, new_n8882, new_n1468);
nand_4 g08498(new_n8884, new_n8883, new_n1247);
nand_4 g08499(new_n8885, new_n8884, new_n1474);
nand_4 g08500(new_n8886, new_n8885, new_n592);
nand_4 g08501(new_n8887, new_n8886, new_n585);
nand_4 g08502(new_n8888, new_n8887, new_n580);
nand_4 g08503(new_n8889, new_n8888, new_n600);
nand_4 g08504(new_n8890, new_n8889, new_n606);
nand_4 g08505(new_n8891, new_n8890, new_n612);
nand_4 g08506(new_n8892_1, new_n8891, new_n575);
nand_4 g08507(new_n8893, new_n8892_1, new_n619);
nand_4 g08508(new_n8894, new_n8893, new_n570);
nand_4 g08509(new_n8895, new_n8894, new_n625);
nand_4 g08510(new_n8896, new_n8895, new_n564);
nand_4 g08511(new_n8897, new_n8896, new_n632);
nand_4 g08512(new_n8898, new_n8897, new_n638);
not_3  g08513(new_n8899, new_n8898);
nor_4  g08514(new_n8900, new_n8899, new_n3075);
nor_4  g08515(new_n8901, new_n8900, new_n3074);
nor_4  g08516(new_n8902, new_n8901, new_n3073);
nor_4  g08517(new_n8903, new_n8902, new_n3072);
nor_4  g08518(new_n8904, new_n8903, new_n3071);
nor_4  g08519(new_n8905, new_n8904, new_n3070);
nor_4  g08520(new_n8906, new_n8905, new_n3069);
nor_4  g08521(new_n8907, new_n8906, new_n3068);
nor_4  g08522(new_n8908, new_n8907, new_n3067);
nor_4  g08523(new_n8909_1, new_n8908, new_n3066);
nor_4  g08524(new_n8910, new_n8909_1, new_n3065);
nor_4  g08525(new_n8911, new_n8910, new_n3064);
nor_4  g08526(new_n8912, new_n8911, new_n3063);
nor_4  g08527(new_n8913, new_n8912, new_n3062);
nor_4  g08528(new_n8914, new_n8913, new_n3061);
nor_4  g08529(new_n8915, new_n8914, new_n3354);
nor_4  g08530(new_n8916, new_n8915, new_n3353);
nor_4  g08531(new_n8917, new_n8916, new_n3352);
nor_4  g08532(new_n8918, new_n8917, new_n3351);
nor_4  g08533(new_n8919, new_n8918, new_n3350);
nor_4  g08534(new_n8920, new_n8919, new_n3349);
nor_4  g08535(new_n8921, new_n8920, new_n3348);
nor_4  g08536(new_n8922, new_n8921, new_n720);
nor_4  g08537(new_n8923, new_n8922, new_n501);
nor_4  g08538(new_n8924, new_n8923, new_n728);
nor_4  g08539(new_n8925, new_n8924, new_n495);
nor_4  g08540(new_n8926_1, new_n8925, new_n736);
not_3  g08541(new_n8927, new_n8926_1);
nand_4 g08542(new_n8928, new_n8927, new_n488);
nand_4 g08543(new_n8929, new_n8928, new_n743);
nand_4 g08544(new_n8930, new_n8929, new_n482);
nand_4 g08545(new_n8931, new_n8930, new_n751);
nand_4 g08546(new_n8932, new_n8931, new_n758);
nand_4 g08547(new_n8933, new_n8932, new_n765);
nand_4 g08548(new_n8934, new_n8933, n9544);
nor_4  g08549(n8471, new_n8934, new_n473);
nand_4 g08550(new_n8936, new_n2160, new_n1321);
nand_4 g08551(new_n8937, new_n8936, new_n2158);
nand_4 g08552(new_n8938, new_n8937, new_n2155);
nand_4 g08553(new_n8939, new_n8938, new_n2151);
nand_4 g08554(new_n8940, new_n8939, new_n2147);
nand_4 g08555(new_n8941, new_n8940, new_n1810);
nand_4 g08556(new_n8942, new_n8941, new_n1806);
nand_4 g08557(new_n8943, new_n8942, new_n1802);
nand_4 g08558(new_n8944, new_n8943, new_n1798);
nand_4 g08559(new_n8945, new_n8944, new_n1820);
nand_4 g08560(new_n8946, new_n8945, new_n1794);
nand_4 g08561(new_n8947, new_n8946, new_n1825);
nand_4 g08562(new_n8948, new_n8947, new_n1789);
nand_4 g08563(new_n8949, new_n8948, new_n1785);
nand_4 g08564(new_n8950, new_n8949, new_n1780);
nand_4 g08565(new_n8951, new_n8950, new_n1777);
nand_4 g08566(new_n8952, new_n8951, new_n1774);
nand_4 g08567(new_n8953, new_n8952, new_n1834);
nand_4 g08568(new_n8954, new_n8953, new_n1769);
nand_4 g08569(new_n8955, new_n8954, new_n1766);
nand_4 g08570(new_n8956, new_n8955, new_n1762);
nand_4 g08571(new_n8957, new_n8956, new_n1758);
nand_4 g08572(new_n8958, new_n8957, new_n1754);
nand_4 g08573(new_n8959, new_n8958, new_n1751);
nand_4 g08574(new_n8960, new_n8959, new_n1748);
nand_4 g08575(new_n8961, new_n8960, new_n1746);
nand_4 g08576(new_n8962, new_n8961, new_n1742);
nand_4 g08577(new_n8963, new_n8962, new_n1738);
nand_4 g08578(new_n8964, new_n8963, new_n1736);
nand_4 g08579(new_n8965, new_n8964, new_n1732);
nand_4 g08580(new_n8966, new_n8965, new_n1729);
nand_4 g08581(new_n8967, new_n8966, new_n1726);
nand_4 g08582(new_n8968, new_n8967, new_n1724);
nand_4 g08583(new_n8969, new_n8968, new_n1721);
nand_4 g08584(new_n8970, new_n8969, new_n1718);
nand_4 g08585(new_n8971, new_n8970, new_n1715);
nand_4 g08586(new_n8972, new_n8971, new_n1711);
nand_4 g08587(new_n8973, new_n8972, new_n1708);
nand_4 g08588(new_n8974, new_n8973, new_n1705);
nand_4 g08589(new_n8975, new_n8974, new_n1703);
nand_4 g08590(new_n8976, new_n8975, new_n1860);
nand_4 g08591(new_n8977, new_n8976, new_n1864);
nand_4 g08592(new_n8978, new_n8977, new_n1699);
nand_4 g08593(new_n8979, new_n8978, new_n1697);
nand_4 g08594(new_n8980, new_n8979, new_n1871);
not_3  g08595(new_n8981, new_n8980);
nor_4  g08596(new_n8982, new_n8981, new_n2132);
nor_4  g08597(new_n8983, new_n8982, new_n1691);
nor_4  g08598(new_n8984, new_n8983, new_n1879);
nor_4  g08599(new_n8985, new_n8984, new_n1883);
nor_4  g08600(new_n8986, new_n8985, new_n1687);
nor_4  g08601(new_n8987, new_n8986, new_n1683);
nor_4  g08602(new_n8988, new_n8987, new_n1679);
nor_4  g08603(new_n8989, new_n8988, new_n1675);
nor_4  g08604(new_n8990, new_n8989, new_n1891);
nor_4  g08605(new_n8991, new_n8990, new_n1670);
nor_4  g08606(new_n8992, new_n8991, new_n1666);
nor_4  g08607(new_n8993, new_n8992, new_n1662);
nor_4  g08608(new_n8994, new_n8993, new_n1658);
nor_4  g08609(new_n8995, new_n8994, new_n1653);
nor_4  g08610(new_n8996, new_n8995, new_n1649);
nor_4  g08611(new_n8997_1, new_n8996, new_n1645);
nor_4  g08612(new_n8998, new_n8997_1, new_n1641);
nor_4  g08613(new_n8999, new_n8998, new_n1637_1);
nor_4  g08614(new_n9000, new_n8999, new_n1633);
nor_4  g08615(new_n9001, new_n9000, new_n1629);
nor_4  g08616(new_n9002, new_n9001, new_n1628);
nor_4  g08617(new_n9003, new_n9002, new_n1627);
nor_4  g08618(new_n9004, new_n9003, new_n1626);
nor_4  g08619(new_n9005, new_n9004, new_n4700);
not_3  g08620(new_n9006, new_n9005);
nand_4 g08621(new_n9007, new_n9006, new_n1357);
nand_4 g08622(new_n9008, new_n9007, new_n1354);
nand_4 g08623(new_n9009, new_n9008, new_n1352);
nand_4 g08624(new_n9010, new_n9009, new_n1350);
nand_4 g08625(new_n9011, new_n9010, new_n1347_1);
nand_4 g08626(new_n9012, new_n9011, new_n1344);
nand_4 g08627(new_n9013, new_n9012, new_n1341);
nand_4 g08628(new_n9014, new_n9013, new_n1338);
nand_4 g08629(new_n9015, new_n9014, new_n1395);
nand_4 g08630(new_n9016, new_n9015, new_n1335);
nand_4 g08631(new_n9017, new_n9016, new_n1332);
nand_4 g08632(new_n9018, new_n9017, new_n1328);
nand_4 g08633(new_n9019, new_n9018, new_n1403);
nand_4 g08634(new_n9020, new_n9019, new_n1325);
nand_4 g08635(new_n9021, new_n9020, new_n1410);
nand_4 g08636(new_n9022, new_n9021, n5786);
nor_4  g08637(n8604, new_n9022, new_n453);
nand_4 g08638(new_n9024, new_n2157, new_n831);
nand_4 g08639(new_n9025, new_n9024, new_n444);
nand_4 g08640(new_n9026_1, new_n9025, new_n439);
nand_4 g08641(new_n9027, new_n9026_1, new_n841);
nand_4 g08642(new_n9028, new_n9027, new_n434);
nand_4 g08643(new_n9029, new_n9028, new_n429);
nand_4 g08644(new_n9030, new_n9029, new_n424);
nand_4 g08645(new_n9031, new_n9030, new_n850);
nand_4 g08646(new_n9032, new_n9031, new_n856);
nand_4 g08647(new_n9033, new_n9032, new_n863);
nand_4 g08648(new_n9034, new_n9033, new_n419);
nand_4 g08649(new_n9035, new_n9034, new_n869);
nand_4 g08650(new_n9036, new_n9035, new_n875);
nand_4 g08651(new_n9037, new_n9036, new_n881);
nand_4 g08652(new_n9038, new_n9037, new_n413);
nand_4 g08653(new_n9039, new_n9038, new_n889);
nand_4 g08654(new_n9040, new_n9039, new_n896);
nand_4 g08655(new_n9041, new_n9040, new_n901);
nand_4 g08656(new_n9042, new_n9041, new_n408);
nand_4 g08657(new_n9043, new_n9042, new_n908);
nand_4 g08658(new_n9044, new_n9043, new_n403);
nand_4 g08659(new_n9045, new_n9044, new_n398);
nand_4 g08660(new_n9046, new_n9045, new_n393);
nand_4 g08661(new_n9047, new_n9046, new_n916);
nand_4 g08662(new_n9048, new_n9047, new_n1123);
nand_4 g08663(new_n9049, new_n9048, new_n1164);
nand_4 g08664(new_n9050, new_n9049, new_n1120);
nand_4 g08665(new_n9051, new_n9050, new_n1169);
nand_4 g08666(new_n9052, new_n9051, new_n1116);
nand_4 g08667(new_n9053, new_n9052, new_n1111);
nand_4 g08668(new_n9054, new_n9053, new_n1106);
nand_4 g08669(new_n9055, new_n9054, new_n1178);
nand_4 g08670(new_n9056, new_n9055, new_n1183);
nand_4 g08671(new_n9057, new_n9056, new_n1102);
nand_4 g08672(new_n9058, new_n9057, new_n1099);
nand_4 g08673(new_n9059, new_n9058, new_n1191);
nand_4 g08674(new_n9060, new_n9059, new_n1095);
nand_4 g08675(new_n9061, new_n9060, new_n1091);
nand_4 g08676(new_n9062, new_n9061, new_n1088);
nand_4 g08677(new_n9063, new_n9062, new_n1084);
nand_4 g08678(new_n9064, new_n9063, new_n1079);
nand_4 g08679(new_n9065, new_n9064, new_n1074);
nand_4 g08680(new_n9066, new_n9065, new_n1070);
nand_4 g08681(new_n9067, new_n9066, new_n1064);
nand_4 g08682(new_n9068, new_n9067, new_n1061);
nand_4 g08683(new_n9069, new_n9068, new_n1055);
nand_4 g08684(new_n9070, new_n9069, new_n1050);
nand_4 g08685(new_n9071, new_n9070, new_n1045);
nand_4 g08686(new_n9072, new_n9071, new_n1041);
nand_4 g08687(new_n9073, new_n9072, new_n1036);
nand_4 g08688(new_n9074, new_n9073, new_n1031);
not_3  g08689(new_n9075, new_n9074);
nor_4  g08690(new_n9076, new_n9075, new_n1026);
nor_4  g08691(new_n9077, new_n9076, new_n1021);
nor_4  g08692(new_n9078, new_n9077, new_n1016);
nor_4  g08693(new_n9079, new_n9078, new_n1011);
nor_4  g08694(new_n9080, new_n9079, new_n1216);
nor_4  g08695(new_n9081, new_n9080, new_n1006);
nor_4  g08696(new_n9082, new_n9081, new_n1001);
nor_4  g08697(new_n9083, new_n9082, new_n995);
nor_4  g08698(new_n9084, new_n9083, new_n990);
nor_4  g08699(new_n9085, new_n9084, new_n985);
nor_4  g08700(new_n9086, new_n9085, new_n979);
nor_4  g08701(new_n9087, new_n9086, new_n974);
nor_4  g08702(new_n9088, new_n9087, new_n968);
nor_4  g08703(new_n9089, new_n9088, new_n965);
nor_4  g08704(new_n9090, new_n9089, new_n961);
nor_4  g08705(new_n9091, new_n9090, new_n958);
nor_4  g08706(new_n9092, new_n9091, new_n953);
nor_4  g08707(new_n9093, new_n9092, new_n3536);
nor_4  g08708(new_n9094, new_n9093, new_n3535);
nor_4  g08709(new_n9095, new_n9094, new_n3534);
nor_4  g08710(new_n9096_1, new_n9095, new_n2520);
nor_4  g08711(new_n9097, new_n9096_1, new_n2519);
nor_4  g08712(new_n9098, new_n9097, new_n2518);
nor_4  g08713(new_n9099, new_n9098, new_n2517);
nor_4  g08714(new_n9100, new_n9099, new_n2516);
nor_4  g08715(new_n9101, new_n9100, new_n2515);
nor_4  g08716(new_n9102, new_n9101, new_n2514);
not_3  g08717(new_n9103, new_n9102);
nand_4 g08718(new_n9104, new_n9103, new_n2183);
nand_4 g08719(new_n9105, new_n9104, new_n2179);
nand_4 g08720(new_n9106, new_n9105, new_n2175_1);
nand_4 g08721(new_n9107, new_n9106, new_n2171);
nand_4 g08722(new_n9108, new_n9107, new_n2168);
nand_4 g08723(new_n9109, new_n9108, new_n2165);
nand_4 g08724(new_n9110_1, new_n9109, n9589);
nor_4  g08725(n8909, new_n9110_1, new_n2159);
not_3  g08726(new_n9112, new_n532);
nand_4 g08727(new_n9113, new_n1882, new_n9112);
nand_4 g08728(new_n9114, new_n9113, new_n1686);
nand_4 g08729(new_n9115, new_n9114, new_n1682);
nand_4 g08730(new_n9116, new_n9115, new_n1678);
nand_4 g08731(new_n9117, new_n9116, new_n1674);
nand_4 g08732(new_n9118, new_n9117, new_n1890);
nand_4 g08733(new_n9119, new_n9118, new_n1669);
nand_4 g08734(new_n9120, new_n9119, new_n1665);
nand_4 g08735(new_n9121, new_n9120, new_n1661);
nand_4 g08736(new_n9122, new_n9121, new_n1657);
nand_4 g08737(new_n9123, new_n9122, new_n1652);
nand_4 g08738(new_n9124, new_n9123, new_n1648);
nand_4 g08739(new_n9125, new_n9124, new_n1644);
nand_4 g08740(new_n9126, new_n9125, new_n1640);
nand_4 g08741(new_n9127, new_n9126, new_n1636);
nand_4 g08742(new_n9128, new_n9127, new_n1632);
nand_4 g08743(new_n9129, new_n9128, new_n1378);
nand_4 g08744(new_n9130, new_n9129, new_n1372);
nand_4 g08745(new_n9131, new_n9130, new_n1367);
nand_4 g08746(new_n9132, new_n9131, new_n1363);
nand_4 g08747(new_n9133, new_n9132, new_n1360);
nand_4 g08748(new_n9134, new_n9133, new_n1357);
nand_4 g08749(new_n9135, new_n9134, new_n1354);
nand_4 g08750(new_n9136, new_n9135, new_n1352);
nand_4 g08751(new_n9137, new_n9136, new_n1350);
nand_4 g08752(new_n9138, new_n9137, new_n1347_1);
nand_4 g08753(new_n9139, new_n9138, new_n1344);
nand_4 g08754(new_n9140, new_n9139, new_n1341);
nand_4 g08755(new_n9141, new_n9140, new_n1338);
nand_4 g08756(new_n9142, new_n9141, new_n1395);
nand_4 g08757(new_n9143, new_n9142, new_n1335);
nand_4 g08758(new_n9144, new_n9143, new_n1332);
nand_4 g08759(new_n9145, new_n9144, new_n1328);
nand_4 g08760(new_n9146, new_n9145, new_n1403);
nand_4 g08761(new_n9147, new_n9146, new_n1325);
nand_4 g08762(new_n9148, new_n9147, new_n1410);
nand_4 g08763(new_n9149, new_n9148, new_n1413);
nand_4 g08764(new_n9150, new_n9149, new_n1322);
nand_4 g08765(new_n9151, new_n9150, new_n1317);
nand_4 g08766(new_n9152, new_n9151, new_n1315);
nand_4 g08767(new_n9153, new_n9152, new_n1419);
nand_4 g08768(new_n9154_1, new_n9153, new_n1310);
nand_4 g08769(new_n9155, new_n9154_1, new_n1305);
nand_4 g08770(new_n9156, new_n9155, new_n1427);
nand_4 g08771(new_n9157, new_n9156, new_n1431);
nand_4 g08772(new_n9158, new_n9157, new_n1302);
nand_4 g08773(new_n9159, new_n9158, new_n1298);
nand_4 g08774(new_n9160, new_n9159, new_n1295);
nand_4 g08775(new_n9161, new_n9160, new_n1291);
nand_4 g08776(new_n9162, new_n9161, new_n1288);
nand_4 g08777(new_n9163, new_n9162, new_n1284);
not_3  g08778(new_n9164, new_n9163);
nor_4  g08779(new_n9165, new_n9164, new_n1281);
nor_4  g08780(new_n9166, new_n9165, new_n1276);
nor_4  g08781(new_n9167, new_n9166, new_n1446);
nor_4  g08782(new_n9168, new_n9167, new_n1271);
nor_4  g08783(new_n9169, new_n9168, new_n1266);
nor_4  g08784(new_n9170, new_n9169, new_n1261);
nor_4  g08785(new_n9171, new_n9170, new_n1257);
nor_4  g08786(new_n9172, new_n9171, new_n1252);
nor_4  g08787(new_n9173, new_n9172, new_n1458);
nor_4  g08788(new_n9174, new_n9173, new_n1463);
nor_4  g08789(new_n9175, new_n9174, new_n1469);
nor_4  g08790(new_n9176, new_n9175, new_n1248);
nor_4  g08791(new_n9177, new_n9176, new_n1475);
nor_4  g08792(new_n9178, new_n9177, new_n1244);
nor_4  g08793(new_n9179, new_n9178, new_n1243);
nor_4  g08794(new_n9180, new_n9179, new_n1242);
nor_4  g08795(new_n9181, new_n9180, new_n1241);
nor_4  g08796(new_n9182, new_n9181, new_n1240);
nor_4  g08797(new_n9183, new_n9182, new_n1239);
nor_4  g08798(new_n9184, new_n9183, new_n3082);
nor_4  g08799(new_n9185, new_n9184, new_n3081);
nor_4  g08800(new_n9186_1, new_n9185, new_n3080);
nor_4  g08801(new_n9187, new_n9186_1, new_n3079);
nor_4  g08802(new_n9188, new_n9187, new_n3078);
nor_4  g08803(new_n9189, new_n9188, new_n3077);
nor_4  g08804(new_n9190, new_n9189, new_n3076);
nor_4  g08805(new_n9191, new_n9190, new_n3075);
not_3  g08806(new_n9192, new_n9191);
nand_4 g08807(new_n9193, new_n9192, new_n554);
nand_4 g08808(new_n9194, new_n9193, new_n646);
nand_4 g08809(new_n9195, new_n9194, new_n652);
nand_4 g08810(new_n9196, new_n9195, new_n549);
nand_4 g08811(new_n9197, new_n9196, new_n544);
nand_4 g08812(new_n9198, new_n9197, new_n660);
nand_4 g08813(new_n9199, new_n9198, n6680);
nor_4  g08814(n9096, new_n9199, new_n536);
not_3  g08815(new_n9201, new_n1444);
nand_4 g08816(new_n9202, new_n9201, new_n887);
nand_4 g08817(new_n9203, new_n9202, new_n1772);
nand_4 g08818(new_n9204, new_n9203, new_n1834);
nand_4 g08819(new_n9205, new_n9204, new_n1769);
nand_4 g08820(new_n9206, new_n9205, new_n1766);
nand_4 g08821(new_n9207, new_n9206, new_n1762);
nand_4 g08822(new_n9208, new_n9207, new_n1758);
nand_4 g08823(new_n9209, new_n9208, new_n1754);
nand_4 g08824(new_n9210, new_n9209, new_n1751);
nand_4 g08825(new_n9211, new_n9210, new_n1748);
nand_4 g08826(new_n9212, new_n9211, new_n1746);
nand_4 g08827(new_n9213, new_n9212, new_n1742);
nand_4 g08828(new_n9214, new_n9213, new_n1738);
nand_4 g08829(new_n9215, new_n9214, new_n1736);
nand_4 g08830(new_n9216, new_n9215, new_n1732);
nand_4 g08831(new_n9217, new_n9216, new_n1729);
nand_4 g08832(new_n9218, new_n9217, new_n1726);
nand_4 g08833(new_n9219, new_n9218, new_n1724);
nand_4 g08834(new_n9220, new_n9219, new_n1721);
nand_4 g08835(new_n9221, new_n9220, new_n1718);
nand_4 g08836(new_n9222, new_n9221, new_n1715);
nand_4 g08837(new_n9223, new_n9222, new_n1711);
nand_4 g08838(new_n9224, new_n9223, new_n1708);
nand_4 g08839(new_n9225, new_n9224, new_n1705);
nand_4 g08840(new_n9226, new_n9225, new_n1703);
nand_4 g08841(new_n9227, new_n9226, new_n1860);
nand_4 g08842(new_n9228, new_n9227, new_n1864);
nand_4 g08843(new_n9229, new_n9228, new_n1699);
nand_4 g08844(new_n9230, new_n9229, new_n1697);
nand_4 g08845(new_n9231, new_n9230, new_n1871);
nand_4 g08846(new_n9232, new_n9231, new_n1694);
nand_4 g08847(new_n9233, new_n9232, new_n1690);
nand_4 g08848(new_n9234, new_n9233, new_n1878);
nand_4 g08849(new_n9235, new_n9234, new_n1882);
nand_4 g08850(new_n9236, new_n9235, new_n1686);
nand_4 g08851(new_n9237, new_n9236, new_n1682);
nand_4 g08852(new_n9238, new_n9237, new_n1678);
nand_4 g08853(new_n9239, new_n9238, new_n1674);
nand_4 g08854(new_n9240, new_n9239, new_n1890);
nand_4 g08855(new_n9241, new_n9240, new_n1669);
nand_4 g08856(new_n9242, new_n9241, new_n1665);
nand_4 g08857(new_n9243, new_n9242, new_n1661);
nand_4 g08858(new_n9244, new_n9243, new_n1657);
nand_4 g08859(new_n9245, new_n9244, new_n1652);
nand_4 g08860(new_n9246, new_n9245, new_n1648);
nand_4 g08861(new_n9247, new_n9246, new_n1644);
nand_4 g08862(new_n9248, new_n9247, new_n1640);
nand_4 g08863(new_n9249, new_n9248, new_n1636);
nand_4 g08864(new_n9250, new_n9249, new_n1632);
nand_4 g08865(new_n9251, new_n9250, new_n1378);
nand_4 g08866(new_n9252_1, new_n9251, new_n1372);
not_3  g08867(new_n9253, new_n9252_1);
nor_4  g08868(new_n9254, new_n9253, new_n1627);
nor_4  g08869(new_n9255, new_n9254, new_n1626);
nor_4  g08870(new_n9256, new_n9255, new_n4700);
nor_4  g08871(new_n9257, new_n9256, new_n4699);
nor_4  g08872(new_n9258, new_n9257, new_n3722);
nor_4  g08873(new_n9259, new_n9258, new_n3721);
nor_4  g08874(new_n9260, new_n9259, new_n3720);
nor_4  g08875(new_n9261, new_n9260, new_n3719);
nor_4  g08876(new_n9262, new_n9261, new_n3718);
nor_4  g08877(new_n9263, new_n9262, new_n3717);
nor_4  g08878(new_n9264, new_n9263, new_n3716);
nor_4  g08879(new_n9265, new_n9264, new_n2611);
nor_4  g08880(new_n9266, new_n9265, new_n2610);
nor_4  g08881(new_n9267, new_n9266, new_n2609);
nor_4  g08882(new_n9268, new_n9267, new_n2413);
nor_4  g08883(new_n9269, new_n9268, new_n2412);
nor_4  g08884(new_n9270, new_n9269, new_n2411);
nor_4  g08885(new_n9271, new_n9270, new_n2410);
nor_4  g08886(new_n9272, new_n9271, new_n2409);
nor_4  g08887(new_n9273, new_n9272, new_n2408);
nor_4  g08888(new_n9274, new_n9273, new_n2407_1);
nor_4  g08889(new_n9275, new_n9274, new_n2406);
nor_4  g08890(new_n9276, new_n9275, new_n2405);
nor_4  g08891(new_n9277, new_n9276, new_n2404);
nor_4  g08892(new_n9278, new_n9277, new_n2403);
not_3  g08893(new_n9279, new_n9278);
nand_4 g08894(new_n9280, new_n9279, new_n1427);
nand_4 g08895(new_n9281, new_n9280, new_n1431);
nand_4 g08896(new_n9282, new_n9281, new_n1302);
nand_4 g08897(new_n9283, new_n9282, new_n1298);
nand_4 g08898(new_n9284, new_n9283, new_n1295);
nand_4 g08899(new_n9285, new_n9284, new_n1291);
nand_4 g08900(new_n9286, new_n9285, new_n1288);
nand_4 g08901(new_n9287, new_n9286, new_n1284);
nand_4 g08902(new_n9288, new_n9287, new_n1280);
nand_4 g08903(new_n9289, new_n9288, n8439);
nor_4  g08904(n9342, new_n9289, new_n1272);
not_3  g08905(new_n9291, new_n680);
nand_4 g08906(new_n9292, new_n9291, new_n676);
nand_4 g08907(new_n9293, new_n9292, new_n1672);
nand_4 g08908(new_n9294, new_n9293, new_n1890);
nand_4 g08909(new_n9295, new_n9294, new_n1669);
nand_4 g08910(new_n9296, new_n9295, new_n1665);
nand_4 g08911(new_n9297, new_n9296, new_n1661);
nand_4 g08912(new_n9298, new_n9297, new_n1657);
nand_4 g08913(new_n9299, new_n9298, new_n1652);
nand_4 g08914(new_n9300, new_n9299, new_n1648);
nand_4 g08915(new_n9301, new_n9300, new_n1644);
nand_4 g08916(new_n9302, new_n9301, new_n1640);
nand_4 g08917(new_n9303, new_n9302, new_n1636);
nand_4 g08918(new_n9304, new_n9303, new_n1632);
nand_4 g08919(new_n9305, new_n9304, new_n1378);
nand_4 g08920(new_n9306, new_n9305, new_n1372);
nand_4 g08921(new_n9307, new_n9306, new_n1367);
nand_4 g08922(new_n9308, new_n9307, new_n1363);
nand_4 g08923(new_n9309, new_n9308, new_n1360);
nand_4 g08924(new_n9310, new_n9309, new_n1357);
nand_4 g08925(new_n9311, new_n9310, new_n1354);
nand_4 g08926(new_n9312, new_n9311, new_n1352);
nand_4 g08927(new_n9313, new_n9312, new_n1350);
nand_4 g08928(new_n9314_1, new_n9313, new_n1347_1);
nand_4 g08929(new_n9315, new_n9314_1, new_n1344);
nand_4 g08930(new_n9316, new_n9315, new_n1341);
nand_4 g08931(new_n9317, new_n9316, new_n1338);
nand_4 g08932(new_n9318, new_n9317, new_n1395);
nand_4 g08933(new_n9319, new_n9318, new_n1335);
nand_4 g08934(new_n9320, new_n9319, new_n1332);
nand_4 g08935(new_n9321, new_n9320, new_n1328);
nand_4 g08936(new_n9322, new_n9321, new_n1403);
nand_4 g08937(new_n9323, new_n9322, new_n1325);
nand_4 g08938(new_n9324, new_n9323, new_n1410);
nand_4 g08939(new_n9325, new_n9324, new_n1413);
nand_4 g08940(new_n9326, new_n9325, new_n1322);
nand_4 g08941(new_n9327, new_n9326, new_n1317);
nand_4 g08942(new_n9328, new_n9327, new_n1315);
nand_4 g08943(new_n9329, new_n9328, new_n1419);
nand_4 g08944(new_n9330, new_n9329, new_n1310);
nand_4 g08945(new_n9331, new_n9330, new_n1305);
nand_4 g08946(new_n9332, new_n9331, new_n1427);
nand_4 g08947(new_n9333, new_n9332, new_n1431);
nand_4 g08948(new_n9334, new_n9333, new_n1302);
nand_4 g08949(new_n9335, new_n9334, new_n1298);
nand_4 g08950(new_n9336, new_n9335, new_n1295);
nand_4 g08951(new_n9337, new_n9336, new_n1291);
not_3  g08952(new_n9338, new_n9337);
nor_4  g08953(new_n9339, new_n9338, new_n2396);
nor_4  g08954(new_n9340, new_n9339, new_n2395);
nor_4  g08955(new_n9341, new_n9340, new_n1281);
nor_4  g08956(new_n9342_1, new_n9341, new_n1276);
nor_4  g08957(new_n9343, new_n9342_1, new_n1446);
nor_4  g08958(new_n9344, new_n9343, new_n1271);
nor_4  g08959(new_n9345, new_n9344, new_n1266);
nor_4  g08960(new_n9346, new_n9345, new_n1261);
nor_4  g08961(new_n9347, new_n9346, new_n1257);
nor_4  g08962(new_n9348, new_n9347, new_n1252);
nor_4  g08963(new_n9349, new_n9348, new_n1458);
nor_4  g08964(new_n9350, new_n9349, new_n1463);
nor_4  g08965(new_n9351, new_n9350, new_n1469);
nor_4  g08966(new_n9352, new_n9351, new_n1248);
nor_4  g08967(new_n9353, new_n9352, new_n1475);
nor_4  g08968(new_n9354, new_n9353, new_n1244);
nor_4  g08969(new_n9355, new_n9354, new_n1243);
nor_4  g08970(new_n9356, new_n9355, new_n1242);
nor_4  g08971(new_n9357, new_n9356, new_n1241);
nor_4  g08972(new_n9358, new_n9357, new_n1240);
nor_4  g08973(new_n9359, new_n9358, new_n1239);
nor_4  g08974(new_n9360, new_n9359, new_n3082);
nor_4  g08975(new_n9361, new_n9360, new_n3081);
nor_4  g08976(new_n9362, new_n9361, new_n3080);
not_3  g08977(new_n9363, new_n9362);
nand_4 g08978(new_n9364, new_n9363, new_n625);
nand_4 g08979(new_n9365, new_n9364, new_n564);
nand_4 g08980(new_n9366, new_n9365, new_n632);
nand_4 g08981(new_n9367, new_n9366, new_n638);
nand_4 g08982(new_n9368, new_n9367, new_n559);
nand_4 g08983(new_n9369, new_n9368, new_n554);
nand_4 g08984(new_n9370, new_n9369, new_n646);
nand_4 g08985(new_n9371, new_n9370, new_n652);
nand_4 g08986(new_n9372, new_n9371, new_n549);
nand_4 g08987(new_n9373, new_n9372, new_n544);
nand_4 g08988(new_n9374, new_n9373, new_n660);
nand_4 g08989(new_n9375, new_n9374, new_n539);
nand_4 g08990(new_n9376, new_n9375, new_n534);
nand_4 g08991(new_n9377, new_n9376, new_n529);
nand_4 g08992(new_n9378, new_n9377, new_n668);
nand_4 g08993(new_n9379, new_n9378, n12614);
nor_4  g08994(n9437, new_n9379, new_n671);
nand_4 g08995(new_n9381, new_n1778, new_n1279);
nand_4 g08996(new_n9382, new_n9381, new_n1777);
nand_4 g08997(new_n9383, new_n9382, new_n1774);
nand_4 g08998(new_n9384, new_n9383, new_n1834);
nand_4 g08999(new_n9385, new_n9384, new_n1769);
nand_4 g09000(new_n9386, new_n9385, new_n1766);
nand_4 g09001(new_n9387, new_n9386, new_n1762);
nand_4 g09002(new_n9388, new_n9387, new_n1758);
nand_4 g09003(new_n9389, new_n9388, new_n1754);
nand_4 g09004(new_n9390, new_n9389, new_n1751);
nand_4 g09005(new_n9391, new_n9390, new_n1748);
nand_4 g09006(new_n9392, new_n9391, new_n1746);
nand_4 g09007(new_n9393, new_n9392, new_n1742);
nand_4 g09008(new_n9394, new_n9393, new_n1738);
nand_4 g09009(new_n9395, new_n9394, new_n1736);
nand_4 g09010(new_n9396, new_n9395, new_n1732);
nand_4 g09011(new_n9397, new_n9396, new_n1729);
nand_4 g09012(new_n9398, new_n9397, new_n1726);
nand_4 g09013(new_n9399, new_n9398, new_n1724);
nand_4 g09014(new_n9400, new_n9399, new_n1721);
nand_4 g09015(new_n9401, new_n9400, new_n1718);
nand_4 g09016(new_n9402, new_n9401, new_n1715);
nand_4 g09017(new_n9403, new_n9402, new_n1711);
nand_4 g09018(new_n9404, new_n9403, new_n1708);
nand_4 g09019(new_n9405, new_n9404, new_n1705);
nand_4 g09020(new_n9406, new_n9405, new_n1703);
nand_4 g09021(new_n9407, new_n9406, new_n1860);
nand_4 g09022(new_n9408, new_n9407, new_n1864);
nand_4 g09023(new_n9409, new_n9408, new_n1699);
nand_4 g09024(new_n9410, new_n9409, new_n1697);
nand_4 g09025(new_n9411, new_n9410, new_n1871);
nand_4 g09026(new_n9412, new_n9411, new_n1694);
nand_4 g09027(new_n9413, new_n9412, new_n1690);
nand_4 g09028(new_n9414, new_n9413, new_n1878);
nand_4 g09029(new_n9415, new_n9414, new_n1882);
nand_4 g09030(new_n9416, new_n9415, new_n1686);
nand_4 g09031(new_n9417, new_n9416, new_n1682);
nand_4 g09032(new_n9418, new_n9417, new_n1678);
nand_4 g09033(new_n9419, new_n9418, new_n1674);
nand_4 g09034(new_n9420, new_n9419, new_n1890);
nand_4 g09035(new_n9421, new_n9420, new_n1669);
nand_4 g09036(new_n9422, new_n9421, new_n1665);
nand_4 g09037(new_n9423, new_n9422, new_n1661);
nand_4 g09038(new_n9424, new_n9423, new_n1657);
nand_4 g09039(new_n9425, new_n9424, new_n1652);
nand_4 g09040(new_n9426, new_n9425, new_n1648);
nand_4 g09041(new_n9427, new_n9426, new_n1644);
nand_4 g09042(new_n9428, new_n9427, new_n1640);
nand_4 g09043(new_n9429, new_n9428, new_n1636);
nand_4 g09044(new_n9430, new_n9429, new_n1632);
nand_4 g09045(new_n9431, new_n9430, new_n1378);
not_3  g09046(new_n9432, new_n9431);
nor_4  g09047(new_n9433, new_n9432, new_n1628);
nor_4  g09048(new_n9434, new_n9433, new_n1627);
nor_4  g09049(new_n9435, new_n9434, new_n1626);
nor_4  g09050(new_n9436, new_n9435, new_n4700);
nor_4  g09051(new_n9437_1, new_n9436, new_n4699);
nor_4  g09052(new_n9438, new_n9437_1, new_n3722);
nor_4  g09053(new_n9439, new_n9438, new_n3721);
nor_4  g09054(new_n9440, new_n9439, new_n3720);
nor_4  g09055(new_n9441, new_n9440, new_n3719);
nor_4  g09056(new_n9442, new_n9441, new_n3718);
nor_4  g09057(new_n9443, new_n9442, new_n3717);
nor_4  g09058(new_n9444, new_n9443, new_n3716);
nor_4  g09059(new_n9445, new_n9444, new_n2611);
nor_4  g09060(new_n9446, new_n9445, new_n2610);
nor_4  g09061(new_n9447_1, new_n9446, new_n2609);
nor_4  g09062(new_n9448, new_n9447_1, new_n2413);
nor_4  g09063(new_n9449, new_n9448, new_n2412);
nor_4  g09064(new_n9450, new_n9449, new_n2411);
nor_4  g09065(new_n9451, new_n9450, new_n2410);
nor_4  g09066(new_n9452, new_n9451, new_n2409);
nor_4  g09067(new_n9453, new_n9452, new_n2408);
nor_4  g09068(new_n9454, new_n9453, new_n2407_1);
nor_4  g09069(new_n9455, new_n9454, new_n2406);
nor_4  g09070(new_n9456, new_n9455, new_n2405);
nor_4  g09071(new_n9457, new_n9456, new_n2404);
nor_4  g09072(new_n9458, new_n9457, new_n2403);
nor_4  g09073(new_n9459, new_n9458, new_n2402);
not_3  g09074(new_n9460, new_n9459);
nand_4 g09075(new_n9461, new_n9460, new_n1431);
nand_4 g09076(new_n9462, new_n9461, new_n1302);
nand_4 g09077(new_n9463, new_n9462, new_n1298);
nand_4 g09078(new_n9464, new_n9463, new_n1295);
nand_4 g09079(new_n9465, new_n9464, new_n1291);
nand_4 g09080(new_n9466, new_n9465, new_n1288);
nand_4 g09081(new_n9467, new_n9466, n12782);
nor_4  g09082(n9447, new_n9467, new_n866);
not_3  g09083(new_n9469, new_n1100);
nand_4 g09084(new_n9470, new_n9469, new_n570);
nand_4 g09085(new_n9471, new_n9470, new_n625);
nand_4 g09086(new_n9472, new_n9471, new_n564);
nand_4 g09087(new_n9473, new_n9472, new_n632);
nand_4 g09088(new_n9474, new_n9473, new_n638);
nand_4 g09089(new_n9475, new_n9474, new_n559);
nand_4 g09090(new_n9476, new_n9475, new_n554);
nand_4 g09091(new_n9477, new_n9476, new_n646);
nand_4 g09092(new_n9478, new_n9477, new_n652);
nand_4 g09093(new_n9479, new_n9478, new_n549);
nand_4 g09094(new_n9480, new_n9479, new_n544);
nand_4 g09095(new_n9481, new_n9480, new_n660);
nand_4 g09096(new_n9482, new_n9481, new_n539);
nand_4 g09097(new_n9483, new_n9482, new_n534);
nand_4 g09098(new_n9484, new_n9483, new_n529);
nand_4 g09099(new_n9485, new_n9484, new_n668);
nand_4 g09100(new_n9486, new_n9485, new_n674_1);
nand_4 g09101(new_n9487, new_n9486, new_n681);
nand_4 g09102(new_n9488, new_n9487, new_n523);
nand_4 g09103(new_n9489, new_n9488, new_n687);
nand_4 g09104(new_n9490, new_n9489, new_n693);
nand_4 g09105(new_n9491, new_n9490, new_n699);
nand_4 g09106(new_n9492, new_n9491, new_n517);
nand_4 g09107(new_n9493, new_n9492, new_n705);
nand_4 g09108(new_n9494, new_n9493, new_n511);
nand_4 g09109(new_n9495, new_n9494, new_n711);
nand_4 g09110(new_n9496, new_n9495, new_n506);
nand_4 g09111(new_n9497, new_n9496, new_n719);
nand_4 g09112(new_n9498, new_n9497, new_n500);
nand_4 g09113(new_n9499, new_n9498, new_n727);
nand_4 g09114(new_n9500, new_n9499, new_n494);
nand_4 g09115(new_n9501, new_n9500, new_n735);
nand_4 g09116(new_n9502, new_n9501, new_n488);
nand_4 g09117(new_n9503, new_n9502, new_n743);
nand_4 g09118(new_n9504, new_n9503, new_n482);
nand_4 g09119(new_n9505, new_n9504, new_n751);
nand_4 g09120(new_n9506, new_n9505, new_n758);
nand_4 g09121(new_n9507, new_n9506, new_n765);
nand_4 g09122(new_n9508, new_n9507, new_n476);
nand_4 g09123(new_n9509, new_n9508, new_n773);
nand_4 g09124(new_n9510, new_n9509, new_n780);
nand_4 g09125(new_n9511, new_n9510, new_n787);
nand_4 g09126(new_n9512, new_n9511, new_n470);
nand_4 g09127(new_n9513, new_n9512, new_n795);
nand_4 g09128(new_n9514, new_n9513, new_n803);
nand_4 g09129(new_n9515, new_n9514, new_n809);
nand_4 g09130(new_n9516, new_n9515, new_n465);
nand_4 g09131(new_n9517, new_n9516, new_n818);
nand_4 g09132(new_n9518, new_n9517, new_n460);
nand_4 g09133(new_n9519, new_n9518, new_n455);
nand_4 g09134(new_n9520, new_n9519, new_n449);
not_3  g09135(new_n9521, new_n9520);
nor_4  g09136(new_n9522, new_n9521, new_n2038);
nor_4  g09137(new_n9523, new_n9522, new_n2037);
nor_4  g09138(new_n9524, new_n9523, new_n2036);
nor_4  g09139(new_n9525, new_n9524, new_n2035);
nor_4  g09140(new_n9526, new_n9525, new_n2034);
nor_4  g09141(new_n9527, new_n9526, new_n2033);
nor_4  g09142(new_n9528, new_n9527, new_n2032);
nor_4  g09143(new_n9529, new_n9528, new_n2031);
nor_4  g09144(new_n9530, new_n9529, new_n2030);
nor_4  g09145(new_n9531, new_n9530, new_n2029);
nor_4  g09146(new_n9532, new_n9531, new_n2028);
nor_4  g09147(new_n9533, new_n9532, new_n2027_1);
nor_4  g09148(new_n9534, new_n9533, new_n2026);
nor_4  g09149(new_n9535, new_n9534, new_n2025);
nor_4  g09150(new_n9536, new_n9535, new_n2024);
nor_4  g09151(new_n9537, new_n9536, new_n2023);
nor_4  g09152(new_n9538, new_n9537, new_n2022);
nor_4  g09153(new_n9539, new_n9538, new_n2021);
nor_4  g09154(new_n9540, new_n9539, new_n2020);
nor_4  g09155(new_n9541, new_n9540, new_n2019);
nor_4  g09156(new_n9542, new_n9541, new_n1537);
nor_4  g09157(new_n9543_1, new_n9542, new_n1536);
nor_4  g09158(new_n9544_1, new_n9543_1, new_n1535);
nor_4  g09159(new_n9545, new_n9544_1, new_n1534);
nor_4  g09160(new_n9546, new_n9545, new_n1533);
nor_4  g09161(new_n9547, new_n9546, new_n1532);
nor_4  g09162(new_n9548, new_n9547, new_n1531);
not_3  g09163(new_n9549, new_n9548);
nand_4 g09164(new_n9550, new_n9549, new_n1120);
nand_4 g09165(new_n9551, new_n9550, new_n1169);
nand_4 g09166(new_n9552, new_n9551, new_n1116);
nand_4 g09167(new_n9553, new_n9552, new_n1111);
nand_4 g09168(new_n9554, new_n9553, new_n1106);
nand_4 g09169(new_n9555_1, new_n9554, new_n1178);
nand_4 g09170(new_n9556, new_n9555_1, n4172);
nor_4  g09171(n9570, new_n9556, new_n1719);
nand_4 g09172(new_n9558, new_n1292, new_n1291);
nand_4 g09173(new_n9559, new_n9558, new_n1288);
nand_4 g09174(new_n9560, new_n9559, new_n1284);
nand_4 g09175(new_n9561, new_n9560, new_n1280);
nand_4 g09176(new_n9562, new_n9561, new_n1275);
nand_4 g09177(new_n9563, new_n9562, new_n1445);
nand_4 g09178(new_n9564, new_n9563, new_n1270);
nand_4 g09179(new_n9565, new_n9564, new_n1265_1);
nand_4 g09180(new_n9566, new_n9565, new_n1260);
nand_4 g09181(new_n9567, new_n9566, new_n1256);
nand_4 g09182(new_n9568, new_n9567, new_n1251);
nand_4 g09183(new_n9569, new_n9568, new_n1457);
nand_4 g09184(new_n9570_1, new_n9569, new_n1462);
nand_4 g09185(new_n9571, new_n9570_1, new_n1468);
nand_4 g09186(new_n9572, new_n9571, new_n1247);
nand_4 g09187(new_n9573, new_n9572, new_n1474);
nand_4 g09188(new_n9574, new_n9573, new_n592);
nand_4 g09189(new_n9575, new_n9574, new_n585);
nand_4 g09190(new_n9576, new_n9575, new_n580);
nand_4 g09191(new_n9577, new_n9576, new_n600);
nand_4 g09192(new_n9578, new_n9577, new_n606);
nand_4 g09193(new_n9579, new_n9578, new_n612);
nand_4 g09194(new_n9580, new_n9579, new_n575);
nand_4 g09195(new_n9581, new_n9580, new_n619);
nand_4 g09196(new_n9582, new_n9581, new_n570);
nand_4 g09197(new_n9583, new_n9582, new_n625);
nand_4 g09198(new_n9584, new_n9583, new_n564);
nand_4 g09199(new_n9585, new_n9584, new_n632);
nand_4 g09200(new_n9586, new_n9585, new_n638);
nand_4 g09201(new_n9587, new_n9586, new_n559);
nand_4 g09202(new_n9588, new_n9587, new_n554);
nand_4 g09203(new_n9589_1, new_n9588, new_n646);
nand_4 g09204(new_n9590, new_n9589_1, new_n652);
nand_4 g09205(new_n9591, new_n9590, new_n549);
nand_4 g09206(new_n9592, new_n9591, new_n544);
not_3  g09207(new_n9593, new_n9592);
nor_4  g09208(new_n9594, new_n9593, new_n3069);
nor_4  g09209(new_n9595, new_n9594, new_n3068);
nor_4  g09210(new_n9596, new_n9595, new_n3067);
nor_4  g09211(new_n9597, new_n9596, new_n3066);
nor_4  g09212(new_n9598, new_n9597, new_n3065);
nor_4  g09213(new_n9599, new_n9598, new_n3064);
nor_4  g09214(new_n9600, new_n9599, new_n3063);
nor_4  g09215(new_n9601, new_n9600, new_n3062);
nor_4  g09216(new_n9602, new_n9601, new_n3061);
nor_4  g09217(new_n9603, new_n9602, new_n3354);
nor_4  g09218(new_n9604, new_n9603, new_n3353);
nor_4  g09219(new_n9605, new_n9604, new_n3352);
nor_4  g09220(new_n9606, new_n9605, new_n3351);
nor_4  g09221(new_n9607, new_n9606, new_n3350);
nor_4  g09222(new_n9608, new_n9607, new_n3349);
nor_4  g09223(new_n9609, new_n9608, new_n3348);
nor_4  g09224(new_n9610, new_n9609, new_n720);
nor_4  g09225(new_n9611, new_n9610, new_n501);
nor_4  g09226(new_n9612, new_n9611, new_n728);
not_3  g09227(new_n9613, new_n9612);
nand_4 g09228(new_n9614, new_n9613, new_n494);
nand_4 g09229(new_n9615, new_n9614, new_n735);
nand_4 g09230(new_n9616, new_n9615, new_n488);
nand_4 g09231(new_n9617, new_n9616, new_n743);
nand_4 g09232(new_n9618, new_n9617, new_n482);
nand_4 g09233(new_n9619, new_n9618, new_n751);
nand_4 g09234(new_n9620, new_n9619, new_n758);
nand_4 g09235(new_n9621, new_n9620, new_n765);
nand_4 g09236(new_n9622, new_n9621, new_n476);
nand_4 g09237(new_n9623, new_n9622, new_n773);
nand_4 g09238(new_n9624, new_n9623, new_n780);
nand_4 g09239(new_n9625, new_n9624, new_n787);
nand_4 g09240(new_n9626, new_n9625, new_n470);
nand_4 g09241(new_n9627, new_n9626, new_n795);
nand_4 g09242(new_n9628, new_n9627, new_n803);
nand_4 g09243(new_n9629, new_n9628, new_n809);
nand_4 g09244(new_n9630, new_n9629, new_n465);
nand_4 g09245(new_n9631, new_n9630, new_n818);
nand_4 g09246(new_n9632, new_n9631, new_n460);
nand_4 g09247(new_n9633, new_n9632, new_n455);
nand_4 g09248(new_n9634, new_n9633, new_n449);
nand_4 g09249(new_n9635, new_n9634, new_n827);
nand_4 g09250(new_n9636, new_n9635, new_n833);
nand_4 g09251(new_n9637, new_n9636, new_n444);
nand_4 g09252(new_n9638, new_n9637, new_n439);
nand_4 g09253(new_n9639, new_n9638, new_n841);
nand_4 g09254(new_n9640, new_n9639, new_n434);
nand_4 g09255(new_n9641, new_n9640, new_n429);
nand_4 g09256(new_n9642, new_n9641, new_n424);
nand_4 g09257(new_n9643, new_n9642, new_n850);
nand_4 g09258(new_n9644, new_n9643, n13511);
nor_4  g09259(n9665, new_n9644, new_n853);
nand_4 g09260(new_n9646, new_n1073, new_n650_1);
nand_4 g09261(new_n9647, new_n9646, new_n549);
nand_4 g09262(new_n9648, new_n9647, new_n544);
nand_4 g09263(new_n9649, new_n9648, new_n660);
nand_4 g09264(new_n9650, new_n9649, new_n539);
nand_4 g09265(new_n9651, new_n9650, new_n534);
nand_4 g09266(new_n9652, new_n9651, new_n529);
nand_4 g09267(new_n9653, new_n9652, new_n668);
nand_4 g09268(new_n9654, new_n9653, new_n674_1);
nand_4 g09269(new_n9655, new_n9654, new_n681);
nand_4 g09270(new_n9656, new_n9655, new_n523);
nand_4 g09271(new_n9657, new_n9656, new_n687);
nand_4 g09272(new_n9658, new_n9657, new_n693);
nand_4 g09273(new_n9659, new_n9658, new_n699);
nand_4 g09274(new_n9660, new_n9659, new_n517);
nand_4 g09275(new_n9661, new_n9660, new_n705);
nand_4 g09276(new_n9662, new_n9661, new_n511);
nand_4 g09277(new_n9663, new_n9662, new_n711);
nand_4 g09278(new_n9664, new_n9663, new_n506);
nand_4 g09279(new_n9665_1, new_n9664, new_n719);
nand_4 g09280(new_n9666, new_n9665_1, new_n500);
nand_4 g09281(new_n9667, new_n9666, new_n727);
nand_4 g09282(new_n9668, new_n9667, new_n494);
nand_4 g09283(new_n9669, new_n9668, new_n735);
nand_4 g09284(new_n9670, new_n9669, new_n488);
nand_4 g09285(new_n9671, new_n9670, new_n743);
nand_4 g09286(new_n9672, new_n9671, new_n482);
nand_4 g09287(new_n9673, new_n9672, new_n751);
nand_4 g09288(new_n9674, new_n9673, new_n758);
nand_4 g09289(new_n9675, new_n9674, new_n765);
nand_4 g09290(new_n9676, new_n9675, new_n476);
nand_4 g09291(new_n9677, new_n9676, new_n773);
nand_4 g09292(new_n9678, new_n9677, new_n780);
nand_4 g09293(new_n9679, new_n9678, new_n787);
nand_4 g09294(new_n9680, new_n9679, new_n470);
nand_4 g09295(new_n9681, new_n9680, new_n795);
nand_4 g09296(new_n9682, new_n9681, new_n803);
nand_4 g09297(new_n9683, new_n9682, new_n809);
nand_4 g09298(new_n9684, new_n9683, new_n465);
nand_4 g09299(new_n9685, new_n9684, new_n818);
nand_4 g09300(new_n9686, new_n9685, new_n460);
nand_4 g09301(new_n9687, new_n9686, new_n455);
nand_4 g09302(new_n9688, new_n9687, new_n449);
nand_4 g09303(new_n9689, new_n9688, new_n827);
nand_4 g09304(new_n9690, new_n9689, new_n833);
nand_4 g09305(new_n9691, new_n9690, new_n444);
not_3  g09306(new_n9692, new_n9691);
nor_4  g09307(new_n9693, new_n9692, new_n2035);
nor_4  g09308(new_n9694, new_n9693, new_n2034);
nor_4  g09309(new_n9695, new_n9694, new_n2033);
nor_4  g09310(new_n9696, new_n9695, new_n2032);
nor_4  g09311(new_n9697, new_n9696, new_n2031);
nor_4  g09312(new_n9698, new_n9697, new_n2030);
nor_4  g09313(new_n9699, new_n9698, new_n2029);
nor_4  g09314(new_n9700, new_n9699, new_n2028);
nor_4  g09315(new_n9701, new_n9700, new_n2027_1);
nor_4  g09316(new_n9702, new_n9701, new_n2026);
nor_4  g09317(new_n9703, new_n9702, new_n2025);
nor_4  g09318(new_n9704, new_n9703, new_n2024);
nor_4  g09319(new_n9705, new_n9704, new_n2023);
nor_4  g09320(new_n9706, new_n9705, new_n2022);
nor_4  g09321(new_n9707, new_n9706, new_n2021);
nor_4  g09322(new_n9708, new_n9707, new_n2020);
nor_4  g09323(new_n9709, new_n9708, new_n2019);
nor_4  g09324(new_n9710, new_n9709, new_n1537);
nor_4  g09325(new_n9711, new_n9710, new_n1536);
nor_4  g09326(new_n9712, new_n9711, new_n1535);
nor_4  g09327(new_n9713, new_n9712, new_n1534);
nor_4  g09328(new_n9714, new_n9713, new_n1533);
nor_4  g09329(new_n9715, new_n9714, new_n1532);
nor_4  g09330(new_n9716, new_n9715, new_n1531);
not_3  g09331(new_n9717_1, new_n9716);
nand_4 g09332(new_n9718, new_n9717_1, new_n1120);
nand_4 g09333(new_n9719, new_n9718, new_n1169);
nand_4 g09334(new_n9720, new_n9719, new_n1116);
nand_4 g09335(new_n9721, new_n9720, new_n1111);
nand_4 g09336(new_n9722, new_n9721, new_n1106);
nand_4 g09337(new_n9723, new_n9722, new_n1178);
nand_4 g09338(new_n9724, new_n9723, new_n1183);
nand_4 g09339(new_n9725, new_n9724, new_n1102);
nand_4 g09340(new_n9726, new_n9725, new_n1099);
nand_4 g09341(new_n9727, new_n9726, new_n1191);
nand_4 g09342(new_n9728, new_n9727, new_n1095);
nand_4 g09343(new_n9729, new_n9728, new_n1091);
nand_4 g09344(new_n9730, new_n9729, new_n1088);
nand_4 g09345(new_n9731, new_n9730, new_n1084);
nand_4 g09346(new_n9732, new_n9731, n6873);
nor_4  g09347(n9717, new_n9732, new_n1862);
nand_4 g09348(new_n9734, new_n1889, new_n1018);
nand_4 g09349(new_n9735, new_n9734, new_n1015);
nand_4 g09350(new_n9736, new_n9735, new_n1010);
nand_4 g09351(new_n9737, new_n9736, new_n1215);
nand_4 g09352(new_n9738, new_n9737, new_n1005);
nand_4 g09353(new_n9739, new_n9738, new_n1000);
nand_4 g09354(new_n9740, new_n9739, new_n994);
nand_4 g09355(new_n9741, new_n9740, new_n989);
nand_4 g09356(new_n9742, new_n9741, new_n984);
nand_4 g09357(new_n9743, new_n9742, new_n978);
nand_4 g09358(new_n9744, new_n9743, new_n973);
nand_4 g09359(new_n9745, new_n9744, new_n967);
nand_4 g09360(new_n9746, new_n9745, new_n964);
nand_4 g09361(new_n9747, new_n9746, new_n960);
nand_4 g09362(new_n9748, new_n9747, new_n957);
nand_4 g09363(new_n9749, new_n9748, new_n952);
nand_4 g09364(new_n9750, new_n9749, new_n948_1);
nand_4 g09365(new_n9751, new_n9750, new_n943);
nand_4 g09366(new_n9752, new_n9751, new_n938);
nand_4 g09367(new_n9753, new_n9752, new_n934);
nand_4 g09368(new_n9754, new_n9753, new_n929);
nand_4 g09369(new_n9755, new_n9754, new_n925);
nand_4 g09370(new_n9756, new_n9755, new_n2194);
nand_4 g09371(new_n9757, new_n9756, new_n2191);
nand_4 g09372(new_n9758, new_n9757, new_n2190);
nand_4 g09373(new_n9759, new_n9758, new_n2186);
nand_4 g09374(new_n9760, new_n9759, new_n2183);
nand_4 g09375(new_n9761, new_n9760, new_n2179);
nand_4 g09376(new_n9762, new_n9761, new_n2175_1);
nand_4 g09377(new_n9763, new_n9762, new_n2171);
nand_4 g09378(new_n9764, new_n9763, new_n2168);
nand_4 g09379(new_n9765, new_n9764, new_n2165);
nand_4 g09380(new_n9766, new_n9765, new_n2162);
nand_4 g09381(new_n9767, new_n9766, new_n2158);
nand_4 g09382(new_n9768, new_n9767, new_n2155);
nand_4 g09383(new_n9769, new_n9768, new_n2151);
nand_4 g09384(new_n9770, new_n9769, new_n2147);
nand_4 g09385(new_n9771, new_n9770, new_n1810);
nand_4 g09386(new_n9772, new_n9771, new_n1806);
nand_4 g09387(new_n9773, new_n9772, new_n1802);
nand_4 g09388(new_n9774, new_n9773, new_n1798);
nand_4 g09389(new_n9775, new_n9774, new_n1820);
not_3  g09390(new_n9776, new_n9775);
nor_4  g09391(new_n9777, new_n9776, new_n2304);
nor_4  g09392(new_n9778, new_n9777, new_n2303);
nor_4  g09393(new_n9779, new_n9778, new_n2302);
nor_4  g09394(new_n9780, new_n9779, new_n2301);
nor_4  g09395(new_n9781, new_n9780, new_n2300);
nor_4  g09396(new_n9782, new_n9781, new_n2299);
nor_4  g09397(new_n9783, new_n9782, new_n2298);
nor_4  g09398(new_n9784, new_n9783, new_n2297);
nor_4  g09399(new_n9785, new_n9784, new_n2296);
nor_4  g09400(new_n9786, new_n9785, new_n2295);
nor_4  g09401(new_n9787, new_n9786, new_n2294);
nor_4  g09402(new_n9788, new_n9787, new_n2293);
nor_4  g09403(new_n9789, new_n9788, new_n2292);
nor_4  g09404(new_n9790, new_n9789, new_n2291);
nor_4  g09405(new_n9791, new_n9790, new_n2290);
nor_4  g09406(new_n9792, new_n9791, new_n2289);
nor_4  g09407(new_n9793, new_n9792, new_n2288);
nor_4  g09408(new_n9794, new_n9793, new_n2287);
nor_4  g09409(new_n9795, new_n9794, new_n2286);
nor_4  g09410(new_n9796, new_n9795, new_n2285);
nor_4  g09411(new_n9797, new_n9796, new_n2284);
nor_4  g09412(new_n9798, new_n9797, new_n2283);
not_3  g09413(new_n9799, new_n9798);
nand_4 g09414(new_n9800, new_n9799, new_n1724);
nand_4 g09415(new_n9801, new_n9800, new_n1721);
nand_4 g09416(new_n9802, new_n9801, new_n1718);
nand_4 g09417(new_n9803, new_n9802, new_n1715);
nand_4 g09418(new_n9804, new_n9803, new_n1711);
nand_4 g09419(new_n9805, new_n9804, new_n1708);
nand_4 g09420(new_n9806, new_n9805, new_n1705);
nand_4 g09421(new_n9807, new_n9806, new_n1703);
nand_4 g09422(new_n9808, new_n9807, new_n1860);
nand_4 g09423(new_n9809, new_n9808, new_n1864);
nand_4 g09424(new_n9810, new_n9809, new_n1699);
nand_4 g09425(new_n9811, new_n9810, new_n1697);
nand_4 g09426(new_n9812, new_n9811, new_n1871);
nand_4 g09427(new_n9813, new_n9812, new_n1694);
nand_4 g09428(new_n9814, new_n9813, new_n1690);
nand_4 g09429(new_n9815, new_n9814, new_n1878);
nand_4 g09430(new_n9816, new_n9815, new_n1882);
nand_4 g09431(new_n9817, new_n9816, new_n1686);
nand_4 g09432(new_n9818, new_n9817, new_n1682);
nand_4 g09433(new_n9819, new_n9818, new_n1678);
nand_4 g09434(new_n9820, new_n9819, n4154);
nor_4  g09435(n10515, new_n9820, new_n1671);
nand_4 g09436(new_n9822, new_n896, new_n886);
nand_4 g09437(new_n9823, new_n9822, new_n901);
nand_4 g09438(new_n9824, new_n9823, new_n408);
nand_4 g09439(new_n9825, new_n9824, new_n908);
nand_4 g09440(new_n9826, new_n9825, new_n403);
nand_4 g09441(new_n9827, new_n9826, new_n398);
nand_4 g09442(new_n9828, new_n9827, new_n393);
nand_4 g09443(new_n9829, new_n9828, new_n916);
nand_4 g09444(new_n9830_1, new_n9829, new_n1123);
nand_4 g09445(new_n9831, new_n9830_1, new_n1164);
nand_4 g09446(new_n9832, new_n9831, new_n1120);
nand_4 g09447(new_n9833, new_n9832, new_n1169);
nand_4 g09448(new_n9834, new_n9833, new_n1116);
nand_4 g09449(new_n9835, new_n9834, new_n1111);
nand_4 g09450(new_n9836, new_n9835, new_n1106);
nand_4 g09451(new_n9837, new_n9836, new_n1178);
nand_4 g09452(new_n9838, new_n9837, new_n1183);
nand_4 g09453(new_n9839, new_n9838, new_n1102);
nand_4 g09454(new_n9840, new_n9839, new_n1099);
nand_4 g09455(new_n9841, new_n9840, new_n1191);
nand_4 g09456(new_n9842, new_n9841, new_n1095);
nand_4 g09457(new_n9843, new_n9842, new_n1091);
nand_4 g09458(new_n9844, new_n9843, new_n1088);
nand_4 g09459(new_n9845, new_n9844, new_n1084);
nand_4 g09460(new_n9846, new_n9845, new_n1079);
nand_4 g09461(new_n9847, new_n9846, new_n1074);
nand_4 g09462(new_n9848, new_n9847, new_n1070);
nand_4 g09463(new_n9849, new_n9848, new_n1064);
nand_4 g09464(new_n9850, new_n9849, new_n1061);
nand_4 g09465(new_n9851, new_n9850, new_n1055);
nand_4 g09466(new_n9852, new_n9851, new_n1050);
nand_4 g09467(new_n9853, new_n9852, new_n1045);
nand_4 g09468(new_n9854, new_n9853, new_n1041);
nand_4 g09469(new_n9855, new_n9854, new_n1036);
nand_4 g09470(new_n9856, new_n9855, new_n1031);
nand_4 g09471(new_n9857, new_n9856, new_n1025);
nand_4 g09472(new_n9858, new_n9857, new_n1020);
nand_4 g09473(new_n9859, new_n9858, new_n1015);
nand_4 g09474(new_n9860, new_n9859, new_n1010);
nand_4 g09475(new_n9861, new_n9860, new_n1215);
nand_4 g09476(new_n9862, new_n9861, new_n1005);
nand_4 g09477(new_n9863, new_n9862, new_n1000);
nand_4 g09478(new_n9864, new_n9863, new_n994);
nand_4 g09479(new_n9865, new_n9864, new_n989);
nand_4 g09480(new_n9866, new_n9865, new_n984);
nand_4 g09481(new_n9867, new_n9866, new_n978);
nand_4 g09482(new_n9868, new_n9867, new_n973);
nand_4 g09483(new_n9869, new_n9868, new_n967);
nand_4 g09484(new_n9870, new_n9869, new_n964);
nand_4 g09485(new_n9871, new_n9870, new_n960);
nand_4 g09486(new_n9872, new_n9871, new_n957);
not_3  g09487(new_n9873, new_n9872);
nor_4  g09488(new_n9874, new_n9873, new_n953);
nor_4  g09489(new_n9875, new_n9874, new_n3536);
nor_4  g09490(new_n9876, new_n9875, new_n3535);
nor_4  g09491(new_n9877, new_n9876, new_n3534);
nor_4  g09492(new_n9878, new_n9877, new_n2520);
nor_4  g09493(new_n9879, new_n9878, new_n2519);
nor_4  g09494(new_n9880, new_n9879, new_n2518);
nor_4  g09495(new_n9881, new_n9880, new_n2517);
nor_4  g09496(new_n9882, new_n9881, new_n2516);
nor_4  g09497(new_n9883, new_n9882, new_n2515);
nor_4  g09498(new_n9884, new_n9883, new_n2514);
nor_4  g09499(new_n9885, new_n9884, new_n2513);
nor_4  g09500(new_n9886, new_n9885, new_n2512);
nor_4  g09501(new_n9887, new_n9886, new_n2511);
nor_4  g09502(new_n9888, new_n9887, new_n2510);
nor_4  g09503(new_n9889, new_n9888, new_n2509);
nor_4  g09504(new_n9890, new_n9889, new_n2508);
nor_4  g09505(new_n9891, new_n9890, new_n2507);
nor_4  g09506(new_n9892, new_n9891, new_n2506);
nor_4  g09507(new_n9893_1, new_n9892, new_n2505);
nor_4  g09508(new_n9894, new_n9893_1, new_n2504);
nor_4  g09509(new_n9895, new_n9894, new_n2503);
nor_4  g09510(new_n9896, new_n9895, new_n2502);
nor_4  g09511(new_n9897, new_n9896, new_n2790);
nor_4  g09512(new_n9898, new_n9897, new_n2789);
nor_4  g09513(new_n9899, new_n9898, new_n2788);
nor_4  g09514(new_n9900, new_n9899, new_n2305);
not_3  g09515(new_n9901, new_n9900);
nand_4 g09516(new_n9902, new_n9901, new_n1794);
nand_4 g09517(new_n9903, new_n9902, new_n1825);
nand_4 g09518(new_n9904, new_n9903, new_n1789);
nand_4 g09519(new_n9905, new_n9904, new_n1785);
nand_4 g09520(new_n9906, new_n9905, new_n1780);
nand_4 g09521(new_n9907, new_n9906, new_n1777);
nand_4 g09522(new_n9908, new_n9907, n3910);
nor_4  g09523(n10591, new_n9908, new_n1771);
nand_4 g09524(new_n9910, new_n1336, new_n786);
nand_4 g09525(new_n9911, new_n9910, new_n1395);
nand_4 g09526(new_n9912, new_n9911, new_n1335);
nand_4 g09527(new_n9913, new_n9912, new_n1332);
nand_4 g09528(new_n9914, new_n9913, new_n1328);
nand_4 g09529(new_n9915, new_n9914, new_n1403);
nand_4 g09530(new_n9916, new_n9915, new_n1325);
nand_4 g09531(new_n9917, new_n9916, new_n1410);
nand_4 g09532(new_n9918, new_n9917, new_n1413);
nand_4 g09533(new_n9919, new_n9918, new_n1322);
nand_4 g09534(new_n9920, new_n9919, new_n1317);
nand_4 g09535(new_n9921_1, new_n9920, new_n1315);
nand_4 g09536(new_n9922, new_n9921_1, new_n1419);
nand_4 g09537(new_n9923, new_n9922, new_n1310);
nand_4 g09538(new_n9924, new_n9923, new_n1305);
nand_4 g09539(new_n9925, new_n9924, new_n1427);
nand_4 g09540(new_n9926, new_n9925, new_n1431);
nand_4 g09541(new_n9927, new_n9926, new_n1302);
nand_4 g09542(new_n9928, new_n9927, new_n1298);
nand_4 g09543(new_n9929, new_n9928, new_n1295);
nand_4 g09544(new_n9930, new_n9929, new_n1291);
nand_4 g09545(new_n9931, new_n9930, new_n1288);
nand_4 g09546(new_n9932, new_n9931, new_n1284);
nand_4 g09547(new_n9933, new_n9932, new_n1280);
nand_4 g09548(new_n9934, new_n9933, new_n1275);
nand_4 g09549(new_n9935, new_n9934, new_n1445);
nand_4 g09550(new_n9936_1, new_n9935, new_n1270);
nand_4 g09551(new_n9937, new_n9936_1, new_n1265_1);
nand_4 g09552(new_n9938, new_n9937, new_n1260);
nand_4 g09553(new_n9939, new_n9938, new_n1256);
nand_4 g09554(new_n9940, new_n9939, new_n1251);
nand_4 g09555(new_n9941, new_n9940, new_n1457);
nand_4 g09556(new_n9942, new_n9941, new_n1462);
nand_4 g09557(new_n9943, new_n9942, new_n1468);
nand_4 g09558(new_n9944, new_n9943, new_n1247);
nand_4 g09559(new_n9945, new_n9944, new_n1474);
nand_4 g09560(new_n9946, new_n9945, new_n592);
nand_4 g09561(new_n9947, new_n9946, new_n585);
nand_4 g09562(new_n9948, new_n9947, new_n580);
nand_4 g09563(new_n9949, new_n9948, new_n600);
nand_4 g09564(new_n9950, new_n9949, new_n606);
nand_4 g09565(new_n9951, new_n9950, new_n612);
nand_4 g09566(new_n9952, new_n9951, new_n575);
nand_4 g09567(new_n9953, new_n9952, new_n619);
nand_4 g09568(new_n9954, new_n9953, new_n570);
nand_4 g09569(new_n9955, new_n9954, new_n625);
not_3  g09570(new_n9956, new_n9955);
nor_4  g09571(new_n9957, new_n9956, new_n3078);
nor_4  g09572(new_n9958, new_n9957, new_n3077);
nor_4  g09573(new_n9959, new_n9958, new_n3076);
nor_4  g09574(new_n9960, new_n9959, new_n3075);
nor_4  g09575(new_n9961, new_n9960, new_n3074);
nor_4  g09576(new_n9962, new_n9961, new_n3073);
nor_4  g09577(new_n9963, new_n9962, new_n3072);
nor_4  g09578(new_n9964, new_n9963, new_n3071);
nor_4  g09579(new_n9965, new_n9964, new_n3070);
nor_4  g09580(new_n9966, new_n9965, new_n3069);
nor_4  g09581(new_n9967, new_n9966, new_n3068);
nor_4  g09582(new_n9968, new_n9967, new_n3067);
nor_4  g09583(new_n9969, new_n9968, new_n3066);
nor_4  g09584(new_n9970, new_n9969, new_n3065);
nor_4  g09585(new_n9971, new_n9970, new_n3064);
nor_4  g09586(new_n9972, new_n9971, new_n3063);
nor_4  g09587(new_n9973, new_n9972, new_n3062);
nor_4  g09588(new_n9974, new_n9973, new_n3061);
nor_4  g09589(new_n9975, new_n9974, new_n3354);
nor_4  g09590(new_n9976, new_n9975, new_n3353);
nor_4  g09591(new_n9977_1, new_n9976, new_n3352);
nor_4  g09592(new_n9978, new_n9977_1, new_n3351);
nor_4  g09593(new_n9979, new_n9978, new_n3350);
nor_4  g09594(new_n9980, new_n9979, new_n3349);
not_3  g09595(new_n9981, new_n9980);
nand_4 g09596(new_n9982, new_n9981, new_n506);
nand_4 g09597(new_n9983, new_n9982, new_n719);
nand_4 g09598(new_n9984, new_n9983, new_n500);
nand_4 g09599(new_n9985, new_n9984, new_n727);
nand_4 g09600(new_n9986, new_n9985, new_n494);
nand_4 g09601(new_n9987, new_n9986, new_n735);
nand_4 g09602(new_n9988, new_n9987, new_n488);
nand_4 g09603(new_n9989, new_n9988, new_n743);
nand_4 g09604(new_n9990, new_n9989, new_n482);
nand_4 g09605(new_n9991, new_n9990, new_n751);
nand_4 g09606(new_n9992, new_n9991, new_n758);
nand_4 g09607(new_n9993, new_n9992, new_n765);
nand_4 g09608(new_n9994, new_n9993, new_n476);
nand_4 g09609(new_n9995, new_n9994, new_n773);
nand_4 g09610(new_n9996, new_n9995, n10378);
nor_4  g09611(n10791, new_n9996, new_n777);
nand_4 g09612(new_n9998, new_n1776_1, new_n411_1);
nand_4 g09613(new_n9999, new_n9998, new_n889);
nand_4 g09614(new_n10000, new_n9999, new_n896);
nand_4 g09615(new_n10001, new_n10000, new_n901);
nand_4 g09616(new_n10002, new_n10001, new_n408);
nand_4 g09617(new_n10003, new_n10002, new_n908);
nand_4 g09618(new_n10004, new_n10003, new_n403);
nand_4 g09619(new_n10005, new_n10004, new_n398);
nand_4 g09620(new_n10006, new_n10005, new_n393);
nand_4 g09621(new_n10007, new_n10006, new_n916);
nand_4 g09622(new_n10008, new_n10007, new_n1123);
nand_4 g09623(new_n10009, new_n10008, new_n1164);
nand_4 g09624(new_n10010, new_n10009, new_n1120);
nand_4 g09625(new_n10011, new_n10010, new_n1169);
nand_4 g09626(new_n10012, new_n10011, new_n1116);
nand_4 g09627(new_n10013, new_n10012, new_n1111);
nand_4 g09628(new_n10014, new_n10013, new_n1106);
nand_4 g09629(new_n10015, new_n10014, new_n1178);
nand_4 g09630(new_n10016, new_n10015, new_n1183);
nand_4 g09631(new_n10017, new_n10016, new_n1102);
nand_4 g09632(new_n10018, new_n10017, new_n1099);
nand_4 g09633(new_n10019, new_n10018, new_n1191);
nand_4 g09634(new_n10020, new_n10019, new_n1095);
nand_4 g09635(new_n10021, new_n10020, new_n1091);
nand_4 g09636(new_n10022, new_n10021, new_n1088);
nand_4 g09637(new_n10023, new_n10022, new_n1084);
nand_4 g09638(new_n10024, new_n10023, new_n1079);
nand_4 g09639(new_n10025, new_n10024, new_n1074);
nand_4 g09640(new_n10026, new_n10025, new_n1070);
nand_4 g09641(new_n10027, new_n10026, new_n1064);
nand_4 g09642(new_n10028, new_n10027, new_n1061);
nand_4 g09643(new_n10029, new_n10028, new_n1055);
nand_4 g09644(new_n10030, new_n10029, new_n1050);
nand_4 g09645(new_n10031, new_n10030, new_n1045);
nand_4 g09646(new_n10032, new_n10031, new_n1041);
nand_4 g09647(new_n10033, new_n10032, new_n1036);
nand_4 g09648(new_n10034, new_n10033, new_n1031);
nand_4 g09649(new_n10035, new_n10034, new_n1025);
nand_4 g09650(new_n10036, new_n10035, new_n1020);
nand_4 g09651(new_n10037, new_n10036, new_n1015);
nand_4 g09652(new_n10038, new_n10037, new_n1010);
nand_4 g09653(new_n10039, new_n10038, new_n1215);
nand_4 g09654(new_n10040, new_n10039, new_n1005);
nand_4 g09655(new_n10041, new_n10040, new_n1000);
nand_4 g09656(new_n10042, new_n10041, new_n994);
nand_4 g09657(new_n10043, new_n10042, new_n989);
not_3  g09658(new_n10044, new_n10043);
nor_4  g09659(new_n10045, new_n10044, new_n985);
nor_4  g09660(new_n10046, new_n10045, new_n979);
nor_4  g09661(new_n10047, new_n10046, new_n974);
nor_4  g09662(new_n10048, new_n10047, new_n968);
nor_4  g09663(new_n10049, new_n10048, new_n965);
nor_4  g09664(new_n10050_1, new_n10049, new_n961);
nor_4  g09665(new_n10051_1, new_n10050_1, new_n958);
nor_4  g09666(new_n10052, new_n10051_1, new_n953);
nor_4  g09667(new_n10053, new_n10052, new_n3536);
nor_4  g09668(new_n10054, new_n10053, new_n3535);
nor_4  g09669(new_n10055, new_n10054, new_n3534);
nor_4  g09670(new_n10056, new_n10055, new_n2520);
nor_4  g09671(new_n10057, new_n10056, new_n2519);
nor_4  g09672(new_n10058, new_n10057, new_n2518);
nor_4  g09673(new_n10059, new_n10058, new_n2517);
nor_4  g09674(new_n10060, new_n10059, new_n2516);
nor_4  g09675(new_n10061_1, new_n10060, new_n2515);
nor_4  g09676(new_n10062, new_n10061_1, new_n2514);
nor_4  g09677(new_n10063, new_n10062, new_n2513);
nor_4  g09678(new_n10064, new_n10063, new_n2512);
nor_4  g09679(new_n10065, new_n10064, new_n2511);
nor_4  g09680(new_n10066, new_n10065, new_n2510);
nor_4  g09681(new_n10067, new_n10066, new_n2509);
nor_4  g09682(new_n10068, new_n10067, new_n2508);
not_3  g09683(new_n10069, new_n10068);
nand_4 g09684(new_n10070, new_n10069, new_n2162);
nand_4 g09685(new_n10071, new_n10070, new_n2158);
nand_4 g09686(new_n10072, new_n10071, new_n2155);
nand_4 g09687(new_n10073, new_n10072, new_n2151);
nand_4 g09688(new_n10074, new_n10073, new_n2147);
nand_4 g09689(new_n10075, new_n10074, new_n1810);
nand_4 g09690(new_n10076, new_n10075, new_n1806);
nand_4 g09691(new_n10077, new_n10076, new_n1802);
nand_4 g09692(new_n10078, new_n10077, new_n1798);
nand_4 g09693(new_n10079, new_n10078, new_n1820);
nand_4 g09694(new_n10080_1, new_n10079, new_n1794);
nand_4 g09695(new_n10081, new_n10080_1, new_n1825);
nand_4 g09696(new_n10082, new_n10081, new_n1789);
nand_4 g09697(new_n10083, new_n10082, new_n1785);
nand_4 g09698(new_n10084, new_n10083, n13186);
nor_4  g09699(n10802, new_n10084, new_n1277);
not_3  g09700(new_n10086, new_n1801);
nand_4 g09701(new_n10087, new_n10086, new_n1300);
nand_4 g09702(new_n10088, new_n10087, new_n422);
nand_4 g09703(new_n10089, new_n10088, new_n850);
nand_4 g09704(new_n10090, new_n10089, new_n856);
nand_4 g09705(new_n10091, new_n10090, new_n863);
nand_4 g09706(new_n10092, new_n10091, new_n419);
nand_4 g09707(new_n10093, new_n10092, new_n869);
nand_4 g09708(new_n10094, new_n10093, new_n875);
nand_4 g09709(new_n10095, new_n10094, new_n881);
nand_4 g09710(new_n10096, new_n10095, new_n413);
nand_4 g09711(new_n10097, new_n10096, new_n889);
nand_4 g09712(new_n10098, new_n10097, new_n896);
nand_4 g09713(new_n10099, new_n10098, new_n901);
nand_4 g09714(new_n10100, new_n10099, new_n408);
nand_4 g09715(new_n10101, new_n10100, new_n908);
nand_4 g09716(new_n10102, new_n10101, new_n403);
nand_4 g09717(new_n10103, new_n10102, new_n398);
nand_4 g09718(new_n10104, new_n10103, new_n393);
nand_4 g09719(new_n10105, new_n10104, new_n916);
nand_4 g09720(new_n10106, new_n10105, new_n1123);
nand_4 g09721(new_n10107, new_n10106, new_n1164);
nand_4 g09722(new_n10108, new_n10107, new_n1120);
nand_4 g09723(new_n10109, new_n10108, new_n1169);
nand_4 g09724(new_n10110, new_n10109, new_n1116);
nand_4 g09725(new_n10111, new_n10110, new_n1111);
nand_4 g09726(new_n10112_1, new_n10111, new_n1106);
nand_4 g09727(new_n10113, new_n10112_1, new_n1178);
nand_4 g09728(new_n10114, new_n10113, new_n1183);
nand_4 g09729(new_n10115, new_n10114, new_n1102);
nand_4 g09730(new_n10116, new_n10115, new_n1099);
nand_4 g09731(new_n10117, new_n10116, new_n1191);
nand_4 g09732(new_n10118, new_n10117, new_n1095);
nand_4 g09733(new_n10119, new_n10118, new_n1091);
nand_4 g09734(new_n10120, new_n10119, new_n1088);
nand_4 g09735(new_n10121, new_n10120, new_n1084);
nand_4 g09736(new_n10122, new_n10121, new_n1079);
nand_4 g09737(new_n10123, new_n10122, new_n1074);
nand_4 g09738(new_n10124, new_n10123, new_n1070);
nand_4 g09739(new_n10125, new_n10124, new_n1064);
nand_4 g09740(new_n10126, new_n10125, new_n1061);
nand_4 g09741(new_n10127, new_n10126, new_n1055);
nand_4 g09742(new_n10128, new_n10127, new_n1050);
nand_4 g09743(new_n10129, new_n10128, new_n1045);
nand_4 g09744(new_n10130, new_n10129, new_n1041);
nand_4 g09745(new_n10131, new_n10130, new_n1036);
nand_4 g09746(new_n10132, new_n10131, new_n1031);
not_3  g09747(new_n10133, new_n10132);
nor_4  g09748(new_n10134, new_n10133, new_n1026);
nor_4  g09749(new_n10135, new_n10134, new_n1021);
nor_4  g09750(new_n10136, new_n10135, new_n1016);
nor_4  g09751(new_n10137, new_n10136, new_n1011);
nor_4  g09752(new_n10138, new_n10137, new_n1216);
nor_4  g09753(new_n10139, new_n10138, new_n1006);
nor_4  g09754(new_n10140, new_n10139, new_n1001);
nor_4  g09755(new_n10141, new_n10140, new_n995);
nor_4  g09756(new_n10142, new_n10141, new_n990);
nor_4  g09757(new_n10143, new_n10142, new_n985);
nor_4  g09758(new_n10144, new_n10143, new_n979);
nor_4  g09759(new_n10145, new_n10144, new_n974);
nor_4  g09760(new_n10146, new_n10145, new_n968);
nor_4  g09761(new_n10147_1, new_n10146, new_n965);
nor_4  g09762(new_n10148, new_n10147_1, new_n961);
nor_4  g09763(new_n10149, new_n10148, new_n958);
nor_4  g09764(new_n10150, new_n10149, new_n953);
nor_4  g09765(new_n10151, new_n10150, new_n3536);
nor_4  g09766(new_n10152, new_n10151, new_n3535);
nor_4  g09767(new_n10153, new_n10152, new_n3534);
nor_4  g09768(new_n10154, new_n10153, new_n2520);
nor_4  g09769(new_n10155, new_n10154, new_n2519);
nor_4  g09770(new_n10156, new_n10155, new_n2518);
nor_4  g09771(new_n10157, new_n10156, new_n2517);
not_3  g09772(new_n10158, new_n10157);
nand_4 g09773(new_n10159, new_n10158, new_n2191);
nand_4 g09774(new_n10160, new_n10159, new_n2190);
nand_4 g09775(new_n10161, new_n10160, new_n2186);
nand_4 g09776(new_n10162, new_n10161, new_n2183);
nand_4 g09777(new_n10163, new_n10162, new_n2179);
nand_4 g09778(new_n10164, new_n10163, new_n2175_1);
nand_4 g09779(new_n10165, new_n10164, new_n2171);
nand_4 g09780(new_n10166, new_n10165, new_n2168);
nand_4 g09781(new_n10167, new_n10166, new_n2165);
nand_4 g09782(new_n10168, new_n10167, new_n2162);
nand_4 g09783(new_n10169, new_n10168, new_n2158);
nand_4 g09784(new_n10170, new_n10169, new_n2155);
nand_4 g09785(new_n10171, new_n10170, new_n2151);
nand_4 g09786(new_n10172, new_n10171, new_n2147);
nand_4 g09787(new_n10173, new_n10172, new_n1810);
nand_4 g09788(new_n10174, new_n10173, n7667);
nor_4  g09789(n10915, new_n10174, new_n1803);
nand_4 g09790(new_n10176, new_n1763_1, new_n1762);
nand_4 g09791(new_n10177, new_n10176, new_n1758);
nand_4 g09792(new_n10178, new_n10177, new_n1754);
nand_4 g09793(new_n10179, new_n10178, new_n1751);
nand_4 g09794(new_n10180, new_n10179, new_n1748);
nand_4 g09795(new_n10181, new_n10180, new_n1746);
nand_4 g09796(new_n10182, new_n10181, new_n1742);
nand_4 g09797(new_n10183, new_n10182, new_n1738);
nand_4 g09798(new_n10184, new_n10183, new_n1736);
nand_4 g09799(new_n10185, new_n10184, new_n1732);
nand_4 g09800(new_n10186, new_n10185, new_n1729);
nand_4 g09801(new_n10187, new_n10186, new_n1726);
nand_4 g09802(new_n10188, new_n10187, new_n1724);
nand_4 g09803(new_n10189, new_n10188, new_n1721);
nand_4 g09804(new_n10190, new_n10189, new_n1718);
nand_4 g09805(new_n10191, new_n10190, new_n1715);
nand_4 g09806(new_n10192, new_n10191, new_n1711);
nand_4 g09807(new_n10193, new_n10192, new_n1708);
nand_4 g09808(new_n10194, new_n10193, new_n1705);
nand_4 g09809(new_n10195, new_n10194, new_n1703);
nand_4 g09810(new_n10196, new_n10195, new_n1860);
nand_4 g09811(new_n10197, new_n10196, new_n1864);
nand_4 g09812(new_n10198, new_n10197, new_n1699);
nand_4 g09813(new_n10199, new_n10198, new_n1697);
nand_4 g09814(new_n10200, new_n10199, new_n1871);
nand_4 g09815(new_n10201, new_n10200, new_n1694);
nand_4 g09816(new_n10202, new_n10201, new_n1690);
nand_4 g09817(new_n10203, new_n10202, new_n1878);
nand_4 g09818(new_n10204, new_n10203, new_n1882);
nand_4 g09819(new_n10205, new_n10204, new_n1686);
nand_4 g09820(new_n10206, new_n10205, new_n1682);
nand_4 g09821(new_n10207, new_n10206, new_n1678);
nand_4 g09822(new_n10208, new_n10207, new_n1674);
nand_4 g09823(new_n10209, new_n10208, new_n1890);
nand_4 g09824(new_n10210, new_n10209, new_n1669);
not_3  g09825(new_n10211, new_n10210);
nor_4  g09826(new_n10212, new_n10211, new_n1666);
nor_4  g09827(new_n10213, new_n10212, new_n1662);
nor_4  g09828(new_n10214, new_n10213, new_n1658);
nor_4  g09829(new_n10215, new_n10214, new_n1653);
nor_4  g09830(new_n10216, new_n10215, new_n1649);
nor_4  g09831(new_n10217, new_n10216, new_n1645);
nor_4  g09832(new_n10218, new_n10217, new_n1641);
nor_4  g09833(new_n10219, new_n10218, new_n1637_1);
nor_4  g09834(new_n10220, new_n10219, new_n1633);
nor_4  g09835(new_n10221, new_n10220, new_n1629);
nor_4  g09836(new_n10222, new_n10221, new_n1628);
nor_4  g09837(new_n10223, new_n10222, new_n1627);
nor_4  g09838(new_n10224, new_n10223, new_n1626);
nor_4  g09839(new_n10225, new_n10224, new_n4700);
nor_4  g09840(new_n10226, new_n10225, new_n4699);
nor_4  g09841(new_n10227, new_n10226, new_n3722);
nor_4  g09842(new_n10228, new_n10227, new_n3721);
nor_4  g09843(new_n10229, new_n10228, new_n3720);
nor_4  g09844(new_n10230, new_n10229, new_n3719);
not_3  g09845(new_n10231, new_n10230);
nand_4 g09846(new_n10232, new_n10231, new_n1344);
nand_4 g09847(new_n10233, new_n10232, new_n1341);
nand_4 g09848(new_n10234, new_n10233, new_n1338);
nand_4 g09849(new_n10235, new_n10234, new_n1395);
nand_4 g09850(new_n10236, new_n10235, new_n1335);
nand_4 g09851(new_n10237, new_n10236, new_n1332);
nand_4 g09852(new_n10238, new_n10237, new_n1328);
nand_4 g09853(new_n10239, new_n10238, new_n1403);
nand_4 g09854(new_n10240, new_n10239, new_n1325);
nand_4 g09855(new_n10241, new_n10240, new_n1410);
nand_4 g09856(new_n10242, new_n10241, new_n1413);
nand_4 g09857(new_n10243, new_n10242, new_n1322);
nand_4 g09858(new_n10244, new_n10243, new_n1317);
nand_4 g09859(new_n10245, new_n10244, new_n1315);
nand_4 g09860(new_n10246, new_n10245, new_n1419);
nand_4 g09861(new_n10247, new_n10246, new_n1310);
nand_4 g09862(new_n10248, new_n10247, new_n1305);
nand_4 g09863(new_n10249, new_n10248, new_n1427);
nand_4 g09864(new_n10250, new_n10249, new_n1431);
nand_4 g09865(new_n10251, new_n10250, new_n1302);
nand_4 g09866(new_n10252, new_n10251, new_n1298);
nand_4 g09867(new_n10253, new_n10252, new_n1295);
nand_4 g09868(new_n10254, new_n10253, new_n1291);
nand_4 g09869(new_n10255_1, new_n10254, new_n1288);
nand_4 g09870(new_n10256, new_n10255_1, new_n1284);
nand_4 g09871(new_n10257, new_n10256, new_n1280);
nand_4 g09872(new_n10258, new_n10257, new_n1275);
nand_4 g09873(new_n10259, new_n10258, new_n1445);
nand_4 g09874(new_n10260, new_n10259, new_n1270);
nand_4 g09875(new_n10261, new_n10260, new_n1265_1);
nand_4 g09876(new_n10262, new_n10261, n8649);
nor_4  g09877(n11122, new_n10262, new_n898);
nand_4 g09878(new_n10264, new_n1273, new_n880);
nand_4 g09879(new_n10265, new_n10264, new_n1445);
nand_4 g09880(new_n10266, new_n10265, new_n1270);
nand_4 g09881(new_n10267, new_n10266, new_n1265_1);
nand_4 g09882(new_n10268, new_n10267, new_n1260);
nand_4 g09883(new_n10269, new_n10268, new_n1256);
nand_4 g09884(new_n10270, new_n10269, new_n1251);
nand_4 g09885(new_n10271, new_n10270, new_n1457);
nand_4 g09886(new_n10272, new_n10271, new_n1462);
nand_4 g09887(new_n10273, new_n10272, new_n1468);
nand_4 g09888(new_n10274, new_n10273, new_n1247);
nand_4 g09889(new_n10275, new_n10274, new_n1474);
nand_4 g09890(new_n10276, new_n10275, new_n592);
nand_4 g09891(new_n10277, new_n10276, new_n585);
nand_4 g09892(new_n10278_1, new_n10277, new_n580);
nand_4 g09893(new_n10279, new_n10278_1, new_n600);
nand_4 g09894(new_n10280, new_n10279, new_n606);
nand_4 g09895(new_n10281, new_n10280, new_n612);
nand_4 g09896(new_n10282, new_n10281, new_n575);
nand_4 g09897(new_n10283_1, new_n10282, new_n619);
nand_4 g09898(new_n10284, new_n10283_1, new_n570);
nand_4 g09899(new_n10285, new_n10284, new_n625);
nand_4 g09900(new_n10286, new_n10285, new_n564);
nand_4 g09901(new_n10287, new_n10286, new_n632);
nand_4 g09902(new_n10288, new_n10287, new_n638);
nand_4 g09903(new_n10289, new_n10288, new_n559);
nand_4 g09904(new_n10290, new_n10289, new_n554);
nand_4 g09905(new_n10291, new_n10290, new_n646);
nand_4 g09906(new_n10292, new_n10291, new_n652);
nand_4 g09907(new_n10293, new_n10292, new_n549);
nand_4 g09908(new_n10294, new_n10293, new_n544);
nand_4 g09909(new_n10295, new_n10294, new_n660);
nand_4 g09910(new_n10296, new_n10295, new_n539);
nand_4 g09911(new_n10297, new_n10296, new_n534);
nand_4 g09912(new_n10298, new_n10297, new_n529);
nand_4 g09913(new_n10299, new_n10298, new_n668);
nand_4 g09914(new_n10300, new_n10299, new_n674_1);
nand_4 g09915(new_n10301, new_n10300, new_n681);
nand_4 g09916(new_n10302, new_n10301, new_n523);
nand_4 g09917(new_n10303, new_n10302, new_n687);
nand_4 g09918(new_n10304, new_n10303, new_n693);
nand_4 g09919(new_n10305, new_n10304, new_n699);
nand_4 g09920(new_n10306, new_n10305, new_n517);
nand_4 g09921(new_n10307, new_n10306, new_n705);
nand_4 g09922(new_n10308, new_n10307, new_n511);
nand_4 g09923(new_n10309, new_n10308, new_n711);
nand_4 g09924(new_n10310, new_n10309, new_n506);
nand_4 g09925(new_n10311, new_n10310, new_n719);
nand_4 g09926(new_n10312, new_n10311, new_n500);
nand_4 g09927(new_n10313, new_n10312, new_n727);
not_3  g09928(new_n10314, new_n10313);
nor_4  g09929(new_n10315, new_n10314, new_n495);
nor_4  g09930(new_n10316, new_n10315, new_n736);
nor_4  g09931(new_n10317, new_n10316, new_n489);
nor_4  g09932(new_n10318, new_n10317, new_n744);
nor_4  g09933(new_n10319, new_n10318, new_n483);
nor_4  g09934(new_n10320, new_n10319, new_n752);
nor_4  g09935(new_n10321, new_n10320, new_n759);
nor_4  g09936(new_n10322, new_n10321, new_n766);
nor_4  g09937(new_n10323, new_n10322, new_n477);
nor_4  g09938(new_n10324, new_n10323, new_n774);
nor_4  g09939(new_n10325, new_n10324, new_n781);
nor_4  g09940(new_n10326, new_n10325, new_n788);
nor_4  g09941(new_n10327, new_n10326, new_n471);
nor_4  g09942(new_n10328, new_n10327, new_n796);
nor_4  g09943(new_n10329, new_n10328, new_n804);
nor_4  g09944(new_n10330, new_n10329, new_n810);
nor_4  g09945(new_n10331, new_n10330, new_n2043);
nor_4  g09946(new_n10332, new_n10331, new_n2042);
nor_4  g09947(new_n10333, new_n10332, new_n2041);
nor_4  g09948(new_n10334, new_n10333, new_n2040);
nor_4  g09949(new_n10335, new_n10334, new_n2039);
nor_4  g09950(new_n10336, new_n10335, new_n2038);
nor_4  g09951(new_n10337, new_n10336, new_n2037);
nor_4  g09952(new_n10338, new_n10337, new_n2036);
nor_4  g09953(new_n10339, new_n10338, new_n2035);
not_3  g09954(new_n10340, new_n10339);
nand_4 g09955(new_n10341, new_n10340, new_n841);
nand_4 g09956(new_n10342, new_n10341, new_n434);
nand_4 g09957(new_n10343, new_n10342, new_n429);
nand_4 g09958(new_n10344, new_n10343, new_n424);
nand_4 g09959(new_n10345, new_n10344, new_n850);
nand_4 g09960(new_n10346, new_n10345, new_n856);
nand_4 g09961(new_n10347, new_n10346, new_n863);
nand_4 g09962(new_n10348, new_n10347, new_n419);
nand_4 g09963(new_n10349, new_n10348, new_n869);
nand_4 g09964(new_n10350, new_n10349, n7748);
nor_4  g09965(n11393, new_n10350, new_n1782);
nand_4 g09966(new_n10352, new_n860, new_n419);
nand_4 g09967(new_n10353, new_n10352, new_n869);
nand_4 g09968(new_n10354, new_n10353, new_n875);
nand_4 g09969(new_n10355, new_n10354, new_n881);
nand_4 g09970(new_n10356, new_n10355, new_n413);
nand_4 g09971(new_n10357, new_n10356, new_n889);
nand_4 g09972(new_n10358, new_n10357, new_n896);
nand_4 g09973(new_n10359, new_n10358, new_n901);
nand_4 g09974(new_n10360, new_n10359, new_n408);
nand_4 g09975(new_n10361, new_n10360, new_n908);
nand_4 g09976(new_n10362, new_n10361, new_n403);
nand_4 g09977(new_n10363, new_n10362, new_n398);
nand_4 g09978(new_n10364, new_n10363, new_n393);
nand_4 g09979(new_n10365, new_n10364, new_n916);
nand_4 g09980(new_n10366, new_n10365, new_n1123);
nand_4 g09981(new_n10367, new_n10366, new_n1164);
nand_4 g09982(new_n10368, new_n10367, new_n1120);
nand_4 g09983(new_n10369, new_n10368, new_n1169);
nand_4 g09984(new_n10370, new_n10369, new_n1116);
nand_4 g09985(new_n10371, new_n10370, new_n1111);
nand_4 g09986(new_n10372, new_n10371, new_n1106);
nand_4 g09987(new_n10373, new_n10372, new_n1178);
nand_4 g09988(new_n10374, new_n10373, new_n1183);
nand_4 g09989(new_n10375, new_n10374, new_n1102);
nand_4 g09990(new_n10376, new_n10375, new_n1099);
nand_4 g09991(new_n10377, new_n10376, new_n1191);
nand_4 g09992(new_n10378_1, new_n10377, new_n1095);
nand_4 g09993(new_n10379, new_n10378_1, new_n1091);
nand_4 g09994(new_n10380, new_n10379, new_n1088);
nand_4 g09995(new_n10381, new_n10380, new_n1084);
nand_4 g09996(new_n10382, new_n10381, new_n1079);
nand_4 g09997(new_n10383, new_n10382, new_n1074);
nand_4 g09998(new_n10384, new_n10383, new_n1070);
nand_4 g09999(new_n10385, new_n10384, new_n1064);
nand_4 g10000(new_n10386, new_n10385, new_n1061);
nand_4 g10001(new_n10387, new_n10386, new_n1055);
nand_4 g10002(new_n10388, new_n10387, new_n1050);
nand_4 g10003(new_n10389, new_n10388, new_n1045);
nand_4 g10004(new_n10390, new_n10389, new_n1041);
nand_4 g10005(new_n10391, new_n10390, new_n1036);
nand_4 g10006(new_n10392, new_n10391, new_n1031);
nand_4 g10007(new_n10393, new_n10392, new_n1025);
nand_4 g10008(new_n10394, new_n10393, new_n1020);
nand_4 g10009(new_n10395, new_n10394, new_n1015);
nand_4 g10010(new_n10396, new_n10395, new_n1010);
nand_4 g10011(new_n10397, new_n10396, new_n1215);
nand_4 g10012(new_n10398, new_n10397, new_n1005);
nand_4 g10013(new_n10399, new_n10398, new_n1000);
nand_4 g10014(new_n10400, new_n10399, new_n994);
nand_4 g10015(new_n10401, new_n10400, new_n989);
nand_4 g10016(new_n10402, new_n10401, new_n984);
not_3  g10017(new_n10403, new_n10402);
nor_4  g10018(new_n10404, new_n10403, new_n979);
nor_4  g10019(new_n10405, new_n10404, new_n974);
nor_4  g10020(new_n10406, new_n10405, new_n968);
nor_4  g10021(new_n10407_1, new_n10406, new_n965);
nor_4  g10022(new_n10408, new_n10407_1, new_n961);
nor_4  g10023(new_n10409, new_n10408, new_n958);
nor_4  g10024(new_n10410, new_n10409, new_n953);
nor_4  g10025(new_n10411, new_n10410, new_n3536);
nor_4  g10026(new_n10412, new_n10411, new_n3535);
nor_4  g10027(new_n10413, new_n10412, new_n3534);
nor_4  g10028(new_n10414, new_n10413, new_n2520);
nor_4  g10029(new_n10415, new_n10414, new_n2519);
nor_4  g10030(new_n10416, new_n10415, new_n2518);
nor_4  g10031(new_n10417, new_n10416, new_n2517);
nor_4  g10032(new_n10418, new_n10417, new_n2516);
nor_4  g10033(new_n10419, new_n10418, new_n2515);
nor_4  g10034(new_n10420, new_n10419, new_n2514);
nor_4  g10035(new_n10421, new_n10420, new_n2513);
nor_4  g10036(new_n10422, new_n10421, new_n2512);
nor_4  g10037(new_n10423, new_n10422, new_n2511);
nor_4  g10038(new_n10424, new_n10423, new_n2510);
nor_4  g10039(new_n10425, new_n10424, new_n2509);
nor_4  g10040(new_n10426_1, new_n10425, new_n2508);
nor_4  g10041(new_n10427, new_n10426_1, new_n2507);
nor_4  g10042(new_n10428, new_n10427, new_n2506);
nor_4  g10043(new_n10429, new_n10428, new_n2505);
nor_4  g10044(new_n10430, new_n10429, new_n2504);
not_3  g10045(new_n10431, new_n10430);
nand_4 g10046(new_n10432, new_n10431, new_n2147);
nand_4 g10047(new_n10433, new_n10432, new_n1810);
nand_4 g10048(new_n10434, new_n10433, new_n1806);
nand_4 g10049(new_n10435, new_n10434, new_n1802);
nand_4 g10050(new_n10436, new_n10435, new_n1798);
nand_4 g10051(new_n10437, new_n10436, new_n1820);
nand_4 g10052(new_n10438, new_n10437, n13364);
nor_4  g10053(n11463, new_n10438, new_n1791);
nand_4 g10054(new_n10440, new_n966, new_n492);
nand_4 g10055(new_n10441, new_n10440, new_n735);
nand_4 g10056(new_n10442, new_n10441, new_n488);
nand_4 g10057(new_n10443, new_n10442, new_n743);
nand_4 g10058(new_n10444, new_n10443, new_n482);
nand_4 g10059(new_n10445, new_n10444, new_n751);
nand_4 g10060(new_n10446_1, new_n10445, new_n758);
nand_4 g10061(new_n10447, new_n10446_1, new_n765);
nand_4 g10062(new_n10448, new_n10447, new_n476);
nand_4 g10063(new_n10449, new_n10448, new_n773);
nand_4 g10064(new_n10450, new_n10449, new_n780);
nand_4 g10065(new_n10451, new_n10450, new_n787);
nand_4 g10066(new_n10452, new_n10451, new_n470);
nand_4 g10067(new_n10453, new_n10452, new_n795);
nand_4 g10068(new_n10454, new_n10453, new_n803);
nand_4 g10069(new_n10455, new_n10454, new_n809);
nand_4 g10070(new_n10456, new_n10455, new_n465);
nand_4 g10071(new_n10457, new_n10456, new_n818);
nand_4 g10072(new_n10458, new_n10457, new_n460);
nand_4 g10073(new_n10459, new_n10458, new_n455);
nand_4 g10074(new_n10460, new_n10459, new_n449);
nand_4 g10075(new_n10461, new_n10460, new_n827);
nand_4 g10076(new_n10462, new_n10461, new_n833);
nand_4 g10077(new_n10463, new_n10462, new_n444);
nand_4 g10078(new_n10464, new_n10463, new_n439);
nand_4 g10079(new_n10465, new_n10464, new_n841);
nand_4 g10080(new_n10466_1, new_n10465, new_n434);
nand_4 g10081(new_n10467, new_n10466_1, new_n429);
nand_4 g10082(new_n10468, new_n10467, new_n424);
nand_4 g10083(new_n10469, new_n10468, new_n850);
nand_4 g10084(new_n10470_1, new_n10469, new_n856);
nand_4 g10085(new_n10471, new_n10470_1, new_n863);
nand_4 g10086(new_n10472, new_n10471, new_n419);
nand_4 g10087(new_n10473, new_n10472, new_n869);
nand_4 g10088(new_n10474, new_n10473, new_n875);
nand_4 g10089(new_n10475, new_n10474, new_n881);
nand_4 g10090(new_n10476, new_n10475, new_n413);
nand_4 g10091(new_n10477, new_n10476, new_n889);
nand_4 g10092(new_n10478, new_n10477, new_n896);
nand_4 g10093(new_n10479, new_n10478, new_n901);
nand_4 g10094(new_n10480, new_n10479, new_n408);
nand_4 g10095(new_n10481, new_n10480, new_n908);
nand_4 g10096(new_n10482, new_n10481, new_n403);
nand_4 g10097(new_n10483, new_n10482, new_n398);
nand_4 g10098(new_n10484, new_n10483, new_n393);
nand_4 g10099(new_n10485, new_n10484, new_n916);
not_3  g10100(new_n10486, new_n10485);
nor_4  g10101(new_n10487, new_n10486, new_n1532);
nor_4  g10102(new_n10488, new_n10487, new_n1531);
nor_4  g10103(new_n10489, new_n10488, new_n1530);
nor_4  g10104(new_n10490, new_n10489, new_n1529);
nor_4  g10105(new_n10491, new_n10490, new_n1528);
nor_4  g10106(new_n10492, new_n10491, new_n1527);
nor_4  g10107(new_n10493, new_n10492, new_n1526);
nor_4  g10108(new_n10494, new_n10493, new_n1525);
nor_4  g10109(new_n10495, new_n10494, new_n1524);
nor_4  g10110(new_n10496, new_n10495, new_n1523);
nor_4  g10111(new_n10497, new_n10496, new_n1522);
nor_4  g10112(new_n10498, new_n10497, new_n1521);
nor_4  g10113(new_n10499, new_n10498, new_n1520);
nor_4  g10114(new_n10500, new_n10499, new_n1519);
nor_4  g10115(new_n10501, new_n10500, new_n1518);
nor_4  g10116(new_n10502, new_n10501, new_n1517);
nor_4  g10117(new_n10503, new_n10502, new_n1516);
nor_4  g10118(new_n10504, new_n10503, new_n1075);
nor_4  g10119(new_n10505, new_n10504, new_n1071);
nor_4  g10120(new_n10506, new_n10505, new_n1065);
nor_4  g10121(new_n10507, new_n10506, new_n1062);
nor_4  g10122(new_n10508, new_n10507, new_n1056);
nor_4  g10123(new_n10509, new_n10508, new_n1051);
nor_4  g10124(new_n10510, new_n10509, new_n1046);
not_3  g10125(new_n10511, new_n10510);
nand_4 g10126(new_n10512, new_n10511, new_n1041);
nand_4 g10127(new_n10513, new_n10512, new_n1036);
nand_4 g10128(new_n10514, new_n10513, new_n1031);
nand_4 g10129(new_n10515_1, new_n10514, new_n1025);
nand_4 g10130(new_n10516, new_n10515_1, new_n1020);
nand_4 g10131(new_n10517, new_n10516, new_n1015);
nand_4 g10132(new_n10518, new_n10517, new_n1010);
nand_4 g10133(new_n10519, new_n10518, new_n1215);
nand_4 g10134(new_n10520, new_n10519, new_n1005);
nand_4 g10135(new_n10521, new_n10520, new_n1000);
nand_4 g10136(new_n10522, new_n10521, new_n994);
nand_4 g10137(new_n10523, new_n10522, new_n989);
nand_4 g10138(new_n10524, new_n10523, new_n984);
nand_4 g10139(new_n10525, new_n10524, new_n978);
nand_4 g10140(new_n10526, new_n10525, n6436);
nor_4  g10141(n11534, new_n10526, new_n970);
nand_4 g10142(new_n10528, new_n1282, new_n868);
nand_4 g10143(new_n10529, new_n10528, new_n1280);
nand_4 g10144(new_n10530, new_n10529, new_n1275);
nand_4 g10145(new_n10531, new_n10530, new_n1445);
nand_4 g10146(new_n10532, new_n10531, new_n1270);
nand_4 g10147(new_n10533, new_n10532, new_n1265_1);
nand_4 g10148(new_n10534, new_n10533, new_n1260);
nand_4 g10149(new_n10535, new_n10534, new_n1256);
nand_4 g10150(new_n10536, new_n10535, new_n1251);
nand_4 g10151(new_n10537, new_n10536, new_n1457);
nand_4 g10152(new_n10538, new_n10537, new_n1462);
nand_4 g10153(new_n10539, new_n10538, new_n1468);
nand_4 g10154(new_n10540, new_n10539, new_n1247);
nand_4 g10155(new_n10541, new_n10540, new_n1474);
nand_4 g10156(new_n10542, new_n10541, new_n592);
nand_4 g10157(new_n10543, new_n10542, new_n585);
nand_4 g10158(new_n10544, new_n10543, new_n580);
nand_4 g10159(new_n10545, new_n10544, new_n600);
nand_4 g10160(new_n10546, new_n10545, new_n606);
nand_4 g10161(new_n10547, new_n10546, new_n612);
nand_4 g10162(new_n10548, new_n10547, new_n575);
nand_4 g10163(new_n10549, new_n10548, new_n619);
nand_4 g10164(new_n10550, new_n10549, new_n570);
nand_4 g10165(new_n10551, new_n10550, new_n625);
nand_4 g10166(new_n10552, new_n10551, new_n564);
nand_4 g10167(new_n10553, new_n10552, new_n632);
nand_4 g10168(new_n10554, new_n10553, new_n638);
nand_4 g10169(new_n10555, new_n10554, new_n559);
nand_4 g10170(new_n10556, new_n10555, new_n554);
nand_4 g10171(new_n10557, new_n10556, new_n646);
nand_4 g10172(new_n10558, new_n10557, new_n652);
nand_4 g10173(new_n10559, new_n10558, new_n549);
nand_4 g10174(new_n10560, new_n10559, new_n544);
nand_4 g10175(new_n10561, new_n10560, new_n660);
nand_4 g10176(new_n10562, new_n10561, new_n539);
nand_4 g10177(new_n10563, new_n10562, new_n534);
nand_4 g10178(new_n10564, new_n10563, new_n529);
nand_4 g10179(new_n10565, new_n10564, new_n668);
nand_4 g10180(new_n10566, new_n10565, new_n674_1);
nand_4 g10181(new_n10567, new_n10566, new_n681);
nand_4 g10182(new_n10568, new_n10567, new_n523);
nand_4 g10183(new_n10569, new_n10568, new_n687);
nand_4 g10184(new_n10570, new_n10569, new_n693);
nand_4 g10185(new_n10571, new_n10570, new_n699);
nand_4 g10186(new_n10572, new_n10571, new_n517);
nand_4 g10187(new_n10573_1, new_n10572, new_n705);
nand_4 g10188(new_n10574, new_n10573_1, new_n511);
nand_4 g10189(new_n10575, new_n10574, new_n711);
nand_4 g10190(new_n10576, new_n10575, new_n506);
nand_4 g10191(new_n10577, new_n10576, new_n719);
nand_4 g10192(new_n10578, new_n10577, new_n500);
not_3  g10193(new_n10579, new_n10578);
nor_4  g10194(new_n10580, new_n10579, new_n728);
nor_4  g10195(new_n10581, new_n10580, new_n495);
nor_4  g10196(new_n10582, new_n10581, new_n736);
nor_4  g10197(new_n10583, new_n10582, new_n489);
nor_4  g10198(new_n10584, new_n10583, new_n744);
nor_4  g10199(new_n10585, new_n10584, new_n483);
nor_4  g10200(new_n10586, new_n10585, new_n752);
nor_4  g10201(new_n10587, new_n10586, new_n759);
nor_4  g10202(new_n10588, new_n10587, new_n766);
nor_4  g10203(new_n10589, new_n10588, new_n477);
nor_4  g10204(new_n10590, new_n10589, new_n774);
nor_4  g10205(new_n10591_1, new_n10590, new_n781);
nor_4  g10206(new_n10592, new_n10591_1, new_n788);
nor_4  g10207(new_n10593, new_n10592, new_n471);
nor_4  g10208(new_n10594, new_n10593, new_n796);
nor_4  g10209(new_n10595, new_n10594, new_n804);
nor_4  g10210(new_n10596, new_n10595, new_n810);
nor_4  g10211(new_n10597, new_n10596, new_n2043);
nor_4  g10212(new_n10598, new_n10597, new_n2042);
nor_4  g10213(new_n10599, new_n10598, new_n2041);
nor_4  g10214(new_n10600, new_n10599, new_n2040);
nor_4  g10215(new_n10601, new_n10600, new_n2039);
nor_4  g10216(new_n10602, new_n10601, new_n2038);
nor_4  g10217(new_n10603, new_n10602, new_n2037);
nor_4  g10218(new_n10604, new_n10603, new_n2036);
nor_4  g10219(new_n10605, new_n10604, new_n2035);
nor_4  g10220(new_n10606, new_n10605, new_n2034);
not_3  g10221(new_n10607, new_n10606);
nand_4 g10222(new_n10608, new_n10607, new_n434);
nand_4 g10223(new_n10609, new_n10608, new_n429);
nand_4 g10224(new_n10610, new_n10609, new_n424);
nand_4 g10225(new_n10611, new_n10610, new_n850);
nand_4 g10226(new_n10612, new_n10611, new_n856);
nand_4 g10227(new_n10613, new_n10612, new_n863);
nand_4 g10228(new_n10614, new_n10613, n9186);
nor_4  g10229(n11627, new_n10614, new_n415);
not_3  g10230(new_n10616, new_n509);
nand_4 g10231(new_n10617, new_n1642, new_n710);
nand_4 g10232(new_n10618, new_n10617, new_n1640);
nand_4 g10233(new_n10619, new_n10618, new_n1636);
nand_4 g10234(new_n10620, new_n10619, new_n1632);
nand_4 g10235(new_n10621, new_n10620, new_n1378);
nand_4 g10236(new_n10622, new_n10621, new_n1372);
nand_4 g10237(new_n10623, new_n10622, new_n1367);
nand_4 g10238(new_n10624, new_n10623, new_n1363);
nand_4 g10239(new_n10625, new_n10624, new_n1360);
nand_4 g10240(new_n10626, new_n10625, new_n1357);
nand_4 g10241(new_n10627, new_n10626, new_n1354);
nand_4 g10242(new_n10628, new_n10627, new_n1352);
nand_4 g10243(new_n10629, new_n10628, new_n1350);
nand_4 g10244(new_n10630_1, new_n10629, new_n1347_1);
nand_4 g10245(new_n10631, new_n10630_1, new_n1344);
nand_4 g10246(new_n10632, new_n10631, new_n1341);
nand_4 g10247(new_n10633, new_n10632, new_n1338);
nand_4 g10248(new_n10634, new_n10633, new_n1395);
nand_4 g10249(new_n10635, new_n10634, new_n1335);
nand_4 g10250(new_n10636, new_n10635, new_n1332);
nand_4 g10251(new_n10637, new_n10636, new_n1328);
nand_4 g10252(new_n10638, new_n10637, new_n1403);
nand_4 g10253(new_n10639, new_n10638, new_n1325);
nand_4 g10254(new_n10640, new_n10639, new_n1410);
nand_4 g10255(new_n10641, new_n10640, new_n1413);
nand_4 g10256(new_n10642, new_n10641, new_n1322);
nand_4 g10257(new_n10643, new_n10642, new_n1317);
nand_4 g10258(new_n10644, new_n10643, new_n1315);
nand_4 g10259(new_n10645, new_n10644, new_n1419);
nand_4 g10260(new_n10646, new_n10645, new_n1310);
nand_4 g10261(new_n10647, new_n10646, new_n1305);
nand_4 g10262(new_n10648, new_n10647, new_n1427);
nand_4 g10263(new_n10649, new_n10648, new_n1431);
nand_4 g10264(new_n10650, new_n10649, new_n1302);
nand_4 g10265(new_n10651, new_n10650, new_n1298);
nand_4 g10266(new_n10652, new_n10651, new_n1295);
nand_4 g10267(new_n10653, new_n10652, new_n1291);
nand_4 g10268(new_n10654, new_n10653, new_n1288);
nand_4 g10269(new_n10655, new_n10654, new_n1284);
nand_4 g10270(new_n10656, new_n10655, new_n1280);
nand_4 g10271(new_n10657, new_n10656, new_n1275);
nand_4 g10272(new_n10658, new_n10657, new_n1445);
nand_4 g10273(new_n10659, new_n10658, new_n1270);
nand_4 g10274(new_n10660, new_n10659, new_n1265_1);
nand_4 g10275(new_n10661, new_n10660, new_n1260);
nand_4 g10276(new_n10662, new_n10661, new_n1256);
nand_4 g10277(new_n10663, new_n10662, new_n1251);
nand_4 g10278(new_n10664, new_n10663, new_n1457);
nand_4 g10279(new_n10665, new_n10664, new_n1462);
nand_4 g10280(new_n10666, new_n10665, new_n1468);
nand_4 g10281(new_n10667, new_n10666, new_n1247);
not_3  g10282(new_n10668, new_n10667);
nor_4  g10283(new_n10669, new_n10668, new_n1475);
nor_4  g10284(new_n10670, new_n10669, new_n1244);
nor_4  g10285(new_n10671, new_n10670, new_n1243);
nor_4  g10286(new_n10672, new_n10671, new_n1242);
nor_4  g10287(new_n10673, new_n10672, new_n1241);
nor_4  g10288(new_n10674, new_n10673, new_n1240);
nor_4  g10289(new_n10675, new_n10674, new_n1239);
nor_4  g10290(new_n10676, new_n10675, new_n3082);
nor_4  g10291(new_n10677, new_n10676, new_n3081);
nor_4  g10292(new_n10678, new_n10677, new_n3080);
nor_4  g10293(new_n10679, new_n10678, new_n3079);
nor_4  g10294(new_n10680, new_n10679, new_n3078);
nor_4  g10295(new_n10681, new_n10680, new_n3077);
nor_4  g10296(new_n10682, new_n10681, new_n3076);
nor_4  g10297(new_n10683, new_n10682, new_n3075);
nor_4  g10298(new_n10684, new_n10683, new_n3074);
nor_4  g10299(new_n10685, new_n10684, new_n3073);
nor_4  g10300(new_n10686, new_n10685, new_n3072);
nor_4  g10301(new_n10687, new_n10686, new_n3071);
nor_4  g10302(new_n10688, new_n10687, new_n3070);
nor_4  g10303(new_n10689, new_n10688, new_n3069);
nor_4  g10304(new_n10690, new_n10689, new_n3068);
nor_4  g10305(new_n10691, new_n10690, new_n3067);
nor_4  g10306(new_n10692, new_n10691, new_n3066);
nor_4  g10307(new_n10693, new_n10692, new_n3065);
nor_4  g10308(new_n10694, new_n10693, new_n3064);
nor_4  g10309(new_n10695, new_n10694, new_n3063);
not_3  g10310(new_n10696, new_n10695);
nand_4 g10311(new_n10697, new_n10696, new_n523);
nand_4 g10312(new_n10698, new_n10697, new_n687);
nand_4 g10313(new_n10699, new_n10698, new_n693);
nand_4 g10314(new_n10700, new_n10699, new_n699);
nand_4 g10315(new_n10701, new_n10700, new_n517);
nand_4 g10316(new_n10702, new_n10701, new_n705);
nand_4 g10317(new_n10703, new_n10702, n13814);
nor_4  g10318(n11664, new_n10703, new_n10616);
not_3  g10319(new_n10705, new_n1869);
nand_4 g10320(new_n10706, new_n1693, new_n1059);
nand_4 g10321(new_n10707, new_n10706, new_n1055);
nand_4 g10322(new_n10708, new_n10707, new_n1050);
nand_4 g10323(new_n10709, new_n10708, new_n1045);
nand_4 g10324(new_n10710, new_n10709, new_n1041);
nand_4 g10325(new_n10711, new_n10710, new_n1036);
nand_4 g10326(new_n10712, new_n10711, new_n1031);
nand_4 g10327(new_n10713, new_n10712, new_n1025);
nand_4 g10328(new_n10714, new_n10713, new_n1020);
nand_4 g10329(new_n10715, new_n10714, new_n1015);
nand_4 g10330(new_n10716, new_n10715, new_n1010);
nand_4 g10331(new_n10717, new_n10716, new_n1215);
nand_4 g10332(new_n10718, new_n10717, new_n1005);
nand_4 g10333(new_n10719, new_n10718, new_n1000);
nand_4 g10334(new_n10720, new_n10719, new_n994);
nand_4 g10335(new_n10721, new_n10720, new_n989);
nand_4 g10336(new_n10722, new_n10721, new_n984);
nand_4 g10337(new_n10723, new_n10722, new_n978);
nand_4 g10338(new_n10724, new_n10723, new_n973);
nand_4 g10339(new_n10725, new_n10724, new_n967);
nand_4 g10340(new_n10726, new_n10725, new_n964);
nand_4 g10341(new_n10727, new_n10726, new_n960);
nand_4 g10342(new_n10728, new_n10727, new_n957);
nand_4 g10343(new_n10729, new_n10728, new_n952);
nand_4 g10344(new_n10730, new_n10729, new_n948_1);
nand_4 g10345(new_n10731, new_n10730, new_n943);
nand_4 g10346(new_n10732, new_n10731, new_n938);
nand_4 g10347(new_n10733, new_n10732, new_n934);
nand_4 g10348(new_n10734, new_n10733, new_n929);
nand_4 g10349(new_n10735, new_n10734, new_n925);
nand_4 g10350(new_n10736_1, new_n10735, new_n2194);
nand_4 g10351(new_n10737, new_n10736_1, new_n2191);
nand_4 g10352(new_n10738, new_n10737, new_n2190);
nand_4 g10353(new_n10739, new_n10738, new_n2186);
nand_4 g10354(new_n10740, new_n10739, new_n2183);
nand_4 g10355(new_n10741, new_n10740, new_n2179);
nand_4 g10356(new_n10742, new_n10741, new_n2175_1);
nand_4 g10357(new_n10743, new_n10742, new_n2171);
nand_4 g10358(new_n10744, new_n10743, new_n2168);
nand_4 g10359(new_n10745, new_n10744, new_n2165);
nand_4 g10360(new_n10746, new_n10745, new_n2162);
nand_4 g10361(new_n10747, new_n10746, new_n2158);
not_3  g10362(new_n10748, new_n10747);
nor_4  g10363(new_n10749, new_n10748, new_n2505);
nor_4  g10364(new_n10750_1, new_n10749, new_n2504);
nor_4  g10365(new_n10751, new_n10750_1, new_n2503);
nor_4  g10366(new_n10752, new_n10751, new_n2502);
nor_4  g10367(new_n10753, new_n10752, new_n2790);
nor_4  g10368(new_n10754, new_n10753, new_n2789);
nor_4  g10369(new_n10755, new_n10754, new_n2788);
nor_4  g10370(new_n10756, new_n10755, new_n2305);
nor_4  g10371(new_n10757, new_n10756, new_n2304);
nor_4  g10372(new_n10758, new_n10757, new_n2303);
nor_4  g10373(new_n10759, new_n10758, new_n2302);
nor_4  g10374(new_n10760, new_n10759, new_n2301);
nor_4  g10375(new_n10761, new_n10760, new_n2300);
nor_4  g10376(new_n10762, new_n10761, new_n2299);
nor_4  g10377(new_n10763, new_n10762, new_n2298);
nor_4  g10378(new_n10764, new_n10763, new_n2297);
nor_4  g10379(new_n10765_1, new_n10764, new_n2296);
nor_4  g10380(new_n10766, new_n10765_1, new_n2295);
nor_4  g10381(new_n10767, new_n10766, new_n2294);
nor_4  g10382(new_n10768, new_n10767, new_n2293);
nor_4  g10383(new_n10769, new_n10768, new_n2292);
nor_4  g10384(new_n10770, new_n10769, new_n2291);
not_3  g10385(new_n10771, new_n10770);
nand_4 g10386(new_n10772, new_n10771, new_n1748);
nand_4 g10387(new_n10773, new_n10772, new_n1746);
nand_4 g10388(new_n10774, new_n10773, new_n1742);
nand_4 g10389(new_n10775, new_n10774, new_n1738);
nand_4 g10390(new_n10776, new_n10775, new_n1736);
nand_4 g10391(new_n10777, new_n10776, new_n1732);
nand_4 g10392(new_n10778, new_n10777, new_n1729);
nand_4 g10393(new_n10779, new_n10778, new_n1726);
nand_4 g10394(new_n10780, new_n10779, new_n1724);
nand_4 g10395(new_n10781, new_n10780, new_n1721);
nand_4 g10396(new_n10782, new_n10781, new_n1718);
nand_4 g10397(new_n10783, new_n10782, new_n1715);
nand_4 g10398(new_n10784, new_n10783, new_n1711);
nand_4 g10399(new_n10785, new_n10784, new_n1708);
nand_4 g10400(new_n10786, new_n10785, new_n1705);
nand_4 g10401(new_n10787, new_n10786, new_n1703);
nand_4 g10402(new_n10788, new_n10787, new_n1860);
nand_4 g10403(new_n10789, new_n10788, new_n1864);
nand_4 g10404(new_n10790, new_n10789, new_n1699);
nand_4 g10405(new_n10791_1, new_n10790, new_n1697);
nand_4 g10406(new_n10792, new_n10791_1, n8746);
nor_4  g10407(n11822, new_n10792, new_n10705);
not_3  g10408(new_n10794, new_n703);
nand_4 g10409(new_n10795, new_n1652, new_n10794);
nand_4 g10410(new_n10796, new_n10795, new_n1648);
nand_4 g10411(new_n10797, new_n10796, new_n1644);
nand_4 g10412(new_n10798, new_n10797, new_n1640);
nand_4 g10413(new_n10799, new_n10798, new_n1636);
nand_4 g10414(new_n10800, new_n10799, new_n1632);
nand_4 g10415(new_n10801, new_n10800, new_n1378);
nand_4 g10416(new_n10802_1, new_n10801, new_n1372);
nand_4 g10417(new_n10803, new_n10802_1, new_n1367);
nand_4 g10418(new_n10804, new_n10803, new_n1363);
nand_4 g10419(new_n10805, new_n10804, new_n1360);
nand_4 g10420(new_n10806, new_n10805, new_n1357);
nand_4 g10421(new_n10807, new_n10806, new_n1354);
nand_4 g10422(new_n10808, new_n10807, new_n1352);
nand_4 g10423(new_n10809, new_n10808, new_n1350);
nand_4 g10424(new_n10810, new_n10809, new_n1347_1);
nand_4 g10425(new_n10811, new_n10810, new_n1344);
nand_4 g10426(new_n10812, new_n10811, new_n1341);
nand_4 g10427(new_n10813, new_n10812, new_n1338);
nand_4 g10428(new_n10814, new_n10813, new_n1395);
nand_4 g10429(new_n10815, new_n10814, new_n1335);
nand_4 g10430(new_n10816, new_n10815, new_n1332);
nand_4 g10431(new_n10817, new_n10816, new_n1328);
nand_4 g10432(new_n10818, new_n10817, new_n1403);
nand_4 g10433(new_n10819, new_n10818, new_n1325);
nand_4 g10434(new_n10820, new_n10819, new_n1410);
nand_4 g10435(new_n10821, new_n10820, new_n1413);
nand_4 g10436(new_n10822, new_n10821, new_n1322);
nand_4 g10437(new_n10823, new_n10822, new_n1317);
nand_4 g10438(new_n10824, new_n10823, new_n1315);
nand_4 g10439(new_n10825, new_n10824, new_n1419);
nand_4 g10440(new_n10826, new_n10825, new_n1310);
nand_4 g10441(new_n10827, new_n10826, new_n1305);
nand_4 g10442(new_n10828, new_n10827, new_n1427);
nand_4 g10443(new_n10829, new_n10828, new_n1431);
nand_4 g10444(new_n10830, new_n10829, new_n1302);
nand_4 g10445(new_n10831, new_n10830, new_n1298);
nand_4 g10446(new_n10832, new_n10831, new_n1295);
nand_4 g10447(new_n10833, new_n10832, new_n1291);
nand_4 g10448(new_n10834, new_n10833, new_n1288);
nand_4 g10449(new_n10835, new_n10834, new_n1284);
nand_4 g10450(new_n10836, new_n10835, new_n1280);
nand_4 g10451(new_n10837, new_n10836, new_n1275);
nand_4 g10452(new_n10838, new_n10837, new_n1445);
nand_4 g10453(new_n10839, new_n10838, new_n1270);
nand_4 g10454(new_n10840, new_n10839, new_n1265_1);
not_3  g10455(new_n10841, new_n10840);
nor_4  g10456(new_n10842, new_n10841, new_n1261);
nor_4  g10457(new_n10843, new_n10842, new_n1257);
nor_4  g10458(new_n10844, new_n10843, new_n1252);
nor_4  g10459(new_n10845, new_n10844, new_n1458);
nor_4  g10460(new_n10846, new_n10845, new_n1463);
nor_4  g10461(new_n10847, new_n10846, new_n1469);
nor_4  g10462(new_n10848, new_n10847, new_n1248);
nor_4  g10463(new_n10849, new_n10848, new_n1475);
nor_4  g10464(new_n10850, new_n10849, new_n1244);
nor_4  g10465(new_n10851, new_n10850, new_n1243);
nor_4  g10466(new_n10852, new_n10851, new_n1242);
nor_4  g10467(new_n10853, new_n10852, new_n1241);
nor_4  g10468(new_n10854, new_n10853, new_n1240);
nor_4  g10469(new_n10855, new_n10854, new_n1239);
nor_4  g10470(new_n10856, new_n10855, new_n3082);
nor_4  g10471(new_n10857, new_n10856, new_n3081);
nor_4  g10472(new_n10858, new_n10857, new_n3080);
nor_4  g10473(new_n10859, new_n10858, new_n3079);
nor_4  g10474(new_n10860, new_n10859, new_n3078);
nor_4  g10475(new_n10861, new_n10860, new_n3077);
nor_4  g10476(new_n10862_1, new_n10861, new_n3076);
nor_4  g10477(new_n10863, new_n10862_1, new_n3075);
nor_4  g10478(new_n10864, new_n10863, new_n3074);
nor_4  g10479(new_n10865, new_n10864, new_n3073);
not_3  g10480(new_n10866, new_n10865);
nand_4 g10481(new_n10867, new_n10866, new_n652);
nand_4 g10482(new_n10868, new_n10867, new_n549);
nand_4 g10483(new_n10869, new_n10868, new_n544);
nand_4 g10484(new_n10870, new_n10869, new_n660);
nand_4 g10485(new_n10871, new_n10870, new_n539);
nand_4 g10486(new_n10872, new_n10871, new_n534);
nand_4 g10487(new_n10873, new_n10872, new_n529);
nand_4 g10488(new_n10874, new_n10873, new_n668);
nand_4 g10489(new_n10875, new_n10874, new_n674_1);
nand_4 g10490(new_n10876, new_n10875, new_n681);
nand_4 g10491(new_n10877, new_n10876, new_n523);
nand_4 g10492(new_n10878, new_n10877, new_n687);
nand_4 g10493(new_n10879, new_n10878, new_n693);
nand_4 g10494(new_n10880, new_n10879, new_n699);
nand_4 g10495(new_n10881, new_n10880, n203);
nor_4  g10496(n11847, new_n10881, new_n513);
nand_4 g10497(new_n10883, new_n1688, new_n659);
nand_4 g10498(new_n10884, new_n10883, new_n1878);
nand_4 g10499(new_n10885, new_n10884, new_n1882);
nand_4 g10500(new_n10886, new_n10885, new_n1686);
nand_4 g10501(new_n10887, new_n10886, new_n1682);
nand_4 g10502(new_n10888, new_n10887, new_n1678);
nand_4 g10503(new_n10889, new_n10888, new_n1674);
nand_4 g10504(new_n10890, new_n10889, new_n1890);
nand_4 g10505(new_n10891, new_n10890, new_n1669);
nand_4 g10506(new_n10892, new_n10891, new_n1665);
nand_4 g10507(new_n10893, new_n10892, new_n1661);
nand_4 g10508(new_n10894, new_n10893, new_n1657);
nand_4 g10509(new_n10895, new_n10894, new_n1652);
nand_4 g10510(new_n10896, new_n10895, new_n1648);
nand_4 g10511(new_n10897, new_n10896, new_n1644);
nand_4 g10512(new_n10898, new_n10897, new_n1640);
nand_4 g10513(new_n10899, new_n10898, new_n1636);
nand_4 g10514(new_n10900, new_n10899, new_n1632);
nand_4 g10515(new_n10901, new_n10900, new_n1378);
nand_4 g10516(new_n10902, new_n10901, new_n1372);
nand_4 g10517(new_n10903, new_n10902, new_n1367);
nand_4 g10518(new_n10904, new_n10903, new_n1363);
nand_4 g10519(new_n10905, new_n10904, new_n1360);
nand_4 g10520(new_n10906, new_n10905, new_n1357);
nand_4 g10521(new_n10907, new_n10906, new_n1354);
nand_4 g10522(new_n10908, new_n10907, new_n1352);
nand_4 g10523(new_n10909, new_n10908, new_n1350);
nand_4 g10524(new_n10910, new_n10909, new_n1347_1);
nand_4 g10525(new_n10911, new_n10910, new_n1344);
nand_4 g10526(new_n10912_1, new_n10911, new_n1341);
nand_4 g10527(new_n10913, new_n10912_1, new_n1338);
nand_4 g10528(new_n10914, new_n10913, new_n1395);
nand_4 g10529(new_n10915_1, new_n10914, new_n1335);
nand_4 g10530(new_n10916, new_n10915_1, new_n1332);
nand_4 g10531(new_n10917, new_n10916, new_n1328);
nand_4 g10532(new_n10918, new_n10917, new_n1403);
nand_4 g10533(new_n10919, new_n10918, new_n1325);
nand_4 g10534(new_n10920, new_n10919, new_n1410);
nand_4 g10535(new_n10921, new_n10920, new_n1413);
nand_4 g10536(new_n10922, new_n10921, new_n1322);
nand_4 g10537(new_n10923, new_n10922, new_n1317);
nand_4 g10538(new_n10924, new_n10923, new_n1315);
nand_4 g10539(new_n10925, new_n10924, new_n1419);
nand_4 g10540(new_n10926, new_n10925, new_n1310);
nand_4 g10541(new_n10927, new_n10926, new_n1305);
nand_4 g10542(new_n10928, new_n10927, new_n1427);
nand_4 g10543(new_n10929, new_n10928, new_n1431);
nand_4 g10544(new_n10930, new_n10929, new_n1302);
nand_4 g10545(new_n10931, new_n10930, new_n1298);
nand_4 g10546(new_n10932, new_n10931, new_n1295);
nand_4 g10547(new_n10933, new_n10932, new_n1291);
not_3  g10548(new_n10934, new_n10933);
nor_4  g10549(new_n10935, new_n10934, new_n2396);
nor_4  g10550(new_n10936, new_n10935, new_n2395);
nor_4  g10551(new_n10937, new_n10936, new_n1281);
nor_4  g10552(new_n10938, new_n10937, new_n1276);
nor_4  g10553(new_n10939, new_n10938, new_n1446);
nor_4  g10554(new_n10940, new_n10939, new_n1271);
nor_4  g10555(new_n10941, new_n10940, new_n1266);
nor_4  g10556(new_n10942, new_n10941, new_n1261);
nor_4  g10557(new_n10943, new_n10942, new_n1257);
nor_4  g10558(new_n10944, new_n10943, new_n1252);
nor_4  g10559(new_n10945_1, new_n10944, new_n1458);
nor_4  g10560(new_n10946, new_n10945_1, new_n1463);
nor_4  g10561(new_n10947, new_n10946, new_n1469);
nor_4  g10562(new_n10948, new_n10947, new_n1248);
nor_4  g10563(new_n10949, new_n10948, new_n1475);
nor_4  g10564(new_n10950, new_n10949, new_n1244);
nor_4  g10565(new_n10951, new_n10950, new_n1243);
nor_4  g10566(new_n10952, new_n10951, new_n1242);
nor_4  g10567(new_n10953, new_n10952, new_n1241);
nor_4  g10568(new_n10954, new_n10953, new_n1240);
nor_4  g10569(new_n10955, new_n10954, new_n1239);
nor_4  g10570(new_n10956, new_n10955, new_n3082);
nor_4  g10571(new_n10957, new_n10956, new_n3081);
nor_4  g10572(new_n10958, new_n10957, new_n3080);
nor_4  g10573(new_n10959, new_n10958, new_n3079);
nor_4  g10574(new_n10960, new_n10959, new_n3078);
nor_4  g10575(new_n10961, new_n10960, new_n3077);
not_3  g10576(new_n10962, new_n10961);
nand_4 g10577(new_n10963, new_n10962, new_n638);
nand_4 g10578(new_n10964, new_n10963, new_n559);
nand_4 g10579(new_n10965, new_n10964, new_n554);
nand_4 g10580(new_n10966, new_n10965, new_n646);
nand_4 g10581(new_n10967, new_n10966, new_n652);
nand_4 g10582(new_n10968, new_n10967, new_n549);
nand_4 g10583(new_n10969, new_n10968, n8550);
nor_4  g10584(n12032, new_n10969, new_n541);
nand_4 g10585(new_n10971, new_n1722, new_n611);
nand_4 g10586(new_n10972, new_n10971, new_n1721);
nand_4 g10587(new_n10973, new_n10972, new_n1718);
nand_4 g10588(new_n10974, new_n10973, new_n1715);
nand_4 g10589(new_n10975, new_n10974, new_n1711);
nand_4 g10590(new_n10976, new_n10975, new_n1708);
nand_4 g10591(new_n10977, new_n10976, new_n1705);
nand_4 g10592(new_n10978, new_n10977, new_n1703);
nand_4 g10593(new_n10979, new_n10978, new_n1860);
nand_4 g10594(new_n10980, new_n10979, new_n1864);
nand_4 g10595(new_n10981, new_n10980, new_n1699);
nand_4 g10596(new_n10982, new_n10981, new_n1697);
nand_4 g10597(new_n10983, new_n10982, new_n1871);
nand_4 g10598(new_n10984, new_n10983, new_n1694);
nand_4 g10599(new_n10985, new_n10984, new_n1690);
nand_4 g10600(new_n10986, new_n10985, new_n1878);
nand_4 g10601(new_n10987, new_n10986, new_n1882);
nand_4 g10602(new_n10988, new_n10987, new_n1686);
nand_4 g10603(new_n10989, new_n10988, new_n1682);
nand_4 g10604(new_n10990, new_n10989, new_n1678);
nand_4 g10605(new_n10991, new_n10990, new_n1674);
nand_4 g10606(new_n10992, new_n10991, new_n1890);
nand_4 g10607(new_n10993, new_n10992, new_n1669);
nand_4 g10608(new_n10994, new_n10993, new_n1665);
nand_4 g10609(new_n10995, new_n10994, new_n1661);
nand_4 g10610(new_n10996, new_n10995, new_n1657);
nand_4 g10611(new_n10997, new_n10996, new_n1652);
nand_4 g10612(new_n10998, new_n10997, new_n1648);
nand_4 g10613(new_n10999, new_n10998, new_n1644);
nand_4 g10614(new_n11000, new_n10999, new_n1640);
nand_4 g10615(new_n11001, new_n11000, new_n1636);
nand_4 g10616(new_n11002, new_n11001, new_n1632);
nand_4 g10617(new_n11003, new_n11002, new_n1378);
nand_4 g10618(new_n11004, new_n11003, new_n1372);
nand_4 g10619(new_n11005, new_n11004, new_n1367);
nand_4 g10620(new_n11006, new_n11005, new_n1363);
nand_4 g10621(new_n11007, new_n11006, new_n1360);
nand_4 g10622(new_n11008, new_n11007, new_n1357);
nand_4 g10623(new_n11009, new_n11008, new_n1354);
nand_4 g10624(new_n11010, new_n11009, new_n1352);
nand_4 g10625(new_n11011, new_n11010, new_n1350);
nand_4 g10626(new_n11012, new_n11011, new_n1347_1);
nand_4 g10627(new_n11013, new_n11012, new_n1344);
nand_4 g10628(new_n11014, new_n11013, new_n1341);
nand_4 g10629(new_n11015, new_n11014, new_n1338);
nand_4 g10630(new_n11016, new_n11015, new_n1395);
nand_4 g10631(new_n11017, new_n11016, new_n1335);
nand_4 g10632(new_n11018, new_n11017, new_n1332);
nand_4 g10633(new_n11019, new_n11018, new_n1328);
nand_4 g10634(new_n11020, new_n11019, new_n1403);
nand_4 g10635(new_n11021, new_n11020, new_n1325);
not_3  g10636(new_n11022, new_n11021);
nor_4  g10637(new_n11023, new_n11022, new_n2410);
nor_4  g10638(new_n11024, new_n11023, new_n2409);
nor_4  g10639(new_n11025, new_n11024, new_n2408);
nor_4  g10640(new_n11026, new_n11025, new_n2407_1);
nor_4  g10641(new_n11027, new_n11026, new_n2406);
nor_4  g10642(new_n11028, new_n11027, new_n2405);
nor_4  g10643(new_n11029, new_n11028, new_n2404);
nor_4  g10644(new_n11030, new_n11029, new_n2403);
nor_4  g10645(new_n11031, new_n11030, new_n2402);
nor_4  g10646(new_n11032, new_n11031, new_n2401);
nor_4  g10647(new_n11033, new_n11032, new_n2400);
nor_4  g10648(new_n11034, new_n11033, new_n2399);
nor_4  g10649(new_n11035, new_n11034, new_n2398);
nor_4  g10650(new_n11036, new_n11035, new_n2397);
nor_4  g10651(new_n11037, new_n11036, new_n2396);
nor_4  g10652(new_n11038, new_n11037, new_n2395);
nor_4  g10653(new_n11039, new_n11038, new_n1281);
nor_4  g10654(new_n11040, new_n11039, new_n1276);
nor_4  g10655(new_n11041, new_n11040, new_n1446);
nor_4  g10656(new_n11042, new_n11041, new_n1271);
nor_4  g10657(new_n11043, new_n11042, new_n1266);
nor_4  g10658(new_n11044, new_n11043, new_n1261);
nor_4  g10659(new_n11045, new_n11044, new_n1257);
nor_4  g10660(new_n11046, new_n11045, new_n1252);
nor_4  g10661(new_n11047, new_n11046, new_n1458);
nor_4  g10662(new_n11048, new_n11047, new_n1463);
nor_4  g10663(new_n11049, new_n11048, new_n1469);
not_3  g10664(new_n11050, new_n11049);
nand_4 g10665(new_n11051, new_n11050, new_n1247);
nand_4 g10666(new_n11052, new_n11051, new_n1474);
nand_4 g10667(new_n11053, new_n11052, new_n592);
nand_4 g10668(new_n11054, new_n11053, new_n585);
nand_4 g10669(new_n11055, new_n11054, new_n580);
nand_4 g10670(new_n11056, new_n11055, new_n600);
nand_4 g10671(new_n11057, new_n11056, n7354);
nor_4  g10672(n12166, new_n11057, new_n603);
nand_4 g10673(new_n11059, new_n1108, new_n1106);
nand_4 g10674(new_n11060, new_n11059, new_n1178);
nand_4 g10675(new_n11061, new_n11060, new_n1183);
nand_4 g10676(new_n11062, new_n11061, new_n1102);
nand_4 g10677(new_n11063, new_n11062, new_n1099);
nand_4 g10678(new_n11064, new_n11063, new_n1191);
nand_4 g10679(new_n11065, new_n11064, new_n1095);
nand_4 g10680(new_n11066, new_n11065, new_n1091);
nand_4 g10681(new_n11067, new_n11066, new_n1088);
nand_4 g10682(new_n11068, new_n11067, new_n1084);
nand_4 g10683(new_n11069, new_n11068, new_n1079);
nand_4 g10684(new_n11070, new_n11069, new_n1074);
nand_4 g10685(new_n11071, new_n11070, new_n1070);
nand_4 g10686(new_n11072, new_n11071, new_n1064);
nand_4 g10687(new_n11073, new_n11072, new_n1061);
nand_4 g10688(new_n11074, new_n11073, new_n1055);
nand_4 g10689(new_n11075, new_n11074, new_n1050);
nand_4 g10690(new_n11076, new_n11075, new_n1045);
nand_4 g10691(new_n11077, new_n11076, new_n1041);
nand_4 g10692(new_n11078, new_n11077, new_n1036);
nand_4 g10693(new_n11079, new_n11078, new_n1031);
nand_4 g10694(new_n11080, new_n11079, new_n1025);
nand_4 g10695(new_n11081, new_n11080, new_n1020);
nand_4 g10696(new_n11082, new_n11081, new_n1015);
nand_4 g10697(new_n11083, new_n11082, new_n1010);
nand_4 g10698(new_n11084, new_n11083, new_n1215);
nand_4 g10699(new_n11085, new_n11084, new_n1005);
nand_4 g10700(new_n11086, new_n11085, new_n1000);
nand_4 g10701(new_n11087, new_n11086, new_n994);
nand_4 g10702(new_n11088, new_n11087, new_n989);
nand_4 g10703(new_n11089, new_n11088, new_n984);
nand_4 g10704(new_n11090, new_n11089, new_n978);
nand_4 g10705(new_n11091, new_n11090, new_n973);
nand_4 g10706(new_n11092, new_n11091, new_n967);
nand_4 g10707(new_n11093, new_n11092, new_n964);
nand_4 g10708(new_n11094, new_n11093, new_n960);
nand_4 g10709(new_n11095, new_n11094, new_n957);
nand_4 g10710(new_n11096, new_n11095, new_n952);
nand_4 g10711(new_n11097, new_n11096, new_n948_1);
nand_4 g10712(new_n11098, new_n11097, new_n943);
nand_4 g10713(new_n11099, new_n11098, new_n938);
nand_4 g10714(new_n11100, new_n11099, new_n934);
nand_4 g10715(new_n11101, new_n11100, new_n929);
nand_4 g10716(new_n11102, new_n11101, new_n925);
nand_4 g10717(new_n11103, new_n11102, new_n2194);
nand_4 g10718(new_n11104, new_n11103, new_n2191);
not_3  g10719(new_n11105, new_n11104);
nor_4  g10720(new_n11106, new_n11105, new_n2515);
nor_4  g10721(new_n11107, new_n11106, new_n2514);
nor_4  g10722(new_n11108, new_n11107, new_n2513);
nor_4  g10723(new_n11109, new_n11108, new_n2512);
nor_4  g10724(new_n11110, new_n11109, new_n2511);
nor_4  g10725(new_n11111, new_n11110, new_n2510);
nor_4  g10726(new_n11112, new_n11111, new_n2509);
nor_4  g10727(new_n11113, new_n11112, new_n2508);
nor_4  g10728(new_n11114, new_n11113, new_n2507);
nor_4  g10729(new_n11115, new_n11114, new_n2506);
nor_4  g10730(new_n11116, new_n11115, new_n2505);
nor_4  g10731(new_n11117, new_n11116, new_n2504);
nor_4  g10732(new_n11118, new_n11117, new_n2503);
nor_4  g10733(new_n11119, new_n11118, new_n2502);
nor_4  g10734(new_n11120, new_n11119, new_n2790);
nor_4  g10735(new_n11121, new_n11120, new_n2789);
nor_4  g10736(new_n11122_1, new_n11121, new_n2788);
nor_4  g10737(new_n11123, new_n11122_1, new_n2305);
nor_4  g10738(new_n11124, new_n11123, new_n2304);
nor_4  g10739(new_n11125, new_n11124, new_n2303);
nor_4  g10740(new_n11126, new_n11125, new_n2302);
nor_4  g10741(new_n11127, new_n11126, new_n2301);
nor_4  g10742(new_n11128, new_n11127, new_n2300);
nor_4  g10743(new_n11129, new_n11128, new_n2299);
not_3  g10744(new_n11130, new_n11129);
nand_4 g10745(new_n11131, new_n11130, new_n1774);
nand_4 g10746(new_n11132, new_n11131, new_n1834);
nand_4 g10747(new_n11133, new_n11132, new_n1769);
nand_4 g10748(new_n11134, new_n11133, new_n1766);
nand_4 g10749(new_n11135, new_n11134, new_n1762);
nand_4 g10750(new_n11136, new_n11135, new_n1758);
nand_4 g10751(new_n11137, new_n11136, new_n1754);
nand_4 g10752(new_n11138, new_n11137, new_n1751);
nand_4 g10753(new_n11139, new_n11138, new_n1748);
nand_4 g10754(new_n11140, new_n11139, new_n1746);
nand_4 g10755(new_n11141, new_n11140, new_n1742);
nand_4 g10756(new_n11142, new_n11141, new_n1738);
nand_4 g10757(new_n11143_1, new_n11142, new_n1736);
nand_4 g10758(new_n11144, new_n11143_1, new_n1732);
nand_4 g10759(new_n11145, new_n11144, n13102);
nor_4  g10760(n12232, new_n11145, new_n597);
nand_4 g10761(new_n11147, new_n1296, new_n849);
nand_4 g10762(new_n11148, new_n11147, new_n1295);
nand_4 g10763(new_n11149, new_n11148, new_n1291);
nand_4 g10764(new_n11150, new_n11149, new_n1288);
nand_4 g10765(new_n11151, new_n11150, new_n1284);
nand_4 g10766(new_n11152, new_n11151, new_n1280);
nand_4 g10767(new_n11153, new_n11152, new_n1275);
nand_4 g10768(new_n11154, new_n11153, new_n1445);
nand_4 g10769(new_n11155, new_n11154, new_n1270);
nand_4 g10770(new_n11156, new_n11155, new_n1265_1);
nand_4 g10771(new_n11157, new_n11156, new_n1260);
nand_4 g10772(new_n11158_1, new_n11157, new_n1256);
nand_4 g10773(new_n11159, new_n11158_1, new_n1251);
nand_4 g10774(new_n11160, new_n11159, new_n1457);
nand_4 g10775(new_n11161, new_n11160, new_n1462);
nand_4 g10776(new_n11162, new_n11161, new_n1468);
nand_4 g10777(new_n11163, new_n11162, new_n1247);
nand_4 g10778(new_n11164, new_n11163, new_n1474);
nand_4 g10779(new_n11165, new_n11164, new_n592);
nand_4 g10780(new_n11166, new_n11165, new_n585);
nand_4 g10781(new_n11167, new_n11166, new_n580);
nand_4 g10782(new_n11168, new_n11167, new_n600);
nand_4 g10783(new_n11169, new_n11168, new_n606);
nand_4 g10784(new_n11170, new_n11169, new_n612);
nand_4 g10785(new_n11171, new_n11170, new_n575);
nand_4 g10786(new_n11172, new_n11171, new_n619);
nand_4 g10787(new_n11173, new_n11172, new_n570);
nand_4 g10788(new_n11174, new_n11173, new_n625);
nand_4 g10789(new_n11175, new_n11174, new_n564);
nand_4 g10790(new_n11176, new_n11175, new_n632);
nand_4 g10791(new_n11177, new_n11176, new_n638);
nand_4 g10792(new_n11178, new_n11177, new_n559);
nand_4 g10793(new_n11179, new_n11178, new_n554);
nand_4 g10794(new_n11180, new_n11179, new_n646);
nand_4 g10795(new_n11181, new_n11180, new_n652);
nand_4 g10796(new_n11182, new_n11181, new_n549);
nand_4 g10797(new_n11183, new_n11182, new_n544);
nand_4 g10798(new_n11184, new_n11183, new_n660);
nand_4 g10799(new_n11185, new_n11184, new_n539);
nand_4 g10800(new_n11186, new_n11185, new_n534);
nand_4 g10801(new_n11187, new_n11186, new_n529);
nand_4 g10802(new_n11188, new_n11187, new_n668);
nand_4 g10803(new_n11189, new_n11188, new_n674_1);
nand_4 g10804(new_n11190, new_n11189, new_n681);
nand_4 g10805(new_n11191, new_n11190, new_n523);
nand_4 g10806(new_n11192, new_n11191, new_n687);
not_3  g10807(new_n11193, new_n11192);
nor_4  g10808(new_n11194, new_n11193, new_n3354);
nor_4  g10809(new_n11195, new_n11194, new_n3353);
nor_4  g10810(new_n11196, new_n11195, new_n3352);
nor_4  g10811(new_n11197, new_n11196, new_n3351);
nor_4  g10812(new_n11198, new_n11197, new_n3350);
nor_4  g10813(new_n11199, new_n11198, new_n3349);
nor_4  g10814(new_n11200, new_n11199, new_n3348);
nor_4  g10815(new_n11201, new_n11200, new_n720);
nor_4  g10816(new_n11202, new_n11201, new_n501);
nor_4  g10817(new_n11203, new_n11202, new_n728);
nor_4  g10818(new_n11204, new_n11203, new_n495);
nor_4  g10819(new_n11205, new_n11204, new_n736);
nor_4  g10820(new_n11206, new_n11205, new_n489);
nor_4  g10821(new_n11207, new_n11206, new_n744);
nor_4  g10822(new_n11208, new_n11207, new_n483);
nor_4  g10823(new_n11209, new_n11208, new_n752);
nor_4  g10824(new_n11210, new_n11209, new_n759);
nor_4  g10825(new_n11211, new_n11210, new_n766);
nor_4  g10826(new_n11212, new_n11211, new_n477);
nor_4  g10827(new_n11213, new_n11212, new_n774);
nor_4  g10828(new_n11214, new_n11213, new_n781);
nor_4  g10829(new_n11215, new_n11214, new_n788);
nor_4  g10830(new_n11216, new_n11215, new_n471);
nor_4  g10831(new_n11217, new_n11216, new_n796);
not_3  g10832(new_n11218, new_n11217);
nand_4 g10833(new_n11219, new_n11218, new_n803);
nand_4 g10834(new_n11220, new_n11219, new_n809);
nand_4 g10835(new_n11221, new_n11220, new_n465);
nand_4 g10836(new_n11222, new_n11221, new_n818);
nand_4 g10837(new_n11223, new_n11222, new_n460);
nand_4 g10838(new_n11224, new_n11223, new_n455);
nand_4 g10839(new_n11225, new_n11224, new_n449);
nand_4 g10840(new_n11226, new_n11225, new_n827);
nand_4 g10841(new_n11227, new_n11226, new_n833);
nand_4 g10842(new_n11228, new_n11227, new_n444);
nand_4 g10843(new_n11229, new_n11228, new_n439);
nand_4 g10844(new_n11230, new_n11229, new_n841);
nand_4 g10845(new_n11231, new_n11230, new_n434);
nand_4 g10846(new_n11232, new_n11231, new_n429);
nand_4 g10847(new_n11233, new_n11232, n14464);
nor_4  g10848(n12355, new_n11233, new_n421);
nand_4 g10849(new_n11235, new_n1737, new_n1118);
nand_4 g10850(new_n11236, new_n11235, new_n1169);
nand_4 g10851(new_n11237, new_n11236, new_n1116);
nand_4 g10852(new_n11238, new_n11237, new_n1111);
nand_4 g10853(new_n11239, new_n11238, new_n1106);
nand_4 g10854(new_n11240, new_n11239, new_n1178);
nand_4 g10855(new_n11241, new_n11240, new_n1183);
nand_4 g10856(new_n11242, new_n11241, new_n1102);
nand_4 g10857(new_n11243, new_n11242, new_n1099);
nand_4 g10858(new_n11244, new_n11243, new_n1191);
nand_4 g10859(new_n11245, new_n11244, new_n1095);
nand_4 g10860(new_n11246, new_n11245, new_n1091);
nand_4 g10861(new_n11247, new_n11246, new_n1088);
nand_4 g10862(new_n11248, new_n11247, new_n1084);
nand_4 g10863(new_n11249, new_n11248, new_n1079);
nand_4 g10864(new_n11250, new_n11249, new_n1074);
nand_4 g10865(new_n11251, new_n11250, new_n1070);
nand_4 g10866(new_n11252, new_n11251, new_n1064);
nand_4 g10867(new_n11253, new_n11252, new_n1061);
nand_4 g10868(new_n11254, new_n11253, new_n1055);
nand_4 g10869(new_n11255, new_n11254, new_n1050);
nand_4 g10870(new_n11256, new_n11255, new_n1045);
nand_4 g10871(new_n11257, new_n11256, new_n1041);
nand_4 g10872(new_n11258, new_n11257, new_n1036);
nand_4 g10873(new_n11259, new_n11258, new_n1031);
nand_4 g10874(new_n11260, new_n11259, new_n1025);
nand_4 g10875(new_n11261, new_n11260, new_n1020);
nand_4 g10876(new_n11262, new_n11261, new_n1015);
nand_4 g10877(new_n11263, new_n11262, new_n1010);
nand_4 g10878(new_n11264, new_n11263, new_n1215);
nand_4 g10879(new_n11265, new_n11264, new_n1005);
nand_4 g10880(new_n11266, new_n11265, new_n1000);
nand_4 g10881(new_n11267, new_n11266, new_n994);
nand_4 g10882(new_n11268, new_n11267, new_n989);
nand_4 g10883(new_n11269_1, new_n11268, new_n984);
nand_4 g10884(new_n11270, new_n11269_1, new_n978);
nand_4 g10885(new_n11271, new_n11270, new_n973);
nand_4 g10886(new_n11272, new_n11271, new_n967);
nand_4 g10887(new_n11273, new_n11272, new_n964);
nand_4 g10888(new_n11274, new_n11273, new_n960);
nand_4 g10889(new_n11275, new_n11274, new_n957);
nand_4 g10890(new_n11276, new_n11275, new_n952);
nand_4 g10891(new_n11277, new_n11276, new_n948_1);
nand_4 g10892(new_n11278, new_n11277, new_n943);
nand_4 g10893(new_n11279, new_n11278, new_n938);
nand_4 g10894(new_n11280, new_n11279, new_n934);
nand_4 g10895(new_n11281, new_n11280, new_n929);
nand_4 g10896(new_n11282, new_n11281, new_n925);
nand_4 g10897(new_n11283, new_n11282, new_n2194);
nand_4 g10898(new_n11284, new_n11283, new_n2191);
nand_4 g10899(new_n11285, new_n11284, new_n2190);
not_3  g10900(new_n11286, new_n11285);
nor_4  g10901(new_n11287, new_n11286, new_n2514);
nor_4  g10902(new_n11288, new_n11287, new_n2513);
nor_4  g10903(new_n11289, new_n11288, new_n2512);
nor_4  g10904(new_n11290, new_n11289, new_n2511);
nor_4  g10905(new_n11291, new_n11290, new_n2510);
nor_4  g10906(new_n11292, new_n11291, new_n2509);
nor_4  g10907(new_n11293, new_n11292, new_n2508);
nor_4  g10908(new_n11294, new_n11293, new_n2507);
nor_4  g10909(new_n11295, new_n11294, new_n2506);
nor_4  g10910(new_n11296, new_n11295, new_n2505);
nor_4  g10911(new_n11297, new_n11296, new_n2504);
nor_4  g10912(new_n11298, new_n11297, new_n2503);
nor_4  g10913(new_n11299, new_n11298, new_n2502);
nor_4  g10914(new_n11300, new_n11299, new_n2790);
nor_4  g10915(new_n11301, new_n11300, new_n2789);
nor_4  g10916(new_n11302, new_n11301, new_n2788);
nor_4  g10917(new_n11303, new_n11302, new_n2305);
nor_4  g10918(new_n11304, new_n11303, new_n2304);
nor_4  g10919(new_n11305, new_n11304, new_n2303);
nor_4  g10920(new_n11306, new_n11305, new_n2302);
nor_4  g10921(new_n11307, new_n11306, new_n2301);
nor_4  g10922(new_n11308, new_n11307, new_n2300);
nor_4  g10923(new_n11309, new_n11308, new_n2299);
nor_4  g10924(new_n11310, new_n11309, new_n2298);
nor_4  g10925(new_n11311, new_n11310, new_n2297);
nor_4  g10926(new_n11312, new_n11311, new_n2296);
nor_4  g10927(new_n11313, new_n11312, new_n2295);
not_3  g10928(new_n11314, new_n11313);
nand_4 g10929(new_n11315, new_n11314, new_n1762);
nand_4 g10930(new_n11316, new_n11315, new_n1758);
nand_4 g10931(new_n11317, new_n11316, new_n1754);
nand_4 g10932(new_n11318, new_n11317, new_n1751);
nand_4 g10933(new_n11319, new_n11318, new_n1748);
nand_4 g10934(new_n11320, new_n11319, new_n1746);
nand_4 g10935(new_n11321, new_n11320, n2201);
nor_4  g10936(n12535, new_n11321, new_n1739_1);
not_3  g10937(new_n11323, new_n1663);
nand_4 g10938(new_n11324, new_n11323, new_n1010);
nand_4 g10939(new_n11325, new_n11324, new_n1215);
nand_4 g10940(new_n11326, new_n11325, new_n1005);
nand_4 g10941(new_n11327, new_n11326, new_n1000);
nand_4 g10942(new_n11328, new_n11327, new_n994);
nand_4 g10943(new_n11329, new_n11328, new_n989);
nand_4 g10944(new_n11330, new_n11329, new_n984);
nand_4 g10945(new_n11331, new_n11330, new_n978);
nand_4 g10946(new_n11332, new_n11331, new_n973);
nand_4 g10947(new_n11333, new_n11332, new_n967);
nand_4 g10948(new_n11334, new_n11333, new_n964);
nand_4 g10949(new_n11335, new_n11334, new_n960);
nand_4 g10950(new_n11336, new_n11335, new_n957);
nand_4 g10951(new_n11337, new_n11336, new_n952);
nand_4 g10952(new_n11338, new_n11337, new_n948_1);
nand_4 g10953(new_n11339, new_n11338, new_n943);
nand_4 g10954(new_n11340, new_n11339, new_n938);
nand_4 g10955(new_n11341, new_n11340, new_n934);
nand_4 g10956(new_n11342, new_n11341, new_n929);
nand_4 g10957(new_n11343, new_n11342, new_n925);
nand_4 g10958(new_n11344, new_n11343, new_n2194);
nand_4 g10959(new_n11345_1, new_n11344, new_n2191);
nand_4 g10960(new_n11346, new_n11345_1, new_n2190);
nand_4 g10961(new_n11347, new_n11346, new_n2186);
nand_4 g10962(new_n11348, new_n11347, new_n2183);
nand_4 g10963(new_n11349, new_n11348, new_n2179);
nand_4 g10964(new_n11350, new_n11349, new_n2175_1);
nand_4 g10965(new_n11351, new_n11350, new_n2171);
nand_4 g10966(new_n11352, new_n11351, new_n2168);
nand_4 g10967(new_n11353, new_n11352, new_n2165);
nand_4 g10968(new_n11354, new_n11353, new_n2162);
nand_4 g10969(new_n11355, new_n11354, new_n2158);
nand_4 g10970(new_n11356, new_n11355, new_n2155);
nand_4 g10971(new_n11357, new_n11356, new_n2151);
nand_4 g10972(new_n11358, new_n11357, new_n2147);
nand_4 g10973(new_n11359, new_n11358, new_n1810);
nand_4 g10974(new_n11360, new_n11359, new_n1806);
nand_4 g10975(new_n11361, new_n11360, new_n1802);
nand_4 g10976(new_n11362, new_n11361, new_n1798);
nand_4 g10977(new_n11363, new_n11362, new_n1820);
nand_4 g10978(new_n11364, new_n11363, new_n1794);
nand_4 g10979(new_n11365, new_n11364, new_n1825);
nand_4 g10980(new_n11366, new_n11365, new_n1789);
nand_4 g10981(new_n11367, new_n11366, new_n1785);
nand_4 g10982(new_n11368, new_n11367, new_n1780);
nand_4 g10983(new_n11369, new_n11368, new_n1777);
nand_4 g10984(new_n11370, new_n11369, new_n1774);
nand_4 g10985(new_n11371, new_n11370, new_n1834);
nand_4 g10986(new_n11372, new_n11371, new_n1769);
nand_4 g10987(new_n11373, new_n11372, new_n1766);
nand_4 g10988(new_n11374, new_n11373, new_n1762);
not_3  g10989(new_n11375, new_n11374);
nor_4  g10990(new_n11376, new_n11375, new_n2293);
nor_4  g10991(new_n11377, new_n11376, new_n2292);
nor_4  g10992(new_n11378, new_n11377, new_n2291);
nor_4  g10993(new_n11379, new_n11378, new_n2290);
nor_4  g10994(new_n11380, new_n11379, new_n2289);
nor_4  g10995(new_n11381, new_n11380, new_n2288);
nor_4  g10996(new_n11382, new_n11381, new_n2287);
nor_4  g10997(new_n11383, new_n11382, new_n2286);
nor_4  g10998(new_n11384, new_n11383, new_n2285);
nor_4  g10999(new_n11385, new_n11384, new_n2284);
nor_4  g11000(new_n11386, new_n11385, new_n2283);
nor_4  g11001(new_n11387, new_n11386, new_n2145);
nor_4  g11002(new_n11388, new_n11387, new_n2144);
nor_4  g11003(new_n11389, new_n11388, new_n2143);
nor_4  g11004(new_n11390, new_n11389, new_n2142);
nor_4  g11005(new_n11391, new_n11390, new_n2141);
nor_4  g11006(new_n11392, new_n11391, new_n2140);
nor_4  g11007(new_n11393_1, new_n11392, new_n2139);
nor_4  g11008(new_n11394, new_n11393_1, new_n2138);
nor_4  g11009(new_n11395, new_n11394, new_n2137);
nor_4  g11010(new_n11396, new_n11395, new_n2136);
nor_4  g11011(new_n11397, new_n11396, new_n2135);
nor_4  g11012(new_n11398, new_n11397, new_n2134);
nor_4  g11013(new_n11399, new_n11398, new_n2133);
nor_4  g11014(new_n11400, new_n11399, new_n2132);
nor_4  g11015(new_n11401, new_n11400, new_n1691);
nor_4  g11016(new_n11402, new_n11401, new_n1879);
not_3  g11017(new_n11403, new_n11402);
nand_4 g11018(new_n11404_1, new_n11403, new_n1882);
nand_4 g11019(new_n11405, new_n11404_1, new_n1686);
nand_4 g11020(new_n11406, new_n11405, new_n1682);
nand_4 g11021(new_n11407, new_n11406, new_n1678);
nand_4 g11022(new_n11408, new_n11407, new_n1674);
nand_4 g11023(new_n11409, new_n11408, new_n1890);
nand_4 g11024(new_n11410, new_n11409, n3893);
nor_4  g11025(n12989, new_n11410, new_n684);
nand_4 g11026(new_n11412, new_n977_1, new_n498_1);
nand_4 g11027(new_n11413, new_n11412, new_n727);
nand_4 g11028(new_n11414, new_n11413, new_n494);
nand_4 g11029(new_n11415, new_n11414, new_n735);
nand_4 g11030(new_n11416, new_n11415, new_n488);
nand_4 g11031(new_n11417, new_n11416, new_n743);
nand_4 g11032(new_n11418, new_n11417, new_n482);
nand_4 g11033(new_n11419, new_n11418, new_n751);
nand_4 g11034(new_n11420, new_n11419, new_n758);
nand_4 g11035(new_n11421, new_n11420, new_n765);
nand_4 g11036(new_n11422, new_n11421, new_n476);
nand_4 g11037(new_n11423, new_n11422, new_n773);
nand_4 g11038(new_n11424, new_n11423, new_n780);
nand_4 g11039(new_n11425, new_n11424, new_n787);
nand_4 g11040(new_n11426, new_n11425, new_n470);
nand_4 g11041(new_n11427, new_n11426, new_n795);
nand_4 g11042(new_n11428, new_n11427, new_n803);
nand_4 g11043(new_n11429, new_n11428, new_n809);
nand_4 g11044(new_n11430, new_n11429, new_n465);
nand_4 g11045(new_n11431, new_n11430, new_n818);
nand_4 g11046(new_n11432, new_n11431, new_n460);
nand_4 g11047(new_n11433, new_n11432, new_n455);
nand_4 g11048(new_n11434, new_n11433, new_n449);
nand_4 g11049(new_n11435, new_n11434, new_n827);
nand_4 g11050(new_n11436, new_n11435, new_n833);
nand_4 g11051(new_n11437, new_n11436, new_n444);
nand_4 g11052(new_n11438, new_n11437, new_n439);
nand_4 g11053(new_n11439, new_n11438, new_n841);
nand_4 g11054(new_n11440, new_n11439, new_n434);
nand_4 g11055(new_n11441, new_n11440, new_n429);
nand_4 g11056(new_n11442, new_n11441, new_n424);
nand_4 g11057(new_n11443, new_n11442, new_n850);
nand_4 g11058(new_n11444, new_n11443, new_n856);
nand_4 g11059(new_n11445, new_n11444, new_n863);
nand_4 g11060(new_n11446, new_n11445, new_n419);
nand_4 g11061(new_n11447, new_n11446, new_n869);
nand_4 g11062(new_n11448, new_n11447, new_n875);
nand_4 g11063(new_n11449, new_n11448, new_n881);
nand_4 g11064(new_n11450, new_n11449, new_n413);
nand_4 g11065(new_n11451, new_n11450, new_n889);
nand_4 g11066(new_n11452, new_n11451, new_n896);
nand_4 g11067(new_n11453, new_n11452, new_n901);
nand_4 g11068(new_n11454, new_n11453, new_n408);
nand_4 g11069(new_n11455, new_n11454, new_n908);
nand_4 g11070(new_n11456, new_n11455, new_n403);
nand_4 g11071(new_n11457, new_n11456, new_n398);
nand_4 g11072(new_n11458, new_n11457, new_n393);
nand_4 g11073(new_n11459, new_n11458, new_n916);
nand_4 g11074(new_n11460, new_n11459, new_n1123);
nand_4 g11075(new_n11461, new_n11460, new_n1164);
not_3  g11076(new_n11462, new_n11461);
nor_4  g11077(new_n11463_1, new_n11462, new_n1530);
nor_4  g11078(new_n11464, new_n11463_1, new_n1529);
nor_4  g11079(new_n11465, new_n11464, new_n1528);
nor_4  g11080(new_n11466, new_n11465, new_n1527);
nor_4  g11081(new_n11467, new_n11466, new_n1526);
nor_4  g11082(new_n11468, new_n11467, new_n1525);
nor_4  g11083(new_n11469, new_n11468, new_n1524);
nor_4  g11084(new_n11470, new_n11469, new_n1523);
nor_4  g11085(new_n11471, new_n11470, new_n1522);
nor_4  g11086(new_n11472, new_n11471, new_n1521);
nor_4  g11087(new_n11473, new_n11472, new_n1520);
nor_4  g11088(new_n11474, new_n11473, new_n1519);
nor_4  g11089(new_n11475, new_n11474, new_n1518);
nor_4  g11090(new_n11476, new_n11475, new_n1517);
nor_4  g11091(new_n11477, new_n11476, new_n1516);
nor_4  g11092(new_n11478, new_n11477, new_n1075);
nor_4  g11093(new_n11479, new_n11478, new_n1071);
nor_4  g11094(new_n11480, new_n11479, new_n1065);
nor_4  g11095(new_n11481, new_n11480, new_n1062);
nor_4  g11096(new_n11482, new_n11481, new_n1056);
nor_4  g11097(new_n11483, new_n11482, new_n1051);
nor_4  g11098(new_n11484, new_n11483, new_n1046);
nor_4  g11099(new_n11485, new_n11484, new_n1042);
nor_4  g11100(new_n11486, new_n11485, new_n1037);
nor_4  g11101(new_n11487, new_n11486, new_n1032);
not_3  g11102(new_n11488, new_n11487);
nand_4 g11103(new_n11489, new_n11488, new_n1025);
nand_4 g11104(new_n11490, new_n11489, new_n1020);
nand_4 g11105(new_n11491, new_n11490, new_n1015);
nand_4 g11106(new_n11492, new_n11491, new_n1010);
nand_4 g11107(new_n11493, new_n11492, new_n1215);
nand_4 g11108(new_n11494, new_n11493, new_n1005);
nand_4 g11109(new_n11495, new_n11494, new_n1000);
nand_4 g11110(new_n11496, new_n11495, new_n994);
nand_4 g11111(new_n11497, new_n11496, new_n989);
nand_4 g11112(new_n11498, new_n11497, n10061);
nor_4  g11113(n13010, new_n11498, new_n981);
nand_4 g11114(new_n11500, new_n931, new_n929);
nand_4 g11115(new_n11501, new_n11500, new_n925);
nand_4 g11116(new_n11502, new_n11501, new_n2194);
nand_4 g11117(new_n11503, new_n11502, new_n2191);
nand_4 g11118(new_n11504, new_n11503, new_n2190);
nand_4 g11119(new_n11505, new_n11504, new_n2186);
nand_4 g11120(new_n11506, new_n11505, new_n2183);
nand_4 g11121(new_n11507, new_n11506, new_n2179);
nand_4 g11122(new_n11508, new_n11507, new_n2175_1);
nand_4 g11123(new_n11509, new_n11508, new_n2171);
nand_4 g11124(new_n11510, new_n11509, new_n2168);
nand_4 g11125(new_n11511, new_n11510, new_n2165);
nand_4 g11126(new_n11512, new_n11511, new_n2162);
nand_4 g11127(new_n11513, new_n11512, new_n2158);
nand_4 g11128(new_n11514, new_n11513, new_n2155);
nand_4 g11129(new_n11515, new_n11514, new_n2151);
nand_4 g11130(new_n11516, new_n11515, new_n2147);
nand_4 g11131(new_n11517, new_n11516, new_n1810);
nand_4 g11132(new_n11518, new_n11517, new_n1806);
nand_4 g11133(new_n11519, new_n11518, new_n1802);
nand_4 g11134(new_n11520, new_n11519, new_n1798);
nand_4 g11135(new_n11521, new_n11520, new_n1820);
nand_4 g11136(new_n11522, new_n11521, new_n1794);
nand_4 g11137(new_n11523, new_n11522, new_n1825);
nand_4 g11138(new_n11524, new_n11523, new_n1789);
nand_4 g11139(new_n11525, new_n11524, new_n1785);
nand_4 g11140(new_n11526, new_n11525, new_n1780);
nand_4 g11141(new_n11527, new_n11526, new_n1777);
nand_4 g11142(new_n11528, new_n11527, new_n1774);
nand_4 g11143(new_n11529_1, new_n11528, new_n1834);
nand_4 g11144(new_n11530, new_n11529_1, new_n1769);
nand_4 g11145(new_n11531, new_n11530, new_n1766);
nand_4 g11146(new_n11532, new_n11531, new_n1762);
nand_4 g11147(new_n11533, new_n11532, new_n1758);
nand_4 g11148(new_n11534_1, new_n11533, new_n1754);
not_3  g11149(new_n11535, new_n11534_1);
nor_4  g11150(new_n11536, new_n11535, new_n2291);
nor_4  g11151(new_n11537, new_n11536, new_n2290);
nor_4  g11152(new_n11538, new_n11537, new_n2289);
nor_4  g11153(new_n11539, new_n11538, new_n2288);
nor_4  g11154(new_n11540, new_n11539, new_n2287);
nor_4  g11155(new_n11541, new_n11540, new_n2286);
nor_4  g11156(new_n11542, new_n11541, new_n2285);
nor_4  g11157(new_n11543, new_n11542, new_n2284);
nor_4  g11158(new_n11544, new_n11543, new_n2283);
nor_4  g11159(new_n11545, new_n11544, new_n2145);
nor_4  g11160(new_n11546, new_n11545, new_n2144);
nor_4  g11161(new_n11547, new_n11546, new_n2143);
nor_4  g11162(new_n11548, new_n11547, new_n2142);
nor_4  g11163(new_n11549, new_n11548, new_n2141);
nor_4  g11164(new_n11550, new_n11549, new_n2140);
nor_4  g11165(new_n11551, new_n11550, new_n2139);
nor_4  g11166(new_n11552, new_n11551, new_n2138);
nor_4  g11167(new_n11553, new_n11552, new_n2137);
nor_4  g11168(new_n11554, new_n11553, new_n2136);
not_3  g11169(new_n11555, new_n11554);
nand_4 g11170(new_n11556, new_n11555, new_n1699);
nand_4 g11171(new_n11557, new_n11556, new_n1697);
nand_4 g11172(new_n11558, new_n11557, new_n1871);
nand_4 g11173(new_n11559, new_n11558, new_n1694);
nand_4 g11174(new_n11560, new_n11559, new_n1690);
nand_4 g11175(new_n11561, new_n11560, new_n1878);
nand_4 g11176(new_n11562, new_n11561, new_n1882);
nand_4 g11177(new_n11563, new_n11562, new_n1686);
nand_4 g11178(new_n11564, new_n11563, new_n1682);
nand_4 g11179(new_n11565, new_n11564, new_n1678);
nand_4 g11180(new_n11566, new_n11565, new_n1674);
nand_4 g11181(new_n11567, new_n11566, new_n1890);
nand_4 g11182(new_n11568, new_n11567, new_n1669);
nand_4 g11183(new_n11569, new_n11568, new_n1665);
nand_4 g11184(new_n11570, new_n11569, new_n1661);
nand_4 g11185(new_n11571, new_n11570, new_n1657);
nand_4 g11186(new_n11572, new_n11571, new_n1652);
nand_4 g11187(new_n11573, new_n11572, new_n1648);
nand_4 g11188(new_n11574, new_n11573, new_n1644);
nand_4 g11189(new_n11575, new_n11574, new_n1640);
nand_4 g11190(new_n11576, new_n11575, new_n1636);
nand_4 g11191(new_n11577, new_n11576, new_n1632);
nand_4 g11192(new_n11578, new_n11577, new_n1378);
nand_4 g11193(new_n11579, new_n11578, new_n1372);
nand_4 g11194(new_n11580, new_n11579, new_n1367);
nand_4 g11195(new_n11581, new_n11580, new_n1363);
nand_4 g11196(new_n11582, new_n11581, new_n1360);
nand_4 g11197(new_n11583, new_n11582, new_n1357);
nand_4 g11198(new_n11584, new_n11583, new_n1354);
nand_4 g11199(new_n11585, new_n11584, new_n1352);
nand_4 g11200(new_n11586, new_n11585, n12321);
nor_4  g11201(n13045, new_n11586, new_n762);
nand_4 g11202(new_n11588, new_n951, new_n480);
nand_4 g11203(new_n11589, new_n11588, new_n751);
nand_4 g11204(new_n11590_1, new_n11589, new_n758);
nand_4 g11205(new_n11591, new_n11590_1, new_n765);
nand_4 g11206(new_n11592, new_n11591, new_n476);
nand_4 g11207(new_n11593, new_n11592, new_n773);
nand_4 g11208(new_n11594, new_n11593, new_n780);
nand_4 g11209(new_n11595, new_n11594, new_n787);
nand_4 g11210(new_n11596, new_n11595, new_n470);
nand_4 g11211(new_n11597, new_n11596, new_n795);
nand_4 g11212(new_n11598, new_n11597, new_n803);
nand_4 g11213(new_n11599, new_n11598, new_n809);
nand_4 g11214(new_n11600, new_n11599, new_n465);
nand_4 g11215(new_n11601, new_n11600, new_n818);
nand_4 g11216(new_n11602, new_n11601, new_n460);
nand_4 g11217(new_n11603, new_n11602, new_n455);
nand_4 g11218(new_n11604, new_n11603, new_n449);
nand_4 g11219(new_n11605_1, new_n11604, new_n827);
nand_4 g11220(new_n11606, new_n11605_1, new_n833);
nand_4 g11221(new_n11607, new_n11606, new_n444);
nand_4 g11222(new_n11608, new_n11607, new_n439);
nand_4 g11223(new_n11609, new_n11608, new_n841);
nand_4 g11224(new_n11610, new_n11609, new_n434);
nand_4 g11225(new_n11611, new_n11610, new_n429);
nand_4 g11226(new_n11612, new_n11611, new_n424);
nand_4 g11227(new_n11613, new_n11612, new_n850);
nand_4 g11228(new_n11614, new_n11613, new_n856);
nand_4 g11229(new_n11615, new_n11614, new_n863);
nand_4 g11230(new_n11616, new_n11615, new_n419);
nand_4 g11231(new_n11617, new_n11616, new_n869);
nand_4 g11232(new_n11618, new_n11617, new_n875);
nand_4 g11233(new_n11619, new_n11618, new_n881);
nand_4 g11234(new_n11620, new_n11619, new_n413);
nand_4 g11235(new_n11621, new_n11620, new_n889);
nand_4 g11236(new_n11622, new_n11621, new_n896);
nand_4 g11237(new_n11623, new_n11622, new_n901);
nand_4 g11238(new_n11624, new_n11623, new_n408);
nand_4 g11239(new_n11625, new_n11624, new_n908);
nand_4 g11240(new_n11626, new_n11625, new_n403);
nand_4 g11241(new_n11627_1, new_n11626, new_n398);
nand_4 g11242(new_n11628, new_n11627_1, new_n393);
nand_4 g11243(new_n11629, new_n11628, new_n916);
nand_4 g11244(new_n11630, new_n11629, new_n1123);
nand_4 g11245(new_n11631, new_n11630, new_n1164);
nand_4 g11246(new_n11632, new_n11631, new_n1120);
not_3  g11247(new_n11633, new_n11632);
nor_4  g11248(new_n11634, new_n11633, new_n1529);
nor_4  g11249(new_n11635, new_n11634, new_n1528);
nor_4  g11250(new_n11636, new_n11635, new_n1527);
nor_4  g11251(new_n11637, new_n11636, new_n1526);
nor_4  g11252(new_n11638, new_n11637, new_n1525);
nor_4  g11253(new_n11639, new_n11638, new_n1524);
nor_4  g11254(new_n11640, new_n11639, new_n1523);
nor_4  g11255(new_n11641, new_n11640, new_n1522);
nor_4  g11256(new_n11642, new_n11641, new_n1521);
nor_4  g11257(new_n11643, new_n11642, new_n1520);
nor_4  g11258(new_n11644, new_n11643, new_n1519);
nor_4  g11259(new_n11645, new_n11644, new_n1518);
nor_4  g11260(new_n11646, new_n11645, new_n1517);
nor_4  g11261(new_n11647, new_n11646, new_n1516);
nor_4  g11262(new_n11648, new_n11647, new_n1075);
nor_4  g11263(new_n11649, new_n11648, new_n1071);
nor_4  g11264(new_n11650, new_n11649, new_n1065);
nor_4  g11265(new_n11651, new_n11650, new_n1062);
nor_4  g11266(new_n11652, new_n11651, new_n1056);
nor_4  g11267(new_n11653, new_n11652, new_n1051);
nor_4  g11268(new_n11654, new_n11653, new_n1046);
nor_4  g11269(new_n11655, new_n11654, new_n1042);
nor_4  g11270(new_n11656, new_n11655, new_n1037);
nor_4  g11271(new_n11657, new_n11656, new_n1032);
not_3  g11272(new_n11658, new_n11657);
nand_4 g11273(new_n11659, new_n11658, new_n1025);
nand_4 g11274(new_n11660, new_n11659, new_n1020);
nand_4 g11275(new_n11661, new_n11660, new_n1015);
nand_4 g11276(new_n11662, new_n11661, new_n1010);
nand_4 g11277(new_n11663, new_n11662, new_n1215);
nand_4 g11278(new_n11664_1, new_n11663, new_n1005);
nand_4 g11279(new_n11665, new_n11664_1, new_n1000);
nand_4 g11280(new_n11666_1, new_n11665, new_n994);
nand_4 g11281(new_n11667, new_n11666_1, new_n989);
nand_4 g11282(new_n11668, new_n11667, new_n984);
nand_4 g11283(new_n11669, new_n11668, new_n978);
nand_4 g11284(new_n11670, new_n11669, new_n973);
nand_4 g11285(new_n11671, new_n11670, new_n967);
nand_4 g11286(new_n11672, new_n11671, new_n964);
nand_4 g11287(new_n11673, new_n11672, new_n960);
nand_4 g11288(new_n11674, new_n11673, n10470);
nor_4  g11289(n13114, new_n11674, new_n955);
nand_4 g11290(new_n11676, new_n2192, new_n1340);
nand_4 g11291(new_n11677, new_n11676, new_n2191);
nand_4 g11292(new_n11678, new_n11677, new_n2190);
nand_4 g11293(new_n11679, new_n11678, new_n2186);
nand_4 g11294(new_n11680, new_n11679, new_n2183);
nand_4 g11295(new_n11681, new_n11680, new_n2179);
nand_4 g11296(new_n11682, new_n11681, new_n2175_1);
nand_4 g11297(new_n11683, new_n11682, new_n2171);
nand_4 g11298(new_n11684, new_n11683, new_n2168);
nand_4 g11299(new_n11685, new_n11684, new_n2165);
nand_4 g11300(new_n11686, new_n11685, new_n2162);
nand_4 g11301(new_n11687, new_n11686, new_n2158);
nand_4 g11302(new_n11688, new_n11687, new_n2155);
nand_4 g11303(new_n11689, new_n11688, new_n2151);
nand_4 g11304(new_n11690, new_n11689, new_n2147);
nand_4 g11305(new_n11691, new_n11690, new_n1810);
nand_4 g11306(new_n11692, new_n11691, new_n1806);
nand_4 g11307(new_n11693, new_n11692, new_n1802);
nand_4 g11308(new_n11694, new_n11693, new_n1798);
nand_4 g11309(new_n11695, new_n11694, new_n1820);
nand_4 g11310(new_n11696, new_n11695, new_n1794);
nand_4 g11311(new_n11697, new_n11696, new_n1825);
nand_4 g11312(new_n11698, new_n11697, new_n1789);
nand_4 g11313(new_n11699, new_n11698, new_n1785);
nand_4 g11314(new_n11700, new_n11699, new_n1780);
nand_4 g11315(new_n11701, new_n11700, new_n1777);
nand_4 g11316(new_n11702, new_n11701, new_n1774);
nand_4 g11317(new_n11703, new_n11702, new_n1834);
nand_4 g11318(new_n11704, new_n11703, new_n1769);
nand_4 g11319(new_n11705, new_n11704, new_n1766);
nand_4 g11320(new_n11706, new_n11705, new_n1762);
nand_4 g11321(new_n11707, new_n11706, new_n1758);
nand_4 g11322(new_n11708, new_n11707, new_n1754);
nand_4 g11323(new_n11709, new_n11708, new_n1751);
nand_4 g11324(new_n11710, new_n11709, new_n1748);
nand_4 g11325(new_n11711, new_n11710, new_n1746);
nand_4 g11326(new_n11712, new_n11711, new_n1742);
nand_4 g11327(new_n11713, new_n11712, new_n1738);
nand_4 g11328(new_n11714, new_n11713, new_n1736);
nand_4 g11329(new_n11715, new_n11714, new_n1732);
nand_4 g11330(new_n11716, new_n11715, new_n1729);
nand_4 g11331(new_n11717, new_n11716, new_n1726);
nand_4 g11332(new_n11718, new_n11717, new_n1724);
nand_4 g11333(new_n11719, new_n11718, new_n1721);
nand_4 g11334(new_n11720, new_n11719, new_n1718);
nand_4 g11335(new_n11721, new_n11720, new_n1715);
nand_4 g11336(new_n11722, new_n11721, new_n1711);
nand_4 g11337(new_n11723, new_n11722, new_n1708);
nand_4 g11338(new_n11724, new_n11723, new_n1705);
nand_4 g11339(new_n11725, new_n11724, new_n1703);
nand_4 g11340(new_n11726, new_n11725, new_n1860);
not_3  g11341(new_n11727, new_n11726);
nor_4  g11342(new_n11728, new_n11727, new_n2136);
nor_4  g11343(new_n11729, new_n11728, new_n2135);
nor_4  g11344(new_n11730, new_n11729, new_n2134);
nor_4  g11345(new_n11731, new_n11730, new_n2133);
nor_4  g11346(new_n11732, new_n11731, new_n2132);
nor_4  g11347(new_n11733, new_n11732, new_n1691);
nor_4  g11348(new_n11734, new_n11733, new_n1879);
nor_4  g11349(new_n11735, new_n11734, new_n1883);
nor_4  g11350(new_n11736, new_n11735, new_n1687);
nor_4  g11351(new_n11737, new_n11736, new_n1683);
nor_4  g11352(new_n11738, new_n11737, new_n1679);
nor_4  g11353(new_n11739, new_n11738, new_n1675);
nor_4  g11354(new_n11740, new_n11739, new_n1891);
nor_4  g11355(new_n11741, new_n11740, new_n1670);
nor_4  g11356(new_n11742, new_n11741, new_n1666);
nor_4  g11357(new_n11743, new_n11742, new_n1662);
nor_4  g11358(new_n11744, new_n11743, new_n1658);
nor_4  g11359(new_n11745, new_n11744, new_n1653);
nor_4  g11360(new_n11746, new_n11745, new_n1649);
nor_4  g11361(new_n11747, new_n11746, new_n1645);
nor_4  g11362(new_n11748, new_n11747, new_n1641);
nor_4  g11363(new_n11749, new_n11748, new_n1637_1);
nor_4  g11364(new_n11750, new_n11749, new_n1633);
nor_4  g11365(new_n11751, new_n11750, new_n1629);
nor_4  g11366(new_n11752, new_n11751, new_n1628);
nor_4  g11367(new_n11753, new_n11752, new_n1627);
nor_4  g11368(new_n11754, new_n11753, new_n1626);
not_3  g11369(new_n11755, new_n11754);
nand_4 g11370(new_n11756_1, new_n11755, new_n1360);
nand_4 g11371(new_n11757, new_n11756_1, new_n1357);
nand_4 g11372(new_n11758, new_n11757, new_n1354);
nand_4 g11373(new_n11759, new_n11758, new_n1352);
nand_4 g11374(new_n11760, new_n11759, new_n1350);
nand_4 g11375(new_n11761, new_n11760, new_n1347_1);
nand_4 g11376(new_n11762, new_n11761, n4147);
nor_4  g11377(n13141, new_n11762, new_n770);
nand_4 g11378(new_n11764, new_n1767, new_n1264);
nand_4 g11379(new_n11765, new_n11764, new_n1766);
nand_4 g11380(new_n11766, new_n11765, new_n1762);
nand_4 g11381(new_n11767, new_n11766, new_n1758);
nand_4 g11382(new_n11768, new_n11767, new_n1754);
nand_4 g11383(new_n11769, new_n11768, new_n1751);
nand_4 g11384(new_n11770, new_n11769, new_n1748);
nand_4 g11385(new_n11771, new_n11770, new_n1746);
nand_4 g11386(new_n11772, new_n11771, new_n1742);
nand_4 g11387(new_n11773, new_n11772, new_n1738);
nand_4 g11388(new_n11774, new_n11773, new_n1736);
nand_4 g11389(new_n11775, new_n11774, new_n1732);
nand_4 g11390(new_n11776_1, new_n11775, new_n1729);
nand_4 g11391(new_n11777, new_n11776_1, new_n1726);
nand_4 g11392(new_n11778, new_n11777, new_n1724);
nand_4 g11393(new_n11779, new_n11778, new_n1721);
nand_4 g11394(new_n11780, new_n11779, new_n1718);
nand_4 g11395(new_n11781, new_n11780, new_n1715);
nand_4 g11396(new_n11782, new_n11781, new_n1711);
nand_4 g11397(new_n11783, new_n11782, new_n1708);
nand_4 g11398(new_n11784, new_n11783, new_n1705);
nand_4 g11399(new_n11785, new_n11784, new_n1703);
nand_4 g11400(new_n11786, new_n11785, new_n1860);
nand_4 g11401(new_n11787, new_n11786, new_n1864);
nand_4 g11402(new_n11788, new_n11787, new_n1699);
nand_4 g11403(new_n11789, new_n11788, new_n1697);
nand_4 g11404(new_n11790, new_n11789, new_n1871);
nand_4 g11405(new_n11791, new_n11790, new_n1694);
nand_4 g11406(new_n11792, new_n11791, new_n1690);
nand_4 g11407(new_n11793, new_n11792, new_n1878);
nand_4 g11408(new_n11794, new_n11793, new_n1882);
nand_4 g11409(new_n11795, new_n11794, new_n1686);
nand_4 g11410(new_n11796, new_n11795, new_n1682);
nand_4 g11411(new_n11797, new_n11796, new_n1678);
nand_4 g11412(new_n11798, new_n11797, new_n1674);
nand_4 g11413(new_n11799, new_n11798, new_n1890);
nand_4 g11414(new_n11800, new_n11799, new_n1669);
nand_4 g11415(new_n11801, new_n11800, new_n1665);
nand_4 g11416(new_n11802, new_n11801, new_n1661);
nand_4 g11417(new_n11803, new_n11802, new_n1657);
nand_4 g11418(new_n11804, new_n11803, new_n1652);
nand_4 g11419(new_n11805, new_n11804, new_n1648);
nand_4 g11420(new_n11806, new_n11805, new_n1644);
nand_4 g11421(new_n11807, new_n11806, new_n1640);
nand_4 g11422(new_n11808, new_n11807, new_n1636);
nand_4 g11423(new_n11809, new_n11808, new_n1632);
not_3  g11424(new_n11810, new_n11809);
nor_4  g11425(new_n11811, new_n11810, new_n1629);
nor_4  g11426(new_n11812, new_n11811, new_n1628);
nor_4  g11427(new_n11813, new_n11812, new_n1627);
nor_4  g11428(new_n11814, new_n11813, new_n1626);
nor_4  g11429(new_n11815, new_n11814, new_n4700);
nor_4  g11430(new_n11816, new_n11815, new_n4699);
nor_4  g11431(new_n11817, new_n11816, new_n3722);
nor_4  g11432(new_n11818, new_n11817, new_n3721);
nor_4  g11433(new_n11819, new_n11818, new_n3720);
nor_4  g11434(new_n11820, new_n11819, new_n3719);
nor_4  g11435(new_n11821, new_n11820, new_n3718);
nor_4  g11436(new_n11822_1, new_n11821, new_n3717);
nor_4  g11437(new_n11823, new_n11822_1, new_n3716);
nor_4  g11438(new_n11824, new_n11823, new_n2611);
nor_4  g11439(new_n11825, new_n11824, new_n2610);
nor_4  g11440(new_n11826, new_n11825, new_n2609);
nor_4  g11441(new_n11827, new_n11826, new_n2413);
nor_4  g11442(new_n11828, new_n11827, new_n2412);
nor_4  g11443(new_n11829, new_n11828, new_n2411);
nor_4  g11444(new_n11830, new_n11829, new_n2410);
nor_4  g11445(new_n11831, new_n11830, new_n2409);
nor_4  g11446(new_n11832, new_n11831, new_n2408);
nor_4  g11447(new_n11833, new_n11832, new_n2407_1);
nor_4  g11448(new_n11834, new_n11833, new_n2406);
not_3  g11449(new_n11835, new_n11834);
nand_4 g11450(new_n11836, new_n11835, new_n1419);
nand_4 g11451(new_n11837, new_n11836, new_n1310);
nand_4 g11452(new_n11838, new_n11837, new_n1305);
nand_4 g11453(new_n11839, new_n11838, new_n1427);
nand_4 g11454(new_n11840, new_n11839, new_n1431);
nand_4 g11455(new_n11841, new_n11840, new_n1302);
nand_4 g11456(new_n11842_1, new_n11841, new_n1298);
nand_4 g11457(new_n11843, new_n11842_1, new_n1295);
nand_4 g11458(new_n11844, new_n11843, new_n1291);
nand_4 g11459(new_n11845, new_n11844, new_n1288);
nand_4 g11460(new_n11846, new_n11845, new_n1284);
nand_4 g11461(new_n11847_1, new_n11846, new_n1280);
nand_4 g11462(new_n11848, new_n11847_1, new_n1275);
nand_4 g11463(new_n11849, new_n11848, new_n1445);
nand_4 g11464(new_n11850, new_n11849, n5467);
nor_4  g11465(n13316, new_n11850, new_n1268_1);
not_3  g11466(new_n11852, new_n1190);
nand_4 g11467(new_n11853, new_n11852, new_n1187);
nand_4 g11468(new_n11854_1, new_n11853, new_n562);
nand_4 g11469(new_n11855, new_n11854_1, new_n632);
nand_4 g11470(new_n11856, new_n11855, new_n638);
nand_4 g11471(new_n11857, new_n11856, new_n559);
nand_4 g11472(new_n11858, new_n11857, new_n554);
nand_4 g11473(new_n11859, new_n11858, new_n646);
nand_4 g11474(new_n11860, new_n11859, new_n652);
nand_4 g11475(new_n11861, new_n11860, new_n549);
nand_4 g11476(new_n11862, new_n11861, new_n544);
nand_4 g11477(new_n11863, new_n11862, new_n660);
nand_4 g11478(new_n11864, new_n11863, new_n539);
nand_4 g11479(new_n11865, new_n11864, new_n534);
nand_4 g11480(new_n11866, new_n11865, new_n529);
nand_4 g11481(new_n11867, new_n11866, new_n668);
nand_4 g11482(new_n11868, new_n11867, new_n674_1);
nand_4 g11483(new_n11869, new_n11868, new_n681);
nand_4 g11484(new_n11870, new_n11869, new_n523);
nand_4 g11485(new_n11871, new_n11870, new_n687);
nand_4 g11486(new_n11872, new_n11871, new_n693);
nand_4 g11487(new_n11873, new_n11872, new_n699);
nand_4 g11488(new_n11874, new_n11873, new_n517);
nand_4 g11489(new_n11875_1, new_n11874, new_n705);
nand_4 g11490(new_n11876, new_n11875_1, new_n511);
nand_4 g11491(new_n11877, new_n11876, new_n711);
nand_4 g11492(new_n11878, new_n11877, new_n506);
nand_4 g11493(new_n11879, new_n11878, new_n719);
nand_4 g11494(new_n11880, new_n11879, new_n500);
nand_4 g11495(new_n11881, new_n11880, new_n727);
nand_4 g11496(new_n11882, new_n11881, new_n494);
nand_4 g11497(new_n11883, new_n11882, new_n735);
nand_4 g11498(new_n11884, new_n11883, new_n488);
nand_4 g11499(new_n11885, new_n11884, new_n743);
nand_4 g11500(new_n11886, new_n11885, new_n482);
nand_4 g11501(new_n11887, new_n11886, new_n751);
nand_4 g11502(new_n11888, new_n11887, new_n758);
nand_4 g11503(new_n11889, new_n11888, new_n765);
nand_4 g11504(new_n11890, new_n11889, new_n476);
nand_4 g11505(new_n11891, new_n11890, new_n773);
nand_4 g11506(new_n11892, new_n11891, new_n780);
nand_4 g11507(new_n11893, new_n11892, new_n787);
nand_4 g11508(new_n11894, new_n11893, new_n470);
nand_4 g11509(new_n11895, new_n11894, new_n795);
nand_4 g11510(new_n11896, new_n11895, new_n803);
nand_4 g11511(new_n11897, new_n11896, new_n809);
nand_4 g11512(new_n11898, new_n11897, new_n465);
not_3  g11513(new_n11899, new_n11898);
nor_4  g11514(new_n11900, new_n11899, new_n2042);
nor_4  g11515(new_n11901, new_n11900, new_n2041);
nor_4  g11516(new_n11902_1, new_n11901, new_n2040);
nor_4  g11517(new_n11903, new_n11902_1, new_n2039);
nor_4  g11518(new_n11904, new_n11903, new_n2038);
nor_4  g11519(new_n11905, new_n11904, new_n2037);
nor_4  g11520(new_n11906, new_n11905, new_n2036);
nor_4  g11521(new_n11907, new_n11906, new_n2035);
nor_4  g11522(new_n11908, new_n11907, new_n2034);
nor_4  g11523(new_n11909, new_n11908, new_n2033);
nor_4  g11524(new_n11910, new_n11909, new_n2032);
nor_4  g11525(new_n11911, new_n11910, new_n2031);
nor_4  g11526(new_n11912, new_n11911, new_n2030);
nor_4  g11527(new_n11913, new_n11912, new_n2029);
nor_4  g11528(new_n11914, new_n11913, new_n2028);
nor_4  g11529(new_n11915, new_n11914, new_n2027_1);
nor_4  g11530(new_n11916, new_n11915, new_n2026);
nor_4  g11531(new_n11917, new_n11916, new_n2025);
nor_4  g11532(new_n11918, new_n11917, new_n2024);
nor_4  g11533(new_n11919, new_n11918, new_n2023);
nor_4  g11534(new_n11920, new_n11919, new_n2022);
nor_4  g11535(new_n11921, new_n11920, new_n2021);
nor_4  g11536(new_n11922, new_n11921, new_n2020);
nor_4  g11537(new_n11923, new_n11922, new_n2019);
not_3  g11538(new_n11924, new_n11923);
nand_4 g11539(new_n11925, new_n11924, new_n908);
nand_4 g11540(new_n11926, new_n11925, new_n403);
nand_4 g11541(new_n11927, new_n11926, new_n398);
nand_4 g11542(new_n11928, new_n11927, new_n393);
nand_4 g11543(new_n11929, new_n11928, new_n916);
nand_4 g11544(new_n11930_1, new_n11929, new_n1123);
nand_4 g11545(new_n11931, new_n11930_1, new_n1164);
nand_4 g11546(new_n11932, new_n11931, new_n1120);
nand_4 g11547(new_n11933_1, new_n11932, new_n1169);
nand_4 g11548(new_n11934, new_n11933_1, new_n1116);
nand_4 g11549(new_n11935, new_n11934, new_n1111);
nand_4 g11550(new_n11936, new_n11935, new_n1106);
nand_4 g11551(new_n11937, new_n11936, new_n1178);
nand_4 g11552(new_n11938, new_n11937, new_n1183);
nand_4 g11553(new_n11939, new_n11938, new_n1102);
nand_4 g11554(new_n11940, new_n11939, n9110);
nor_4  g11555(n13577, new_n11940, new_n1096);
nand_4 g11556(new_n11942, new_n1249, new_n907);
nand_4 g11557(new_n11943, new_n11942, new_n1457);
nand_4 g11558(new_n11944, new_n11943, new_n1462);
nand_4 g11559(new_n11945, new_n11944, new_n1468);
nand_4 g11560(new_n11946, new_n11945, new_n1247);
nand_4 g11561(new_n11947, new_n11946, new_n1474);
nand_4 g11562(new_n11948, new_n11947, new_n592);
nand_4 g11563(new_n11949, new_n11948, new_n585);
nand_4 g11564(new_n11950, new_n11949, new_n580);
nand_4 g11565(new_n11951, new_n11950, new_n600);
nand_4 g11566(new_n11952, new_n11951, new_n606);
nand_4 g11567(new_n11953, new_n11952, new_n612);
nand_4 g11568(new_n11954, new_n11953, new_n575);
nand_4 g11569(new_n11955, new_n11954, new_n619);
nand_4 g11570(new_n11956, new_n11955, new_n570);
nand_4 g11571(new_n11957, new_n11956, new_n625);
nand_4 g11572(new_n11958, new_n11957, new_n564);
nand_4 g11573(new_n11959, new_n11958, new_n632);
nand_4 g11574(new_n11960, new_n11959, new_n638);
nand_4 g11575(new_n11961_1, new_n11960, new_n559);
nand_4 g11576(new_n11962, new_n11961_1, new_n554);
nand_4 g11577(new_n11963, new_n11962, new_n646);
nand_4 g11578(new_n11964, new_n11963, new_n652);
nand_4 g11579(new_n11965, new_n11964, new_n549);
nand_4 g11580(new_n11966, new_n11965, new_n544);
nand_4 g11581(new_n11967, new_n11966, new_n660);
nand_4 g11582(new_n11968, new_n11967, new_n539);
nand_4 g11583(new_n11969, new_n11968, new_n534);
nand_4 g11584(new_n11970, new_n11969, new_n529);
nand_4 g11585(new_n11971, new_n11970, new_n668);
nand_4 g11586(new_n11972, new_n11971, new_n674_1);
nand_4 g11587(new_n11973, new_n11972, new_n681);
nand_4 g11588(new_n11974, new_n11973, new_n523);
nand_4 g11589(new_n11975, new_n11974, new_n687);
nand_4 g11590(new_n11976, new_n11975, new_n693);
nand_4 g11591(new_n11977, new_n11976, new_n699);
nand_4 g11592(new_n11978, new_n11977, new_n517);
nand_4 g11593(new_n11979, new_n11978, new_n705);
nand_4 g11594(new_n11980, new_n11979, new_n511);
nand_4 g11595(new_n11981, new_n11980, new_n711);
nand_4 g11596(new_n11982, new_n11981, new_n506);
nand_4 g11597(new_n11983, new_n11982, new_n719);
nand_4 g11598(new_n11984, new_n11983, new_n500);
nand_4 g11599(new_n11985, new_n11984, new_n727);
nand_4 g11600(new_n11986, new_n11985, new_n494);
nand_4 g11601(new_n11987, new_n11986, new_n735);
nand_4 g11602(new_n11988, new_n11987, new_n488);
nand_4 g11603(new_n11989, new_n11988, new_n743);
nand_4 g11604(new_n11990, new_n11989, new_n482);
nand_4 g11605(new_n11991, new_n11990, new_n751);
nand_4 g11606(new_n11992, new_n11991, new_n758);
not_3  g11607(new_n11993, new_n11992);
nor_4  g11608(new_n11994, new_n11993, new_n766);
nor_4  g11609(new_n11995, new_n11994, new_n477);
nor_4  g11610(new_n11996, new_n11995, new_n774);
nor_4  g11611(new_n11997, new_n11996, new_n781);
nor_4  g11612(new_n11998, new_n11997, new_n788);
nor_4  g11613(new_n11999, new_n11998, new_n471);
nor_4  g11614(new_n12000, new_n11999, new_n796);
nor_4  g11615(new_n12001, new_n12000, new_n804);
nor_4  g11616(new_n12002, new_n12001, new_n810);
nor_4  g11617(new_n12003, new_n12002, new_n2043);
nor_4  g11618(new_n12004, new_n12003, new_n2042);
nor_4  g11619(new_n12005, new_n12004, new_n2041);
nor_4  g11620(new_n12006, new_n12005, new_n2040);
nor_4  g11621(new_n12007, new_n12006, new_n2039);
nor_4  g11622(new_n12008, new_n12007, new_n2038);
nor_4  g11623(new_n12009_1, new_n12008, new_n2037);
nor_4  g11624(new_n12010, new_n12009_1, new_n2036);
nor_4  g11625(new_n12011, new_n12010, new_n2035);
nor_4  g11626(new_n12012_1, new_n12011, new_n2034);
nor_4  g11627(new_n12013, new_n12012_1, new_n2033);
nor_4  g11628(new_n12014, new_n12013, new_n2032);
nor_4  g11629(new_n12015, new_n12014, new_n2031);
nor_4  g11630(new_n12016, new_n12015, new_n2030);
nor_4  g11631(new_n12017, new_n12016, new_n2029);
nor_4  g11632(new_n12018, new_n12017, new_n2028);
nor_4  g11633(new_n12019, new_n12018, new_n2027_1);
nor_4  g11634(new_n12020, new_n12019, new_n2026);
not_3  g11635(new_n12021, new_n12020);
nand_4 g11636(new_n12022, new_n12021, new_n875);
nand_4 g11637(new_n12023, new_n12022, new_n881);
nand_4 g11638(new_n12024, new_n12023, new_n413);
nand_4 g11639(new_n12025_1, new_n12024, new_n889);
nand_4 g11640(new_n12026, new_n12025_1, new_n896);
nand_4 g11641(new_n12027, new_n12026, new_n901);
nand_4 g11642(new_n12028, new_n12027, n12927);
nor_4  g11643(n13639, new_n12028, new_n405);
nand_4 g11644(new_n12030, new_n1258, new_n900);
nand_4 g11645(new_n12031, new_n12030, new_n1256);
nand_4 g11646(new_n12032_1, new_n12031, new_n1251);
nand_4 g11647(new_n12033, new_n12032_1, new_n1457);
nand_4 g11648(new_n12034, new_n12033, new_n1462);
nand_4 g11649(new_n12035, new_n12034, new_n1468);
nand_4 g11650(new_n12036, new_n12035, new_n1247);
nand_4 g11651(new_n12037, new_n12036, new_n1474);
nand_4 g11652(new_n12038, new_n12037, new_n592);
nand_4 g11653(new_n12039, new_n12038, new_n585);
nand_4 g11654(new_n12040, new_n12039, new_n580);
nand_4 g11655(new_n12041, new_n12040, new_n600);
nand_4 g11656(new_n12042, new_n12041, new_n606);
nand_4 g11657(new_n12043, new_n12042, new_n612);
nand_4 g11658(new_n12044, new_n12043, new_n575);
nand_4 g11659(new_n12045, new_n12044, new_n619);
nand_4 g11660(new_n12046, new_n12045, new_n570);
nand_4 g11661(new_n12047, new_n12046, new_n625);
nand_4 g11662(new_n12048, new_n12047, new_n564);
nand_4 g11663(new_n12049, new_n12048, new_n632);
nand_4 g11664(new_n12050, new_n12049, new_n638);
nand_4 g11665(new_n12051, new_n12050, new_n559);
nand_4 g11666(new_n12052, new_n12051, new_n554);
nand_4 g11667(new_n12053, new_n12052, new_n646);
nand_4 g11668(new_n12054, new_n12053, new_n652);
nand_4 g11669(new_n12055, new_n12054, new_n549);
nand_4 g11670(new_n12056, new_n12055, new_n544);
nand_4 g11671(new_n12057, new_n12056, new_n660);
nand_4 g11672(new_n12058, new_n12057, new_n539);
nand_4 g11673(new_n12059, new_n12058, new_n534);
nand_4 g11674(new_n12060, new_n12059, new_n529);
nand_4 g11675(new_n12061, new_n12060, new_n668);
nand_4 g11676(new_n12062, new_n12061, new_n674_1);
nand_4 g11677(new_n12063, new_n12062, new_n681);
nand_4 g11678(new_n12064, new_n12063, new_n523);
nand_4 g11679(new_n12065, new_n12064, new_n687);
nand_4 g11680(new_n12066, new_n12065, new_n693);
nand_4 g11681(new_n12067, new_n12066, new_n699);
nand_4 g11682(new_n12068, new_n12067, new_n517);
nand_4 g11683(new_n12069, new_n12068, new_n705);
nand_4 g11684(new_n12070, new_n12069, new_n511);
nand_4 g11685(new_n12071, new_n12070, new_n711);
nand_4 g11686(new_n12072, new_n12071, new_n506);
nand_4 g11687(new_n12073, new_n12072, new_n719);
nand_4 g11688(new_n12074, new_n12073, new_n500);
nand_4 g11689(new_n12075, new_n12074, new_n727);
not_3  g11690(new_n12076, new_n12075);
nor_4  g11691(new_n12077, new_n12076, new_n495);
nor_4  g11692(new_n12078, new_n12077, new_n736);
nor_4  g11693(new_n12079, new_n12078, new_n489);
nor_4  g11694(new_n12080, new_n12079, new_n744);
nor_4  g11695(new_n12081, new_n12080, new_n483);
nor_4  g11696(new_n12082, new_n12081, new_n752);
nor_4  g11697(new_n12083, new_n12082, new_n759);
nor_4  g11698(new_n12084, new_n12083, new_n766);
nor_4  g11699(new_n12085, new_n12084, new_n477);
nor_4  g11700(new_n12086, new_n12085, new_n774);
nor_4  g11701(new_n12087, new_n12086, new_n781);
nor_4  g11702(new_n12088, new_n12087, new_n788);
nor_4  g11703(new_n12089, new_n12088, new_n471);
nor_4  g11704(new_n12090, new_n12089, new_n796);
nor_4  g11705(new_n12091, new_n12090, new_n804);
nor_4  g11706(new_n12092, new_n12091, new_n810);
nor_4  g11707(new_n12093, new_n12092, new_n2043);
nor_4  g11708(new_n12094, new_n12093, new_n2042);
nor_4  g11709(new_n12095, new_n12094, new_n2041);
nor_4  g11710(new_n12096, new_n12095, new_n2040);
nor_4  g11711(new_n12097, new_n12096, new_n2039);
nor_4  g11712(new_n12098, new_n12097, new_n2038);
nor_4  g11713(new_n12099, new_n12098, new_n2037);
nor_4  g11714(new_n12100, new_n12099, new_n2036);
not_3  g11715(new_n12101, new_n12100);
nand_4 g11716(new_n12102, new_n12101, new_n439);
nand_4 g11717(new_n12103, new_n12102, new_n841);
nand_4 g11718(new_n12104, new_n12103, new_n434);
nand_4 g11719(new_n12105, new_n12104, new_n429);
nand_4 g11720(new_n12106, new_n12105, new_n424);
nand_4 g11721(new_n12107, new_n12106, new_n850);
nand_4 g11722(new_n12108, new_n12107, new_n856);
nand_4 g11723(new_n12109, new_n12108, new_n863);
nand_4 g11724(new_n12110, new_n12109, new_n419);
nand_4 g11725(new_n12111, new_n12110, new_n869);
nand_4 g11726(new_n12112, new_n12111, new_n875);
nand_4 g11727(new_n12113, new_n12112, new_n881);
nand_4 g11728(new_n12114, new_n12113, new_n413);
nand_4 g11729(new_n12115, new_n12114, new_n889);
nand_4 g11730(new_n12116, new_n12115, n7282);
nor_4  g11731(n13658, new_n12116, new_n892);
not_3  g11732(new_n12118, n13231);
not_3  g11733(new_n12119, new_n1714);
nand_4 g11734(new_n12120, new_n12119, new_n12118);
nand_4 g11735(new_n12121, new_n12120, new_n1097);
nand_4 g11736(new_n12122, new_n12121, new_n1191);
nand_4 g11737(new_n12123, new_n12122, new_n1095);
nand_4 g11738(new_n12124, new_n12123, new_n1091);
nand_4 g11739(new_n12125, new_n12124, new_n1088);
nand_4 g11740(new_n12126, new_n12125, new_n1084);
nand_4 g11741(new_n12127, new_n12126, new_n1079);
nand_4 g11742(new_n12128, new_n12127, new_n1074);
nand_4 g11743(new_n12129, new_n12128, new_n1070);
nand_4 g11744(new_n12130, new_n12129, new_n1064);
nand_4 g11745(new_n12131, new_n12130, new_n1061);
nand_4 g11746(new_n12132, new_n12131, new_n1055);
nand_4 g11747(new_n12133, new_n12132, new_n1050);
nand_4 g11748(new_n12134, new_n12133, new_n1045);
nand_4 g11749(new_n12135, new_n12134, new_n1041);
nand_4 g11750(new_n12136, new_n12135, new_n1036);
nand_4 g11751(new_n12137, new_n12136, new_n1031);
nand_4 g11752(new_n12138, new_n12137, new_n1025);
nand_4 g11753(new_n12139, new_n12138, new_n1020);
nand_4 g11754(new_n12140, new_n12139, new_n1015);
nand_4 g11755(new_n12141, new_n12140, new_n1010);
nand_4 g11756(new_n12142_1, new_n12141, new_n1215);
nand_4 g11757(new_n12143, new_n12142_1, new_n1005);
nand_4 g11758(new_n12144, new_n12143, new_n1000);
nand_4 g11759(new_n12145, new_n12144, new_n994);
nand_4 g11760(new_n12146, new_n12145, new_n989);
nand_4 g11761(new_n12147, new_n12146, new_n984);
nand_4 g11762(new_n12148, new_n12147, new_n978);
nand_4 g11763(new_n12149, new_n12148, new_n973);
nand_4 g11764(new_n12150, new_n12149, new_n967);
nand_4 g11765(new_n12151, new_n12150, new_n964);
nand_4 g11766(new_n12152, new_n12151, new_n960);
nand_4 g11767(new_n12153, new_n12152, new_n957);
nand_4 g11768(new_n12154, new_n12153, new_n952);
nand_4 g11769(new_n12155, new_n12154, new_n948_1);
nand_4 g11770(new_n12156, new_n12155, new_n943);
nand_4 g11771(new_n12157, new_n12156, new_n938);
nand_4 g11772(new_n12158, new_n12157, new_n934);
nand_4 g11773(new_n12159, new_n12158, new_n929);
nand_4 g11774(new_n12160, new_n12159, new_n925);
nand_4 g11775(new_n12161, new_n12160, new_n2194);
nand_4 g11776(new_n12162, new_n12161, new_n2191);
nand_4 g11777(new_n12163, new_n12162, new_n2190);
nand_4 g11778(new_n12164, new_n12163, new_n2186);
nand_4 g11779(new_n12165, new_n12164, new_n2183);
nand_4 g11780(new_n12166_1, new_n12165, new_n2179);
nand_4 g11781(new_n12167, new_n12166_1, new_n2175_1);
nand_4 g11782(new_n12168, new_n12167, new_n2171);
nand_4 g11783(new_n12169, new_n12168, new_n2168);
nand_4 g11784(new_n12170, new_n12169, new_n2165);
not_3  g11785(new_n12171, new_n12170);
nor_4  g11786(new_n12172, new_n12171, new_n2507);
nor_4  g11787(new_n12173, new_n12172, new_n2506);
nor_4  g11788(new_n12174, new_n12173, new_n2505);
nor_4  g11789(new_n12175, new_n12174, new_n2504);
nor_4  g11790(new_n12176, new_n12175, new_n2503);
nor_4  g11791(new_n12177, new_n12176, new_n2502);
nor_4  g11792(new_n12178, new_n12177, new_n2790);
nor_4  g11793(new_n12179, new_n12178, new_n2789);
nor_4  g11794(new_n12180, new_n12179, new_n2788);
nor_4  g11795(new_n12181, new_n12180, new_n2305);
nor_4  g11796(new_n12182, new_n12181, new_n2304);
nor_4  g11797(new_n12183, new_n12182, new_n2303);
nor_4  g11798(new_n12184, new_n12183, new_n2302);
nor_4  g11799(new_n12185, new_n12184, new_n2301);
nor_4  g11800(new_n12186, new_n12185, new_n2300);
nor_4  g11801(new_n12187, new_n12186, new_n2299);
nor_4  g11802(new_n12188, new_n12187, new_n2298);
nor_4  g11803(new_n12189, new_n12188, new_n2297);
nor_4  g11804(new_n12190, new_n12189, new_n2296);
nor_4  g11805(new_n12191, new_n12190, new_n2295);
nor_4  g11806(new_n12192, new_n12191, new_n2294);
nor_4  g11807(new_n12193, new_n12192, new_n2293);
nor_4  g11808(new_n12194, new_n12193, new_n2292);
nor_4  g11809(new_n12195, new_n12194, new_n2291);
nor_4  g11810(new_n12196, new_n12195, new_n2290);
not_3  g11811(new_n12197, new_n12196);
nand_4 g11812(new_n12198, new_n12197, new_n1746);
nand_4 g11813(new_n12199, new_n12198, new_n1742);
nand_4 g11814(new_n12200, new_n12199, new_n1738);
nand_4 g11815(new_n12201, new_n12200, new_n1736);
nand_4 g11816(new_n12202, new_n12201, new_n1732);
nand_4 g11817(new_n12203, new_n12202, new_n1729);
nand_4 g11818(new_n12204, new_n12203, new_n1726);
nand_4 g11819(new_n12205, new_n12204, new_n1724);
nand_4 g11820(new_n12206, new_n12205, new_n1721);
nand_4 g11821(new_n12207, new_n12206, n74);
nor_4  g11822(n13693, new_n12207, new_n616);
not_3  g11823(new_n12209, new_n2173);
nand_4 g11824(new_n12210, new_n2170, new_n458);
nand_4 g11825(new_n12211, new_n12210, new_n455);
nand_4 g11826(new_n12212, new_n12211, new_n449);
nand_4 g11827(new_n12213, new_n12212, new_n827);
nand_4 g11828(new_n12214, new_n12213, new_n833);
nand_4 g11829(new_n12215, new_n12214, new_n444);
nand_4 g11830(new_n12216, new_n12215, new_n439);
nand_4 g11831(new_n12217, new_n12216, new_n841);
nand_4 g11832(new_n12218_1, new_n12217, new_n434);
nand_4 g11833(new_n12219, new_n12218_1, new_n429);
nand_4 g11834(new_n12220, new_n12219, new_n424);
nand_4 g11835(new_n12221, new_n12220, new_n850);
nand_4 g11836(new_n12222, new_n12221, new_n856);
nand_4 g11837(new_n12223, new_n12222, new_n863);
nand_4 g11838(new_n12224, new_n12223, new_n419);
nand_4 g11839(new_n12225, new_n12224, new_n869);
nand_4 g11840(new_n12226, new_n12225, new_n875);
nand_4 g11841(new_n12227, new_n12226, new_n881);
nand_4 g11842(new_n12228, new_n12227, new_n413);
nand_4 g11843(new_n12229, new_n12228, new_n889);
nand_4 g11844(new_n12230, new_n12229, new_n896);
nand_4 g11845(new_n12231, new_n12230, new_n901);
nand_4 g11846(new_n12232_1, new_n12231, new_n408);
nand_4 g11847(new_n12233, new_n12232_1, new_n908);
nand_4 g11848(new_n12234, new_n12233, new_n403);
nand_4 g11849(new_n12235, new_n12234, new_n398);
nand_4 g11850(new_n12236, new_n12235, new_n393);
nand_4 g11851(new_n12237, new_n12236, new_n916);
nand_4 g11852(new_n12238, new_n12237, new_n1123);
nand_4 g11853(new_n12239, new_n12238, new_n1164);
nand_4 g11854(new_n12240, new_n12239, new_n1120);
nand_4 g11855(new_n12241, new_n12240, new_n1169);
nand_4 g11856(new_n12242, new_n12241, new_n1116);
nand_4 g11857(new_n12243, new_n12242, new_n1111);
nand_4 g11858(new_n12244, new_n12243, new_n1106);
nand_4 g11859(new_n12245, new_n12244, new_n1178);
nand_4 g11860(new_n12246, new_n12245, new_n1183);
nand_4 g11861(new_n12247, new_n12246, new_n1102);
nand_4 g11862(new_n12248, new_n12247, new_n1099);
nand_4 g11863(new_n12249, new_n12248, new_n1191);
nand_4 g11864(new_n12250, new_n12249, new_n1095);
nand_4 g11865(new_n12251, new_n12250, new_n1091);
nand_4 g11866(new_n12252, new_n12251, new_n1088);
nand_4 g11867(new_n12253, new_n12252, new_n1084);
nand_4 g11868(new_n12254, new_n12253, new_n1079);
nand_4 g11869(new_n12255, new_n12254, new_n1074);
nand_4 g11870(new_n12256, new_n12255, new_n1070);
nand_4 g11871(new_n12257, new_n12256, new_n1064);
nand_4 g11872(new_n12258, new_n12257, new_n1061);
nand_4 g11873(new_n12259, new_n12258, new_n1055);
nand_4 g11874(new_n12260, new_n12259, new_n1050);
not_3  g11875(new_n12261, new_n12260);
nor_4  g11876(new_n12262, new_n12261, new_n1046);
nor_4  g11877(new_n12263, new_n12262, new_n1042);
nor_4  g11878(new_n12264, new_n12263, new_n1037);
nor_4  g11879(new_n12265, new_n12264, new_n1032);
nor_4  g11880(new_n12266, new_n12265, new_n1026);
nor_4  g11881(new_n12267, new_n12266, new_n1021);
nor_4  g11882(new_n12268, new_n12267, new_n1016);
nor_4  g11883(new_n12269, new_n12268, new_n1011);
nor_4  g11884(new_n12270_1, new_n12269, new_n1216);
nor_4  g11885(new_n12271, new_n12270_1, new_n1006);
nor_4  g11886(new_n12272, new_n12271, new_n1001);
nor_4  g11887(new_n12273, new_n12272, new_n995);
nor_4  g11888(new_n12274, new_n12273, new_n990);
nor_4  g11889(new_n12275, new_n12274, new_n985);
nor_4  g11890(new_n12276, new_n12275, new_n979);
nor_4  g11891(new_n12277, new_n12276, new_n974);
nor_4  g11892(new_n12278, new_n12277, new_n968);
nor_4  g11893(new_n12279, new_n12278, new_n965);
nor_4  g11894(new_n12280, new_n12279, new_n961);
nor_4  g11895(new_n12281, new_n12280, new_n958);
nor_4  g11896(new_n12282, new_n12281, new_n953);
nor_4  g11897(new_n12283, new_n12282, new_n3536);
nor_4  g11898(new_n12284, new_n12283, new_n3535);
nor_4  g11899(new_n12285, new_n12284, new_n3534);
nor_4  g11900(new_n12286, new_n12285, new_n2520);
nor_4  g11901(new_n12287, new_n12286, new_n2519);
nor_4  g11902(new_n12288, new_n12287, new_n2518);
not_3  g11903(new_n12289, new_n12288);
nand_4 g11904(new_n12290, new_n12289, new_n2194);
nand_4 g11905(new_n12291, new_n12290, new_n2191);
nand_4 g11906(new_n12292, new_n12291, new_n2190);
nand_4 g11907(new_n12293, new_n12292, new_n2186);
nand_4 g11908(new_n12294, new_n12293, new_n2183);
nand_4 g11909(new_n12295, new_n12294, new_n2179);
nand_4 g11910(new_n12296, new_n12295, n9921);
nor_4  g11911(n13760, new_n12296, new_n12209);
nand_4 g11912(new_n12298, new_n1081, new_n1079);
nand_4 g11913(new_n12299, new_n12298, new_n1074);
nand_4 g11914(new_n12300, new_n12299, new_n1070);
nand_4 g11915(new_n12301, new_n12300, new_n1064);
nand_4 g11916(new_n12302, new_n12301, new_n1061);
nand_4 g11917(new_n12303, new_n12302, new_n1055);
nand_4 g11918(new_n12304, new_n12303, new_n1050);
nand_4 g11919(new_n12305, new_n12304, new_n1045);
nand_4 g11920(new_n12306, new_n12305, new_n1041);
nand_4 g11921(new_n12307, new_n12306, new_n1036);
nand_4 g11922(new_n12308, new_n12307, new_n1031);
nand_4 g11923(new_n12309, new_n12308, new_n1025);
nand_4 g11924(new_n12310, new_n12309, new_n1020);
nand_4 g11925(new_n12311, new_n12310, new_n1015);
nand_4 g11926(new_n12312, new_n12311, new_n1010);
nand_4 g11927(new_n12313, new_n12312, new_n1215);
nand_4 g11928(new_n12314, new_n12313, new_n1005);
nand_4 g11929(new_n12315, new_n12314, new_n1000);
nand_4 g11930(new_n12316, new_n12315, new_n994);
nand_4 g11931(new_n12317, new_n12316, new_n989);
nand_4 g11932(new_n12318, new_n12317, new_n984);
nand_4 g11933(new_n12319, new_n12318, new_n978);
nand_4 g11934(new_n12320, new_n12319, new_n973);
nand_4 g11935(new_n12321_1, new_n12320, new_n967);
nand_4 g11936(new_n12322, new_n12321_1, new_n964);
nand_4 g11937(new_n12323, new_n12322, new_n960);
nand_4 g11938(new_n12324, new_n12323, new_n957);
nand_4 g11939(new_n12325, new_n12324, new_n952);
nand_4 g11940(new_n12326, new_n12325, new_n948_1);
nand_4 g11941(new_n12327, new_n12326, new_n943);
nand_4 g11942(new_n12328, new_n12327, new_n938);
nand_4 g11943(new_n12329, new_n12328, new_n934);
nand_4 g11944(new_n12330, new_n12329, new_n929);
nand_4 g11945(new_n12331, new_n12330, new_n925);
nand_4 g11946(new_n12332, new_n12331, new_n2194);
not_3  g11947(new_n12333, new_n12332);
nor_4  g11948(new_n12334, new_n12333, new_n2516);
nor_4  g11949(new_n12335, new_n12334, new_n2515);
nor_4  g11950(new_n12336_1, new_n12335, new_n2514);
nor_4  g11951(new_n12337, new_n12336_1, new_n2513);
nor_4  g11952(new_n12338, new_n12337, new_n2512);
nor_4  g11953(new_n12339, new_n12338, new_n2511);
nor_4  g11954(new_n12340, new_n12339, new_n2510);
nor_4  g11955(new_n12341, new_n12340, new_n2509);
nor_4  g11956(new_n12342, new_n12341, new_n2508);
nor_4  g11957(new_n12343, new_n12342, new_n2507);
nor_4  g11958(new_n12344, new_n12343, new_n2506);
nor_4  g11959(new_n12345, new_n12344, new_n2505);
nor_4  g11960(new_n12346, new_n12345, new_n2504);
nor_4  g11961(new_n12347, new_n12346, new_n2503);
nor_4  g11962(new_n12348, new_n12347, new_n2502);
nor_4  g11963(new_n12349, new_n12348, new_n2790);
nor_4  g11964(new_n12350, new_n12349, new_n2789);
nor_4  g11965(new_n12351, new_n12350, new_n2788);
nor_4  g11966(new_n12352, new_n12351, new_n2305);
not_3  g11967(new_n12353, new_n12352);
nand_4 g11968(new_n12354, new_n12353, new_n1794);
nand_4 g11969(new_n12355_1, new_n12354, new_n1825);
nand_4 g11970(new_n12356, new_n12355_1, new_n1789);
nand_4 g11971(new_n12357, new_n12356, new_n1785);
nand_4 g11972(new_n12358, new_n12357, new_n1780);
nand_4 g11973(new_n12359, new_n12358, new_n1777);
nand_4 g11974(new_n12360, new_n12359, new_n1774);
nand_4 g11975(new_n12361, new_n12360, new_n1834);
nand_4 g11976(new_n12362, new_n12361, new_n1769);
nand_4 g11977(new_n12363, new_n12362, new_n1766);
nand_4 g11978(new_n12364, new_n12363, new_n1762);
nand_4 g11979(new_n12365, new_n12364, new_n1758);
nand_4 g11980(new_n12366, new_n12365, new_n1754);
nand_4 g11981(new_n12367, new_n12366, new_n1751);
nand_4 g11982(new_n12368, new_n12367, new_n1748);
nand_4 g11983(new_n12369, new_n12368, new_n1746);
nand_4 g11984(new_n12370, new_n12369, new_n1742);
nand_4 g11985(new_n12371, new_n12370, new_n1738);
nand_4 g11986(new_n12372, new_n12371, new_n1736);
nand_4 g11987(new_n12373, new_n12372, new_n1732);
nand_4 g11988(new_n12374, new_n12373, new_n1729);
nand_4 g11989(new_n12375, new_n12374, new_n1726);
nand_4 g11990(new_n12376, new_n12375, new_n1724);
nand_4 g11991(new_n12377, new_n12376, new_n1721);
nand_4 g11992(new_n12378, new_n12377, new_n1718);
nand_4 g11993(new_n12379, new_n12378, new_n1715);
nand_4 g11994(new_n12380, new_n12379, new_n1711);
nand_4 g11995(new_n12381, new_n12380, new_n1708);
nand_4 g11996(new_n12382, new_n12381, new_n1705);
nand_4 g11997(new_n12383, new_n12382, new_n1703);
nand_4 g11998(new_n12384, new_n12383, n3367);
nor_4  g11999(n13853, new_n12384, new_n556);
not_3  g12000(new_n12386, n7450);
not_3  g12001(new_n12387, new_n942);
nand_4 g12002(new_n12388, new_n12387, new_n12386);
nand_4 g12003(new_n12389, new_n12388, new_n756);
nand_4 g12004(new_n12390, new_n12389, new_n765);
nand_4 g12005(new_n12391, new_n12390, new_n476);
nand_4 g12006(new_n12392, new_n12391, new_n773);
nand_4 g12007(new_n12393, new_n12392, new_n780);
nand_4 g12008(new_n12394, new_n12393, new_n787);
nand_4 g12009(new_n12395, new_n12394, new_n470);
nand_4 g12010(new_n12396, new_n12395, new_n795);
nand_4 g12011(new_n12397, new_n12396, new_n803);
nand_4 g12012(new_n12398, new_n12397, new_n809);
nand_4 g12013(new_n12399, new_n12398, new_n465);
nand_4 g12014(new_n12400, new_n12399, new_n818);
nand_4 g12015(new_n12401, new_n12400, new_n460);
nand_4 g12016(new_n12402, new_n12401, new_n455);
nand_4 g12017(new_n12403, new_n12402, new_n449);
nand_4 g12018(new_n12404, new_n12403, new_n827);
nand_4 g12019(new_n12405, new_n12404, new_n833);
nand_4 g12020(new_n12406, new_n12405, new_n444);
nand_4 g12021(new_n12407, new_n12406, new_n439);
nand_4 g12022(new_n12408, new_n12407, new_n841);
nand_4 g12023(new_n12409, new_n12408, new_n434);
nand_4 g12024(new_n12410, new_n12409, new_n429);
nand_4 g12025(new_n12411, new_n12410, new_n424);
nand_4 g12026(new_n12412, new_n12411, new_n850);
nand_4 g12027(new_n12413, new_n12412, new_n856);
nand_4 g12028(new_n12414, new_n12413, new_n863);
nand_4 g12029(new_n12415, new_n12414, new_n419);
nand_4 g12030(new_n12416, new_n12415, new_n869);
nand_4 g12031(new_n12417, new_n12416, new_n875);
nand_4 g12032(new_n12418, new_n12417, new_n881);
nand_4 g12033(new_n12419, new_n12418, new_n413);
nand_4 g12034(new_n12420, new_n12419, new_n889);
nand_4 g12035(new_n12421, new_n12420, new_n896);
nand_4 g12036(new_n12422, new_n12421, new_n901);
nand_4 g12037(new_n12423, new_n12422, new_n408);
nand_4 g12038(new_n12424, new_n12423, new_n908);
nand_4 g12039(new_n12425, new_n12424, new_n403);
nand_4 g12040(new_n12426, new_n12425, new_n398);
nand_4 g12041(new_n12427, new_n12426, new_n393);
nand_4 g12042(new_n12428, new_n12427, new_n916);
nand_4 g12043(new_n12429, new_n12428, new_n1123);
nand_4 g12044(new_n12430, new_n12429, new_n1164);
nand_4 g12045(new_n12431, new_n12430, new_n1120);
nand_4 g12046(new_n12432, new_n12431, new_n1169);
nand_4 g12047(new_n12433, new_n12432, new_n1116);
not_3  g12048(new_n12434, new_n12433);
nor_4  g12049(new_n12435, new_n12434, new_n1527);
nor_4  g12050(new_n12436, new_n12435, new_n1526);
nor_4  g12051(new_n12437, new_n12436, new_n1525);
nor_4  g12052(new_n12438, new_n12437, new_n1524);
nor_4  g12053(new_n12439, new_n12438, new_n1523);
nor_4  g12054(new_n12440, new_n12439, new_n1522);
nor_4  g12055(new_n12441, new_n12440, new_n1521);
nor_4  g12056(new_n12442, new_n12441, new_n1520);
nor_4  g12057(new_n12443, new_n12442, new_n1519);
nor_4  g12058(new_n12444, new_n12443, new_n1518);
nor_4  g12059(new_n12445, new_n12444, new_n1517);
nor_4  g12060(new_n12446, new_n12445, new_n1516);
nor_4  g12061(new_n12447, new_n12446, new_n1075);
nor_4  g12062(new_n12448, new_n12447, new_n1071);
nor_4  g12063(new_n12449, new_n12448, new_n1065);
nor_4  g12064(new_n12450, new_n12449, new_n1062);
nor_4  g12065(new_n12451, new_n12450, new_n1056);
nor_4  g12066(new_n12452, new_n12451, new_n1051);
nor_4  g12067(new_n12453, new_n12452, new_n1046);
nor_4  g12068(new_n12454, new_n12453, new_n1042);
nor_4  g12069(new_n12455, new_n12454, new_n1037);
nor_4  g12070(new_n12456, new_n12455, new_n1032);
nor_4  g12071(new_n12457, new_n12456, new_n1026);
nor_4  g12072(new_n12458, new_n12457, new_n1021);
not_3  g12073(new_n12459, new_n12458);
nand_4 g12074(new_n12460, new_n12459, new_n1015);
nand_4 g12075(new_n12461, new_n12460, new_n1010);
nand_4 g12076(new_n12462, new_n12461, new_n1215);
nand_4 g12077(new_n12463, new_n12462, new_n1005);
nand_4 g12078(new_n12464, new_n12463, new_n1000);
nand_4 g12079(new_n12465, new_n12464, new_n994);
nand_4 g12080(new_n12466, new_n12465, new_n989);
nand_4 g12081(new_n12467, new_n12466, new_n984);
nand_4 g12082(new_n12468, new_n12467, new_n978);
nand_4 g12083(new_n12469, new_n12468, new_n973);
nand_4 g12084(new_n12470, new_n12469, new_n967);
nand_4 g12085(new_n12471, new_n12470, new_n964);
nand_4 g12086(new_n12472, new_n12471, new_n960);
nand_4 g12087(new_n12473, new_n12472, new_n957);
nand_4 g12088(new_n12474, new_n12473, new_n952);
nand_4 g12089(new_n12475, new_n12474, n7972);
nor_4  g12090(n13870, new_n12475, new_n945);
nand_4 g12091(new_n12477, new_n1369, new_n1367);
nand_4 g12092(new_n12478, new_n12477, new_n1363);
nand_4 g12093(new_n12479, new_n12478, new_n1360);
nand_4 g12094(new_n12480, new_n12479, new_n1357);
nand_4 g12095(new_n12481, new_n12480, new_n1354);
nand_4 g12096(new_n12482, new_n12481, new_n1352);
nand_4 g12097(new_n12483, new_n12482, new_n1350);
nand_4 g12098(new_n12484, new_n12483, new_n1347_1);
nand_4 g12099(new_n12485, new_n12484, new_n1344);
nand_4 g12100(new_n12486, new_n12485, new_n1341);
nand_4 g12101(new_n12487, new_n12486, new_n1338);
nand_4 g12102(new_n12488, new_n12487, new_n1395);
nand_4 g12103(new_n12489, new_n12488, new_n1335);
nand_4 g12104(new_n12490, new_n12489, new_n1332);
nand_4 g12105(new_n12491, new_n12490, new_n1328);
nand_4 g12106(new_n12492, new_n12491, new_n1403);
nand_4 g12107(new_n12493, new_n12492, new_n1325);
nand_4 g12108(new_n12494, new_n12493, new_n1410);
nand_4 g12109(new_n12495, new_n12494, new_n1413);
nand_4 g12110(new_n12496, new_n12495, new_n1322);
nand_4 g12111(new_n12497, new_n12496, new_n1317);
nand_4 g12112(new_n12498, new_n12497, new_n1315);
nand_4 g12113(new_n12499, new_n12498, new_n1419);
nand_4 g12114(new_n12500, new_n12499, new_n1310);
nand_4 g12115(new_n12501, new_n12500, new_n1305);
nand_4 g12116(new_n12502, new_n12501, new_n1427);
nand_4 g12117(new_n12503, new_n12502, new_n1431);
nand_4 g12118(new_n12504, new_n12503, new_n1302);
nand_4 g12119(new_n12505, new_n12504, new_n1298);
nand_4 g12120(new_n12506, new_n12505, new_n1295);
nand_4 g12121(new_n12507, new_n12506, new_n1291);
nand_4 g12122(new_n12508, new_n12507, new_n1288);
nand_4 g12123(new_n12509, new_n12508, new_n1284);
nand_4 g12124(new_n12510, new_n12509, new_n1280);
nand_4 g12125(new_n12511, new_n12510, new_n1275);
nand_4 g12126(new_n12512, new_n12511, new_n1445);
nand_4 g12127(new_n12513, new_n12512, new_n1270);
nand_4 g12128(new_n12514, new_n12513, new_n1265_1);
nand_4 g12129(new_n12515, new_n12514, new_n1260);
nand_4 g12130(new_n12516, new_n12515, new_n1256);
nand_4 g12131(new_n12517, new_n12516, new_n1251);
nand_4 g12132(new_n12518, new_n12517, new_n1457);
nand_4 g12133(new_n12519, new_n12518, new_n1462);
nand_4 g12134(new_n12520, new_n12519, new_n1468);
nand_4 g12135(new_n12521, new_n12520, new_n1247);
nand_4 g12136(new_n12522, new_n12521, new_n1474);
nand_4 g12137(new_n12523, new_n12522, new_n592);
nand_4 g12138(new_n12524, new_n12523, new_n585);
nand_4 g12139(new_n12525, new_n12524, new_n580);
nand_4 g12140(new_n12526, new_n12525, new_n600);
nand_4 g12141(new_n12527, new_n12526, new_n606);
not_3  g12142(new_n12528, new_n12527);
nor_4  g12143(new_n12529, new_n12528, new_n1239);
nor_4  g12144(new_n12530, new_n12529, new_n3082);
nor_4  g12145(new_n12531, new_n12530, new_n3081);
nor_4  g12146(new_n12532, new_n12531, new_n3080);
nor_4  g12147(new_n12533, new_n12532, new_n3079);
nor_4  g12148(new_n12534, new_n12533, new_n3078);
nor_4  g12149(new_n12535_1, new_n12534, new_n3077);
nor_4  g12150(new_n12536, new_n12535_1, new_n3076);
nor_4  g12151(new_n12537, new_n12536, new_n3075);
nor_4  g12152(new_n12538, new_n12537, new_n3074);
nor_4  g12153(new_n12539, new_n12538, new_n3073);
nor_4  g12154(new_n12540, new_n12539, new_n3072);
nor_4  g12155(new_n12541, new_n12540, new_n3071);
nor_4  g12156(new_n12542, new_n12541, new_n3070);
nor_4  g12157(new_n12543, new_n12542, new_n3069);
nor_4  g12158(new_n12544, new_n12543, new_n3068);
nor_4  g12159(new_n12545, new_n12544, new_n3067);
nor_4  g12160(new_n12546, new_n12545, new_n3066);
nor_4  g12161(new_n12547, new_n12546, new_n3065);
nor_4  g12162(new_n12548, new_n12547, new_n3064);
nor_4  g12163(new_n12549, new_n12548, new_n3063);
nor_4  g12164(new_n12550, new_n12549, new_n3062);
nor_4  g12165(new_n12551, new_n12550, new_n3061);
nor_4  g12166(new_n12552, new_n12551, new_n3354);
nor_4  g12167(new_n12553, new_n12552, new_n3353);
nor_4  g12168(new_n12554, new_n12553, new_n3352);
nor_4  g12169(new_n12555, new_n12554, new_n3351);
not_3  g12170(new_n12556, new_n12555);
nand_4 g12171(new_n12557, new_n12556, new_n511);
nand_4 g12172(new_n12558, new_n12557, new_n711);
nand_4 g12173(new_n12559, new_n12558, new_n506);
nand_4 g12174(new_n12560, new_n12559, new_n719);
nand_4 g12175(new_n12561, new_n12560, new_n500);
nand_4 g12176(new_n12562, new_n12561, new_n727);
nand_4 g12177(new_n12563, new_n12562, n11158);
nor_4  g12178(n13953, new_n12563, new_n491);
nand_4 g12179(new_n12565, new_n1858, new_n558);
nand_4 g12180(new_n12566, new_n12565, new_n1864);
nand_4 g12181(new_n12567, new_n12566, new_n1699);
nand_4 g12182(new_n12568, new_n12567, new_n1697);
nand_4 g12183(new_n12569, new_n12568, new_n1871);
nand_4 g12184(new_n12570, new_n12569, new_n1694);
nand_4 g12185(new_n12571, new_n12570, new_n1690);
nand_4 g12186(new_n12572, new_n12571, new_n1878);
nand_4 g12187(new_n12573_1, new_n12572, new_n1882);
nand_4 g12188(new_n12574, new_n12573_1, new_n1686);
nand_4 g12189(new_n12575, new_n12574, new_n1682);
nand_4 g12190(new_n12576, new_n12575, new_n1678);
nand_4 g12191(new_n12577, new_n12576, new_n1674);
nand_4 g12192(new_n12578, new_n12577, new_n1890);
nand_4 g12193(new_n12579, new_n12578, new_n1669);
nand_4 g12194(new_n12580, new_n12579, new_n1665);
nand_4 g12195(new_n12581, new_n12580, new_n1661);
nand_4 g12196(new_n12582, new_n12581, new_n1657);
nand_4 g12197(new_n12583, new_n12582, new_n1652);
nand_4 g12198(new_n12584, new_n12583, new_n1648);
nand_4 g12199(new_n12585, new_n12584, new_n1644);
nand_4 g12200(new_n12586, new_n12585, new_n1640);
nand_4 g12201(new_n12587, new_n12586, new_n1636);
nand_4 g12202(new_n12588, new_n12587, new_n1632);
nand_4 g12203(new_n12589, new_n12588, new_n1378);
nand_4 g12204(new_n12590, new_n12589, new_n1372);
nand_4 g12205(new_n12591, new_n12590, new_n1367);
nand_4 g12206(new_n12592, new_n12591, new_n1363);
nand_4 g12207(new_n12593, new_n12592, new_n1360);
nand_4 g12208(new_n12594, new_n12593, new_n1357);
nand_4 g12209(new_n12595, new_n12594, new_n1354);
nand_4 g12210(new_n12596, new_n12595, new_n1352);
nand_4 g12211(new_n12597, new_n12596, new_n1350);
nand_4 g12212(new_n12598, new_n12597, new_n1347_1);
nand_4 g12213(new_n12599, new_n12598, new_n1344);
nand_4 g12214(new_n12600, new_n12599, new_n1341);
nand_4 g12215(new_n12601, new_n12600, new_n1338);
nand_4 g12216(new_n12602, new_n12601, new_n1395);
nand_4 g12217(new_n12603, new_n12602, new_n1335);
nand_4 g12218(new_n12604, new_n12603, new_n1332);
nand_4 g12219(new_n12605, new_n12604, new_n1328);
nand_4 g12220(new_n12606, new_n12605, new_n1403);
nand_4 g12221(new_n12607, new_n12606, new_n1325);
nand_4 g12222(new_n12608, new_n12607, new_n1410);
nand_4 g12223(new_n12609, new_n12608, new_n1413);
nand_4 g12224(new_n12610, new_n12609, new_n1322);
nand_4 g12225(new_n12611, new_n12610, new_n1317);
nand_4 g12226(new_n12612, new_n12611, new_n1315);
nand_4 g12227(new_n12613, new_n12612, new_n1419);
nand_4 g12228(new_n12614_1, new_n12613, new_n1310);
nand_4 g12229(new_n12615, new_n12614_1, new_n1305);
not_3  g12230(new_n12616, new_n12615);
nor_4  g12231(new_n12617, new_n12616, new_n2402);
nor_4  g12232(new_n12618, new_n12617, new_n2401);
nor_4  g12233(new_n12619, new_n12618, new_n2400);
nor_4  g12234(new_n12620, new_n12619, new_n2399);
nor_4  g12235(new_n12621, new_n12620, new_n2398);
nor_4  g12236(new_n12622, new_n12621, new_n2397);
nor_4  g12237(new_n12623, new_n12622, new_n2396);
nor_4  g12238(new_n12624, new_n12623, new_n2395);
nor_4  g12239(new_n12625, new_n12624, new_n1281);
nor_4  g12240(new_n12626, new_n12625, new_n1276);
nor_4  g12241(new_n12627, new_n12626, new_n1446);
nor_4  g12242(new_n12628, new_n12627, new_n1271);
nor_4  g12243(new_n12629, new_n12628, new_n1266);
nor_4  g12244(new_n12630, new_n12629, new_n1261);
nor_4  g12245(new_n12631, new_n12630, new_n1257);
nor_4  g12246(new_n12632, new_n12631, new_n1252);
nor_4  g12247(new_n12633, new_n12632, new_n1458);
nor_4  g12248(new_n12634, new_n12633, new_n1463);
nor_4  g12249(new_n12635, new_n12634, new_n1469);
nor_4  g12250(new_n12636, new_n12635, new_n1248);
nor_4  g12251(new_n12637, new_n12636, new_n1475);
nor_4  g12252(new_n12638, new_n12637, new_n1244);
nor_4  g12253(new_n12639, new_n12638, new_n1243);
nor_4  g12254(new_n12640, new_n12639, new_n1242);
nor_4  g12255(new_n12641, new_n12640, new_n1241);
nor_4  g12256(new_n12642, new_n12641, new_n1240);
nor_4  g12257(new_n12643, new_n12642, new_n1239);
not_3  g12258(new_n12644, new_n12643);
nand_4 g12259(new_n12645, new_n12644, new_n575);
nand_4 g12260(new_n12646, new_n12645, new_n619);
nand_4 g12261(new_n12647, new_n12646, new_n570);
nand_4 g12262(new_n12648, new_n12647, new_n625);
nand_4 g12263(new_n12649, new_n12648, new_n564);
nand_4 g12264(new_n12650, new_n12649, new_n632);
nand_4 g12265(new_n12651, new_n12650, n2334);
nor_4  g12266(n13959, new_n12651, new_n635);
not_3  g12267(new_n12653, new_n427_1);
nand_4 g12268(new_n12654, new_n1431, new_n12653);
nand_4 g12269(new_n12655, new_n12654, new_n1302);
nand_4 g12270(new_n12656, new_n12655, new_n1298);
nand_4 g12271(new_n12657, new_n12656, new_n1295);
nand_4 g12272(new_n12658, new_n12657, new_n1291);
nand_4 g12273(new_n12659, new_n12658, new_n1288);
nand_4 g12274(new_n12660, new_n12659, new_n1284);
nand_4 g12275(new_n12661, new_n12660, new_n1280);
nand_4 g12276(new_n12662, new_n12661, new_n1275);
nand_4 g12277(new_n12663, new_n12662, new_n1445);
nand_4 g12278(new_n12664, new_n12663, new_n1270);
nand_4 g12279(new_n12665, new_n12664, new_n1265_1);
nand_4 g12280(new_n12666, new_n12665, new_n1260);
nand_4 g12281(new_n12667, new_n12666, new_n1256);
nand_4 g12282(new_n12668, new_n12667, new_n1251);
nand_4 g12283(new_n12669, new_n12668, new_n1457);
nand_4 g12284(new_n12670, new_n12669, new_n1462);
nand_4 g12285(new_n12671, new_n12670, new_n1468);
nand_4 g12286(new_n12672, new_n12671, new_n1247);
nand_4 g12287(new_n12673, new_n12672, new_n1474);
nand_4 g12288(new_n12674, new_n12673, new_n592);
nand_4 g12289(new_n12675, new_n12674, new_n585);
nand_4 g12290(new_n12676, new_n12675, new_n580);
nand_4 g12291(new_n12677, new_n12676, new_n600);
nand_4 g12292(new_n12678, new_n12677, new_n606);
nand_4 g12293(new_n12679, new_n12678, new_n612);
nand_4 g12294(new_n12680, new_n12679, new_n575);
nand_4 g12295(new_n12681, new_n12680, new_n619);
nand_4 g12296(new_n12682, new_n12681, new_n570);
nand_4 g12297(new_n12683, new_n12682, new_n625);
nand_4 g12298(new_n12684, new_n12683, new_n564);
nand_4 g12299(new_n12685, new_n12684, new_n632);
nand_4 g12300(new_n12686, new_n12685, new_n638);
nand_4 g12301(new_n12687, new_n12686, new_n559);
nand_4 g12302(new_n12688, new_n12687, new_n554);
nand_4 g12303(new_n12689, new_n12688, new_n646);
nand_4 g12304(new_n12690, new_n12689, new_n652);
nand_4 g12305(new_n12691, new_n12690, new_n549);
nand_4 g12306(new_n12692, new_n12691, new_n544);
nand_4 g12307(new_n12693, new_n12692, new_n660);
nand_4 g12308(new_n12694, new_n12693, new_n539);
nand_4 g12309(new_n12695, new_n12694, new_n534);
nand_4 g12310(new_n12696, new_n12695, new_n529);
nand_4 g12311(new_n12697, new_n12696, new_n668);
nand_4 g12312(new_n12698, new_n12697, new_n674_1);
nand_4 g12313(new_n12699, new_n12698, new_n681);
not_3  g12314(new_n12700, new_n12699);
nor_4  g12315(new_n12701, new_n12700, new_n3062);
nor_4  g12316(new_n12702, new_n12701, new_n3061);
nor_4  g12317(new_n12703, new_n12702, new_n3354);
nor_4  g12318(new_n12704, new_n12703, new_n3353);
nor_4  g12319(new_n12705, new_n12704, new_n3352);
nor_4  g12320(new_n12706, new_n12705, new_n3351);
nor_4  g12321(new_n12707, new_n12706, new_n3350);
nor_4  g12322(new_n12708, new_n12707, new_n3349);
nor_4  g12323(new_n12709, new_n12708, new_n3348);
nor_4  g12324(new_n12710, new_n12709, new_n720);
nor_4  g12325(new_n12711, new_n12710, new_n501);
nor_4  g12326(new_n12712, new_n12711, new_n728);
nor_4  g12327(new_n12713, new_n12712, new_n495);
nor_4  g12328(new_n12714, new_n12713, new_n736);
nor_4  g12329(new_n12715, new_n12714, new_n489);
nor_4  g12330(new_n12716, new_n12715, new_n744);
nor_4  g12331(new_n12717, new_n12716, new_n483);
nor_4  g12332(new_n12718, new_n12717, new_n752);
nor_4  g12333(new_n12719, new_n12718, new_n759);
nor_4  g12334(new_n12720, new_n12719, new_n766);
nor_4  g12335(new_n12721, new_n12720, new_n477);
nor_4  g12336(new_n12722, new_n12721, new_n774);
nor_4  g12337(new_n12723, new_n12722, new_n781);
nor_4  g12338(new_n12724, new_n12723, new_n788);
not_3  g12339(new_n12725, new_n12724);
nand_4 g12340(new_n12726, new_n12725, new_n470);
nand_4 g12341(new_n12727, new_n12726, new_n795);
nand_4 g12342(new_n12728, new_n12727, new_n803);
nand_4 g12343(new_n12729, new_n12728, new_n809);
nand_4 g12344(new_n12730, new_n12729, new_n465);
nand_4 g12345(new_n12731, new_n12730, new_n818);
nand_4 g12346(new_n12732, new_n12731, new_n460);
nand_4 g12347(new_n12733, new_n12732, new_n455);
nand_4 g12348(new_n12734, new_n12733, new_n449);
nand_4 g12349(new_n12735, new_n12734, new_n827);
nand_4 g12350(new_n12736, new_n12735, new_n833);
nand_4 g12351(new_n12737, new_n12736, new_n444);
nand_4 g12352(new_n12738, new_n12737, new_n439);
nand_4 g12353(new_n12739, new_n12738, new_n841);
nand_4 g12354(new_n12740, new_n12739, n14303);
nor_4  g12355(n14289, new_n12740, new_n431);
nand_4 g12356(new_n12742, new_n2166_1, new_n1409);
nand_4 g12357(new_n12743, new_n12742, new_n2165);
nand_4 g12358(new_n12744, new_n12743, new_n2162);
nand_4 g12359(new_n12745, new_n12744, new_n2158);
nand_4 g12360(new_n12746, new_n12745, new_n2155);
nand_4 g12361(new_n12747, new_n12746, new_n2151);
nand_4 g12362(new_n12748, new_n12747, new_n2147);
nand_4 g12363(new_n12749, new_n12748, new_n1810);
nand_4 g12364(new_n12750, new_n12749, new_n1806);
nand_4 g12365(new_n12751, new_n12750, new_n1802);
nand_4 g12366(new_n12752, new_n12751, new_n1798);
nand_4 g12367(new_n12753, new_n12752, new_n1820);
nand_4 g12368(new_n12754, new_n12753, new_n1794);
nand_4 g12369(new_n12755, new_n12754, new_n1825);
nand_4 g12370(new_n12756, new_n12755, new_n1789);
nand_4 g12371(new_n12757, new_n12756, new_n1785);
nand_4 g12372(new_n12758, new_n12757, new_n1780);
nand_4 g12373(new_n12759, new_n12758, new_n1777);
nand_4 g12374(new_n12760, new_n12759, new_n1774);
nand_4 g12375(new_n12761, new_n12760, new_n1834);
nand_4 g12376(new_n12762, new_n12761, new_n1769);
nand_4 g12377(new_n12763, new_n12762, new_n1766);
nand_4 g12378(new_n12764, new_n12763, new_n1762);
nand_4 g12379(new_n12765, new_n12764, new_n1758);
nand_4 g12380(new_n12766, new_n12765, new_n1754);
nand_4 g12381(new_n12767, new_n12766, new_n1751);
nand_4 g12382(new_n12768, new_n12767, new_n1748);
nand_4 g12383(new_n12769, new_n12768, new_n1746);
nand_4 g12384(new_n12770, new_n12769, new_n1742);
nand_4 g12385(new_n12771, new_n12770, new_n1738);
nand_4 g12386(new_n12772, new_n12771, new_n1736);
nand_4 g12387(new_n12773, new_n12772, new_n1732);
nand_4 g12388(new_n12774, new_n12773, new_n1729);
nand_4 g12389(new_n12775, new_n12774, new_n1726);
nand_4 g12390(new_n12776, new_n12775, new_n1724);
nand_4 g12391(new_n12777, new_n12776, new_n1721);
nand_4 g12392(new_n12778, new_n12777, new_n1718);
nand_4 g12393(new_n12779, new_n12778, new_n1715);
nand_4 g12394(new_n12780, new_n12779, new_n1711);
nand_4 g12395(new_n12781, new_n12780, new_n1708);
nand_4 g12396(new_n12782_1, new_n12781, new_n1705);
nand_4 g12397(new_n12783, new_n12782_1, new_n1703);
nand_4 g12398(new_n12784, new_n12783, new_n1860);
nand_4 g12399(new_n12785, new_n12784, new_n1864);
nand_4 g12400(new_n12786, new_n12785, new_n1699);
nand_4 g12401(new_n12787, new_n12786, new_n1697);
nand_4 g12402(new_n12788, new_n12787, new_n1871);
nand_4 g12403(new_n12789, new_n12788, new_n1694);
nand_4 g12404(new_n12790, new_n12789, new_n1690);
nand_4 g12405(new_n12791, new_n12790, new_n1878);
nand_4 g12406(new_n12792, new_n12791, new_n1882);
not_3  g12407(new_n12793, new_n12792);
nor_4  g12408(new_n12794, new_n12793, new_n1687);
nor_4  g12409(new_n12795, new_n12794, new_n1683);
nor_4  g12410(new_n12796, new_n12795, new_n1679);
nor_4  g12411(new_n12797, new_n12796, new_n1675);
nor_4  g12412(new_n12798, new_n12797, new_n1891);
nor_4  g12413(new_n12799, new_n12798, new_n1670);
nor_4  g12414(new_n12800, new_n12799, new_n1666);
nor_4  g12415(new_n12801, new_n12800, new_n1662);
nor_4  g12416(new_n12802, new_n12801, new_n1658);
nor_4  g12417(new_n12803, new_n12802, new_n1653);
nor_4  g12418(new_n12804, new_n12803, new_n1649);
nor_4  g12419(new_n12805, new_n12804, new_n1645);
nor_4  g12420(new_n12806, new_n12805, new_n1641);
nor_4  g12421(new_n12807, new_n12806, new_n1637_1);
nor_4  g12422(new_n12808, new_n12807, new_n1633);
nor_4  g12423(new_n12809, new_n12808, new_n1629);
nor_4  g12424(new_n12810, new_n12809, new_n1628);
nor_4  g12425(new_n12811, new_n12810, new_n1627);
nor_4  g12426(new_n12812, new_n12811, new_n1626);
nor_4  g12427(new_n12813, new_n12812, new_n4700);
nor_4  g12428(new_n12814, new_n12813, new_n4699);
nor_4  g12429(new_n12815, new_n12814, new_n3722);
nor_4  g12430(new_n12816, new_n12815, new_n3721);
nor_4  g12431(new_n12817, new_n12816, new_n3720);
nor_4  g12432(new_n12818, new_n12817, new_n3719);
nor_4  g12433(new_n12819, new_n12818, new_n3718);
nor_4  g12434(new_n12820, new_n12819, new_n3717);
not_3  g12435(new_n12821, new_n12820);
nand_4 g12436(new_n12822, new_n12821, new_n1338);
nand_4 g12437(new_n12823, new_n12822, new_n1395);
nand_4 g12438(new_n12824, new_n12823, new_n1335);
nand_4 g12439(new_n12825, new_n12824, new_n1332);
nand_4 g12440(new_n12826, new_n12825, new_n1328);
nand_4 g12441(new_n12827, new_n12826, new_n1403);
nand_4 g12442(new_n12828, new_n12827, n6480);
nor_4  g12443(n14307, new_n12828, new_n815);
nand_4 g12444(new_n12830, new_n1054, new_n537);
nand_4 g12445(new_n12831, new_n12830, new_n534);
nand_4 g12446(new_n12832, new_n12831, new_n529);
nand_4 g12447(new_n12833, new_n12832, new_n668);
nand_4 g12448(new_n12834, new_n12833, new_n674_1);
nand_4 g12449(new_n12835, new_n12834, new_n681);
nand_4 g12450(new_n12836, new_n12835, new_n523);
nand_4 g12451(new_n12837, new_n12836, new_n687);
nand_4 g12452(new_n12838, new_n12837, new_n693);
nand_4 g12453(new_n12839, new_n12838, new_n699);
nand_4 g12454(new_n12840, new_n12839, new_n517);
nand_4 g12455(new_n12841, new_n12840, new_n705);
nand_4 g12456(new_n12842, new_n12841, new_n511);
nand_4 g12457(new_n12843, new_n12842, new_n711);
nand_4 g12458(new_n12844, new_n12843, new_n506);
nand_4 g12459(new_n12845, new_n12844, new_n719);
nand_4 g12460(new_n12846, new_n12845, new_n500);
nand_4 g12461(new_n12847, new_n12846, new_n727);
nand_4 g12462(new_n12848, new_n12847, new_n494);
nand_4 g12463(new_n12849, new_n12848, new_n735);
nand_4 g12464(new_n12850, new_n12849, new_n488);
nand_4 g12465(new_n12851, new_n12850, new_n743);
nand_4 g12466(new_n12852, new_n12851, new_n482);
nand_4 g12467(new_n12853, new_n12852, new_n751);
nand_4 g12468(new_n12854, new_n12853, new_n758);
nand_4 g12469(new_n12855, new_n12854, new_n765);
nand_4 g12470(new_n12856, new_n12855, new_n476);
nand_4 g12471(new_n12857, new_n12856, new_n773);
nand_4 g12472(new_n12858, new_n12857, new_n780);
nand_4 g12473(new_n12859, new_n12858, new_n787);
nand_4 g12474(new_n12860, new_n12859, new_n470);
nand_4 g12475(new_n12861, new_n12860, new_n795);
nand_4 g12476(new_n12862, new_n12861, new_n803);
nand_4 g12477(new_n12863, new_n12862, new_n809);
nand_4 g12478(new_n12864, new_n12863, new_n465);
nand_4 g12479(new_n12865, new_n12864, new_n818);
nand_4 g12480(new_n12866, new_n12865, new_n460);
nand_4 g12481(new_n12867, new_n12866, new_n455);
nand_4 g12482(new_n12868, new_n12867, new_n449);
nand_4 g12483(new_n12869, new_n12868, new_n827);
nand_4 g12484(new_n12870, new_n12869, new_n833);
nand_4 g12485(new_n12871, new_n12870, new_n444);
nand_4 g12486(new_n12872, new_n12871, new_n439);
nand_4 g12487(new_n12873, new_n12872, new_n841);
nand_4 g12488(new_n12874, new_n12873, new_n434);
not_3  g12489(new_n12875, new_n12874);
nor_4  g12490(new_n12876, new_n12875, new_n2032);
nor_4  g12491(new_n12877, new_n12876, new_n2031);
nor_4  g12492(new_n12878, new_n12877, new_n2030);
nor_4  g12493(new_n12879, new_n12878, new_n2029);
nor_4  g12494(new_n12880, new_n12879, new_n2028);
nor_4  g12495(new_n12881, new_n12880, new_n2027_1);
nor_4  g12496(new_n12882, new_n12881, new_n2026);
nor_4  g12497(new_n12883, new_n12882, new_n2025);
nor_4  g12498(new_n12884, new_n12883, new_n2024);
nor_4  g12499(new_n12885_1, new_n12884, new_n2023);
nor_4  g12500(new_n12886, new_n12885_1, new_n2022);
nor_4  g12501(new_n12887, new_n12886, new_n2021);
nor_4  g12502(new_n12888, new_n12887, new_n2020);
nor_4  g12503(new_n12889, new_n12888, new_n2019);
nor_4  g12504(new_n12890, new_n12889, new_n1537);
nor_4  g12505(new_n12891, new_n12890, new_n1536);
nor_4  g12506(new_n12892, new_n12891, new_n1535);
nor_4  g12507(new_n12893, new_n12892, new_n1534);
nor_4  g12508(new_n12894, new_n12893, new_n1533);
nor_4  g12509(new_n12895, new_n12894, new_n1532);
nor_4  g12510(new_n12896, new_n12895, new_n1531);
nor_4  g12511(new_n12897, new_n12896, new_n1530);
nor_4  g12512(new_n12898, new_n12897, new_n1529);
nor_4  g12513(new_n12899, new_n12898, new_n1528);
not_3  g12514(new_n12900, new_n12899);
nand_4 g12515(new_n12901, new_n12900, new_n1111);
nand_4 g12516(new_n12902, new_n12901, new_n1106);
nand_4 g12517(new_n12903, new_n12902, new_n1178);
nand_4 g12518(new_n12904, new_n12903, new_n1183);
nand_4 g12519(new_n12905, new_n12904, new_n1102);
nand_4 g12520(new_n12906, new_n12905, new_n1099);
nand_4 g12521(new_n12907, new_n12906, new_n1191);
nand_4 g12522(new_n12908, new_n12907, new_n1095);
nand_4 g12523(new_n12909, new_n12908, new_n1091);
nand_4 g12524(new_n12910, new_n12909, new_n1088);
nand_4 g12525(new_n12911, new_n12910, new_n1084);
nand_4 g12526(new_n12912, new_n12911, new_n1079);
nand_4 g12527(new_n12913, new_n12912, new_n1074);
nand_4 g12528(new_n12914, new_n12913, new_n1070);
nand_4 g12529(new_n12915, new_n12914, new_n1064);
nand_4 g12530(new_n12916, new_n12915, n5725);
nor_4  g12531(n14330, new_n12916, new_n1058);
nand_4 g12532(new_n12918, new_n678, new_n523);
nand_4 g12533(new_n12919, new_n12918, new_n687);
nand_4 g12534(new_n12920, new_n12919, new_n693);
nand_4 g12535(new_n12921, new_n12920, new_n699);
nand_4 g12536(new_n12922, new_n12921, new_n517);
nand_4 g12537(new_n12923, new_n12922, new_n705);
nand_4 g12538(new_n12924, new_n12923, new_n511);
nand_4 g12539(new_n12925, new_n12924, new_n711);
nand_4 g12540(new_n12926, new_n12925, new_n506);
nand_4 g12541(new_n12927_1, new_n12926, new_n719);
nand_4 g12542(new_n12928, new_n12927_1, new_n500);
nand_4 g12543(new_n12929, new_n12928, new_n727);
nand_4 g12544(new_n12930, new_n12929, new_n494);
nand_4 g12545(new_n12931, new_n12930, new_n735);
nand_4 g12546(new_n12932, new_n12931, new_n488);
nand_4 g12547(new_n12933, new_n12932, new_n743);
nand_4 g12548(new_n12934, new_n12933, new_n482);
nand_4 g12549(new_n12935, new_n12934, new_n751);
nand_4 g12550(new_n12936, new_n12935, new_n758);
nand_4 g12551(new_n12937, new_n12936, new_n765);
nand_4 g12552(new_n12938, new_n12937, new_n476);
nand_4 g12553(new_n12939, new_n12938, new_n773);
nand_4 g12554(new_n12940, new_n12939, new_n780);
nand_4 g12555(new_n12941, new_n12940, new_n787);
nand_4 g12556(new_n12942, new_n12941, new_n470);
nand_4 g12557(new_n12943, new_n12942, new_n795);
nand_4 g12558(new_n12944, new_n12943, new_n803);
nand_4 g12559(new_n12945, new_n12944, new_n809);
nand_4 g12560(new_n12946, new_n12945, new_n465);
nand_4 g12561(new_n12947, new_n12946, new_n818);
nand_4 g12562(new_n12948, new_n12947, new_n460);
nand_4 g12563(new_n12949, new_n12948, new_n455);
nand_4 g12564(new_n12950, new_n12949, new_n449);
nand_4 g12565(new_n12951, new_n12950, new_n827);
nand_4 g12566(new_n12952, new_n12951, new_n833);
nand_4 g12567(new_n12953, new_n12952, new_n444);
nand_4 g12568(new_n12954, new_n12953, new_n439);
nand_4 g12569(new_n12955, new_n12954, new_n841);
nand_4 g12570(new_n12956, new_n12955, new_n434);
nand_4 g12571(new_n12957, new_n12956, new_n429);
nand_4 g12572(new_n12958, new_n12957, new_n424);
nand_4 g12573(new_n12959, new_n12958, new_n850);
nand_4 g12574(new_n12960, new_n12959, new_n856);
nand_4 g12575(new_n12961, new_n12960, new_n863);
nand_4 g12576(new_n12962, new_n12961, new_n419);
nand_4 g12577(new_n12963, new_n12962, new_n869);
nand_4 g12578(new_n12964, new_n12963, new_n875);
nand_4 g12579(new_n12965, new_n12964, new_n881);
nand_4 g12580(new_n12966, new_n12965, new_n413);
nand_4 g12581(new_n12967, new_n12966, new_n889);
nand_4 g12582(new_n12968, new_n12967, new_n896);
not_3  g12583(new_n12969, new_n12968);
nor_4  g12584(new_n12970, new_n12969, new_n2020);
nor_4  g12585(new_n12971, new_n12970, new_n2019);
nor_4  g12586(new_n12972, new_n12971, new_n1537);
nor_4  g12587(new_n12973, new_n12972, new_n1536);
nor_4  g12588(new_n12974, new_n12973, new_n1535);
nor_4  g12589(new_n12975, new_n12974, new_n1534);
nor_4  g12590(new_n12976_1, new_n12975, new_n1533);
nor_4  g12591(new_n12977, new_n12976_1, new_n1532);
nor_4  g12592(new_n12978, new_n12977, new_n1531);
nor_4  g12593(new_n12979, new_n12978, new_n1530);
nor_4  g12594(new_n12980, new_n12979, new_n1529);
nor_4  g12595(new_n12981, new_n12980, new_n1528);
nor_4  g12596(new_n12982, new_n12981, new_n1527);
nor_4  g12597(new_n12983, new_n12982, new_n1526);
nor_4  g12598(new_n12984, new_n12983, new_n1525);
nor_4  g12599(new_n12985, new_n12984, new_n1524);
nor_4  g12600(new_n12986, new_n12985, new_n1523);
nor_4  g12601(new_n12987, new_n12986, new_n1522);
nor_4  g12602(new_n12988, new_n12987, new_n1521);
nor_4  g12603(new_n12989_1, new_n12988, new_n1520);
nor_4  g12604(new_n12990, new_n12989_1, new_n1519);
nor_4  g12605(new_n12991, new_n12990, new_n1518);
nor_4  g12606(new_n12992, new_n12991, new_n1517);
nor_4  g12607(new_n12993, new_n12992, new_n1516);
nor_4  g12608(new_n12994, new_n12993, new_n1075);
nor_4  g12609(new_n12995, new_n12994, new_n1071);
nor_4  g12610(new_n12996, new_n12995, new_n1065);
not_3  g12611(new_n12997, new_n12996);
nand_4 g12612(new_n12998, new_n12997, new_n1061);
nand_4 g12613(new_n12999, new_n12998, new_n1055);
nand_4 g12614(new_n13000_1, new_n12999, new_n1050);
nand_4 g12615(new_n13001, new_n13000_1, new_n1045);
nand_4 g12616(new_n13002, new_n13001, new_n1041);
nand_4 g12617(new_n13003, new_n13002, new_n1036);
nand_4 g12618(new_n13004, new_n13003, n10765);
nor_4  g12619(n14399, new_n13004, new_n1028);
not_3  g12620(new_n13006, new_n644);
nand_4 g12621(new_n13007, new_n1699, new_n13006);
nand_4 g12622(new_n13008, new_n13007, new_n1697);
nand_4 g12623(new_n13009, new_n13008, new_n1871);
nand_4 g12624(new_n13010_1, new_n13009, new_n1694);
nand_4 g12625(new_n13011, new_n13010_1, new_n1690);
nand_4 g12626(new_n13012, new_n13011, new_n1878);
nand_4 g12627(new_n13013, new_n13012, new_n1882);
nand_4 g12628(new_n13014, new_n13013, new_n1686);
nand_4 g12629(new_n13015, new_n13014, new_n1682);
nand_4 g12630(new_n13016, new_n13015, new_n1678);
nand_4 g12631(new_n13017, new_n13016, new_n1674);
nand_4 g12632(new_n13018, new_n13017, new_n1890);
nand_4 g12633(new_n13019, new_n13018, new_n1669);
nand_4 g12634(new_n13020, new_n13019, new_n1665);
nand_4 g12635(new_n13021, new_n13020, new_n1661);
nand_4 g12636(new_n13022, new_n13021, new_n1657);
nand_4 g12637(new_n13023, new_n13022, new_n1652);
nand_4 g12638(new_n13024, new_n13023, new_n1648);
nand_4 g12639(new_n13025, new_n13024, new_n1644);
nand_4 g12640(new_n13026, new_n13025, new_n1640);
nand_4 g12641(new_n13027, new_n13026, new_n1636);
nand_4 g12642(new_n13028, new_n13027, new_n1632);
nand_4 g12643(new_n13029, new_n13028, new_n1378);
nand_4 g12644(new_n13030, new_n13029, new_n1372);
nand_4 g12645(new_n13031, new_n13030, new_n1367);
nand_4 g12646(new_n13032, new_n13031, new_n1363);
nand_4 g12647(new_n13033, new_n13032, new_n1360);
nand_4 g12648(new_n13034, new_n13033, new_n1357);
nand_4 g12649(new_n13035, new_n13034, new_n1354);
nand_4 g12650(new_n13036, new_n13035, new_n1352);
nand_4 g12651(new_n13037, new_n13036, new_n1350);
nand_4 g12652(new_n13038, new_n13037, new_n1347_1);
nand_4 g12653(new_n13039, new_n13038, new_n1344);
nand_4 g12654(new_n13040, new_n13039, new_n1341);
nand_4 g12655(new_n13041, new_n13040, new_n1338);
nand_4 g12656(new_n13042, new_n13041, new_n1395);
nand_4 g12657(new_n13043, new_n13042, new_n1335);
nand_4 g12658(new_n13044, new_n13043, new_n1332);
nand_4 g12659(new_n13045_1, new_n13044, new_n1328);
nand_4 g12660(new_n13046, new_n13045_1, new_n1403);
nand_4 g12661(new_n13047, new_n13046, new_n1325);
nand_4 g12662(new_n13048, new_n13047, new_n1410);
nand_4 g12663(new_n13049, new_n13048, new_n1413);
nand_4 g12664(new_n13050, new_n13049, new_n1322);
nand_4 g12665(new_n13051, new_n13050, new_n1317);
nand_4 g12666(new_n13052, new_n13051, new_n1315);
nand_4 g12667(new_n13053, new_n13052, new_n1419);
nand_4 g12668(new_n13054, new_n13053, new_n1310);
nand_4 g12669(new_n13055, new_n13054, new_n1305);
nand_4 g12670(new_n13056, new_n13055, new_n1427);
nand_4 g12671(new_n13057, new_n13056, new_n1431);
not_3  g12672(new_n13058, new_n13057);
nor_4  g12673(new_n13059, new_n13058, new_n2400);
nor_4  g12674(new_n13060, new_n13059, new_n2399);
nor_4  g12675(new_n13061, new_n13060, new_n2398);
nor_4  g12676(new_n13062, new_n13061, new_n2397);
nor_4  g12677(new_n13063, new_n13062, new_n2396);
nor_4  g12678(new_n13064, new_n13063, new_n2395);
nor_4  g12679(new_n13065, new_n13064, new_n1281);
nor_4  g12680(new_n13066, new_n13065, new_n1276);
nor_4  g12681(new_n13067, new_n13066, new_n1446);
nor_4  g12682(new_n13068, new_n13067, new_n1271);
nor_4  g12683(new_n13069, new_n13068, new_n1266);
nor_4  g12684(new_n13070, new_n13069, new_n1261);
nor_4  g12685(new_n13071, new_n13070, new_n1257);
nor_4  g12686(new_n13072, new_n13071, new_n1252);
nor_4  g12687(new_n13073, new_n13072, new_n1458);
nor_4  g12688(new_n13074, new_n13073, new_n1463);
nor_4  g12689(new_n13075, new_n13074, new_n1469);
nor_4  g12690(new_n13076, new_n13075, new_n1248);
nor_4  g12691(new_n13077, new_n13076, new_n1475);
nor_4  g12692(new_n13078, new_n13077, new_n1244);
nor_4  g12693(new_n13079, new_n13078, new_n1243);
nor_4  g12694(new_n13080, new_n13079, new_n1242);
nor_4  g12695(new_n13081, new_n13080, new_n1241);
nor_4  g12696(new_n13082, new_n13081, new_n1240);
nor_4  g12697(new_n13083, new_n13082, new_n1239);
nor_4  g12698(new_n13084, new_n13083, new_n3082);
nor_4  g12699(new_n13085, new_n13084, new_n3081);
not_3  g12700(new_n13086, new_n13085);
nand_4 g12701(new_n13087, new_n13086, new_n570);
nand_4 g12702(new_n13088, new_n13087, new_n625);
nand_4 g12703(new_n13089, new_n13088, new_n564);
nand_4 g12704(new_n13090, new_n13089, new_n632);
nand_4 g12705(new_n13091, new_n13090, new_n638);
nand_4 g12706(new_n13092, new_n13091, new_n559);
nand_4 g12707(new_n13093_1, new_n13092, n11776);
nor_4  g12708(n14463, new_n13093_1, new_n551);
endmodule


