// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Fri Jun 14 22:42:05 2024

module top_810026173_826291639_946996917_1246901 ( 
    n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213, n223,
    n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414, n424,
    n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649, n653,
    n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788, n801,
    n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764,
    n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156, n174,
    n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299, n317,
    n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457, n460,
    n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547, n549,
    n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648, n665,
    n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773, n790,
    n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888, n891,
    n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989, n991,
    n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103, n1113,
    n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183, n1191,
    n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255, n1260,
    n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347, n1348,
    n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426, n1440,
    n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502, n1507,
    n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633, n1635,
    n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690, n1721,
    n1727, n1729, n1731, n1737, n1746  );
  input  n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213,
    n223, n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414,
    n424, n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649,
    n653, n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788,
    n801, n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764;
  output n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156,
    n174, n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299,
    n317, n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457,
    n460, n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547,
    n549, n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648,
    n665, n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773,
    n790, n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888,
    n891, n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989,
    n991, n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103,
    n1113, n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183,
    n1191, n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255,
    n1260, n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347,
    n1348, n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426,
    n1440, n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502,
    n1507, n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633,
    n1635, n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690,
    n1721, n1727, n1729, n1731, n1737, n1746;
  wire new_n276_1, new_n277_1, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290_1, new_n291, new_n292_1, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299_1, new_n300, new_n301,
    new_n302, new_n303_1, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317_1, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329_1,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347_1, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353_1, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372_1, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378_1, new_n379_1, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387_1, new_n388, new_n389, new_n390,
    new_n391_1, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401_1, new_n402_1, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414_1, new_n415, new_n416_1,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423_1,
    new_n424_1, new_n425, new_n426_1, new_n427, new_n428, new_n429_1,
    new_n430, new_n431, new_n432_1, new_n433_1, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444_1, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452_1, new_n453, new_n454, new_n455, new_n456,
    new_n457_1, new_n458, new_n459, new_n460_1, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469_1,
    new_n470, new_n471, new_n472_1, new_n473, new_n474, new_n475,
    new_n476_1, new_n478, new_n479, new_n480, new_n481, new_n482_1,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488_1, new_n489,
    new_n490, new_n491, new_n492, new_n493_1, new_n494, new_n495, new_n496,
    new_n497, new_n498_1, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510_1,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517_1,
    new_n518, new_n519, new_n520, new_n521, new_n522_1, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532_1, new_n533, new_n534_1, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541_1, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547_1, new_n548, new_n549_1, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555_1, new_n556,
    new_n557_1, new_n558, new_n559_1, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n569_1, new_n571,
    new_n573_1, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585_1, new_n586, new_n587,
    new_n588_1, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n597, new_n598, new_n599_1, new_n600_1, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607_1, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627_1, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638_1, new_n639, new_n640, new_n641, new_n642, new_n643_1,
    new_n644, new_n645, new_n646_1, new_n647_1, new_n648_1, new_n649_1,
    new_n650, new_n651, new_n652, new_n653_1, new_n654, new_n655_1,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665_1, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675_1, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682_1,
    new_n683_1, new_n684_1, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693_1, new_n694,
    new_n695_1, new_n696, new_n697, new_n698, new_n699_1, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712_1, new_n713, new_n714,
    new_n715_1, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724_1, new_n725_1, new_n726, new_n727,
    new_n728, new_n729_1, new_n730, new_n731_1, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738_1, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747_1,
    new_n748_1, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759_1, new_n760,
    new_n761_1, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770_1, new_n771, new_n772, new_n773_1,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788_1,
    new_n789, new_n790_1, new_n791, new_n792_1, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801_1,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813_1, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823_1, new_n824_1, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836_1, new_n837, new_n838, new_n839_1, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846_1, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858_1, new_n859, new_n860, new_n861, new_n862_1,
    new_n863, new_n864, new_n865_1, new_n866, new_n867_1, new_n868,
    new_n869, new_n870_1, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882_1,
    new_n883_1, new_n884, new_n885, new_n886, new_n887, new_n888_1,
    new_n889, new_n890, new_n891_1, new_n892_1, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902_1, new_n903, new_n904, new_n905_1, new_n906_1, new_n908,
    new_n909, new_n910, new_n911, new_n912_1, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927_1, new_n928, new_n929,
    new_n930, new_n931_1, new_n932, new_n933, new_n934, new_n935_1,
    new_n937, new_n938, new_n940, new_n941, new_n942_1, new_n943, new_n945,
    new_n947, new_n950, new_n951, new_n952_1, new_n953_1, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961_1,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968_1,
    new_n969, new_n970, new_n971, new_n972, new_n975, new_n976, new_n977,
    new_n978, new_n979_1, new_n980_1, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989_1, new_n990,
    new_n991_1, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000_1, new_n1001, new_n1002, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012_1,
    new_n1013, new_n1014, new_n1015_1, new_n1016_1, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025_1, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030_1,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062_1, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067_1, new_n1068_1, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1098, new_n1101, new_n1102, new_n1103_1, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113_1, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119_1, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135_1, new_n1136,
    new_n1137, new_n1138_1, new_n1139, new_n1140_1, new_n1141, new_n1142_1,
    new_n1143, new_n1144, new_n1145_1, new_n1146, new_n1147, new_n1148,
    new_n1149_1, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161_1, new_n1162_1, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172_1,
    new_n1173, new_n1174, new_n1175_1, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183_1, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191_1,
    new_n1192, new_n1193, new_n1194_1, new_n1195, new_n1196, new_n1199_1,
    new_n1201_1, new_n1202_1, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222_1, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234_1, new_n1235_1, new_n1236, new_n1237_1,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249_1,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255_1,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260_1, new_n1261,
    new_n1262, new_n1263_1, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277_1, new_n1278_1, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283_1, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296_1, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305_1, new_n1306, new_n1307, new_n1308, new_n1312,
    new_n1313, new_n1314, new_n1315_1, new_n1316, new_n1317, new_n1320,
    new_n1322, new_n1323, new_n1326, new_n1327, new_n1329, new_n1331,
    new_n1332_1, new_n1333, new_n1334, new_n1336, new_n1338_1, new_n1339,
    new_n1340_1, new_n1341_1, new_n1342, new_n1343, new_n1344, new_n1346,
    new_n1347_1, new_n1348_1, new_n1349_1, new_n1350, new_n1351_1,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1360, new_n1363_1, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369_1, new_n1370, new_n1371, new_n1373,
    new_n1375, new_n1378, new_n1379, new_n1380, new_n1381_1, new_n1382,
    new_n1384, new_n1385_1, new_n1389, new_n1391, new_n1392, new_n1393_1,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399_1,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407_1, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422_1, new_n1424,
    new_n1425_1, new_n1426_1, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435_1, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440_1, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453_1, new_n1454,
    new_n1455, new_n1456, new_n1457_1, new_n1458, new_n1459, new_n1460_1,
    new_n1461_1, new_n1462, new_n1463_1, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1470_1, new_n1471, new_n1472, new_n1473,
    new_n1474, new_n1475, new_n1476, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481_1, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1487, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1494, new_n1495_1, new_n1496, new_n1497, new_n1498_1, new_n1499,
    new_n1500, new_n1501_1, new_n1502_1, new_n1503, new_n1504, new_n1505,
    new_n1506, new_n1507_1, new_n1508, new_n1509, new_n1510, new_n1511,
    new_n1512, new_n1513, new_n1514, new_n1515, new_n1516, new_n1517,
    new_n1518, new_n1519, new_n1520, new_n1521, new_n1522, new_n1523,
    new_n1524, new_n1525_1, new_n1526, new_n1527_1, new_n1528, new_n1529,
    new_n1530_1, new_n1531, new_n1532, new_n1533, new_n1534, new_n1535_1,
    new_n1536, new_n1537_1, new_n1538, new_n1539, new_n1540, new_n1541,
    new_n1542, new_n1543, new_n1544_1, new_n1545, new_n1546, new_n1547,
    new_n1548, new_n1549, new_n1550, new_n1551, new_n1552, new_n1553,
    new_n1554, new_n1555, new_n1556_1, new_n1557, new_n1558, new_n1559,
    new_n1560, new_n1561, new_n1562, new_n1563, new_n1564, new_n1565,
    new_n1566, new_n1567, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1572, new_n1573, new_n1574, new_n1575, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580, new_n1581, new_n1582, new_n1583,
    new_n1584, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595_1,
    new_n1596, new_n1597_1, new_n1598, new_n1599, new_n1600_1, new_n1601_1,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613_1,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622_1, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1629_1, new_n1630, new_n1631,
    new_n1633_1, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642_1, new_n1643_1, new_n1644, new_n1645, new_n1650,
    new_n1653, new_n1655, new_n1657_1, new_n1658, new_n1659, new_n1660_1,
    new_n1661, new_n1663, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675_1, new_n1676, new_n1677_1,
    new_n1678_1, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683_1,
    new_n1684, new_n1685, new_n1686_1, new_n1687, new_n1688_1, new_n1689,
    new_n1690_1, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1703, new_n1704,
    new_n1706, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1719, new_n1721_1, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1727_1, new_n1729_1, new_n1731_1, new_n1734,
    new_n1737_1, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743_1,
    new_n1744, new_n1745, new_n1746_1, new_n1748, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757_1,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763_1,
    new_n1764_1, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1784, new_n1785,
    new_n1786, new_n1788, new_n1791, new_n1793, new_n1794, new_n1796,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1805, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1819, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1830, new_n1831, new_n1832, new_n1834, new_n1835,
    new_n1838, new_n1839, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1851,
    new_n1854, new_n1856, new_n1857, new_n1863, new_n1865, new_n1866,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1873, new_n1874,
    new_n1875, new_n1878, new_n1880, new_n1882, new_n1884, new_n1885,
    new_n1887, new_n1888, new_n1890, new_n1892, new_n1896, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1909, new_n1911, new_n1914,
    new_n1917, new_n1923, new_n1924, new_n1927, new_n1928, new_n1929,
    new_n1933, new_n1942;
nor_4  g0000(new_n276_1, n1643, n36);
xor_3  g0001(new_n277_1, n1643, n36);
not_3  g0002(new_n278, new_n277_1);
nor_4  g0003(new_n279, n788, n555);
not_3  g0004(new_n280, new_n279);
xnor_3 g0005(new_n281, n788, n555);
not_3  g0006(new_n282, new_n281);
nor_4  g0007(new_n283, n747, n353);
not_3  g0008(new_n284, new_n283);
nand_4 g0009(new_n285, n747, n353);
not_3  g0010(new_n286, new_n285);
nor_4  g0011(new_n287, new_n286, new_n283);
nor_4  g0012(new_n288, n952, n329);
not_3  g0013(new_n289, new_n288);
nand_4 g0014(new_n290_1, n1145, n931);
xnor_3 g0015(new_n291, n952, n329);
not_3  g0016(new_n292_1, new_n291);
nand_4 g0017(new_n293, new_n292_1, new_n290_1);
nand_4 g0018(new_n294, new_n293, new_n289);
nand_4 g0019(new_n295, new_n294, new_n287);
nand_4 g0020(new_n296, new_n295, new_n284);
nand_4 g0021(new_n297, new_n296, new_n282);
nand_4 g0022(new_n298, new_n297, new_n280);
not_3  g0023(new_n299_1, new_n298);
nor_4  g0024(new_n300, new_n299_1, new_n278);
nor_4  g0025(new_n301, new_n300, new_n276_1);
nand_4 g0026(new_n302, new_n301, n1501);
xnor_3 g0027(new_n303_1, new_n302, n433);
nand_4 g0028(new_n304, n1000, n870);
not_3  g0029(new_n305, n1000);
nand_4 g0030(new_n306, new_n305, n66);
nand_4 g0031(new_n307, new_n306, new_n304);
nand_4 g0032(new_n308, n1000, n585);
nand_4 g0033(new_n309, new_n305, n968);
nand_4 g0034(new_n310, new_n309, new_n308);
nor_4  g0035(new_n311, new_n310, new_n307);
nand_4 g0036(new_n312, n1000, n155);
not_3  g0037(new_n313, new_n312);
not_3  g0038(new_n314, n1435);
nor_4  g0039(new_n315, new_n314, n1000);
nor_4  g0040(new_n316, new_n315, new_n313);
nand_4 g0041(new_n317_1, new_n316, new_n311);
nor_4  g0042(new_n318, n1000, n682);
nor_4  g0043(new_n319, n1678, new_n305);
nor_4  g0044(new_n320, new_n319, new_n318);
not_3  g0045(new_n321, new_n320);
nor_4  g0046(new_n322, new_n321, new_n317_1);
xor_3  g0047(new_n323, n1597, n682);
nor_4  g0048(new_n324, new_n323, n1000);
xnor_3 g0049(new_n325, n1678, n607);
nor_4  g0050(new_n326, new_n325, new_n305);
nor_4  g0051(new_n327, new_n326, new_n324);
xnor_3 g0052(new_n328, new_n327, new_n322);
not_3  g0053(new_n329_1, new_n317_1);
nor_4  g0054(new_n330, new_n320, new_n329_1);
nor_4  g0055(new_n331, new_n330, new_n322);
nor_4  g0056(new_n332, new_n316, new_n311);
nor_4  g0057(new_n333, new_n332, new_n329_1);
not_3  g0058(new_n334, new_n333);
not_3  g0059(new_n335, new_n308);
not_3  g0060(new_n336, n968);
nor_4  g0061(new_n337, n1000, new_n336);
nor_4  g0062(new_n338, new_n337, new_n335);
xnor_3 g0063(new_n339, new_n338, new_n307);
not_3  g0064(new_n340, new_n339);
nand_4 g0065(new_n341, new_n340, n693);
not_3  g0066(new_n342, n693);
nand_4 g0067(new_n343, new_n339, new_n342);
nand_4 g0068(new_n344, new_n338, n1763);
not_3  g0069(new_n345, n1763);
nand_4 g0070(new_n346, new_n310, new_n345);
not_3  g0071(new_n347_1, n1530);
nand_4 g0072(new_n348, n1461, n1000);
not_3  g0073(new_n349, new_n348);
not_3  g0074(new_n350, n347);
nor_4  g0075(new_n351, n1000, new_n350);
nor_4  g0076(new_n352, new_n351, new_n349);
nor_4  g0077(new_n353_1, new_n352, new_n347_1);
nand_4 g0078(new_n354, new_n353_1, new_n346);
nand_4 g0079(new_n355, new_n354, new_n344);
nand_4 g0080(new_n356, new_n355, new_n343);
nand_4 g0081(new_n357, new_n356, new_n341);
nand_4 g0082(new_n358, new_n357, new_n334);
nor_4  g0083(new_n359, new_n358, new_n331);
nand_4 g0084(new_n360, new_n359, new_n328);
nand_4 g0085(new_n361, new_n327, new_n322);
not_3  g0086(new_n362, n682);
nor_4  g0087(new_n363, n1597, n46);
nand_4 g0088(new_n364, new_n363, new_n362);
not_3  g0089(new_n365, new_n364);
not_3  g0090(new_n366, n46);
nor_4  g0091(new_n367, n1597, n682);
nor_4  g0092(new_n368, new_n367, new_n366);
nor_4  g0093(new_n369, new_n368, new_n365);
nor_4  g0094(new_n370, new_n369, n1000);
not_3  g0095(new_n371, n1678);
nand_4 g0096(new_n372_1, n607, n26);
nor_4  g0097(new_n373, new_n372_1, new_n371);
not_3  g0098(new_n374, n26);
nand_4 g0099(new_n375, n1678, n607);
nand_4 g0100(new_n376, new_n375, new_n374);
nand_4 g0101(new_n377, new_n376, n1000);
nor_4  g0102(new_n378_1, new_n377, new_n373);
nor_4  g0103(new_n379_1, new_n378_1, new_n370);
xnor_3 g0104(new_n380, new_n379_1, new_n361);
xnor_3 g0105(new_n381, new_n380, new_n360);
xnor_3 g0106(new_n382, new_n381, new_n303_1);
not_3  g0107(new_n383, new_n382);
xnor_3 g0108(new_n384, new_n359, new_n328);
xnor_3 g0109(new_n385, new_n301, n1501);
nand_4 g0110(new_n386, new_n385, new_n384);
not_3  g0111(new_n387_1, n1501);
xnor_3 g0112(new_n388, new_n301, new_n387_1);
xnor_3 g0113(new_n389, new_n388, new_n384);
xnor_3 g0114(new_n390, new_n358, new_n331);
xnor_3 g0115(new_n391_1, new_n298, new_n277_1);
not_3  g0116(new_n392, new_n391_1);
nor_4  g0117(new_n393, new_n392, new_n390);
xnor_3 g0118(new_n394, new_n357, new_n333);
not_3  g0119(new_n395, new_n394);
xnor_3 g0120(new_n396, new_n296, new_n282);
not_3  g0121(new_n397, new_n396);
nand_4 g0122(new_n398, new_n397, new_n395);
xnor_3 g0123(new_n399, new_n397, new_n394);
xnor_3 g0124(new_n400, new_n294, new_n287);
not_3  g0125(new_n401_1, new_n400);
not_3  g0126(new_n402_1, new_n290_1);
nor_4  g0127(new_n403, n1145, n931);
nor_4  g0128(new_n404, new_n403, new_n402_1);
nand_4 g0129(new_n405, new_n305, n347);
nand_4 g0130(new_n406, new_n405, new_n348);
xnor_3 g0131(new_n407, new_n406, new_n347_1);
nand_4 g0132(new_n408, new_n407, new_n404);
not_3  g0133(new_n409, new_n408);
xnor_3 g0134(new_n410, new_n291, new_n402_1);
nor_4  g0135(new_n411, new_n410, new_n409);
not_3  g0136(new_n412, new_n411);
nor_4  g0137(new_n413, new_n408, new_n291);
nand_4 g0138(new_n414_1, new_n346, new_n344);
xnor_3 g0139(new_n415, new_n414_1, new_n353_1);
nor_4  g0140(new_n416_1, new_n415, new_n413);
not_3  g0141(new_n417, new_n416_1);
nand_4 g0142(new_n418, new_n417, new_n412);
nor_4  g0143(new_n419, new_n418, new_n401_1);
nor_4  g0144(new_n420, new_n416_1, new_n411);
nor_4  g0145(new_n421, new_n420, new_n400);
not_3  g0146(new_n422, new_n355);
nand_4 g0147(new_n423_1, new_n343, new_n341);
xnor_3 g0148(new_n424_1, new_n423_1, new_n422);
nor_4  g0149(new_n425, new_n424_1, new_n421);
nor_4  g0150(new_n426_1, new_n425, new_n419);
nand_4 g0151(new_n427, new_n426_1, new_n399);
nand_4 g0152(new_n428, new_n427, new_n398);
xnor_3 g0153(new_n429_1, new_n392, new_n390);
nor_4  g0154(new_n430, new_n429_1, new_n428);
nor_4  g0155(new_n431, new_n430, new_n393);
nand_4 g0156(new_n432_1, new_n431, new_n389);
nand_4 g0157(new_n433_1, new_n432_1, new_n386);
xor_3  g0158(n19, new_n433_1, new_n383);
not_3  g0159(new_n435, n69);
not_3  g0160(new_n436, n402);
nor_4  g0161(new_n437, n1381, new_n436);
nor_4  g0162(new_n438, new_n437, n870);
not_3  g0163(new_n439, n1381);
nand_4 g0164(new_n440, new_n439, n402);
nor_4  g0165(new_n441, new_n440, n66);
nor_4  g0166(new_n442, new_n441, new_n438);
xnor_3 g0167(new_n443, new_n442, new_n435);
not_3  g0168(new_n444_1, new_n443);
nor_4  g0169(new_n445, new_n437, n585);
nor_4  g0170(new_n446, new_n440, n968);
nor_4  g0171(new_n447, new_n446, new_n445);
nand_4 g0172(new_n448, new_n447, n953);
not_3  g0173(new_n449, n303);
not_3  g0174(new_n450, n1461);
nand_4 g0175(new_n451, new_n440, new_n450);
nand_4 g0176(new_n452_1, new_n437, new_n350);
nand_4 g0177(new_n453, new_n452_1, new_n451);
nor_4  g0178(new_n454, new_n453, new_n449);
not_3  g0179(new_n455, n953);
xnor_3 g0180(new_n456, new_n447, new_n455);
nand_4 g0181(new_n457_1, new_n456, new_n454);
nand_4 g0182(new_n458, new_n457_1, new_n448);
xnor_3 g0183(new_n459, new_n458, new_n444_1);
nor_4  g0184(new_n460_1, new_n459, new_n400);
xnor_3 g0185(new_n461, new_n458, new_n443);
nor_4  g0186(new_n462, new_n461, new_n401_1);
nor_4  g0187(new_n463, new_n462, new_n460_1);
not_3  g0188(new_n464, new_n463);
not_3  g0189(new_n465, new_n404);
xnor_3 g0190(new_n466, new_n453, n303);
not_3  g0191(new_n467, new_n466);
nor_4  g0192(new_n468, new_n467, new_n465);
nor_4  g0193(new_n469_1, new_n468, new_n410);
not_3  g0194(new_n470, new_n469_1);
xnor_3 g0195(new_n471, new_n456, new_n454);
not_3  g0196(new_n472_1, new_n468);
nor_4  g0197(new_n473, new_n472_1, new_n291);
nor_4  g0198(new_n474, new_n473, new_n469_1);
nand_4 g0199(new_n475, new_n474, new_n471);
nand_4 g0200(new_n476_1, new_n475, new_n470);
xor_3  g0201(n33, new_n476_1, new_n464);
not_3  g0202(new_n478, n247);
nor_4  g0203(new_n479, n607, n26);
nand_4 g0204(new_n480, new_n479, new_n478);
xor_3  g0205(new_n481, new_n480, n1642);
nor_4  g0206(new_n482_1, new_n481, new_n439);
not_3  g0207(new_n483, n1527);
nand_4 g0208(new_n484, new_n483, new_n366);
nor_4  g0209(new_n485, new_n484, n379);
not_3  g0210(new_n486, n379);
nor_4  g0211(new_n487, n1527, n46);
nor_4  g0212(new_n488_1, new_n487, new_n486);
nor_4  g0213(new_n489, new_n488_1, new_n436);
not_3  g0214(new_n490, new_n489);
nor_4  g0215(new_n491, new_n490, new_n485);
not_3  g0216(new_n492, n1642);
nor_4  g0217(new_n493_1, new_n492, n1381);
nor_4  g0218(new_n494, new_n493_1, new_n437);
nor_4  g0219(new_n495, new_n494, new_n491);
nor_4  g0220(new_n496, new_n495, new_n482_1);
not_3  g0221(new_n497, new_n496);
xor_3  g0222(new_n498_1, new_n479, new_n478);
nor_4  g0223(new_n499, new_n498_1, new_n439);
nand_4 g0224(new_n500, n1527, n46);
nand_4 g0225(new_n501, new_n500, n402);
nor_4  g0226(new_n502, new_n501, new_n487);
nor_4  g0227(new_n503, n1381, new_n478);
nor_4  g0228(new_n504, new_n503, new_n437);
nor_4  g0229(new_n505, new_n504, new_n502);
nor_4  g0230(new_n506, new_n505, new_n499);
nor_4  g0231(new_n507, new_n437, n1678);
nor_4  g0232(new_n508, new_n440, n682);
nor_4  g0233(new_n509, new_n508, new_n507);
nor_4  g0234(new_n510_1, new_n509, n1643);
not_3  g0235(new_n511, new_n510_1);
xor_3  g0236(new_n512, new_n509, n1643);
not_3  g0237(new_n513, n555);
nor_4  g0238(new_n514, new_n437, n155);
nor_4  g0239(new_n515, new_n440, n1435);
nor_4  g0240(new_n516, new_n515, new_n514);
not_3  g0241(new_n517_1, new_n516);
nor_4  g0242(new_n518, new_n517_1, new_n513);
nor_4  g0243(new_n519, new_n442, n353);
not_3  g0244(new_n520, new_n519);
xor_3  g0245(new_n521, new_n442, n353);
nor_4  g0246(new_n522_1, new_n447, n952);
not_3  g0247(new_n523, new_n522_1);
not_3  g0248(new_n524, n1145);
nor_4  g0249(new_n525, new_n453, new_n524);
not_3  g0250(new_n526, new_n525);
xor_3  g0251(new_n527, new_n447, n952);
nand_4 g0252(new_n528, new_n527, new_n526);
nand_4 g0253(new_n529, new_n528, new_n523);
nand_4 g0254(new_n530, new_n529, new_n521);
nand_4 g0255(new_n531, new_n530, new_n520);
xor_3  g0256(new_n532_1, new_n516, n555);
not_3  g0257(new_n533, new_n532_1);
nor_4  g0258(new_n534_1, new_n533, new_n531);
nor_4  g0259(new_n535, new_n534_1, new_n518);
nand_4 g0260(new_n536, new_n535, new_n512);
nand_4 g0261(new_n537, new_n536, new_n511);
nand_4 g0262(new_n538, n1381, n607);
not_3  g0263(new_n539, new_n538);
nor_4  g0264(new_n540, n1597, new_n436);
nor_4  g0265(new_n541_1, n607, n402);
nor_4  g0266(new_n542, new_n541_1, new_n540);
nor_4  g0267(new_n543, new_n542, n1381);
nor_4  g0268(new_n544, new_n543, new_n539);
not_3  g0269(new_n545, new_n544);
nor_4  g0270(new_n546, new_n545, new_n537);
nand_4 g0271(new_n547_1, n402, n46);
not_3  g0272(new_n548, new_n547_1);
nor_4  g0273(new_n549_1, n402, n26);
nor_4  g0274(new_n550, new_n549_1, new_n548);
nor_4  g0275(new_n551, new_n550, n1381);
not_3  g0276(new_n552, new_n372_1);
nor_4  g0277(new_n553, new_n479, new_n552);
not_3  g0278(new_n554, new_n553);
nor_4  g0279(new_n555_1, new_n554, new_n439);
nor_4  g0280(new_n556, new_n555_1, new_n551);
nand_4 g0281(new_n557_1, new_n556, new_n546);
nor_4  g0282(new_n558, new_n557_1, new_n506);
nor_4  g0283(new_n559_1, new_n558, new_n497);
nand_4 g0284(new_n560, new_n558, new_n497);
not_3  g0285(new_n561, new_n560);
nor_4  g0286(n1731, new_n561, new_n559_1);
not_3  g0287(new_n563, new_n506);
not_3  g0288(new_n564, new_n557_1);
nor_4  g0289(new_n565, new_n564, new_n563);
nor_4  g0290(n1138, new_n565, new_n558);
not_3  g0291(new_n567, new_n556);
not_3  g0292(new_n568, new_n537);
nor_4  g0293(new_n569_1, new_n544, new_n568);
nor_4  g0294(n1727, new_n569_1, new_n546);
not_3  g0295(new_n571, new_n527);
xor_3  g0296(n1457, new_n571, new_n526);
nand_4 g0297(new_n573_1, new_n453, new_n524);
and_4  g0298(n1183, new_n573_1, new_n526);
nor_4  g0299(new_n575, n1183, n1457);
not_3  g0300(new_n576, new_n530);
nor_4  g0301(new_n577, new_n529, new_n521);
nor_4  g0302(new_n578, new_n577, new_n576);
nand_4 g0303(new_n579, new_n578, new_n575);
not_3  g0304(new_n580, new_n531);
nor_4  g0305(new_n581, new_n532_1, new_n580);
nor_4  g0306(n1721, new_n581, new_n534_1);
nor_4  g0307(new_n583, n1721, new_n579);
not_3  g0308(new_n584, new_n536);
nor_4  g0309(new_n585_1, new_n535, new_n512);
nor_4  g0310(new_n586, new_n585_1, new_n584);
nor_4  g0311(new_n587, new_n586, new_n583);
nand_4 g0312(new_n588_1, new_n587, n1727);
nor_4  g0313(new_n589, new_n588_1, new_n567);
nand_4 g0314(new_n590, new_n589, n1138);
not_3  g0315(new_n591, new_n590);
nor_4  g0316(new_n592, new_n591, n1731);
nor_4  g0317(new_n593, new_n590, new_n496);
nor_4  g0318(n44, new_n593, new_n592);
not_3  g0319(new_n595, new_n407);
xor_3  g0320(n55, new_n595, new_n465);
not_3  g0321(new_n597, n1332);
nor_4  g0322(new_n598, n1707, n1643);
not_3  g0323(new_n599_1, new_n598);
xor_3  g0324(new_n600_1, n1707, n1643);
nor_4  g0325(new_n601, n1140, n555);
not_3  g0326(new_n602, new_n601);
xor_3  g0327(new_n603, n1140, n555);
nor_4  g0328(new_n604, n1351, n353);
not_3  g0329(new_n605, new_n604);
xor_3  g0330(new_n606, n1351, n353);
nor_4  g0331(new_n607_1, n952, n729);
nand_4 g0332(new_n608, n1145, n684);
not_3  g0333(new_n609, new_n608);
nand_4 g0334(new_n610, n952, n729);
not_3  g0335(new_n611, new_n610);
nor_4  g0336(new_n612, new_n611, new_n607_1);
not_3  g0337(new_n613, new_n612);
nor_4  g0338(new_n614, new_n613, new_n609);
nor_4  g0339(new_n615, new_n614, new_n607_1);
not_3  g0340(new_n616, new_n615);
nand_4 g0341(new_n617, new_n616, new_n606);
nand_4 g0342(new_n618, new_n617, new_n605);
nand_4 g0343(new_n619, new_n618, new_n603);
nand_4 g0344(new_n620, new_n619, new_n602);
nand_4 g0345(new_n621, new_n620, new_n600_1);
nand_4 g0346(new_n622, new_n621, new_n599_1);
nor_4  g0347(new_n623, new_n622, new_n597);
nand_4 g0348(new_n624, new_n623, n391);
xnor_3 g0349(new_n625, new_n624, n1544);
nand_4 g0350(new_n626, n607, n266);
not_3  g0351(new_n627_1, new_n626);
nor_4  g0352(new_n628, n1597, n266);
nor_4  g0353(new_n629, new_n628, new_n627_1);
not_3  g0354(new_n630, new_n629);
nand_4 g0355(new_n631, n266, n155);
not_3  g0356(new_n632, n266);
nand_4 g0357(new_n633, n1435, new_n632);
nand_4 g0358(new_n634, new_n633, new_n631);
nand_4 g0359(new_n635, n870, n266);
nand_4 g0360(new_n636, new_n632, n66);
nand_4 g0361(new_n637, new_n636, new_n635);
nor_4  g0362(new_n638_1, new_n637, new_n634);
nand_4 g0363(new_n639, n1678, n266);
nand_4 g0364(new_n640, n682, new_n632);
nand_4 g0365(new_n641, new_n640, new_n639);
not_3  g0366(new_n642, new_n641);
nand_4 g0367(new_n643_1, new_n642, new_n638_1);
nor_4  g0368(new_n644, new_n643_1, new_n630);
nor_4  g0369(new_n645, new_n632, n26);
not_3  g0370(new_n646_1, new_n645);
xor_3  g0371(new_n647_1, n1597, n46);
nand_4 g0372(new_n648_1, new_n647_1, new_n632);
nand_4 g0373(new_n649_1, new_n648_1, new_n646_1);
xnor_3 g0374(new_n650, new_n649_1, new_n644);
xnor_3 g0375(new_n651, new_n643_1, new_n629);
xor_3  g0376(new_n652, new_n641, new_n638_1);
xnor_3 g0377(new_n653_1, new_n637, new_n634);
nand_4 g0378(new_n654, new_n653_1, n223);
not_3  g0379(new_n655_1, new_n654);
nor_4  g0380(new_n656, new_n653_1, n223);
nor_4  g0381(new_n657, new_n656, new_n655_1);
not_3  g0382(new_n658, n444);
nor_4  g0383(new_n659, new_n637, new_n658);
not_3  g0384(new_n660, new_n659);
nand_4 g0385(new_n661, n585, n266);
nand_4 g0386(new_n662, n968, new_n632);
nand_4 g0387(new_n663, new_n662, new_n661);
nor_4  g0388(new_n664, new_n663, n472);
not_3  g0389(new_n665_1, n801);
nand_4 g0390(new_n666, n1461, n266);
not_3  g0391(new_n667, new_n666);
nor_4  g0392(new_n668, new_n350, n266);
nor_4  g0393(new_n669, new_n668, new_n667);
nor_4  g0394(new_n670, new_n669, new_n665_1);
not_3  g0395(new_n671, n472);
not_3  g0396(new_n672, new_n661);
nor_4  g0397(new_n673, new_n336, n266);
nor_4  g0398(new_n674, new_n673, new_n672);
xnor_3 g0399(new_n675_1, new_n674, new_n671);
nor_4  g0400(new_n676, new_n675_1, new_n670);
nor_4  g0401(new_n677, new_n676, new_n664);
xnor_3 g0402(new_n678, new_n637, new_n658);
not_3  g0403(new_n679, new_n678);
nand_4 g0404(new_n680, new_n679, new_n677);
nand_4 g0405(new_n681, new_n680, new_n660);
nand_4 g0406(new_n682_1, new_n681, new_n657);
nand_4 g0407(new_n683_1, new_n682_1, new_n654);
nand_4 g0408(new_n684_1, new_n683_1, new_n652);
nor_4  g0409(new_n685, new_n684_1, new_n651);
nand_4 g0410(new_n686, new_n685, new_n650);
not_3  g0411(new_n687, new_n644);
xor_3  g0412(new_n688, n1597, new_n366);
nor_4  g0413(new_n689, new_n688, n266);
nor_4  g0414(new_n690, new_n689, new_n645);
nor_4  g0415(new_n691, new_n690, new_n687);
not_3  g0416(new_n692, n1597);
nand_4 g0417(new_n693_1, new_n487, new_n692);
not_3  g0418(new_n694, new_n693_1);
nor_4  g0419(new_n695_1, new_n363, new_n483);
nor_4  g0420(new_n696, new_n695_1, new_n694);
nand_4 g0421(new_n697, new_n696, new_n632);
not_3  g0422(new_n698, new_n697);
nor_4  g0423(new_n699_1, new_n632, n247);
nor_4  g0424(new_n700, new_n699_1, new_n698);
not_3  g0425(new_n701, new_n700);
nor_4  g0426(new_n702, new_n701, new_n691);
nand_4 g0427(new_n703, new_n649_1, new_n644);
nor_4  g0428(new_n704, new_n700, new_n703);
nor_4  g0429(new_n705, new_n704, new_n702);
xnor_3 g0430(new_n706, new_n705, new_n686);
xnor_3 g0431(new_n707, new_n706, new_n625);
not_3  g0432(new_n708, new_n707);
not_3  g0433(new_n709, n391);
xnor_3 g0434(new_n710, new_n623, new_n709);
xnor_3 g0435(new_n711, new_n649_1, new_n687);
xnor_3 g0436(new_n712_1, new_n685, new_n711);
nor_4  g0437(new_n713, new_n712_1, new_n710);
not_3  g0438(new_n714, new_n713);
xnor_3 g0439(new_n715_1, new_n684_1, new_n651);
not_3  g0440(new_n716, new_n715_1);
xnor_3 g0441(new_n717, new_n622, n1332);
nor_4  g0442(new_n718, new_n717, new_n716);
not_3  g0443(new_n719, new_n718);
xnor_3 g0444(new_n720, new_n717, new_n715_1);
xnor_3 g0445(new_n721, new_n683_1, new_n652);
xnor_3 g0446(new_n722, new_n620, new_n600_1);
not_3  g0447(new_n723, new_n722);
nand_4 g0448(new_n724_1, new_n723, new_n721);
xnor_3 g0449(new_n725_1, new_n722, new_n721);
xnor_3 g0450(new_n726, new_n653_1, n223);
not_3  g0451(new_n727, new_n664);
nand_4 g0452(new_n728, n347, new_n632);
nand_4 g0453(new_n729_1, new_n728, new_n666);
nand_4 g0454(new_n730, new_n729_1, n801);
xnor_3 g0455(new_n731_1, new_n674, n472);
nand_4 g0456(new_n732, new_n731_1, new_n730);
nand_4 g0457(new_n733, new_n732, new_n727);
nor_4  g0458(new_n734, new_n678, new_n733);
nor_4  g0459(new_n735, new_n734, new_n659);
xnor_3 g0460(new_n736, new_n735, new_n726);
xnor_3 g0461(new_n737, new_n618, new_n603);
not_3  g0462(new_n738_1, new_n737);
nand_4 g0463(new_n739, new_n738_1, new_n736);
xnor_3 g0464(new_n740, new_n737, new_n736);
xnor_3 g0465(new_n741, new_n679, new_n677);
xnor_3 g0466(new_n742, new_n615, new_n606);
nand_4 g0467(new_n743, new_n742, new_n741);
nor_4  g0468(new_n744, new_n612, new_n608);
not_3  g0469(new_n745, new_n614);
nor_4  g0470(new_n746, n1145, n684);
nor_4  g0471(new_n747_1, new_n746, new_n609);
nor_4  g0472(new_n748_1, new_n729_1, n801);
nor_4  g0473(new_n749, new_n748_1, new_n670);
nand_4 g0474(new_n750, new_n749, new_n747_1);
nand_4 g0475(new_n751, new_n750, new_n745);
nor_4  g0476(new_n752, new_n751, new_n744);
not_3  g0477(new_n753, new_n752);
xnor_3 g0478(new_n754, new_n731_1, new_n670);
nor_4  g0479(new_n755, new_n750, new_n613);
nor_4  g0480(new_n756, new_n755, new_n752);
nand_4 g0481(new_n757, new_n756, new_n754);
nand_4 g0482(new_n758, new_n757, new_n753);
not_3  g0483(new_n759_1, new_n743);
nor_4  g0484(new_n760, new_n742, new_n741);
nor_4  g0485(new_n761_1, new_n760, new_n759_1);
nand_4 g0486(new_n762, new_n761_1, new_n758);
nand_4 g0487(new_n763, new_n762, new_n743);
nand_4 g0488(new_n764, new_n763, new_n740);
nand_4 g0489(new_n765, new_n764, new_n739);
nand_4 g0490(new_n766, new_n765, new_n725_1);
nand_4 g0491(new_n767, new_n766, new_n724_1);
nand_4 g0492(new_n768, new_n767, new_n720);
nand_4 g0493(new_n769, new_n768, new_n719);
xnor_3 g0494(new_n770_1, new_n685, new_n650);
xnor_3 g0495(new_n771, new_n770_1, new_n710);
nand_4 g0496(new_n772, new_n771, new_n769);
nand_4 g0497(new_n773_1, new_n772, new_n714);
xor_3  g0498(n56, new_n773_1, new_n708);
nor_4  g0499(new_n775, new_n705, new_n686);
nor_4  g0500(new_n776, n1642, new_n632);
not_3  g0501(new_n777, new_n776);
xor_3  g0502(new_n778, new_n693_1, n379);
nand_4 g0503(new_n779, new_n778, new_n632);
nand_4 g0504(new_n780, new_n779, new_n777);
xnor_3 g0505(new_n781, new_n780, new_n704);
nand_4 g0506(new_n782, new_n781, new_n775);
nand_4 g0507(new_n783, new_n780, new_n704);
nor_4  g0508(new_n784, new_n632, n171);
not_3  g0509(new_n785, n1263);
nor_4  g0510(new_n786, new_n693_1, n379);
nor_4  g0511(new_n787, new_n786, new_n785);
nand_4 g0512(new_n788_1, new_n485, new_n785);
nor_4  g0513(new_n789, new_n788_1, n1597);
nor_4  g0514(new_n790_1, new_n789, new_n787);
nand_4 g0515(new_n791, new_n790_1, new_n632);
not_3  g0516(new_n792_1, new_n791);
nor_4  g0517(new_n793, new_n792_1, new_n784);
nor_4  g0518(new_n794, new_n793, new_n783);
nand_4 g0519(new_n795, new_n701, new_n691);
xor_3  g0520(new_n796, new_n693_1, new_n486);
nor_4  g0521(new_n797, new_n796, n266);
nor_4  g0522(new_n798, new_n797, new_n776);
nor_4  g0523(new_n799, new_n798, new_n795);
not_3  g0524(new_n800, new_n793);
nor_4  g0525(new_n801_1, new_n800, new_n799);
nor_4  g0526(new_n802, new_n801_1, new_n794);
nor_4  g0527(new_n803, new_n802, new_n782);
not_3  g0528(new_n804, new_n794);
nor_4  g0529(new_n805, n557, new_n632);
not_3  g0530(new_n806, n1422);
not_3  g0531(new_n807, new_n788_1);
nand_4 g0532(new_n808, new_n807, new_n806);
nor_4  g0533(new_n809, new_n808, n1597);
not_3  g0534(new_n810, new_n789);
nand_4 g0535(new_n811, new_n810, n1422);
not_3  g0536(new_n812, new_n811);
nor_4  g0537(new_n813_1, new_n812, new_n809);
nand_4 g0538(new_n814, new_n813_1, new_n632);
not_3  g0539(new_n815, new_n814);
nor_4  g0540(new_n816, new_n815, new_n805);
xor_3  g0541(new_n817, new_n816, new_n804);
not_3  g0542(new_n818, new_n817);
xor_3  g0543(new_n819, new_n818, new_n803);
not_3  g0544(new_n820, n1544);
nor_4  g0545(new_n821, new_n624, new_n820);
nand_4 g0546(new_n822, new_n821, n649);
not_3  g0547(new_n823_1, new_n822);
xnor_3 g0548(new_n824_1, new_n802, new_n782);
not_3  g0549(new_n825, new_n824_1);
nor_4  g0550(new_n826, new_n825, new_n823_1);
not_3  g0551(new_n827, new_n826);
xor_3  g0552(new_n828, new_n825, new_n823_1);
nor_4  g0553(new_n829, new_n821, n649);
nor_4  g0554(new_n830, new_n829, new_n823_1);
not_3  g0555(new_n831, new_n781);
xnor_3 g0556(new_n832, new_n831, new_n775);
nor_4  g0557(new_n833, new_n832, new_n830);
not_3  g0558(new_n834, new_n833);
xnor_3 g0559(new_n835, new_n832, new_n830);
not_3  g0560(new_n836_1, new_n835);
xnor_3 g0561(new_n837, new_n700, new_n703);
xnor_3 g0562(new_n838, new_n837, new_n686);
nor_4  g0563(new_n839_1, new_n838, new_n625);
not_3  g0564(new_n840, new_n839_1);
nand_4 g0565(new_n841, new_n773_1, new_n707);
nand_4 g0566(new_n842, new_n841, new_n840);
nand_4 g0567(new_n843, new_n842, new_n836_1);
nand_4 g0568(new_n844, new_n843, new_n834);
nand_4 g0569(new_n845, new_n844, new_n828);
nand_4 g0570(new_n846_1, new_n845, new_n827);
not_3  g0571(new_n847, new_n846_1);
nor_4  g0572(new_n848, new_n847, new_n819);
not_3  g0573(new_n849, new_n819);
nor_4  g0574(new_n850, new_n846_1, new_n849);
nor_4  g0575(n67, new_n850, new_n848);
not_3  g0576(new_n852, new_n390);
xor_3  g0577(new_n853, n1643, n469);
nor_4  g0578(new_n854, n927, n555);
not_3  g0579(new_n855, new_n854);
xor_3  g0580(new_n856, n927, n555);
nor_4  g0581(new_n857, n655, n353);
xnor_3 g0582(new_n858_1, n655, n353);
nor_4  g0583(new_n859, n952, n653);
nand_4 g0584(new_n860, n1764, n1145);
not_3  g0585(new_n861, new_n860);
nand_4 g0586(new_n862_1, n952, n653);
not_3  g0587(new_n863, new_n862_1);
nor_4  g0588(new_n864, new_n863, new_n859);
not_3  g0589(new_n865_1, new_n864);
nor_4  g0590(new_n866, new_n865_1, new_n861);
nor_4  g0591(new_n867_1, new_n866, new_n859);
nor_4  g0592(new_n868, new_n867_1, new_n858_1);
nor_4  g0593(new_n869, new_n868, new_n857);
not_3  g0594(new_n870_1, new_n869);
nand_4 g0595(new_n871, new_n870_1, new_n856);
nand_4 g0596(new_n872, new_n871, new_n855);
xnor_3 g0597(new_n873, new_n872, new_n853);
nand_4 g0598(new_n874, new_n873, new_n852);
not_3  g0599(new_n875, new_n874);
nor_4  g0600(new_n876, new_n873, new_n852);
nor_4  g0601(new_n877, new_n876, new_n875);
xnor_3 g0602(new_n878, new_n870_1, new_n856);
nor_4  g0603(new_n879, new_n878, new_n394);
not_3  g0604(new_n880, new_n878);
nor_4  g0605(new_n881, new_n880, new_n395);
nor_4  g0606(new_n882_1, new_n881, new_n879);
not_3  g0607(new_n883_1, new_n882_1);
nor_4  g0608(new_n884, new_n864, new_n860);
not_3  g0609(new_n885, new_n866);
nor_4  g0610(new_n886, n1764, n1145);
nor_4  g0611(new_n887, new_n886, new_n861);
nand_4 g0612(new_n888_1, new_n887, new_n407);
nand_4 g0613(new_n889, new_n888_1, new_n885);
nor_4  g0614(new_n890, new_n889, new_n884);
not_3  g0615(new_n891_1, new_n890);
not_3  g0616(new_n892_1, new_n415);
nor_4  g0617(new_n893, new_n888_1, new_n865_1);
nor_4  g0618(new_n894, new_n893, new_n890);
nand_4 g0619(new_n895, new_n894, new_n892_1);
nand_4 g0620(new_n896, new_n895, new_n891_1);
xnor_3 g0621(new_n897, new_n867_1, new_n858_1);
not_3  g0622(new_n898, new_n897);
nor_4  g0623(new_n899, new_n898, new_n896);
not_3  g0624(new_n900, new_n899);
not_3  g0625(new_n901, new_n424_1);
xnor_3 g0626(new_n902_1, new_n897, new_n896);
nand_4 g0627(new_n903, new_n902_1, new_n901);
nand_4 g0628(new_n904, new_n903, new_n900);
nor_4  g0629(new_n905_1, new_n904, new_n883_1);
nor_4  g0630(new_n906_1, new_n905_1, new_n879);
xor_3  g0631(n74, new_n906_1, new_n877);
not_3  g0632(new_n908, n171);
nor_4  g0633(new_n909, new_n480, n1642);
xor_3  g0634(new_n910, new_n909, new_n908);
nor_4  g0635(new_n911, new_n910, new_n439);
xor_3  g0636(new_n912_1, new_n485, new_n785);
not_3  g0637(new_n913, new_n912_1);
nor_4  g0638(new_n914, new_n913, new_n436);
nor_4  g0639(new_n915, n402, n171);
nor_4  g0640(new_n916, new_n915, n1381);
not_3  g0641(new_n917, new_n916);
nor_4  g0642(new_n918, new_n917, new_n914);
nor_4  g0643(new_n919, new_n918, new_n911);
nor_4  g0644(new_n920, new_n919, new_n560);
xor_3  g0645(new_n921, new_n788_1, n1422);
not_3  g0646(new_n922, new_n921);
nor_4  g0647(new_n923, new_n922, new_n436);
nor_4  g0648(new_n924, n557, n402);
nor_4  g0649(new_n925, new_n924, n1381);
not_3  g0650(new_n926, new_n925);
nor_4  g0651(new_n927_1, new_n926, new_n923);
nand_4 g0652(new_n928, new_n909, new_n908);
xor_3  g0653(new_n929, new_n928, n557);
nor_4  g0654(new_n930, new_n929, new_n439);
nor_4  g0655(new_n931_1, new_n930, new_n927_1);
not_3  g0656(new_n932, new_n931_1);
nor_4  g0657(new_n933, new_n932, new_n920);
nand_4 g0658(new_n934, new_n932, new_n920);
not_3  g0659(new_n935_1, new_n934);
nor_4  g0660(n156, new_n935_1, new_n933);
not_3  g0661(new_n937, new_n919);
nor_4  g0662(new_n938, new_n937, new_n561);
nor_4  g0663(n1149, new_n938, new_n920);
nand_4 g0664(new_n940, n1149, new_n593);
not_3  g0665(new_n941, new_n940);
nor_4  g0666(new_n942_1, new_n941, n156);
nor_4  g0667(new_n943, new_n940, new_n931_1);
nor_4  g0668(n106, new_n943, new_n942_1);
not_3  g0669(new_n945, new_n588_1);
xor_3  g0670(n1385, new_n556, new_n546);
nor_4  g0671(new_n947, n1385, new_n945);
nor_4  g0672(n126, new_n947, new_n589);
xnor_3 g0673(n135, new_n765, new_n725_1);
nor_4  g0674(new_n950, new_n641, n1643);
xor_3  g0675(new_n951, new_n641, n1643);
not_3  g0676(new_n952_1, new_n634);
nand_4 g0677(new_n953_1, new_n952_1, new_n513);
not_3  g0678(new_n954, n353);
not_3  g0679(new_n955, new_n637);
nand_4 g0680(new_n956, new_n955, new_n954);
xor_3  g0681(new_n957, new_n955, new_n954);
not_3  g0682(new_n958, n952);
nand_4 g0683(new_n959, new_n674, new_n958);
nand_4 g0684(new_n960, new_n729_1, n1145);
xor_3  g0685(new_n961_1, new_n674, new_n958);
nand_4 g0686(new_n962, new_n961_1, new_n960);
nand_4 g0687(new_n963, new_n962, new_n959);
nand_4 g0688(new_n964, new_n963, new_n957);
nand_4 g0689(new_n965, new_n964, new_n956);
xor_3  g0690(new_n966, new_n634, n555);
nand_4 g0691(new_n967, new_n966, new_n965);
nand_4 g0692(new_n968_1, new_n967, new_n953_1);
nand_4 g0693(new_n969, new_n968_1, new_n951);
not_3  g0694(new_n970, new_n969);
nor_4  g0695(new_n971, new_n970, new_n950);
nand_4 g0696(new_n972, new_n971, new_n630);
xor_3  g0697(n145, new_n972, new_n649_1);
xor_3  g0698(n174, new_n404, n347);
xnor_3 g0699(new_n975, new_n388, new_n692);
not_3  g0700(new_n976, new_n975);
nand_4 g0701(new_n977, new_n391_1, n682);
xnor_3 g0702(new_n978, new_n391_1, new_n362);
nand_4 g0703(new_n979_1, new_n396, n1435);
xnor_3 g0704(new_n980_1, new_n396, new_n314);
nand_4 g0705(new_n981, new_n400, n66);
not_3  g0706(new_n982, new_n981);
nor_4  g0707(new_n983, new_n400, n66);
nor_4  g0708(new_n984, new_n983, new_n982);
nor_4  g0709(new_n985, new_n410, n968);
nor_4  g0710(new_n986, new_n465, new_n350);
xnor_3 g0711(new_n987, new_n410, n968);
nor_4  g0712(new_n988, new_n987, new_n986);
nor_4  g0713(new_n989_1, new_n988, new_n985);
nand_4 g0714(new_n990, new_n989_1, new_n984);
nand_4 g0715(new_n991_1, new_n990, new_n981);
nand_4 g0716(new_n992, new_n991_1, new_n980_1);
nand_4 g0717(new_n993, new_n992, new_n979_1);
nand_4 g0718(new_n994, new_n993, new_n978);
nand_4 g0719(new_n995, new_n994, new_n977);
xor_3  g0720(new_n996, new_n995, new_n976);
xor_3  g0721(new_n997, new_n993, new_n978);
not_3  g0722(new_n998, new_n997);
xor_3  g0723(n1426, new_n989_1, new_n984);
xor_3  g0724(new_n1000_1, new_n991_1, new_n980_1);
nor_4  g0725(new_n1001, new_n1000_1, n1426);
nand_4 g0726(new_n1002, new_n1001, new_n998);
xor_3  g0727(n181, new_n1002, new_n996);
nor_4  g0728(new_n1004, new_n421, new_n419);
xor_3  g0729(n208, new_n1004, new_n901);
nor_4  g0730(new_n1006, new_n637, n213);
not_3  g0731(new_n1007, new_n1006);
not_3  g0732(new_n1008, n213);
nor_4  g0733(new_n1009, new_n955, new_n1008);
nor_4  g0734(new_n1010, new_n1009, new_n1006);
nor_4  g0735(new_n1011, new_n663, n1743);
not_3  g0736(new_n1012_1, new_n1011);
not_3  g0737(new_n1013, n600);
nor_4  g0738(new_n1014, new_n669, new_n1013);
not_3  g0739(new_n1015_1, new_n1014);
not_3  g0740(new_n1016_1, n1743);
nor_4  g0741(new_n1017, new_n674, new_n1016_1);
nor_4  g0742(new_n1018, new_n1017, new_n1011);
nand_4 g0743(new_n1019, new_n1018, new_n1015_1);
nand_4 g0744(new_n1020, new_n1019, new_n1012_1);
nand_4 g0745(new_n1021, new_n1020, new_n1010);
nand_4 g0746(new_n1022, new_n1021, new_n1007);
nor_4  g0747(new_n1023, new_n1022, new_n952_1);
nand_4 g0748(new_n1024, new_n1023, new_n641);
xnor_3 g0749(new_n1025_1, new_n1024, new_n630);
nor_4  g0750(new_n1026, n1643, n424);
not_3  g0751(new_n1027, new_n1026);
xor_3  g0752(new_n1028, n1643, n424);
nor_4  g0753(new_n1029, n1363, n555);
not_3  g0754(new_n1030_1, new_n1029);
xor_3  g0755(new_n1031, n1363, n555);
nor_4  g0756(new_n1032, n498, n353);
not_3  g0757(new_n1033, new_n1032);
nand_4 g0758(new_n1034, n498, n353);
not_3  g0759(new_n1035, new_n1034);
nor_4  g0760(new_n1036, new_n1035, new_n1032);
nor_4  g0761(new_n1037, n952, n414);
not_3  g0762(new_n1038, new_n1037);
nand_4 g0763(new_n1039, n1145, n183);
nand_4 g0764(new_n1040, n952, n414);
not_3  g0765(new_n1041, new_n1040);
nor_4  g0766(new_n1042, new_n1041, new_n1037);
nand_4 g0767(new_n1043, new_n1042, new_n1039);
nand_4 g0768(new_n1044, new_n1043, new_n1038);
nand_4 g0769(new_n1045, new_n1044, new_n1036);
nand_4 g0770(new_n1046, new_n1045, new_n1033);
nand_4 g0771(new_n1047, new_n1046, new_n1031);
nand_4 g0772(new_n1048, new_n1047, new_n1030_1);
nand_4 g0773(new_n1049, new_n1048, new_n1028);
nand_4 g0774(new_n1050, new_n1049, new_n1027);
xnor_3 g0775(new_n1051, new_n1050, n17);
xnor_3 g0776(new_n1052, new_n1051, new_n1025_1);
not_3  g0777(new_n1053, new_n1052);
xnor_3 g0778(new_n1054, new_n1023, new_n642);
xnor_3 g0779(new_n1055, new_n1048, new_n1028);
nor_4  g0780(new_n1056, new_n1055, new_n1054);
xnor_3 g0781(new_n1057, new_n1022, new_n952_1);
xnor_3 g0782(new_n1058, new_n1046, new_n1031);
not_3  g0783(new_n1059, new_n1058);
nand_4 g0784(new_n1060, new_n1059, new_n1057);
xnor_3 g0785(new_n1061, new_n1058, new_n1057);
xnor_3 g0786(new_n1062_1, new_n1020, new_n1010);
not_3  g0787(new_n1063, new_n1062_1);
not_3  g0788(new_n1064, new_n1045);
nor_4  g0789(new_n1065, new_n1044, new_n1036);
nor_4  g0790(new_n1066, new_n1065, new_n1064);
nand_4 g0791(new_n1067_1, new_n1066, new_n1063);
nor_4  g0792(new_n1068_1, new_n1042, new_n1039);
not_3  g0793(new_n1069, new_n1039);
nor_4  g0794(new_n1070, n1145, n183);
nor_4  g0795(new_n1071, new_n1070, new_n1069);
nor_4  g0796(new_n1072, new_n729_1, n600);
nor_4  g0797(new_n1073, new_n1072, new_n1014);
nand_4 g0798(new_n1074, new_n1073, new_n1071);
nand_4 g0799(new_n1075, new_n1074, new_n1043);
nor_4  g0800(new_n1076, new_n1075, new_n1068_1);
not_3  g0801(new_n1077, new_n1076);
xnor_3 g0802(new_n1078, new_n1018, new_n1014);
not_3  g0803(new_n1079, new_n1042);
nor_4  g0804(new_n1080, new_n1074, new_n1079);
nor_4  g0805(new_n1081, new_n1080, new_n1076);
nand_4 g0806(new_n1082, new_n1081, new_n1078);
nand_4 g0807(new_n1083, new_n1082, new_n1077);
xnor_3 g0808(new_n1084, new_n1066, new_n1062_1);
nand_4 g0809(new_n1085, new_n1084, new_n1083);
nand_4 g0810(new_n1086, new_n1085, new_n1067_1);
nand_4 g0811(new_n1087, new_n1086, new_n1061);
nand_4 g0812(new_n1088, new_n1087, new_n1060);
not_3  g0813(new_n1089, new_n1054);
not_3  g0814(new_n1090, new_n1028);
xnor_3 g0815(new_n1091, new_n1048, new_n1090);
nor_4  g0816(new_n1092, new_n1091, new_n1089);
nor_4  g0817(new_n1093, new_n1092, new_n1056);
nand_4 g0818(new_n1094, new_n1093, new_n1088);
not_3  g0819(new_n1095, new_n1094);
nor_4  g0820(new_n1096, new_n1095, new_n1056);
xor_3  g0821(n216, new_n1096, new_n1053);
not_3  g0822(new_n1098, new_n1084);
xor_3  g0823(n218, new_n1098, new_n1083);
xnor_3 g0824(n231, new_n844, new_n828);
not_3  g0825(new_n1101, n1747);
not_3  g0826(new_n1102, n738);
not_3  g0827(new_n1103_1, n17);
nor_4  g0828(new_n1104, new_n1050, new_n1103_1);
nand_4 g0829(new_n1105, new_n1104, n961);
nor_4  g0830(new_n1106, new_n1105, new_n1102);
not_3  g0831(new_n1107, new_n1106);
xor_3  g0832(new_n1108, new_n1107, new_n1101);
nor_4  g0833(new_n1109, new_n1024, new_n629);
nand_4 g0834(new_n1110, new_n1109, new_n690);
nor_4  g0835(new_n1111, new_n1110, new_n701);
xnor_3 g0836(new_n1112, new_n1111, new_n780);
xnor_3 g0837(new_n1113_1, new_n1112, new_n1108);
xnor_3 g0838(new_n1114, new_n1105, n738);
xnor_3 g0839(new_n1115, new_n1110, new_n700);
nor_4  g0840(new_n1116, new_n1115, new_n1114);
xnor_3 g0841(new_n1117, new_n1115, new_n1114);
not_3  g0842(new_n1118, n961);
xnor_3 g0843(new_n1119_1, new_n1104, new_n1118);
xnor_3 g0844(new_n1120, new_n1109, new_n649_1);
nor_4  g0845(new_n1121, new_n1120, new_n1119_1);
xnor_3 g0846(new_n1122, new_n1120, new_n1119_1);
nor_4  g0847(new_n1123, new_n1051, new_n1025_1);
nor_4  g0848(new_n1124, new_n1096, new_n1052);
nor_4  g0849(new_n1125, new_n1124, new_n1123);
nor_4  g0850(new_n1126, new_n1125, new_n1122);
nor_4  g0851(new_n1127, new_n1126, new_n1121);
nor_4  g0852(new_n1128, new_n1127, new_n1117);
nor_4  g0853(new_n1129, new_n1128, new_n1116);
xnor_3 g0854(n238, new_n1129, new_n1113_1);
not_3  g0855(new_n1131, n675);
not_3  g0856(new_n1132, n433);
nor_4  g0857(new_n1133, new_n302, new_n1132);
nand_4 g0858(new_n1134, new_n1133, n1537);
nor_4  g0859(new_n1135_1, new_n1134, new_n1131);
xor_3  g0860(new_n1136, new_n1135_1, n1263);
not_3  g0861(new_n1137, new_n1134);
nor_4  g0862(new_n1138_1, new_n1137, n675);
nor_4  g0863(new_n1139, new_n1138_1, new_n1135_1);
not_3  g0864(new_n1140_1, new_n1139);
nor_4  g0865(new_n1141, new_n1140_1, new_n486);
xnor_3 g0866(new_n1142_1, new_n1139, n379);
xnor_3 g0867(new_n1143, new_n1133, n1537);
nor_4  g0868(new_n1144, new_n1143, new_n483);
xnor_3 g0869(new_n1145_1, new_n1143, n1527);
nand_4 g0870(new_n1146, new_n303_1, n46);
nand_4 g0871(new_n1147, new_n388, n1597);
nand_4 g0872(new_n1148, new_n995, new_n975);
nand_4 g0873(new_n1149_1, new_n1148, new_n1147);
xnor_3 g0874(new_n1150, new_n303_1, new_n366);
nand_4 g0875(new_n1151, new_n1150, new_n1149_1);
nand_4 g0876(new_n1152, new_n1151, new_n1146);
nand_4 g0877(new_n1153, new_n1152, new_n1145_1);
not_3  g0878(new_n1154, new_n1153);
nor_4  g0879(new_n1155, new_n1154, new_n1144);
nor_4  g0880(new_n1156, new_n1155, new_n1142_1);
nor_4  g0881(new_n1157, new_n1156, new_n1141);
nand_4 g0882(new_n1158, new_n1157, new_n1136);
not_3  g0883(new_n1159, new_n1158);
nor_4  g0884(new_n1160, new_n1157, new_n1136);
nor_4  g0885(new_n1161_1, new_n1160, new_n1159);
not_3  g0886(new_n1162_1, new_n1161_1);
not_3  g0887(new_n1163, new_n1142_1);
xor_3  g0888(new_n1164, new_n1155, new_n1163);
nor_4  g0889(new_n1165, new_n1152, new_n1145_1);
nor_4  g0890(new_n1166, new_n1165, new_n1154);
not_3  g0891(new_n1167, new_n1166);
nor_4  g0892(new_n1168, new_n1000_1, new_n997);
nand_4 g0893(new_n1169, new_n1168, new_n996);
xnor_3 g0894(new_n1170, new_n1150, new_n1149_1);
not_3  g0895(new_n1171, new_n1170);
nor_4  g0896(new_n1172_1, new_n1171, new_n1169);
nand_4 g0897(new_n1173, new_n1172_1, new_n1167);
nor_4  g0898(new_n1174, new_n1173, n1426);
nand_4 g0899(new_n1175_1, new_n1174, new_n1164);
xnor_3 g0900(n270, new_n1175_1, new_n1162_1);
xnor_3 g0901(new_n1177, new_n721, new_n391_1);
not_3  g0902(new_n1178, new_n1177);
nor_4  g0903(new_n1179, new_n736, new_n397);
nor_4  g0904(new_n1180, new_n741, new_n401_1);
not_3  g0905(new_n1181, new_n410);
nand_4 g0906(new_n1182, new_n749, new_n404);
nand_4 g0907(new_n1183_1, new_n1182, new_n1181);
xnor_3 g0908(new_n1184, new_n669, new_n665_1);
nor_4  g0909(new_n1185, new_n1184, new_n465);
nor_4  g0910(new_n1186, new_n1185, new_n410);
nor_4  g0911(new_n1187, new_n1182, new_n291);
nor_4  g0912(new_n1188, new_n1187, new_n1186);
nand_4 g0913(new_n1189, new_n1188, new_n754);
nand_4 g0914(new_n1190, new_n1189, new_n1183_1);
xnor_3 g0915(new_n1191_1, new_n741, new_n401_1);
nor_4  g0916(new_n1192, new_n1191_1, new_n1190);
nor_4  g0917(new_n1193, new_n1192, new_n1180);
xnor_3 g0918(new_n1194_1, new_n736, new_n397);
nor_4  g0919(new_n1195, new_n1194_1, new_n1193);
nor_4  g0920(new_n1196, new_n1195, new_n1179);
xor_3  g0921(n276, new_n1196, new_n1178);
xor_3  g0922(n290, new_n887, new_n407);
not_3  g0923(new_n1199_1, new_n987);
xor_3  g0924(n292, new_n1199_1, new_n986);
not_3  g0925(new_n1201_1, new_n809);
nor_4  g0926(new_n1202_1, new_n1201_1, n266);
not_3  g0927(new_n1203, new_n1202_1);
nand_4 g0928(new_n1204, new_n1111, new_n798);
nor_4  g0929(new_n1205, new_n1204, new_n800);
nand_4 g0930(new_n1206, new_n1205, new_n816);
xor_3  g0931(new_n1207, new_n1205, new_n816);
nor_4  g0932(new_n1208, new_n1107, new_n1101);
xor_3  g0933(new_n1209, new_n1204, new_n800);
nor_4  g0934(new_n1210, new_n1209, new_n1208);
xnor_3 g0935(new_n1211, new_n1209, new_n1208);
nor_4  g0936(new_n1212, new_n1112, new_n1108);
nor_4  g0937(new_n1213, new_n1129, new_n1113_1);
nor_4  g0938(new_n1214, new_n1213, new_n1212);
nor_4  g0939(new_n1215, new_n1214, new_n1211);
nor_4  g0940(new_n1216, new_n1215, new_n1210);
nand_4 g0941(new_n1217, new_n1216, new_n1207);
nand_4 g0942(new_n1218, new_n1217, new_n1206);
nor_4  g0943(n299, new_n1218, new_n1203);
nand_4 g0944(new_n1220, new_n516, n1341);
xnor_3 g0945(new_n1221, new_n517_1, n1341);
nand_4 g0946(new_n1222_1, new_n442, n69);
nand_4 g0947(new_n1223, new_n458, new_n443);
nand_4 g0948(new_n1224, new_n1223, new_n1222_1);
nand_4 g0949(new_n1225, new_n1224, new_n1221);
nand_4 g0950(new_n1226, new_n1225, new_n1220);
nand_4 g0951(new_n1227, new_n1226, new_n509);
not_3  g0952(new_n1228, new_n1227);
nand_4 g0953(new_n1229, new_n1228, new_n544);
xnor_3 g0954(new_n1230, new_n1229, new_n556);
not_3  g0955(new_n1231, new_n1230);
not_3  g0956(new_n1232, n862);
nor_4  g0957(new_n1233, n1643, n761);
not_3  g0958(new_n1234_1, new_n1233);
xor_3  g0959(new_n1235_1, n1643, n761);
nor_4  g0960(new_n1236, n1172, n555);
not_3  g0961(new_n1237_1, new_n1236);
xor_3  g0962(new_n1238, n1172, n555);
nor_4  g0963(new_n1239, n695, n353);
nand_4 g0964(new_n1240, n695, n353);
not_3  g0965(new_n1241, new_n1240);
nor_4  g0966(new_n1242, new_n1241, new_n1239);
not_3  g0967(new_n1243, new_n1242);
nor_4  g0968(new_n1244, n1296, n952);
nand_4 g0969(new_n1245, n1145, n1062);
not_3  g0970(new_n1246, new_n1245);
not_3  g0971(new_n1247, new_n1244);
nand_4 g0972(new_n1248, n1296, n952);
nand_4 g0973(new_n1249_1, new_n1248, new_n1247);
nor_4  g0974(new_n1250, new_n1249_1, new_n1246);
nor_4  g0975(new_n1251, new_n1250, new_n1244);
nor_4  g0976(new_n1252, new_n1251, new_n1243);
nor_4  g0977(new_n1253, new_n1252, new_n1239);
not_3  g0978(new_n1254, new_n1253);
nand_4 g0979(new_n1255_1, new_n1254, new_n1238);
nand_4 g0980(new_n1256, new_n1255_1, new_n1237_1);
nand_4 g0981(new_n1257, new_n1256, new_n1235_1);
nand_4 g0982(new_n1258, new_n1257, new_n1234_1);
nor_4  g0983(new_n1259, new_n1258, new_n1232);
nor_4  g0984(new_n1260_1, new_n1259, n1222);
not_3  g0985(new_n1261, n1222);
not_3  g0986(new_n1262, new_n1259);
nor_4  g0987(new_n1263_1, new_n1262, new_n1261);
nor_4  g0988(new_n1264, new_n1263_1, new_n1260_1);
xnor_3 g0989(new_n1265, new_n1264, new_n1231);
xnor_3 g0990(new_n1266, new_n1227, new_n545);
xnor_3 g0991(new_n1267, new_n1258, new_n1232);
nand_4 g0992(new_n1268, new_n1267, new_n1266);
not_3  g0993(new_n1269, new_n1268);
xnor_3 g0994(new_n1270, new_n1267, new_n1266);
xnor_3 g0995(new_n1271, new_n1226, new_n509);
not_3  g0996(new_n1272, new_n1271);
xnor_3 g0997(new_n1273, new_n1256, new_n1235_1);
nor_4  g0998(new_n1274, new_n1273, new_n1272);
xnor_3 g0999(new_n1275, new_n1273, new_n1271);
xnor_3 g1000(new_n1276, new_n1224, new_n1221);
xnor_3 g1001(new_n1277_1, new_n1253, new_n1238);
nand_4 g1002(new_n1278_1, new_n1277_1, new_n1276);
not_3  g1003(new_n1279, new_n1221);
xnor_3 g1004(new_n1280, new_n1224, new_n1279);
xnor_3 g1005(new_n1281, new_n1277_1, new_n1280);
not_3  g1006(new_n1282, new_n1251);
nor_4  g1007(new_n1283_1, new_n1282, new_n1242);
nor_4  g1008(new_n1284, new_n1283_1, new_n1252);
nand_4 g1009(new_n1285, new_n1284, new_n461);
xnor_3 g1010(new_n1286, new_n1284, new_n459);
not_3  g1011(new_n1287, new_n1249_1);
nor_4  g1012(new_n1288, new_n1287, new_n1245);
not_3  g1013(new_n1289, new_n1250);
nor_4  g1014(new_n1290, n1145, n1062);
nor_4  g1015(new_n1291, new_n1290, new_n1246);
nand_4 g1016(new_n1292, new_n1291, new_n466);
nand_4 g1017(new_n1293, new_n1292, new_n1289);
nor_4  g1018(new_n1294, new_n1293, new_n1288);
not_3  g1019(new_n1295, new_n1294);
nor_4  g1020(new_n1296_1, new_n1292, new_n1249_1);
nor_4  g1021(new_n1297, new_n1296_1, new_n1294);
nand_4 g1022(new_n1298, new_n1297, new_n471);
nand_4 g1023(new_n1299, new_n1298, new_n1295);
nand_4 g1024(new_n1300, new_n1299, new_n1286);
nand_4 g1025(new_n1301, new_n1300, new_n1285);
nand_4 g1026(new_n1302, new_n1301, new_n1281);
nand_4 g1027(new_n1303, new_n1302, new_n1278_1);
nand_4 g1028(new_n1304, new_n1303, new_n1275);
not_3  g1029(new_n1305_1, new_n1304);
nor_4  g1030(new_n1306, new_n1305_1, new_n1274);
nor_4  g1031(new_n1307, new_n1306, new_n1270);
nor_4  g1032(new_n1308, new_n1307, new_n1269);
xor_3  g1033(n317, new_n1308, new_n1265);
xor_3  g1034(n372, new_n1291, new_n466);
xor_3  g1035(n378, new_n904, new_n882_1);
not_3  g1036(new_n1312, new_n816);
nor_4  g1037(new_n1313, new_n972, new_n649_1);
nand_4 g1038(new_n1314, new_n1313, new_n700);
nor_4  g1039(new_n1315_1, new_n1314, new_n780);
nand_4 g1040(new_n1316, new_n1315_1, new_n793);
nor_4  g1041(new_n1317, new_n1316, new_n1312);
xor_3  g1042(n1425, new_n1317, new_n1202_1);
xor_3  g1043(n1249, new_n1315_1, new_n793);
not_3  g1044(new_n1320, n1249);
xor_3  g1045(n1119, new_n1313, new_n700);
not_3  g1046(new_n1322, n1119);
nand_4 g1047(new_n1323, new_n669, new_n524);
and_4  g1048(n647, new_n1323, new_n960);
not_3  g1049(n1255, n647);
xor_3  g1050(new_n1326, new_n961_1, new_n960);
nand_4 g1051(new_n1327, new_n1326, n1255);
xnor_3 g1052(n1016, new_n963, new_n957);
nor_4  g1053(new_n1329, n1016, new_n1327);
xnor_3 g1054(n1683, new_n966, new_n965);
not_3  g1055(new_n1331, n1683);
nor_4  g1056(new_n1332_1, new_n1331, new_n1329);
nor_4  g1057(new_n1333, new_n968_1, new_n951);
nor_4  g1058(new_n1334, new_n1333, new_n970);
not_3  g1059(n569, new_n1334);
nand_4 g1060(new_n1336, n569, new_n1332_1);
xor_3  g1061(n773, new_n971, new_n630);
not_3  g1062(new_n1338_1, n773);
nor_4  g1063(new_n1339, new_n1338_1, new_n1336);
nand_4 g1064(new_n1340_1, new_n1339, new_n690);
nor_4  g1065(new_n1341_1, new_n1340_1, new_n1322);
nand_4 g1066(new_n1342, new_n1341_1, new_n798);
nor_4  g1067(new_n1343, new_n1342, new_n1320);
nand_4 g1068(new_n1344, new_n1343, new_n816);
xnor_3 g1069(n387, new_n1344, n1425);
nor_4  g1070(new_n1346, new_n1229, new_n567);
nand_4 g1071(new_n1347_1, new_n1346, new_n563);
not_3  g1072(new_n1348_1, new_n1347_1);
nor_4  g1073(new_n1349_1, new_n1346, new_n563);
nor_4  g1074(new_n1350, new_n1349_1, new_n1348_1);
xnor_3 g1075(new_n1351_1, new_n1263_1, n1757);
not_3  g1076(new_n1352, new_n1351_1);
nor_4  g1077(new_n1353, new_n1352, new_n1350);
not_3  g1078(new_n1354, new_n1350);
nor_4  g1079(new_n1355, new_n1351_1, new_n1354);
nor_4  g1080(new_n1356, new_n1355, new_n1353);
nor_4  g1081(new_n1357, new_n1264, new_n1230);
not_3  g1082(new_n1358, new_n1265);
nor_4  g1083(new_n1359, new_n1308, new_n1358);
nor_4  g1084(new_n1360, new_n1359, new_n1357);
xor_3  g1085(n401, new_n1360, new_n1356);
not_3  g1086(n416, new_n578);
xnor_3 g1087(new_n1363_1, new_n898, new_n896);
xor_3  g1088(n423, new_n1363_1, new_n424_1);
nor_4  g1089(new_n1365, new_n1280, new_n396);
nor_4  g1090(new_n1366, new_n1276, new_n397);
nor_4  g1091(new_n1367, new_n1366, new_n1365);
not_3  g1092(new_n1368, new_n1367);
not_3  g1093(new_n1369_1, new_n460_1);
nand_4 g1094(new_n1370, new_n476_1, new_n463);
nand_4 g1095(new_n1371, new_n1370, new_n1369_1);
xor_3  g1096(n426, new_n1371, new_n1368);
not_3  g1097(new_n1373, new_n1344);
xor_3  g1098(n493, new_n1316, new_n1312);
nor_4  g1099(new_n1375, n493, new_n1343);
nor_4  g1100(n429, new_n1375, new_n1373);
xor_3  g1101(n432, new_n1338_1, new_n1336);
xnor_3 g1102(new_n1378, new_n1271, new_n391_1);
not_3  g1103(new_n1379, new_n1378);
not_3  g1104(new_n1380, new_n1365);
nand_4 g1105(new_n1381_1, new_n1371, new_n1367);
nand_4 g1106(new_n1382, new_n1381_1, new_n1380);
xor_3  g1107(n452, new_n1382, new_n1379);
not_3  g1108(new_n1384, new_n996);
nor_4  g1109(new_n1385_1, new_n1002, new_n1384);
xor_3  g1110(n457, new_n1171, new_n1385_1);
xnor_3 g1111(n460, new_n1214, new_n1211);
xor_3  g1112(n476, new_n749, new_n747_1);
not_3  g1113(new_n1389, new_n426_1);
xor_3  g1114(n482, new_n1389, new_n399);
nor_4  g1115(new_n1391, new_n1347_1, new_n496);
xor_3  g1116(new_n1392, new_n1391, new_n937);
xnor_3 g1117(new_n1393_1, new_n1392, new_n1135_1);
xnor_3 g1118(new_n1394, new_n1347_1, new_n496);
not_3  g1119(new_n1395, new_n1394);
nor_4  g1120(new_n1396, new_n1395, new_n1139);
xnor_3 g1121(new_n1397, new_n1394, new_n1140_1);
not_3  g1122(new_n1398, new_n1143);
nor_4  g1123(new_n1399_1, new_n1350, new_n1398);
xnor_3 g1124(new_n1400, new_n1350, new_n1398);
xnor_3 g1125(new_n1401, new_n302, new_n1132);
nor_4  g1126(new_n1402, new_n1231, new_n1401);
not_3  g1127(new_n1403, new_n1402);
not_3  g1128(new_n1404, new_n1266);
nor_4  g1129(new_n1405, new_n1404, new_n388);
not_3  g1130(new_n1406, new_n1405);
nor_4  g1131(new_n1407_1, new_n1266, new_n385);
nor_4  g1132(new_n1408, new_n1407_1, new_n1405);
nand_4 g1133(new_n1409, new_n1271, new_n392);
nand_4 g1134(new_n1410, new_n1382, new_n1378);
nand_4 g1135(new_n1411, new_n1410, new_n1409);
nand_4 g1136(new_n1412, new_n1411, new_n1408);
nand_4 g1137(new_n1413, new_n1412, new_n1406);
not_3  g1138(new_n1414, new_n1413);
nor_4  g1139(new_n1415, new_n1230, new_n303_1);
nor_4  g1140(new_n1416, new_n1415, new_n1402);
nand_4 g1141(new_n1417, new_n1416, new_n1414);
nand_4 g1142(new_n1418, new_n1417, new_n1403);
nor_4  g1143(new_n1419, new_n1418, new_n1400);
nor_4  g1144(new_n1420, new_n1419, new_n1399_1);
nor_4  g1145(new_n1421, new_n1420, new_n1397);
nor_4  g1146(new_n1422_1, new_n1421, new_n1396);
xnor_3 g1147(n510, new_n1422_1, new_n1393_1);
xnor_3 g1148(new_n1424, new_n1139, new_n1112);
nor_4  g1149(new_n1425_1, new_n1398, new_n1115);
not_3  g1150(new_n1426_1, new_n1425_1);
not_3  g1151(new_n1427, new_n1115);
nor_4  g1152(new_n1428, new_n1143, new_n1427);
nor_4  g1153(new_n1429, new_n1428, new_n1425_1);
nor_4  g1154(new_n1430, new_n1120, new_n303_1);
not_3  g1155(new_n1431, new_n1430);
not_3  g1156(new_n1432, new_n1120);
nor_4  g1157(new_n1433, new_n1432, new_n1401);
nor_4  g1158(new_n1434, new_n1433, new_n1430);
nor_4  g1159(new_n1435_1, new_n1025_1, new_n388);
not_3  g1160(new_n1436, new_n1435_1);
not_3  g1161(new_n1437, new_n1025_1);
nor_4  g1162(new_n1438, new_n1437, new_n385);
nor_4  g1163(new_n1439, new_n1438, new_n1435_1);
nor_4  g1164(new_n1440_1, new_n1089, new_n392);
nand_4 g1165(new_n1441, new_n1057, new_n397);
xnor_3 g1166(new_n1442, new_n1057, new_n396);
nor_4  g1167(new_n1443, new_n1062_1, new_n400);
not_3  g1168(new_n1444, new_n1443);
nor_4  g1169(new_n1445, new_n1063, new_n401_1);
nor_4  g1170(new_n1446, new_n1445, new_n1443);
not_3  g1171(new_n1447, new_n1073);
nor_4  g1172(new_n1448, new_n1447, new_n465);
nor_4  g1173(new_n1449, new_n1448, new_n410);
not_3  g1174(new_n1450, new_n1449);
not_3  g1175(new_n1451, new_n1448);
nor_4  g1176(new_n1452, new_n1451, new_n291);
nor_4  g1177(new_n1453_1, new_n1452, new_n1449);
nand_4 g1178(new_n1454, new_n1453_1, new_n1078);
nand_4 g1179(new_n1455, new_n1454, new_n1450);
nand_4 g1180(new_n1456, new_n1455, new_n1446);
nand_4 g1181(new_n1457_1, new_n1456, new_n1444);
nand_4 g1182(new_n1458, new_n1457_1, new_n1442);
nand_4 g1183(new_n1459, new_n1458, new_n1441);
xnor_3 g1184(new_n1460_1, new_n1054, new_n391_1);
nor_4  g1185(new_n1461_1, new_n1460_1, new_n1459);
nor_4  g1186(new_n1462, new_n1461_1, new_n1440_1);
nand_4 g1187(new_n1463_1, new_n1462, new_n1439);
nand_4 g1188(new_n1464, new_n1463_1, new_n1436);
nand_4 g1189(new_n1465, new_n1464, new_n1434);
nand_4 g1190(new_n1466, new_n1465, new_n1431);
nand_4 g1191(new_n1467, new_n1466, new_n1429);
nand_4 g1192(new_n1468, new_n1467, new_n1426_1);
xor_3  g1193(n517, new_n1468, new_n1424);
xnor_3 g1194(new_n1470_1, new_n1140_1, new_n832);
nand_4 g1195(new_n1471, new_n1143, new_n706);
xnor_3 g1196(new_n1472, new_n1143, new_n838);
nand_4 g1197(new_n1473, new_n770_1, new_n1401);
nand_4 g1198(new_n1474, new_n715_1, new_n385);
xnor_3 g1199(new_n1475, new_n715_1, new_n388);
nand_4 g1200(new_n1476, new_n721, new_n392);
nand_4 g1201(new_n1477, new_n1196, new_n1177);
nand_4 g1202(new_n1478, new_n1477, new_n1476);
nand_4 g1203(new_n1479, new_n1478, new_n1475);
nand_4 g1204(new_n1480, new_n1479, new_n1474);
xnor_3 g1205(new_n1481_1, new_n712_1, new_n1401);
nand_4 g1206(new_n1482, new_n1481_1, new_n1480);
nand_4 g1207(new_n1483, new_n1482, new_n1473);
nand_4 g1208(new_n1484, new_n1483, new_n1472);
nand_4 g1209(new_n1485, new_n1484, new_n1471);
xnor_3 g1210(n522, new_n1485, new_n1470_1);
xor_3  g1211(new_n1487, new_n1155, new_n1142_1);
xnor_3 g1212(n532, new_n1173, new_n1487);
not_3  g1213(new_n1489, new_n318);
nor_4  g1214(new_n1490, new_n1201_1, new_n1489);
not_3  g1215(new_n1491, new_n379_1);
nor_4  g1216(new_n1492, new_n1491, new_n361);
xor_3  g1217(new_n1493, new_n373, new_n478);
nand_4 g1218(new_n1494, new_n1493, n1000);
nor_4  g1219(new_n1495_1, new_n693_1, n682);
nand_4 g1220(new_n1496, new_n364, n1527);
not_3  g1221(new_n1497, new_n1496);
nor_4  g1222(new_n1498_1, new_n1497, new_n1495_1);
nand_4 g1223(new_n1499, new_n1498_1, new_n305);
nand_4 g1224(new_n1500, new_n1499, new_n1494);
nand_4 g1225(new_n1501_1, new_n1500, new_n1492);
xor_3  g1226(new_n1502_1, new_n1495_1, n379);
nand_4 g1227(new_n1503, new_n1502_1, new_n305);
nand_4 g1228(new_n1504, new_n373, n247);
xor_3  g1229(new_n1505, new_n1504, new_n492);
nand_4 g1230(new_n1506, new_n1505, n1000);
nand_4 g1231(new_n1507_1, new_n1506, new_n1503);
nor_4  g1232(new_n1508, new_n1507_1, new_n1501_1);
nand_4 g1233(new_n1509, new_n1495_1, new_n486);
nand_4 g1234(new_n1510, new_n1509, n1263);
nor_4  g1235(new_n1511, new_n810, n682);
nor_4  g1236(new_n1512, new_n1511, n1000);
nand_4 g1237(new_n1513, new_n1512, new_n1510);
nor_4  g1238(new_n1514, new_n1504, new_n492);
xor_3  g1239(new_n1515, new_n1514, new_n908);
nand_4 g1240(new_n1516, new_n1515, n1000);
nand_4 g1241(new_n1517, new_n1516, new_n1513);
nand_4 g1242(new_n1518, new_n1517, new_n1508);
nand_4 g1243(new_n1519, new_n1514, n171);
nand_4 g1244(new_n1520, n1000, n557);
nor_4  g1245(new_n1521, new_n1520, new_n1519);
nand_4 g1246(new_n1522, new_n1512, n1422);
not_3  g1247(new_n1523, new_n1520);
nor_4  g1248(new_n1524, new_n1519, new_n305);
nor_4  g1249(new_n1525_1, new_n1524, new_n1523);
nand_4 g1250(new_n1526, new_n1525_1, new_n1522);
nor_4  g1251(new_n1527_1, new_n1526, new_n1490);
nor_4  g1252(new_n1528, new_n1527_1, new_n1521);
nor_4  g1253(new_n1529, new_n1528, new_n1518);
nor_4  g1254(new_n1530_1, new_n1521, new_n1490);
and_4  g1255(new_n1531, new_n1530_1, new_n1529);
nor_4  g1256(new_n1532, new_n1531, new_n1490);
not_3  g1257(new_n1533, new_n1518);
xor_3  g1258(new_n1534, new_n1528, new_n1533);
not_3  g1259(new_n1535_1, new_n1534);
not_3  g1260(new_n1536, new_n322);
xor_3  g1261(new_n1537_1, n1597, new_n362);
nand_4 g1262(new_n1538, new_n1537_1, new_n305);
not_3  g1263(new_n1539, new_n326);
nand_4 g1264(new_n1540, new_n1539, new_n1538);
nor_4  g1265(new_n1541, new_n1540, new_n1536);
nand_4 g1266(new_n1542, new_n379_1, new_n1541);
xor_3  g1267(new_n1543, new_n373, n247);
nor_4  g1268(new_n1544_1, new_n1543, new_n305);
not_3  g1269(new_n1545, new_n1499);
nor_4  g1270(new_n1546, new_n1545, new_n1544_1);
nor_4  g1271(new_n1547, new_n1546, new_n1542);
xor_3  g1272(new_n1548, new_n1495_1, new_n486);
nor_4  g1273(new_n1549, new_n1548, n1000);
xor_3  g1274(new_n1550, new_n1504, n1642);
nor_4  g1275(new_n1551, new_n1550, new_n305);
nor_4  g1276(new_n1552, new_n1551, new_n1549);
nor_4  g1277(new_n1553, new_n1552, new_n1547);
nor_4  g1278(new_n1554, new_n1553, new_n1508);
nor_4  g1279(new_n1555, new_n380, new_n360);
xnor_3 g1280(new_n1556_1, new_n1500, new_n1492);
nand_4 g1281(new_n1557, new_n1556_1, new_n1555);
nor_4  g1282(new_n1558, new_n1557, new_n1554);
xnor_3 g1283(new_n1559, new_n1517, new_n1508);
nand_4 g1284(new_n1560, new_n1559, new_n1558);
nor_4  g1285(new_n1561, new_n1560, new_n1535_1);
nor_4  g1286(new_n1562, new_n1561, new_n1532);
not_3  g1287(new_n1563, new_n1562);
xnor_3 g1288(new_n1564, new_n1560, new_n1534);
not_3  g1289(new_n1565, new_n1564);
not_3  g1290(new_n1566, n277);
not_3  g1291(new_n1567, n1622);
not_3  g1292(new_n1568, n49);
nor_4  g1293(new_n1569, n1643, n469);
not_3  g1294(new_n1570, new_n1569);
nand_4 g1295(new_n1571, new_n872, new_n853);
nand_4 g1296(new_n1572, new_n1571, new_n1570);
nor_4  g1297(new_n1573, new_n1572, new_n1568);
not_3  g1298(new_n1574, new_n1573);
nor_4  g1299(new_n1575, new_n1574, new_n1567);
nand_4 g1300(new_n1576, new_n1575, n906);
nor_4  g1301(new_n1577, new_n1576, new_n1566);
not_3  g1302(new_n1578, new_n1560);
nor_4  g1303(new_n1579, new_n1559, new_n1558);
nor_4  g1304(new_n1580, new_n1579, new_n1578);
nor_4  g1305(new_n1581, new_n1580, new_n1577);
not_3  g1306(new_n1582, new_n1581);
not_3  g1307(new_n1583, new_n1577);
not_3  g1308(new_n1584, new_n1580);
nor_4  g1309(new_n1585, new_n1584, new_n1583);
nor_4  g1310(new_n1586, new_n1585, new_n1581);
not_3  g1311(new_n1587, new_n1576);
nor_4  g1312(new_n1588, new_n1587, n277);
nor_4  g1313(new_n1589, new_n1588, new_n1577);
xnor_3 g1314(new_n1590, new_n1557, new_n1554);
not_3  g1315(new_n1591, new_n1590);
nor_4  g1316(new_n1592, new_n1591, new_n1589);
not_3  g1317(new_n1593, new_n1592);
not_3  g1318(new_n1594, new_n1589);
nor_4  g1319(new_n1595_1, new_n1590, new_n1594);
nor_4  g1320(new_n1596, new_n1595_1, new_n1592);
nor_4  g1321(new_n1597_1, new_n1575, n906);
nor_4  g1322(new_n1598, new_n1597_1, new_n1587);
nor_4  g1323(new_n1599, new_n1500, new_n1492);
nor_4  g1324(new_n1600_1, new_n1599, new_n1547);
xnor_3 g1325(new_n1601_1, new_n1600_1, new_n1555);
nor_4  g1326(new_n1602, new_n1601_1, new_n1598);
not_3  g1327(new_n1603, new_n1602);
xnor_3 g1328(new_n1604, new_n1601_1, new_n1598);
not_3  g1329(new_n1605, new_n1604);
not_3  g1330(new_n1606, new_n381);
nor_4  g1331(new_n1607, new_n1573, n1622);
nor_4  g1332(new_n1608, new_n1607, new_n1575);
nor_4  g1333(new_n1609, new_n1608, new_n1606);
not_3  g1334(new_n1610, new_n1609);
xnor_3 g1335(new_n1611, new_n1608, new_n1606);
not_3  g1336(new_n1612, new_n1611);
xnor_3 g1337(new_n1613_1, new_n1572, new_n1568);
nor_4  g1338(new_n1614, new_n1613_1, new_n384);
not_3  g1339(new_n1615, new_n1614);
xnor_3 g1340(new_n1616, new_n1613_1, new_n384);
not_3  g1341(new_n1617, new_n1616);
nand_4 g1342(new_n1618, new_n906_1, new_n877);
nand_4 g1343(new_n1619, new_n1618, new_n874);
nand_4 g1344(new_n1620, new_n1619, new_n1617);
nand_4 g1345(new_n1621, new_n1620, new_n1615);
not_3  g1346(new_n1622_1, new_n1621);
nand_4 g1347(new_n1623, new_n1622_1, new_n1612);
nand_4 g1348(new_n1624, new_n1623, new_n1610);
nand_4 g1349(new_n1625, new_n1624, new_n1605);
nand_4 g1350(new_n1626, new_n1625, new_n1603);
nand_4 g1351(new_n1627, new_n1626, new_n1596);
nand_4 g1352(new_n1628, new_n1627, new_n1593);
nand_4 g1353(new_n1629_1, new_n1628, new_n1586);
nand_4 g1354(new_n1630, new_n1629_1, new_n1582);
nor_4  g1355(new_n1631, new_n1630, new_n1565);
nor_4  g1356(n534, new_n1631, new_n1563);
not_3  g1357(new_n1633_1, new_n579);
xor_3  g1358(n541, n1721, new_n1633_1);
not_3  g1359(n547, n1426);
nor_4  g1360(new_n1636, new_n1209, new_n1135_1);
xnor_3 g1361(new_n1637, new_n1209, new_n1135_1);
nor_4  g1362(new_n1638, new_n1139, new_n1112);
not_3  g1363(new_n1639, new_n1468);
nor_4  g1364(new_n1640, new_n1639, new_n1424);
nor_4  g1365(new_n1641, new_n1640, new_n1638);
nor_4  g1366(new_n1642_1, new_n1641, new_n1637);
nor_4  g1367(new_n1643_1, new_n1642_1, new_n1636);
nand_4 g1368(new_n1644, new_n1643_1, new_n1207);
nand_4 g1369(new_n1645, new_n1644, new_n1206);
nor_4  g1370(n549, new_n1645, new_n1203);
xnor_3 g1371(n559, new_n1481_1, new_n1480);
xor_3  g1372(n573, new_n1460_1, new_n1459);
xnor_3 g1373(n588, new_n1641, new_n1637);
not_3  g1374(new_n1650, new_n575);
xor_3  g1375(n599, new_n578, new_n1650);
nor_4  g1376(n824, new_n1317, new_n1203);
not_3  g1377(new_n1653, n824);
nor_4  g1378(n627, new_n1373, new_n1653);
not_3  g1379(new_n1655, new_n1207);
xnor_3 g1380(n638, new_n1216, new_n1655);
nor_4  g1381(new_n1657_1, new_n928, n557);
nand_4 g1382(new_n1658, new_n1657_1, n1381);
or_4   g1383(new_n1659, new_n808, new_n440);
nand_4 g1384(new_n1660_1, new_n1659, new_n1658);
nand_4 g1385(new_n1661, new_n1660_1, new_n934);
not_3  g1386(n643, new_n1661);
not_3  g1387(new_n1663, new_n960);
xor_3  g1388(n646, new_n961_1, new_n1663);
xor_3  g1389(n648, new_n1619, new_n1617);
xnor_3 g1390(n665, new_n767, new_n720);
xnor_3 g1391(n683, new_n1127, new_n1117);
nor_4  g1392(new_n1668, new_n1564, new_n1135_1);
not_3  g1393(new_n1669, new_n1668);
not_3  g1394(new_n1670, new_n1135_1);
xnor_3 g1395(new_n1671, new_n1564, new_n1670);
nand_4 g1396(new_n1672, new_n1584, new_n1670);
xnor_3 g1397(new_n1673, new_n1580, new_n1670);
nand_4 g1398(new_n1674, new_n1590, new_n1140_1);
xnor_3 g1399(new_n1675_1, new_n1590, new_n1139);
xnor_3 g1400(new_n1676, new_n1556_1, new_n1555);
nand_4 g1401(new_n1677_1, new_n1676, new_n1143);
xnor_3 g1402(new_n1678_1, new_n1601_1, new_n1143);
nand_4 g1403(new_n1679, new_n381, new_n1401);
nand_4 g1404(new_n1680, new_n433_1, new_n382);
nand_4 g1405(new_n1681, new_n1680, new_n1679);
nand_4 g1406(new_n1682, new_n1681, new_n1678_1);
nand_4 g1407(new_n1683_1, new_n1682, new_n1677_1);
nand_4 g1408(new_n1684, new_n1683_1, new_n1675_1);
nand_4 g1409(new_n1685, new_n1684, new_n1674);
nand_4 g1410(new_n1686_1, new_n1685, new_n1673);
nand_4 g1411(new_n1687, new_n1686_1, new_n1672);
nand_4 g1412(new_n1688_1, new_n1687, new_n1671);
nand_4 g1413(new_n1689, new_n1688_1, new_n1669);
xor_3  g1414(new_n1690_1, new_n1530_1, new_n1529);
xnor_3 g1415(new_n1691, new_n1690_1, new_n1561);
nand_4 g1416(new_n1692, new_n1691, new_n1689);
nor_4  g1417(new_n1693, new_n1691, new_n1135_1);
not_3  g1418(new_n1694, new_n1671);
not_3  g1419(new_n1695, new_n1687);
nor_4  g1420(new_n1696, new_n1695, new_n1694);
nor_4  g1421(new_n1697, new_n1696, new_n1670);
nor_4  g1422(new_n1698, new_n1697, new_n1693);
nand_4 g1423(new_n1699, new_n1698, new_n1692);
xnor_3 g1424(n699, new_n1699, new_n1562);
xor_3  g1425(n712, new_n894, new_n415);
not_3  g1426(n715, new_n586);
not_3  g1427(new_n1703, new_n1340_1);
nor_4  g1428(new_n1704, new_n1339, n145);
nor_4  g1429(n724, new_n1704, new_n1703);
not_3  g1430(new_n1706, n1016);
xor_3  g1431(n725, new_n1706, new_n1327);
xnor_3 g1432(n731, new_n1483, new_n1472);
xnor_3 g1433(n748, new_n1681, new_n1678_1);
xnor_3 g1434(n759, new_n1418, new_n1400);
not_3  g1435(new_n1711, new_n1173);
nand_4 g1436(new_n1712, new_n1711, new_n1164);
nor_4  g1437(new_n1713, new_n1712, new_n1162_1);
nor_4  g1438(new_n1714, new_n1135_1, n1263);
nor_4  g1439(new_n1715, new_n1159, new_n1714);
nor_4  g1440(new_n1716, new_n1715, n1422);
nand_4 g1441(new_n1717, new_n1716, new_n1713);
not_3  g1442(n770, new_n1717);
not_3  g1443(new_n1719, new_n1439);
xor_3  g1444(n790, new_n1462, new_n1719);
xor_3  g1445(new_n1721_1, new_n1135_1, new_n825);
nor_4  g1446(new_n1722, new_n1139, new_n832);
nand_4 g1447(new_n1723, new_n1485, new_n1470_1);
not_3  g1448(new_n1724, new_n1723);
nor_4  g1449(new_n1725, new_n1724, new_n1722);
xor_3  g1450(n792, new_n1725, new_n1721_1);
not_3  g1451(new_n1727_1, new_n1093);
xor_3  g1452(n813, new_n1727_1, new_n1088);
not_3  g1453(new_n1729_1, new_n1286);
xor_3  g1454(n823, new_n1299, new_n1729_1);
not_3  g1455(new_n1731_1, new_n471);
xor_3  g1456(n836, new_n474, new_n1731_1);
xnor_3 g1457(n846, new_n1683_1, new_n1675_1);
not_3  g1458(new_n1734, new_n1270);
xor_3  g1459(n858, new_n1306, new_n1734);
xor_3  g1460(n865, new_n1314, new_n780);
not_3  g1461(new_n1737_1, new_n1429);
xor_3  g1462(n867, new_n1466, new_n1737_1);
not_3  g1463(new_n1739, new_n1391);
nor_4  g1464(new_n1740, new_n1739, new_n919);
not_3  g1465(new_n1741, new_n1740);
xor_3  g1466(new_n1742, new_n1741, new_n931_1);
not_3  g1467(new_n1743_1, new_n1742);
nor_4  g1468(new_n1744, new_n1392, new_n1135_1);
nor_4  g1469(new_n1745, new_n1422_1, new_n1393_1);
nor_4  g1470(new_n1746_1, new_n1745, new_n1744);
xnor_3 g1471(n883, new_n1746_1, new_n1743_1);
not_3  g1472(new_n1748, new_n771);
xor_3  g1473(n888, new_n1748, new_n769);
not_3  g1474(new_n1750, new_n1392);
not_3  g1475(new_n1751, n839);
nand_4 g1476(new_n1752, new_n1263_1, n1757);
nor_4  g1477(new_n1753, new_n1752, new_n1751);
not_3  g1478(new_n1754, new_n1753);
nand_4 g1479(new_n1755, new_n1754, new_n1750);
not_3  g1480(new_n1756, new_n1755);
xnor_3 g1481(new_n1757_1, new_n1753, new_n1392);
not_3  g1482(new_n1758, new_n1752);
nor_4  g1483(new_n1759, new_n1758, n839);
nor_4  g1484(new_n1760, new_n1759, new_n1753);
nor_4  g1485(new_n1761, new_n1760, new_n1395);
not_3  g1486(new_n1762, new_n1760);
nor_4  g1487(new_n1763_1, new_n1762, new_n1394);
nor_4  g1488(new_n1764_1, new_n1763_1, new_n1761);
not_3  g1489(new_n1765, new_n1764_1);
not_3  g1490(new_n1766, new_n1356);
nor_4  g1491(new_n1767, new_n1360, new_n1766);
nor_4  g1492(new_n1768, new_n1767, new_n1353);
nor_4  g1493(new_n1769, new_n1768, new_n1765);
nor_4  g1494(new_n1770, new_n1769, new_n1761);
nor_4  g1495(new_n1771, new_n1770, new_n1757_1);
nor_4  g1496(new_n1772, new_n1771, new_n1756);
nand_4 g1497(new_n1773, new_n1772, new_n1742);
not_3  g1498(new_n1774, new_n1773);
nor_4  g1499(new_n1775, new_n1772, new_n1742);
nor_4  g1500(n891, new_n1775, new_n1774);
not_3  g1501(new_n1777, new_n1660_1);
nor_4  g1502(new_n1778, new_n1741, new_n931_1);
not_3  g1503(new_n1779, new_n1778);
nand_4 g1504(new_n1780, new_n1773, new_n1779);
nor_4  g1505(n892, new_n1780, new_n1777);
xor_3  g1506(n902, new_n1073, new_n1071);
xor_3  g1507(n905, new_n1194_1, new_n1193);
not_3  g1508(new_n1784, new_n1174);
nand_4 g1509(new_n1785, new_n1170, new_n1385_1);
nand_4 g1510(new_n1786, new_n1785, new_n1166);
nand_4 g1511(n912, new_n1786, new_n1784);
nor_4  g1512(new_n1788, n1149, new_n593);
nor_4  g1513(n935, new_n1788, new_n941);
xor_3  g1514(n942, new_n1703, n1119);
not_3  g1515(new_n1791, new_n1122);
xor_3  g1516(n944, new_n1125, new_n1791);
nor_4  g1517(new_n1793, new_n1175_1, new_n1162_1);
nand_4 g1518(new_n1794, new_n1716, new_n1793);
not_3  g1519(n974, new_n1794);
not_3  g1520(new_n1796, new_n389);
xor_3  g1521(n979, new_n431, new_n1796);
not_3  g1522(new_n1798, new_n803);
nor_4  g1523(new_n1799, new_n817, new_n1798);
nor_4  g1524(new_n1800, new_n816, new_n804);
nor_4  g1525(new_n1801, new_n1202_1, new_n1800);
nor_4  g1526(new_n1802, new_n1801, new_n1799);
not_3  g1527(new_n1803, new_n1802);
nor_4  g1528(n980, new_n1803, new_n850);
not_3  g1529(new_n1805, new_n1434);
xor_3  g1530(n989, new_n1464, new_n1805);
xor_3  g1531(n991, new_n1695, new_n1671);
xor_3  g1532(n1005, new_n1768, new_n1764_1);
xnor_3 g1533(n1012, new_n1420, new_n1397);
xor_3  g1534(n1015, new_n1168, new_n1384);
nand_4 g1535(new_n1811, new_n1801, new_n850);
not_3  g1536(new_n1812, new_n850);
nand_4 g1537(new_n1813, new_n1801, new_n1799);
and_4  g1538(new_n1814, new_n1813, new_n1803);
not_3  g1539(new_n1815, new_n1814);
nand_4 g1540(new_n1816, new_n1815, new_n1812);
nand_4 g1541(n1025, new_n1816, new_n1811);
xnor_3 g1542(n1030, new_n1770, new_n1757_1);
not_3  g1543(new_n1819, new_n842);
xor_3  g1544(n1067, new_n1819, new_n836_1);
xnor_3 g1545(n1068, new_n1780, new_n1777);
xor_3  g1546(n1103, new_n586, new_n583);
xor_3  g1547(n1113, new_n467, new_n465);
nor_4  g1548(new_n1824, new_n1173, new_n1487);
nand_4 g1549(new_n1825, new_n1824, new_n1161_1);
not_3  g1550(new_n1826, new_n1715);
nor_4  g1551(new_n1827, new_n1826, new_n806);
nand_4 g1552(new_n1828, new_n1827, new_n1825);
nand_4 g1553(n1135, new_n1828, new_n1717);
nand_4 g1554(new_n1830, new_n1690_1, new_n1631);
not_3  g1555(new_n1831, new_n1631);
nand_4 g1556(new_n1832, new_n1691, new_n1831);
nand_4 g1557(n1142, new_n1832, new_n1830);
not_3  g1558(new_n1834, new_n1689);
xnor_3 g1559(new_n1835, new_n1691, new_n1135_1);
xnor_3 g1560(n1161, new_n1835, new_n1834);
xor_3  g1561(n1162, new_n1170, new_n1169);
not_3  g1562(new_n1838, new_n1342);
nor_4  g1563(new_n1839, n865, new_n1341_1);
nor_4  g1564(n1175, new_n1839, new_n1838);
nor_4  g1565(new_n1841, new_n1135_1, new_n819);
nor_4  g1566(new_n1842, new_n1135_1, new_n824_1);
and_4  g1567(new_n1843, new_n1842, new_n1725);
not_3  g1568(new_n1844, new_n1722);
nand_4 g1569(new_n1845, new_n1723, new_n1844);
nand_4 g1570(new_n1846, new_n1845, new_n1721_1);
nor_4  g1571(new_n1847, new_n1846, new_n819);
nor_4  g1572(new_n1848, new_n1847, new_n1843);
nor_4  g1573(new_n1849, new_n1848, new_n1841);
xnor_3 g1574(n1191, new_n1849, new_n1814);
not_3  g1575(new_n1851, new_n1172_1);
xor_3  g1576(n1194, new_n1851, new_n1167);
xor_3  g1577(n1199, new_n429_1, new_n428);
not_3  g1578(new_n1854, new_n1446);
xor_3  g1579(n1201, new_n1455, new_n1854);
not_3  g1580(new_n1856, new_n962);
nand_4 g1581(new_n1857, new_n1323, new_n1856);
nand_4 g1582(n1202, new_n1857, new_n1327);
xor_3  g1583(n1234, n569, new_n1332_1);
xnor_3 g1584(n1235, new_n1712, new_n1162_1);
not_3  g1585(n1237, n1183);
xnor_3 g1586(n1260, new_n1218, new_n1203);
nor_4  g1587(new_n1863, new_n1838, n1249);
nor_4  g1588(n1277, new_n1863, new_n1343);
nand_4 g1589(new_n1865, new_n1746_1, new_n1742);
nand_4 g1590(new_n1866, new_n1865, new_n1779);
nor_4  g1591(n1278, new_n1866, new_n1777);
nor_4  g1592(new_n1868, new_n415, new_n412);
not_3  g1593(new_n1869, new_n413);
nor_4  g1594(new_n1870, new_n892_1, new_n1869);
nor_4  g1595(new_n1871, new_n1870, new_n418);
nor_4  g1596(n1283, new_n1871, new_n1868);
nor_4  g1597(new_n1873, new_n1784, new_n1487);
nand_4 g1598(new_n1874, new_n1873, new_n1161_1);
nand_4 g1599(new_n1875, new_n1827, new_n1874);
nand_4 g1600(n1305, new_n1875, new_n1794);
xor_3  g1601(n1315, new_n587, n1727);
not_3  g1602(new_n1878, new_n1596);
xor_3  g1603(n1330, new_n1626, new_n1878);
not_3  g1604(new_n1880, new_n1475);
xor_3  g1605(n1338, new_n1478, new_n1880);
not_3  g1606(new_n1882, new_n754);
xor_3  g1607(n1340, new_n756, new_n1882);
not_3  g1608(new_n1884, new_n1630);
nor_4  g1609(new_n1885, new_n1884, new_n1564);
nor_4  g1610(n1347, new_n1885, new_n1631);
nor_4  g1611(new_n1887, new_n1660_1, new_n934);
nor_4  g1612(new_n1888, new_n1887, n643);
not_3  g1613(n1348, new_n1888);
not_3  g1614(new_n1890, new_n1275);
xor_3  g1615(n1349, new_n1303, new_n1890);
nor_4  g1616(new_n1892, new_n1827, new_n1716);
xnor_3 g1617(n1369, new_n1892, new_n1825);
xnor_3 g1618(n1383, new_n1892, new_n1874);
xor_3  g1619(n1393, new_n1622_1, new_n1611);
not_3  g1620(new_n1896, new_n1078);
xor_3  g1621(n1399, new_n1453_1, new_n1896);
xor_3  g1622(n1407, new_n1191_1, new_n1190);
nor_4  g1623(n1440, new_n1661, new_n943);
xor_3  g1624(n1453, new_n1000_1, new_n998);
xor_3  g1625(n1460, new_n1188, new_n1882);
not_3  g1626(new_n1902, new_n1843);
not_3  g1627(new_n1903, new_n1846);
nand_4 g1628(new_n1904, new_n1903, new_n1135_1);
nand_4 g1629(new_n1905, new_n1904, new_n1902);
xnor_3 g1630(n1463, new_n1905, new_n849);
xnor_3 g1631(n1470, new_n1784, new_n1487);
xor_3  g1632(n1481, new_n1447, new_n465);
not_3  g1633(new_n1909, new_n758);
xor_3  g1634(n1495, new_n761_1, new_n1909);
not_3  g1635(new_n1911, new_n1061);
xor_3  g1636(n1498, new_n1086, new_n1911);
xor_3  g1637(n1502, new_n1624, new_n1604);
not_3  g1638(new_n1914, new_n1301);
xor_3  g1639(n1507, new_n1914, new_n1281);
xor_3  g1640(n1525, new_n1331, new_n1329);
not_3  g1641(new_n1917, new_n763);
xor_3  g1642(n1535, new_n1917, new_n740);
not_3  g1643(n1601, new_n1000_1);
xor_3  g1644(n1556, n1601, n1426);
xnor_3 g1645(n1595, new_n1888, new_n943);
xnor_3 g1646(n1600, new_n1457_1, new_n1442);
not_3  g1647(new_n1923, new_n528);
and_4  g1648(new_n1924, new_n573_1, new_n1923);
or_4   g1649(n1613, new_n1924, new_n575);
xor_3  g1650(n1629, new_n1297, new_n1731_1);
nor_4  g1651(new_n1927, new_n1849, new_n1802);
nand_4 g1652(new_n1928, new_n1843, new_n819);
nand_4 g1653(new_n1929, new_n1928, new_n1813);
nor_4  g1654(n1633, new_n1929, new_n1927);
xor_3  g1655(n1635, new_n1001, new_n997);
xor_3  g1656(n1654, new_n1416, new_n1414);
nor_4  g1657(new_n1933, new_n589, n1138);
nor_4  g1658(n1657, new_n1933, new_n591);
xnor_3 g1659(n1660, new_n1866, new_n1777);
xor_3  g1660(n1675, new_n1081, new_n1896);
xnor_3 g1661(n1686, new_n1643_1, new_n1655);
xor_3  g1662(n1688, new_n1184, new_n465);
xnor_3 g1663(n1690, new_n1628, new_n1586);
xnor_3 g1664(n1729, new_n1685, new_n1673);
xnor_3 g1665(n1737, new_n1645, new_n1203);
not_3  g1666(new_n1942, new_n1408);
xor_3  g1667(n1746, new_n1411, new_n1942);
xor_3  g1668(n488, new_n404, n347);
xor_3  g1669(n1677, new_n1199_1, new_n986);
endmodule


