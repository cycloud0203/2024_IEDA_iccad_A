// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Fri Jun 14 22:42:05 2024

module top_810026173_826291639_946996917_1246901 ( 
    n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213, n223,
    n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414, n424,
    n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649, n653,
    n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788, n801,
    n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764,
    n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156, n174,
    n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299, n317,
    n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457, n460,
    n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547, n549,
    n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648, n665,
    n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773, n790,
    n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888, n891,
    n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989, n991,
    n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103, n1113,
    n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183, n1191,
    n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255, n1260,
    n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347, n1348,
    n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426, n1440,
    n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502, n1507,
    n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633, n1635,
    n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690, n1721,
    n1727, n1729, n1731, n1737, n1746  );
  input  n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213,
    n223, n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414,
    n424, n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649,
    n653, n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788,
    n801, n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764;
  output n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156,
    n174, n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299,
    n317, n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457,
    n460, n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547,
    n549, n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648,
    n665, n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773,
    n790, n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888,
    n891, n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989,
    n991, n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103,
    n1113, n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183,
    n1191, n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255,
    n1260, n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347,
    n1348, n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426,
    n1440, n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502,
    n1507, n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633,
    n1635, n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690,
    n1721, n1727, n1729, n1731, n1737, n1746;
  wire new_n276_1, new_n277_1, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290_1, new_n291, new_n292_1, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299_1, new_n300, new_n301,
    new_n302, new_n303_1, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317_1, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329_1,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347_1, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353_1, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372_1, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378_1, new_n379_1, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387_1, new_n388, new_n389, new_n390,
    new_n391_1, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401_1, new_n402_1, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414_1, new_n415, new_n416_1,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423_1,
    new_n424_1, new_n425, new_n426_1, new_n427, new_n428, new_n429_1,
    new_n430, new_n431, new_n432_1, new_n433_1, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444_1, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452_1, new_n453, new_n454, new_n455, new_n456,
    new_n457_1, new_n458, new_n459, new_n460_1, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469_1,
    new_n470, new_n471, new_n472_1, new_n473, new_n474, new_n475,
    new_n476_1, new_n478, new_n479, new_n480, new_n481, new_n482_1,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488_1, new_n489,
    new_n490, new_n491, new_n492, new_n493_1, new_n494, new_n495, new_n496,
    new_n497, new_n498_1, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510_1,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517_1,
    new_n518, new_n519, new_n520, new_n521, new_n522_1, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532_1, new_n533, new_n534_1, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541_1, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547_1, new_n548, new_n549_1, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555_1, new_n556,
    new_n557_1, new_n558, new_n559_1, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n567, new_n568, new_n569_1, new_n571,
    new_n573_1, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585_1, new_n586, new_n587,
    new_n588_1, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n597, new_n598, new_n599_1, new_n600_1, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607_1, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627_1, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638_1, new_n639, new_n640, new_n641, new_n642, new_n643_1,
    new_n644, new_n645, new_n646_1, new_n647_1, new_n648_1, new_n649_1,
    new_n650, new_n651, new_n652, new_n653_1, new_n654, new_n655_1,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665_1, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675_1, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682_1,
    new_n683_1, new_n684_1, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693_1, new_n694,
    new_n695_1, new_n696, new_n697, new_n698, new_n699_1, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712_1, new_n713, new_n714,
    new_n715_1, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724_1, new_n725_1, new_n726, new_n727,
    new_n728, new_n729_1, new_n730, new_n731_1, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738_1, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747_1,
    new_n748_1, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759_1, new_n760,
    new_n761_1, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770_1, new_n771, new_n772, new_n773_1,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788_1,
    new_n789, new_n790_1, new_n791, new_n792_1, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801_1,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813_1, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823_1, new_n824_1, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836_1, new_n837, new_n838, new_n839_1, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846_1, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858_1, new_n859, new_n860, new_n861, new_n862_1,
    new_n863, new_n864, new_n865_1, new_n866, new_n867_1, new_n868,
    new_n869, new_n870_1, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882_1,
    new_n883_1, new_n884, new_n885, new_n886, new_n887, new_n888_1,
    new_n889, new_n890, new_n891_1, new_n892_1, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902_1, new_n903, new_n904, new_n905_1, new_n906_1, new_n908,
    new_n909, new_n910, new_n911, new_n912_1, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927_1, new_n928, new_n929,
    new_n930, new_n931_1, new_n932, new_n933, new_n934, new_n935_1,
    new_n937, new_n938, new_n940, new_n941, new_n942_1, new_n943, new_n945,
    new_n947, new_n950, new_n951, new_n952_1, new_n953_1, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961_1,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968_1,
    new_n969, new_n970, new_n971, new_n972, new_n975, new_n976, new_n977,
    new_n978, new_n979_1, new_n980_1, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989_1, new_n990,
    new_n991_1, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000_1, new_n1001, new_n1002, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012_1,
    new_n1013, new_n1014, new_n1015_1, new_n1016_1, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025_1, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030_1,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062_1, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067_1, new_n1068_1, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1098, new_n1101, new_n1102, new_n1103_1, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113_1, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119_1, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135_1, new_n1136,
    new_n1137, new_n1138_1, new_n1139, new_n1140_1, new_n1141, new_n1142_1,
    new_n1143, new_n1144, new_n1145_1, new_n1146, new_n1147, new_n1148,
    new_n1149_1, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161_1, new_n1162_1, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172_1,
    new_n1173, new_n1174, new_n1175_1, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183_1, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191_1,
    new_n1192, new_n1193, new_n1194_1, new_n1195, new_n1196, new_n1199_1,
    new_n1201_1, new_n1202_1, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1220, new_n1221, new_n1222_1, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234_1, new_n1235_1, new_n1236, new_n1237_1,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249_1,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255_1,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260_1, new_n1261,
    new_n1262, new_n1263_1, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277_1, new_n1278_1, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283_1, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296_1, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305_1, new_n1306, new_n1307, new_n1308, new_n1312,
    new_n1313, new_n1314, new_n1315_1, new_n1316, new_n1317, new_n1320,
    new_n1322, new_n1323, new_n1326, new_n1327, new_n1329, new_n1331,
    new_n1332_1, new_n1333, new_n1334, new_n1336, new_n1338_1, new_n1339,
    new_n1340_1, new_n1341_1, new_n1342, new_n1343, new_n1344, new_n1346,
    new_n1347_1, new_n1348_1, new_n1349_1, new_n1350, new_n1351_1,
    new_n1352, new_n1353, new_n1354, new_n1355, new_n1356, new_n1357,
    new_n1358, new_n1359, new_n1360, new_n1363_1, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369_1, new_n1370, new_n1371, new_n1373,
    new_n1375, new_n1378, new_n1379, new_n1380, new_n1381_1, new_n1382,
    new_n1384, new_n1385_1, new_n1389, new_n1391, new_n1392, new_n1393_1,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399_1,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407_1, new_n1408, new_n1409, new_n1410, new_n1411,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1422_1, new_n1424,
    new_n1425_1, new_n1426_1, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435_1, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440_1, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453_1, new_n1454,
    new_n1455, new_n1456, new_n1457_1, new_n1458, new_n1459, new_n1460_1,
    new_n1461_1, new_n1462, new_n1463_1, new_n1464, new_n1465, new_n1466,
    new_n1467, new_n1468, new_n1470_1, new_n1471, new_n1472, new_n1473,
    new_n1474, new_n1475, new_n1476, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481_1, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1487, new_n1489, new_n1490, new_n1491, new_n1492, new_n1493,
    new_n1494, new_n1495_1, new_n1496, new_n1497, new_n1498_1, new_n1499,
    new_n1500, new_n1501_1, new_n1502_1, new_n1503, new_n1504, new_n1505,
    new_n1506, new_n1507_1, new_n1508, new_n1509, new_n1510, new_n1511,
    new_n1512, new_n1513, new_n1514, new_n1515, new_n1516, new_n1517,
    new_n1518, new_n1519, new_n1520, new_n1521, new_n1522, new_n1523,
    new_n1524, new_n1525_1, new_n1526, new_n1527_1, new_n1528, new_n1529,
    new_n1530_1, new_n1531, new_n1532, new_n1533, new_n1534, new_n1535_1,
    new_n1536, new_n1537_1, new_n1538, new_n1539, new_n1540, new_n1541,
    new_n1542, new_n1543, new_n1544_1, new_n1545, new_n1546, new_n1547,
    new_n1548, new_n1549, new_n1550, new_n1551, new_n1552, new_n1553,
    new_n1554, new_n1555, new_n1556_1, new_n1557, new_n1558, new_n1559,
    new_n1560, new_n1561, new_n1562, new_n1563, new_n1564, new_n1565,
    new_n1566, new_n1567, new_n1568, new_n1569, new_n1570, new_n1571,
    new_n1572, new_n1573, new_n1574, new_n1575, new_n1576, new_n1577,
    new_n1578, new_n1579, new_n1580, new_n1581, new_n1582, new_n1583,
    new_n1584, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595_1,
    new_n1596, new_n1597_1, new_n1598, new_n1599, new_n1600_1, new_n1601_1,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613_1,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622_1, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1629_1, new_n1630, new_n1631,
    new_n1633_1, new_n1636, new_n1637, new_n1638, new_n1639, new_n1640,
    new_n1641, new_n1642_1, new_n1643_1, new_n1644, new_n1645, new_n1650,
    new_n1653, new_n1655, new_n1657_1, new_n1658, new_n1659, new_n1660_1,
    new_n1661, new_n1663, new_n1668, new_n1669, new_n1670, new_n1671,
    new_n1672, new_n1673, new_n1674, new_n1675_1, new_n1676, new_n1677_1,
    new_n1678_1, new_n1679, new_n1680, new_n1681, new_n1682, new_n1683_1,
    new_n1684, new_n1685, new_n1686_1, new_n1687, new_n1688_1, new_n1689,
    new_n1690_1, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1703, new_n1704,
    new_n1706, new_n1711, new_n1712, new_n1713, new_n1714, new_n1715,
    new_n1716, new_n1717, new_n1719, new_n1721_1, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1727_1, new_n1729_1, new_n1731_1, new_n1734,
    new_n1737_1, new_n1739, new_n1740, new_n1741, new_n1742, new_n1743_1,
    new_n1744, new_n1745, new_n1746_1, new_n1748, new_n1750, new_n1751,
    new_n1752, new_n1753, new_n1754, new_n1755, new_n1756, new_n1757_1,
    new_n1758, new_n1759, new_n1760, new_n1761, new_n1762, new_n1763_1,
    new_n1764_1, new_n1765, new_n1766, new_n1767, new_n1768, new_n1769,
    new_n1770, new_n1771, new_n1772, new_n1773, new_n1774, new_n1775,
    new_n1777, new_n1778, new_n1779, new_n1780, new_n1784, new_n1785,
    new_n1786, new_n1788, new_n1791, new_n1793, new_n1794, new_n1796,
    new_n1798, new_n1799, new_n1800, new_n1801, new_n1802, new_n1803,
    new_n1805, new_n1811, new_n1812, new_n1813, new_n1814, new_n1815,
    new_n1816, new_n1819, new_n1824, new_n1825, new_n1826, new_n1827,
    new_n1828, new_n1830, new_n1831, new_n1832, new_n1834, new_n1835,
    new_n1838, new_n1839, new_n1841, new_n1842, new_n1843, new_n1844,
    new_n1845, new_n1846, new_n1847, new_n1848, new_n1849, new_n1851,
    new_n1854, new_n1856, new_n1857, new_n1863, new_n1865, new_n1866,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1873, new_n1874,
    new_n1875, new_n1878, new_n1880, new_n1882, new_n1884, new_n1885,
    new_n1887, new_n1888, new_n1890, new_n1892, new_n1896, new_n1902,
    new_n1903, new_n1904, new_n1905, new_n1909, new_n1911, new_n1914,
    new_n1917, new_n1923, new_n1924, new_n1927, new_n1928, new_n1929,
    new_n1933, new_n1942;
  nor_4  g0000(.A(n1643), .B(n36), .Y(new_n276_1));
  xor_3  g0001(.A(n1643), .B(n36), .Y(new_n277_1));
  not_3  g0002(.A(new_n277_1), .Y(new_n278));
  nor_4  g0003(.A(n788), .B(n555), .Y(new_n279));
  not_3  g0004(.A(new_n279), .Y(new_n280));
  xnor_3 g0005(.A(n788), .B(n555), .Y(new_n281));
  not_3  g0006(.A(new_n281), .Y(new_n282));
  nor_4  g0007(.A(n747), .B(n353), .Y(new_n283));
  not_3  g0008(.A(new_n283), .Y(new_n284));
  nand_4 g0009(.A(n747), .B(n353), .Y(new_n285));
  not_3  g0010(.A(new_n285), .Y(new_n286));
  nor_4  g0011(.A(new_n286), .B(new_n283), .Y(new_n287));
  nor_4  g0012(.A(n952), .B(n329), .Y(new_n288));
  not_3  g0013(.A(new_n288), .Y(new_n289));
  nand_4 g0014(.A(n1145), .B(n931), .Y(new_n290_1));
  xnor_3 g0015(.A(n952), .B(n329), .Y(new_n291));
  not_3  g0016(.A(new_n291), .Y(new_n292_1));
  nand_4 g0017(.A(new_n292_1), .B(new_n290_1), .Y(new_n293));
  nand_4 g0018(.A(new_n293), .B(new_n289), .Y(new_n294));
  nand_4 g0019(.A(new_n294), .B(new_n287), .Y(new_n295));
  nand_4 g0020(.A(new_n295), .B(new_n284), .Y(new_n296));
  nand_4 g0021(.A(new_n296), .B(new_n282), .Y(new_n297));
  nand_4 g0022(.A(new_n297), .B(new_n280), .Y(new_n298));
  not_3  g0023(.A(new_n298), .Y(new_n299_1));
  nor_4  g0024(.A(new_n299_1), .B(new_n278), .Y(new_n300));
  nor_4  g0025(.A(new_n300), .B(new_n276_1), .Y(new_n301));
  nand_4 g0026(.A(new_n301), .B(n1501), .Y(new_n302));
  xnor_3 g0027(.A(new_n302), .B(n433), .Y(new_n303_1));
  nand_4 g0028(.A(n1000), .B(n870), .Y(new_n304));
  not_3  g0029(.A(n1000), .Y(new_n305));
  nand_4 g0030(.A(new_n305), .B(n66), .Y(new_n306));
  nand_4 g0031(.A(new_n306), .B(new_n304), .Y(new_n307));
  nand_4 g0032(.A(n1000), .B(n585), .Y(new_n308));
  nand_4 g0033(.A(new_n305), .B(n968), .Y(new_n309));
  nand_4 g0034(.A(new_n309), .B(new_n308), .Y(new_n310));
  nor_4  g0035(.A(new_n310), .B(new_n307), .Y(new_n311));
  nand_4 g0036(.A(n1000), .B(n155), .Y(new_n312));
  not_3  g0037(.A(new_n312), .Y(new_n313));
  not_3  g0038(.A(n1435), .Y(new_n314));
  nor_4  g0039(.A(new_n314), .B(n1000), .Y(new_n315));
  nor_4  g0040(.A(new_n315), .B(new_n313), .Y(new_n316));
  nand_4 g0041(.A(new_n316), .B(new_n311), .Y(new_n317_1));
  nor_4  g0042(.A(n1000), .B(n682), .Y(new_n318));
  nor_4  g0043(.A(n1678), .B(new_n305), .Y(new_n319));
  nor_4  g0044(.A(new_n319), .B(new_n318), .Y(new_n320));
  not_3  g0045(.A(new_n320), .Y(new_n321));
  nor_4  g0046(.A(new_n321), .B(new_n317_1), .Y(new_n322));
  xor_3  g0047(.A(n1597), .B(n682), .Y(new_n323));
  nor_4  g0048(.A(new_n323), .B(n1000), .Y(new_n324));
  xnor_3 g0049(.A(n1678), .B(n607), .Y(new_n325));
  nor_4  g0050(.A(new_n325), .B(new_n305), .Y(new_n326));
  nor_4  g0051(.A(new_n326), .B(new_n324), .Y(new_n327));
  xnor_3 g0052(.A(new_n327), .B(new_n322), .Y(new_n328));
  not_3  g0053(.A(new_n317_1), .Y(new_n329_1));
  nor_4  g0054(.A(new_n320), .B(new_n329_1), .Y(new_n330));
  nor_4  g0055(.A(new_n330), .B(new_n322), .Y(new_n331));
  nor_4  g0056(.A(new_n316), .B(new_n311), .Y(new_n332));
  nor_4  g0057(.A(new_n332), .B(new_n329_1), .Y(new_n333));
  not_3  g0058(.A(new_n333), .Y(new_n334));
  not_3  g0059(.A(new_n308), .Y(new_n335));
  not_3  g0060(.A(n968), .Y(new_n336));
  nor_4  g0061(.A(n1000), .B(new_n336), .Y(new_n337));
  nor_4  g0062(.A(new_n337), .B(new_n335), .Y(new_n338));
  xnor_3 g0063(.A(new_n338), .B(new_n307), .Y(new_n339));
  not_3  g0064(.A(new_n339), .Y(new_n340));
  nand_4 g0065(.A(new_n340), .B(n693), .Y(new_n341));
  not_3  g0066(.A(n693), .Y(new_n342));
  nand_4 g0067(.A(new_n339), .B(new_n342), .Y(new_n343));
  nand_4 g0068(.A(new_n338), .B(n1763), .Y(new_n344));
  not_3  g0069(.A(n1763), .Y(new_n345));
  nand_4 g0070(.A(new_n310), .B(new_n345), .Y(new_n346));
  not_3  g0071(.A(n1530), .Y(new_n347_1));
  nand_4 g0072(.A(n1461), .B(n1000), .Y(new_n348));
  not_3  g0073(.A(new_n348), .Y(new_n349));
  not_3  g0074(.A(n347), .Y(new_n350));
  nor_4  g0075(.A(n1000), .B(new_n350), .Y(new_n351));
  nor_4  g0076(.A(new_n351), .B(new_n349), .Y(new_n352));
  nor_4  g0077(.A(new_n352), .B(new_n347_1), .Y(new_n353_1));
  nand_4 g0078(.A(new_n353_1), .B(new_n346), .Y(new_n354));
  nand_4 g0079(.A(new_n354), .B(new_n344), .Y(new_n355));
  nand_4 g0080(.A(new_n355), .B(new_n343), .Y(new_n356));
  nand_4 g0081(.A(new_n356), .B(new_n341), .Y(new_n357));
  nand_4 g0082(.A(new_n357), .B(new_n334), .Y(new_n358));
  nor_4  g0083(.A(new_n358), .B(new_n331), .Y(new_n359));
  nand_4 g0084(.A(new_n359), .B(new_n328), .Y(new_n360));
  nand_4 g0085(.A(new_n327), .B(new_n322), .Y(new_n361));
  not_3  g0086(.A(n682), .Y(new_n362));
  nor_4  g0087(.A(n1597), .B(n46), .Y(new_n363));
  nand_4 g0088(.A(new_n363), .B(new_n362), .Y(new_n364));
  not_3  g0089(.A(new_n364), .Y(new_n365));
  not_3  g0090(.A(n46), .Y(new_n366));
  nor_4  g0091(.A(n1597), .B(n682), .Y(new_n367));
  nor_4  g0092(.A(new_n367), .B(new_n366), .Y(new_n368));
  nor_4  g0093(.A(new_n368), .B(new_n365), .Y(new_n369));
  nor_4  g0094(.A(new_n369), .B(n1000), .Y(new_n370));
  not_3  g0095(.A(n1678), .Y(new_n371));
  nand_4 g0096(.A(n607), .B(n26), .Y(new_n372_1));
  nor_4  g0097(.A(new_n372_1), .B(new_n371), .Y(new_n373));
  not_3  g0098(.A(n26), .Y(new_n374));
  nand_4 g0099(.A(n1678), .B(n607), .Y(new_n375));
  nand_4 g0100(.A(new_n375), .B(new_n374), .Y(new_n376));
  nand_4 g0101(.A(new_n376), .B(n1000), .Y(new_n377));
  nor_4  g0102(.A(new_n377), .B(new_n373), .Y(new_n378_1));
  nor_4  g0103(.A(new_n378_1), .B(new_n370), .Y(new_n379_1));
  xnor_3 g0104(.A(new_n379_1), .B(new_n361), .Y(new_n380));
  xnor_3 g0105(.A(new_n380), .B(new_n360), .Y(new_n381));
  xnor_3 g0106(.A(new_n381), .B(new_n303_1), .Y(new_n382));
  not_3  g0107(.A(new_n382), .Y(new_n383));
  xnor_3 g0108(.A(new_n359), .B(new_n328), .Y(new_n384));
  xnor_3 g0109(.A(new_n301), .B(n1501), .Y(new_n385));
  nand_4 g0110(.A(new_n385), .B(new_n384), .Y(new_n386));
  not_3  g0111(.A(n1501), .Y(new_n387_1));
  xnor_3 g0112(.A(new_n301), .B(new_n387_1), .Y(new_n388));
  xnor_3 g0113(.A(new_n388), .B(new_n384), .Y(new_n389));
  xnor_3 g0114(.A(new_n358), .B(new_n331), .Y(new_n390));
  xnor_3 g0115(.A(new_n298), .B(new_n277_1), .Y(new_n391_1));
  not_3  g0116(.A(new_n391_1), .Y(new_n392));
  nor_4  g0117(.A(new_n392), .B(new_n390), .Y(new_n393));
  xnor_3 g0118(.A(new_n357), .B(new_n333), .Y(new_n394));
  not_3  g0119(.A(new_n394), .Y(new_n395));
  xnor_3 g0120(.A(new_n296), .B(new_n282), .Y(new_n396));
  not_3  g0121(.A(new_n396), .Y(new_n397));
  nand_4 g0122(.A(new_n397), .B(new_n395), .Y(new_n398));
  xnor_3 g0123(.A(new_n397), .B(new_n394), .Y(new_n399));
  xnor_3 g0124(.A(new_n294), .B(new_n287), .Y(new_n400));
  not_3  g0125(.A(new_n400), .Y(new_n401_1));
  not_3  g0126(.A(new_n290_1), .Y(new_n402_1));
  nor_4  g0127(.A(n1145), .B(n931), .Y(new_n403));
  nor_4  g0128(.A(new_n403), .B(new_n402_1), .Y(new_n404));
  nand_4 g0129(.A(new_n305), .B(n347), .Y(new_n405));
  nand_4 g0130(.A(new_n405), .B(new_n348), .Y(new_n406));
  xnor_3 g0131(.A(new_n406), .B(new_n347_1), .Y(new_n407));
  nand_4 g0132(.A(new_n407), .B(new_n404), .Y(new_n408));
  not_3  g0133(.A(new_n408), .Y(new_n409));
  xnor_3 g0134(.A(new_n291), .B(new_n402_1), .Y(new_n410));
  nor_4  g0135(.A(new_n410), .B(new_n409), .Y(new_n411));
  not_3  g0136(.A(new_n411), .Y(new_n412));
  nor_4  g0137(.A(new_n408), .B(new_n291), .Y(new_n413));
  nand_4 g0138(.A(new_n346), .B(new_n344), .Y(new_n414_1));
  xnor_3 g0139(.A(new_n414_1), .B(new_n353_1), .Y(new_n415));
  nor_4  g0140(.A(new_n415), .B(new_n413), .Y(new_n416_1));
  not_3  g0141(.A(new_n416_1), .Y(new_n417));
  nand_4 g0142(.A(new_n417), .B(new_n412), .Y(new_n418));
  nor_4  g0143(.A(new_n418), .B(new_n401_1), .Y(new_n419));
  nor_4  g0144(.A(new_n416_1), .B(new_n411), .Y(new_n420));
  nor_4  g0145(.A(new_n420), .B(new_n400), .Y(new_n421));
  not_3  g0146(.A(new_n355), .Y(new_n422));
  nand_4 g0147(.A(new_n343), .B(new_n341), .Y(new_n423_1));
  xnor_3 g0148(.A(new_n423_1), .B(new_n422), .Y(new_n424_1));
  nor_4  g0149(.A(new_n424_1), .B(new_n421), .Y(new_n425));
  nor_4  g0150(.A(new_n425), .B(new_n419), .Y(new_n426_1));
  nand_4 g0151(.A(new_n426_1), .B(new_n399), .Y(new_n427));
  nand_4 g0152(.A(new_n427), .B(new_n398), .Y(new_n428));
  xnor_3 g0153(.A(new_n392), .B(new_n390), .Y(new_n429_1));
  nor_4  g0154(.A(new_n429_1), .B(new_n428), .Y(new_n430));
  nor_4  g0155(.A(new_n430), .B(new_n393), .Y(new_n431));
  nand_4 g0156(.A(new_n431), .B(new_n389), .Y(new_n432_1));
  nand_4 g0157(.A(new_n432_1), .B(new_n386), .Y(new_n433_1));
  xor_3  g0158(.A(new_n433_1), .B(new_n383), .Y(n19));
  not_3  g0159(.A(n69), .Y(new_n435));
  not_3  g0160(.A(n402), .Y(new_n436));
  nor_4  g0161(.A(n1381), .B(new_n436), .Y(new_n437));
  nor_4  g0162(.A(new_n437), .B(n870), .Y(new_n438));
  not_3  g0163(.A(n1381), .Y(new_n439));
  nand_4 g0164(.A(new_n439), .B(n402), .Y(new_n440));
  nor_4  g0165(.A(new_n440), .B(n66), .Y(new_n441));
  nor_4  g0166(.A(new_n441), .B(new_n438), .Y(new_n442));
  xnor_3 g0167(.A(new_n442), .B(new_n435), .Y(new_n443));
  not_3  g0168(.A(new_n443), .Y(new_n444_1));
  nor_4  g0169(.A(new_n437), .B(n585), .Y(new_n445));
  nor_4  g0170(.A(new_n440), .B(n968), .Y(new_n446));
  nor_4  g0171(.A(new_n446), .B(new_n445), .Y(new_n447));
  nand_4 g0172(.A(new_n447), .B(n953), .Y(new_n448));
  not_3  g0173(.A(n303), .Y(new_n449));
  not_3  g0174(.A(n1461), .Y(new_n450));
  nand_4 g0175(.A(new_n440), .B(new_n450), .Y(new_n451));
  nand_4 g0176(.A(new_n437), .B(new_n350), .Y(new_n452_1));
  nand_4 g0177(.A(new_n452_1), .B(new_n451), .Y(new_n453));
  nor_4  g0178(.A(new_n453), .B(new_n449), .Y(new_n454));
  not_3  g0179(.A(n953), .Y(new_n455));
  xnor_3 g0180(.A(new_n447), .B(new_n455), .Y(new_n456));
  nand_4 g0181(.A(new_n456), .B(new_n454), .Y(new_n457_1));
  nand_4 g0182(.A(new_n457_1), .B(new_n448), .Y(new_n458));
  xnor_3 g0183(.A(new_n458), .B(new_n444_1), .Y(new_n459));
  nor_4  g0184(.A(new_n459), .B(new_n400), .Y(new_n460_1));
  xnor_3 g0185(.A(new_n458), .B(new_n443), .Y(new_n461));
  nor_4  g0186(.A(new_n461), .B(new_n401_1), .Y(new_n462));
  nor_4  g0187(.A(new_n462), .B(new_n460_1), .Y(new_n463));
  not_3  g0188(.A(new_n463), .Y(new_n464));
  not_3  g0189(.A(new_n404), .Y(new_n465));
  xnor_3 g0190(.A(new_n453), .B(n303), .Y(new_n466));
  not_3  g0191(.A(new_n466), .Y(new_n467));
  nor_4  g0192(.A(new_n467), .B(new_n465), .Y(new_n468));
  nor_4  g0193(.A(new_n468), .B(new_n410), .Y(new_n469_1));
  not_3  g0194(.A(new_n469_1), .Y(new_n470));
  xnor_3 g0195(.A(new_n456), .B(new_n454), .Y(new_n471));
  not_3  g0196(.A(new_n468), .Y(new_n472_1));
  nor_4  g0197(.A(new_n472_1), .B(new_n291), .Y(new_n473));
  nor_4  g0198(.A(new_n473), .B(new_n469_1), .Y(new_n474));
  nand_4 g0199(.A(new_n474), .B(new_n471), .Y(new_n475));
  nand_4 g0200(.A(new_n475), .B(new_n470), .Y(new_n476_1));
  xor_3  g0201(.A(new_n476_1), .B(new_n464), .Y(n33));
  not_3  g0202(.A(n247), .Y(new_n478));
  nor_4  g0203(.A(n607), .B(n26), .Y(new_n479));
  nand_4 g0204(.A(new_n479), .B(new_n478), .Y(new_n480));
  xor_3  g0205(.A(new_n480), .B(n1642), .Y(new_n481));
  nor_4  g0206(.A(new_n481), .B(new_n439), .Y(new_n482_1));
  not_3  g0207(.A(n1527), .Y(new_n483));
  nand_4 g0208(.A(new_n483), .B(new_n366), .Y(new_n484));
  nor_4  g0209(.A(new_n484), .B(n379), .Y(new_n485));
  not_3  g0210(.A(n379), .Y(new_n486));
  nor_4  g0211(.A(n1527), .B(n46), .Y(new_n487));
  nor_4  g0212(.A(new_n487), .B(new_n486), .Y(new_n488_1));
  nor_4  g0213(.A(new_n488_1), .B(new_n436), .Y(new_n489));
  not_3  g0214(.A(new_n489), .Y(new_n490));
  nor_4  g0215(.A(new_n490), .B(new_n485), .Y(new_n491));
  not_3  g0216(.A(n1642), .Y(new_n492));
  nor_4  g0217(.A(new_n492), .B(n1381), .Y(new_n493_1));
  nor_4  g0218(.A(new_n493_1), .B(new_n437), .Y(new_n494));
  nor_4  g0219(.A(new_n494), .B(new_n491), .Y(new_n495));
  nor_4  g0220(.A(new_n495), .B(new_n482_1), .Y(new_n496));
  not_3  g0221(.A(new_n496), .Y(new_n497));
  xor_3  g0222(.A(new_n479), .B(new_n478), .Y(new_n498_1));
  nor_4  g0223(.A(new_n498_1), .B(new_n439), .Y(new_n499));
  nand_4 g0224(.A(n1527), .B(n46), .Y(new_n500));
  nand_4 g0225(.A(new_n500), .B(n402), .Y(new_n501));
  nor_4  g0226(.A(new_n501), .B(new_n487), .Y(new_n502));
  nor_4  g0227(.A(n1381), .B(new_n478), .Y(new_n503));
  nor_4  g0228(.A(new_n503), .B(new_n437), .Y(new_n504));
  nor_4  g0229(.A(new_n504), .B(new_n502), .Y(new_n505));
  nor_4  g0230(.A(new_n505), .B(new_n499), .Y(new_n506));
  nor_4  g0231(.A(new_n437), .B(n1678), .Y(new_n507));
  nor_4  g0232(.A(new_n440), .B(n682), .Y(new_n508));
  nor_4  g0233(.A(new_n508), .B(new_n507), .Y(new_n509));
  nor_4  g0234(.A(new_n509), .B(n1643), .Y(new_n510_1));
  not_3  g0235(.A(new_n510_1), .Y(new_n511));
  xor_3  g0236(.A(new_n509), .B(n1643), .Y(new_n512));
  not_3  g0237(.A(n555), .Y(new_n513));
  nor_4  g0238(.A(new_n437), .B(n155), .Y(new_n514));
  nor_4  g0239(.A(new_n440), .B(n1435), .Y(new_n515));
  nor_4  g0240(.A(new_n515), .B(new_n514), .Y(new_n516));
  not_3  g0241(.A(new_n516), .Y(new_n517_1));
  nor_4  g0242(.A(new_n517_1), .B(new_n513), .Y(new_n518));
  nor_4  g0243(.A(new_n442), .B(n353), .Y(new_n519));
  not_3  g0244(.A(new_n519), .Y(new_n520));
  xor_3  g0245(.A(new_n442), .B(n353), .Y(new_n521));
  nor_4  g0246(.A(new_n447), .B(n952), .Y(new_n522_1));
  not_3  g0247(.A(new_n522_1), .Y(new_n523));
  not_3  g0248(.A(n1145), .Y(new_n524));
  nor_4  g0249(.A(new_n453), .B(new_n524), .Y(new_n525));
  not_3  g0250(.A(new_n525), .Y(new_n526));
  xor_3  g0251(.A(new_n447), .B(n952), .Y(new_n527));
  nand_4 g0252(.A(new_n527), .B(new_n526), .Y(new_n528));
  nand_4 g0253(.A(new_n528), .B(new_n523), .Y(new_n529));
  nand_4 g0254(.A(new_n529), .B(new_n521), .Y(new_n530));
  nand_4 g0255(.A(new_n530), .B(new_n520), .Y(new_n531));
  xor_3  g0256(.A(new_n516), .B(n555), .Y(new_n532_1));
  not_3  g0257(.A(new_n532_1), .Y(new_n533));
  nor_4  g0258(.A(new_n533), .B(new_n531), .Y(new_n534_1));
  nor_4  g0259(.A(new_n534_1), .B(new_n518), .Y(new_n535));
  nand_4 g0260(.A(new_n535), .B(new_n512), .Y(new_n536));
  nand_4 g0261(.A(new_n536), .B(new_n511), .Y(new_n537));
  nand_4 g0262(.A(n1381), .B(n607), .Y(new_n538));
  not_3  g0263(.A(new_n538), .Y(new_n539));
  nor_4  g0264(.A(n1597), .B(new_n436), .Y(new_n540));
  nor_4  g0265(.A(n607), .B(n402), .Y(new_n541_1));
  nor_4  g0266(.A(new_n541_1), .B(new_n540), .Y(new_n542));
  nor_4  g0267(.A(new_n542), .B(n1381), .Y(new_n543));
  nor_4  g0268(.A(new_n543), .B(new_n539), .Y(new_n544));
  not_3  g0269(.A(new_n544), .Y(new_n545));
  nor_4  g0270(.A(new_n545), .B(new_n537), .Y(new_n546));
  nand_4 g0271(.A(n402), .B(n46), .Y(new_n547_1));
  not_3  g0272(.A(new_n547_1), .Y(new_n548));
  nor_4  g0273(.A(n402), .B(n26), .Y(new_n549_1));
  nor_4  g0274(.A(new_n549_1), .B(new_n548), .Y(new_n550));
  nor_4  g0275(.A(new_n550), .B(n1381), .Y(new_n551));
  not_3  g0276(.A(new_n372_1), .Y(new_n552));
  nor_4  g0277(.A(new_n479), .B(new_n552), .Y(new_n553));
  not_3  g0278(.A(new_n553), .Y(new_n554));
  nor_4  g0279(.A(new_n554), .B(new_n439), .Y(new_n555_1));
  nor_4  g0280(.A(new_n555_1), .B(new_n551), .Y(new_n556));
  nand_4 g0281(.A(new_n556), .B(new_n546), .Y(new_n557_1));
  nor_4  g0282(.A(new_n557_1), .B(new_n506), .Y(new_n558));
  nor_4  g0283(.A(new_n558), .B(new_n497), .Y(new_n559_1));
  nand_4 g0284(.A(new_n558), .B(new_n497), .Y(new_n560));
  not_3  g0285(.A(new_n560), .Y(new_n561));
  nor_4  g0286(.A(new_n561), .B(new_n559_1), .Y(n1731));
  not_3  g0287(.A(new_n506), .Y(new_n563));
  not_3  g0288(.A(new_n557_1), .Y(new_n564));
  nor_4  g0289(.A(new_n564), .B(new_n563), .Y(new_n565));
  nor_4  g0290(.A(new_n565), .B(new_n558), .Y(n1138));
  not_3  g0291(.A(new_n556), .Y(new_n567));
  not_3  g0292(.A(new_n537), .Y(new_n568));
  nor_4  g0293(.A(new_n544), .B(new_n568), .Y(new_n569_1));
  nor_4  g0294(.A(new_n569_1), .B(new_n546), .Y(n1727));
  not_3  g0295(.A(new_n527), .Y(new_n571));
  xor_3  g0296(.A(new_n571), .B(new_n526), .Y(n1457));
  nand_4 g0297(.A(new_n453), .B(new_n524), .Y(new_n573_1));
  and_4  g0298(.A(new_n573_1), .B(new_n526), .Y(n1183));
  nor_4  g0299(.A(n1183), .B(n1457), .Y(new_n575));
  not_3  g0300(.A(new_n530), .Y(new_n576));
  nor_4  g0301(.A(new_n529), .B(new_n521), .Y(new_n577));
  nor_4  g0302(.A(new_n577), .B(new_n576), .Y(new_n578));
  nand_4 g0303(.A(new_n578), .B(new_n575), .Y(new_n579));
  not_3  g0304(.A(new_n531), .Y(new_n580));
  nor_4  g0305(.A(new_n532_1), .B(new_n580), .Y(new_n581));
  nor_4  g0306(.A(new_n581), .B(new_n534_1), .Y(n1721));
  nor_4  g0307(.A(n1721), .B(new_n579), .Y(new_n583));
  not_3  g0308(.A(new_n536), .Y(new_n584));
  nor_4  g0309(.A(new_n535), .B(new_n512), .Y(new_n585_1));
  nor_4  g0310(.A(new_n585_1), .B(new_n584), .Y(new_n586));
  nor_4  g0311(.A(new_n586), .B(new_n583), .Y(new_n587));
  nand_4 g0312(.A(new_n587), .B(n1727), .Y(new_n588_1));
  nor_4  g0313(.A(new_n588_1), .B(new_n567), .Y(new_n589));
  nand_4 g0314(.A(new_n589), .B(n1138), .Y(new_n590));
  not_3  g0315(.A(new_n590), .Y(new_n591));
  nor_4  g0316(.A(new_n591), .B(n1731), .Y(new_n592));
  nor_4  g0317(.A(new_n590), .B(new_n496), .Y(new_n593));
  nor_4  g0318(.A(new_n593), .B(new_n592), .Y(n44));
  not_3  g0319(.A(new_n407), .Y(new_n595));
  xor_3  g0320(.A(new_n595), .B(new_n465), .Y(n55));
  not_3  g0321(.A(n1332), .Y(new_n597));
  nor_4  g0322(.A(n1707), .B(n1643), .Y(new_n598));
  not_3  g0323(.A(new_n598), .Y(new_n599_1));
  xor_3  g0324(.A(n1707), .B(n1643), .Y(new_n600_1));
  nor_4  g0325(.A(n1140), .B(n555), .Y(new_n601));
  not_3  g0326(.A(new_n601), .Y(new_n602));
  xor_3  g0327(.A(n1140), .B(n555), .Y(new_n603));
  nor_4  g0328(.A(n1351), .B(n353), .Y(new_n604));
  not_3  g0329(.A(new_n604), .Y(new_n605));
  xor_3  g0330(.A(n1351), .B(n353), .Y(new_n606));
  nor_4  g0331(.A(n952), .B(n729), .Y(new_n607_1));
  nand_4 g0332(.A(n1145), .B(n684), .Y(new_n608));
  not_3  g0333(.A(new_n608), .Y(new_n609));
  nand_4 g0334(.A(n952), .B(n729), .Y(new_n610));
  not_3  g0335(.A(new_n610), .Y(new_n611));
  nor_4  g0336(.A(new_n611), .B(new_n607_1), .Y(new_n612));
  not_3  g0337(.A(new_n612), .Y(new_n613));
  nor_4  g0338(.A(new_n613), .B(new_n609), .Y(new_n614));
  nor_4  g0339(.A(new_n614), .B(new_n607_1), .Y(new_n615));
  not_3  g0340(.A(new_n615), .Y(new_n616));
  nand_4 g0341(.A(new_n616), .B(new_n606), .Y(new_n617));
  nand_4 g0342(.A(new_n617), .B(new_n605), .Y(new_n618));
  nand_4 g0343(.A(new_n618), .B(new_n603), .Y(new_n619));
  nand_4 g0344(.A(new_n619), .B(new_n602), .Y(new_n620));
  nand_4 g0345(.A(new_n620), .B(new_n600_1), .Y(new_n621));
  nand_4 g0346(.A(new_n621), .B(new_n599_1), .Y(new_n622));
  nor_4  g0347(.A(new_n622), .B(new_n597), .Y(new_n623));
  nand_4 g0348(.A(new_n623), .B(n391), .Y(new_n624));
  xnor_3 g0349(.A(new_n624), .B(n1544), .Y(new_n625));
  nand_4 g0350(.A(n607), .B(n266), .Y(new_n626));
  not_3  g0351(.A(new_n626), .Y(new_n627_1));
  nor_4  g0352(.A(n1597), .B(n266), .Y(new_n628));
  nor_4  g0353(.A(new_n628), .B(new_n627_1), .Y(new_n629));
  not_3  g0354(.A(new_n629), .Y(new_n630));
  nand_4 g0355(.A(n266), .B(n155), .Y(new_n631));
  not_3  g0356(.A(n266), .Y(new_n632));
  nand_4 g0357(.A(n1435), .B(new_n632), .Y(new_n633));
  nand_4 g0358(.A(new_n633), .B(new_n631), .Y(new_n634));
  nand_4 g0359(.A(n870), .B(n266), .Y(new_n635));
  nand_4 g0360(.A(new_n632), .B(n66), .Y(new_n636));
  nand_4 g0361(.A(new_n636), .B(new_n635), .Y(new_n637));
  nor_4  g0362(.A(new_n637), .B(new_n634), .Y(new_n638_1));
  nand_4 g0363(.A(n1678), .B(n266), .Y(new_n639));
  nand_4 g0364(.A(n682), .B(new_n632), .Y(new_n640));
  nand_4 g0365(.A(new_n640), .B(new_n639), .Y(new_n641));
  not_3  g0366(.A(new_n641), .Y(new_n642));
  nand_4 g0367(.A(new_n642), .B(new_n638_1), .Y(new_n643_1));
  nor_4  g0368(.A(new_n643_1), .B(new_n630), .Y(new_n644));
  nor_4  g0369(.A(new_n632), .B(n26), .Y(new_n645));
  not_3  g0370(.A(new_n645), .Y(new_n646_1));
  xor_3  g0371(.A(n1597), .B(n46), .Y(new_n647_1));
  nand_4 g0372(.A(new_n647_1), .B(new_n632), .Y(new_n648_1));
  nand_4 g0373(.A(new_n648_1), .B(new_n646_1), .Y(new_n649_1));
  xnor_3 g0374(.A(new_n649_1), .B(new_n644), .Y(new_n650));
  xnor_3 g0375(.A(new_n643_1), .B(new_n629), .Y(new_n651));
  xor_3  g0376(.A(new_n641), .B(new_n638_1), .Y(new_n652));
  xnor_3 g0377(.A(new_n637), .B(new_n634), .Y(new_n653_1));
  nand_4 g0378(.A(new_n653_1), .B(n223), .Y(new_n654));
  not_3  g0379(.A(new_n654), .Y(new_n655_1));
  nor_4  g0380(.A(new_n653_1), .B(n223), .Y(new_n656));
  nor_4  g0381(.A(new_n656), .B(new_n655_1), .Y(new_n657));
  not_3  g0382(.A(n444), .Y(new_n658));
  nor_4  g0383(.A(new_n637), .B(new_n658), .Y(new_n659));
  not_3  g0384(.A(new_n659), .Y(new_n660));
  nand_4 g0385(.A(n585), .B(n266), .Y(new_n661));
  nand_4 g0386(.A(n968), .B(new_n632), .Y(new_n662));
  nand_4 g0387(.A(new_n662), .B(new_n661), .Y(new_n663));
  nor_4  g0388(.A(new_n663), .B(n472), .Y(new_n664));
  not_3  g0389(.A(n801), .Y(new_n665_1));
  nand_4 g0390(.A(n1461), .B(n266), .Y(new_n666));
  not_3  g0391(.A(new_n666), .Y(new_n667));
  nor_4  g0392(.A(new_n350), .B(n266), .Y(new_n668));
  nor_4  g0393(.A(new_n668), .B(new_n667), .Y(new_n669));
  nor_4  g0394(.A(new_n669), .B(new_n665_1), .Y(new_n670));
  not_3  g0395(.A(n472), .Y(new_n671));
  not_3  g0396(.A(new_n661), .Y(new_n672));
  nor_4  g0397(.A(new_n336), .B(n266), .Y(new_n673));
  nor_4  g0398(.A(new_n673), .B(new_n672), .Y(new_n674));
  xnor_3 g0399(.A(new_n674), .B(new_n671), .Y(new_n675_1));
  nor_4  g0400(.A(new_n675_1), .B(new_n670), .Y(new_n676));
  nor_4  g0401(.A(new_n676), .B(new_n664), .Y(new_n677));
  xnor_3 g0402(.A(new_n637), .B(new_n658), .Y(new_n678));
  not_3  g0403(.A(new_n678), .Y(new_n679));
  nand_4 g0404(.A(new_n679), .B(new_n677), .Y(new_n680));
  nand_4 g0405(.A(new_n680), .B(new_n660), .Y(new_n681));
  nand_4 g0406(.A(new_n681), .B(new_n657), .Y(new_n682_1));
  nand_4 g0407(.A(new_n682_1), .B(new_n654), .Y(new_n683_1));
  nand_4 g0408(.A(new_n683_1), .B(new_n652), .Y(new_n684_1));
  nor_4  g0409(.A(new_n684_1), .B(new_n651), .Y(new_n685));
  nand_4 g0410(.A(new_n685), .B(new_n650), .Y(new_n686));
  not_3  g0411(.A(new_n644), .Y(new_n687));
  xor_3  g0412(.A(n1597), .B(new_n366), .Y(new_n688));
  nor_4  g0413(.A(new_n688), .B(n266), .Y(new_n689));
  nor_4  g0414(.A(new_n689), .B(new_n645), .Y(new_n690));
  nor_4  g0415(.A(new_n690), .B(new_n687), .Y(new_n691));
  not_3  g0416(.A(n1597), .Y(new_n692));
  nand_4 g0417(.A(new_n487), .B(new_n692), .Y(new_n693_1));
  not_3  g0418(.A(new_n693_1), .Y(new_n694));
  nor_4  g0419(.A(new_n363), .B(new_n483), .Y(new_n695_1));
  nor_4  g0420(.A(new_n695_1), .B(new_n694), .Y(new_n696));
  nand_4 g0421(.A(new_n696), .B(new_n632), .Y(new_n697));
  not_3  g0422(.A(new_n697), .Y(new_n698));
  nor_4  g0423(.A(new_n632), .B(n247), .Y(new_n699_1));
  nor_4  g0424(.A(new_n699_1), .B(new_n698), .Y(new_n700));
  not_3  g0425(.A(new_n700), .Y(new_n701));
  nor_4  g0426(.A(new_n701), .B(new_n691), .Y(new_n702));
  nand_4 g0427(.A(new_n649_1), .B(new_n644), .Y(new_n703));
  nor_4  g0428(.A(new_n700), .B(new_n703), .Y(new_n704));
  nor_4  g0429(.A(new_n704), .B(new_n702), .Y(new_n705));
  xnor_3 g0430(.A(new_n705), .B(new_n686), .Y(new_n706));
  xnor_3 g0431(.A(new_n706), .B(new_n625), .Y(new_n707));
  not_3  g0432(.A(new_n707), .Y(new_n708));
  not_3  g0433(.A(n391), .Y(new_n709));
  xnor_3 g0434(.A(new_n623), .B(new_n709), .Y(new_n710));
  xnor_3 g0435(.A(new_n649_1), .B(new_n687), .Y(new_n711));
  xnor_3 g0436(.A(new_n685), .B(new_n711), .Y(new_n712_1));
  nor_4  g0437(.A(new_n712_1), .B(new_n710), .Y(new_n713));
  not_3  g0438(.A(new_n713), .Y(new_n714));
  xnor_3 g0439(.A(new_n684_1), .B(new_n651), .Y(new_n715_1));
  not_3  g0440(.A(new_n715_1), .Y(new_n716));
  xnor_3 g0441(.A(new_n622), .B(n1332), .Y(new_n717));
  nor_4  g0442(.A(new_n717), .B(new_n716), .Y(new_n718));
  not_3  g0443(.A(new_n718), .Y(new_n719));
  xnor_3 g0444(.A(new_n717), .B(new_n715_1), .Y(new_n720));
  xnor_3 g0445(.A(new_n683_1), .B(new_n652), .Y(new_n721));
  xnor_3 g0446(.A(new_n620), .B(new_n600_1), .Y(new_n722));
  not_3  g0447(.A(new_n722), .Y(new_n723));
  nand_4 g0448(.A(new_n723), .B(new_n721), .Y(new_n724_1));
  xnor_3 g0449(.A(new_n722), .B(new_n721), .Y(new_n725_1));
  xnor_3 g0450(.A(new_n653_1), .B(n223), .Y(new_n726));
  not_3  g0451(.A(new_n664), .Y(new_n727));
  nand_4 g0452(.A(n347), .B(new_n632), .Y(new_n728));
  nand_4 g0453(.A(new_n728), .B(new_n666), .Y(new_n729_1));
  nand_4 g0454(.A(new_n729_1), .B(n801), .Y(new_n730));
  xnor_3 g0455(.A(new_n674), .B(n472), .Y(new_n731_1));
  nand_4 g0456(.A(new_n731_1), .B(new_n730), .Y(new_n732));
  nand_4 g0457(.A(new_n732), .B(new_n727), .Y(new_n733));
  nor_4  g0458(.A(new_n678), .B(new_n733), .Y(new_n734));
  nor_4  g0459(.A(new_n734), .B(new_n659), .Y(new_n735));
  xnor_3 g0460(.A(new_n735), .B(new_n726), .Y(new_n736));
  xnor_3 g0461(.A(new_n618), .B(new_n603), .Y(new_n737));
  not_3  g0462(.A(new_n737), .Y(new_n738_1));
  nand_4 g0463(.A(new_n738_1), .B(new_n736), .Y(new_n739));
  xnor_3 g0464(.A(new_n737), .B(new_n736), .Y(new_n740));
  xnor_3 g0465(.A(new_n679), .B(new_n677), .Y(new_n741));
  xnor_3 g0466(.A(new_n615), .B(new_n606), .Y(new_n742));
  nand_4 g0467(.A(new_n742), .B(new_n741), .Y(new_n743));
  nor_4  g0468(.A(new_n612), .B(new_n608), .Y(new_n744));
  not_3  g0469(.A(new_n614), .Y(new_n745));
  nor_4  g0470(.A(n1145), .B(n684), .Y(new_n746));
  nor_4  g0471(.A(new_n746), .B(new_n609), .Y(new_n747_1));
  nor_4  g0472(.A(new_n729_1), .B(n801), .Y(new_n748_1));
  nor_4  g0473(.A(new_n748_1), .B(new_n670), .Y(new_n749));
  nand_4 g0474(.A(new_n749), .B(new_n747_1), .Y(new_n750));
  nand_4 g0475(.A(new_n750), .B(new_n745), .Y(new_n751));
  nor_4  g0476(.A(new_n751), .B(new_n744), .Y(new_n752));
  not_3  g0477(.A(new_n752), .Y(new_n753));
  xnor_3 g0478(.A(new_n731_1), .B(new_n670), .Y(new_n754));
  nor_4  g0479(.A(new_n750), .B(new_n613), .Y(new_n755));
  nor_4  g0480(.A(new_n755), .B(new_n752), .Y(new_n756));
  nand_4 g0481(.A(new_n756), .B(new_n754), .Y(new_n757));
  nand_4 g0482(.A(new_n757), .B(new_n753), .Y(new_n758));
  not_3  g0483(.A(new_n743), .Y(new_n759_1));
  nor_4  g0484(.A(new_n742), .B(new_n741), .Y(new_n760));
  nor_4  g0485(.A(new_n760), .B(new_n759_1), .Y(new_n761_1));
  nand_4 g0486(.A(new_n761_1), .B(new_n758), .Y(new_n762));
  nand_4 g0487(.A(new_n762), .B(new_n743), .Y(new_n763));
  nand_4 g0488(.A(new_n763), .B(new_n740), .Y(new_n764));
  nand_4 g0489(.A(new_n764), .B(new_n739), .Y(new_n765));
  nand_4 g0490(.A(new_n765), .B(new_n725_1), .Y(new_n766));
  nand_4 g0491(.A(new_n766), .B(new_n724_1), .Y(new_n767));
  nand_4 g0492(.A(new_n767), .B(new_n720), .Y(new_n768));
  nand_4 g0493(.A(new_n768), .B(new_n719), .Y(new_n769));
  xnor_3 g0494(.A(new_n685), .B(new_n650), .Y(new_n770_1));
  xnor_3 g0495(.A(new_n770_1), .B(new_n710), .Y(new_n771));
  nand_4 g0496(.A(new_n771), .B(new_n769), .Y(new_n772));
  nand_4 g0497(.A(new_n772), .B(new_n714), .Y(new_n773_1));
  xor_3  g0498(.A(new_n773_1), .B(new_n708), .Y(n56));
  nor_4  g0499(.A(new_n705), .B(new_n686), .Y(new_n775));
  nor_4  g0500(.A(n1642), .B(new_n632), .Y(new_n776));
  not_3  g0501(.A(new_n776), .Y(new_n777));
  xor_3  g0502(.A(new_n693_1), .B(n379), .Y(new_n778));
  nand_4 g0503(.A(new_n778), .B(new_n632), .Y(new_n779));
  nand_4 g0504(.A(new_n779), .B(new_n777), .Y(new_n780));
  xnor_3 g0505(.A(new_n780), .B(new_n704), .Y(new_n781));
  nand_4 g0506(.A(new_n781), .B(new_n775), .Y(new_n782));
  nand_4 g0507(.A(new_n780), .B(new_n704), .Y(new_n783));
  nor_4  g0508(.A(new_n632), .B(n171), .Y(new_n784));
  not_3  g0509(.A(n1263), .Y(new_n785));
  nor_4  g0510(.A(new_n693_1), .B(n379), .Y(new_n786));
  nor_4  g0511(.A(new_n786), .B(new_n785), .Y(new_n787));
  nand_4 g0512(.A(new_n485), .B(new_n785), .Y(new_n788_1));
  nor_4  g0513(.A(new_n788_1), .B(n1597), .Y(new_n789));
  nor_4  g0514(.A(new_n789), .B(new_n787), .Y(new_n790_1));
  nand_4 g0515(.A(new_n790_1), .B(new_n632), .Y(new_n791));
  not_3  g0516(.A(new_n791), .Y(new_n792_1));
  nor_4  g0517(.A(new_n792_1), .B(new_n784), .Y(new_n793));
  nor_4  g0518(.A(new_n793), .B(new_n783), .Y(new_n794));
  nand_4 g0519(.A(new_n701), .B(new_n691), .Y(new_n795));
  xor_3  g0520(.A(new_n693_1), .B(new_n486), .Y(new_n796));
  nor_4  g0521(.A(new_n796), .B(n266), .Y(new_n797));
  nor_4  g0522(.A(new_n797), .B(new_n776), .Y(new_n798));
  nor_4  g0523(.A(new_n798), .B(new_n795), .Y(new_n799));
  not_3  g0524(.A(new_n793), .Y(new_n800));
  nor_4  g0525(.A(new_n800), .B(new_n799), .Y(new_n801_1));
  nor_4  g0526(.A(new_n801_1), .B(new_n794), .Y(new_n802));
  nor_4  g0527(.A(new_n802), .B(new_n782), .Y(new_n803));
  not_3  g0528(.A(new_n794), .Y(new_n804));
  nor_4  g0529(.A(n557), .B(new_n632), .Y(new_n805));
  not_3  g0530(.A(n1422), .Y(new_n806));
  not_3  g0531(.A(new_n788_1), .Y(new_n807));
  nand_4 g0532(.A(new_n807), .B(new_n806), .Y(new_n808));
  nor_4  g0533(.A(new_n808), .B(n1597), .Y(new_n809));
  not_3  g0534(.A(new_n789), .Y(new_n810));
  nand_4 g0535(.A(new_n810), .B(n1422), .Y(new_n811));
  not_3  g0536(.A(new_n811), .Y(new_n812));
  nor_4  g0537(.A(new_n812), .B(new_n809), .Y(new_n813_1));
  nand_4 g0538(.A(new_n813_1), .B(new_n632), .Y(new_n814));
  not_3  g0539(.A(new_n814), .Y(new_n815));
  nor_4  g0540(.A(new_n815), .B(new_n805), .Y(new_n816));
  xor_3  g0541(.A(new_n816), .B(new_n804), .Y(new_n817));
  not_3  g0542(.A(new_n817), .Y(new_n818));
  xor_3  g0543(.A(new_n818), .B(new_n803), .Y(new_n819));
  not_3  g0544(.A(n1544), .Y(new_n820));
  nor_4  g0545(.A(new_n624), .B(new_n820), .Y(new_n821));
  nand_4 g0546(.A(new_n821), .B(n649), .Y(new_n822));
  not_3  g0547(.A(new_n822), .Y(new_n823_1));
  xnor_3 g0548(.A(new_n802), .B(new_n782), .Y(new_n824_1));
  not_3  g0549(.A(new_n824_1), .Y(new_n825));
  nor_4  g0550(.A(new_n825), .B(new_n823_1), .Y(new_n826));
  not_3  g0551(.A(new_n826), .Y(new_n827));
  xor_3  g0552(.A(new_n825), .B(new_n823_1), .Y(new_n828));
  nor_4  g0553(.A(new_n821), .B(n649), .Y(new_n829));
  nor_4  g0554(.A(new_n829), .B(new_n823_1), .Y(new_n830));
  not_3  g0555(.A(new_n781), .Y(new_n831));
  xnor_3 g0556(.A(new_n831), .B(new_n775), .Y(new_n832));
  nor_4  g0557(.A(new_n832), .B(new_n830), .Y(new_n833));
  not_3  g0558(.A(new_n833), .Y(new_n834));
  xnor_3 g0559(.A(new_n832), .B(new_n830), .Y(new_n835));
  not_3  g0560(.A(new_n835), .Y(new_n836_1));
  xnor_3 g0561(.A(new_n700), .B(new_n703), .Y(new_n837));
  xnor_3 g0562(.A(new_n837), .B(new_n686), .Y(new_n838));
  nor_4  g0563(.A(new_n838), .B(new_n625), .Y(new_n839_1));
  not_3  g0564(.A(new_n839_1), .Y(new_n840));
  nand_4 g0565(.A(new_n773_1), .B(new_n707), .Y(new_n841));
  nand_4 g0566(.A(new_n841), .B(new_n840), .Y(new_n842));
  nand_4 g0567(.A(new_n842), .B(new_n836_1), .Y(new_n843));
  nand_4 g0568(.A(new_n843), .B(new_n834), .Y(new_n844));
  nand_4 g0569(.A(new_n844), .B(new_n828), .Y(new_n845));
  nand_4 g0570(.A(new_n845), .B(new_n827), .Y(new_n846_1));
  not_3  g0571(.A(new_n846_1), .Y(new_n847));
  nor_4  g0572(.A(new_n847), .B(new_n819), .Y(new_n848));
  not_3  g0573(.A(new_n819), .Y(new_n849));
  nor_4  g0574(.A(new_n846_1), .B(new_n849), .Y(new_n850));
  nor_4  g0575(.A(new_n850), .B(new_n848), .Y(n67));
  not_3  g0576(.A(new_n390), .Y(new_n852));
  xor_3  g0577(.A(n1643), .B(n469), .Y(new_n853));
  nor_4  g0578(.A(n927), .B(n555), .Y(new_n854));
  not_3  g0579(.A(new_n854), .Y(new_n855));
  xor_3  g0580(.A(n927), .B(n555), .Y(new_n856));
  nor_4  g0581(.A(n655), .B(n353), .Y(new_n857));
  xnor_3 g0582(.A(n655), .B(n353), .Y(new_n858_1));
  nor_4  g0583(.A(n952), .B(n653), .Y(new_n859));
  nand_4 g0584(.A(n1764), .B(n1145), .Y(new_n860));
  not_3  g0585(.A(new_n860), .Y(new_n861));
  nand_4 g0586(.A(n952), .B(n653), .Y(new_n862_1));
  not_3  g0587(.A(new_n862_1), .Y(new_n863));
  nor_4  g0588(.A(new_n863), .B(new_n859), .Y(new_n864));
  not_3  g0589(.A(new_n864), .Y(new_n865_1));
  nor_4  g0590(.A(new_n865_1), .B(new_n861), .Y(new_n866));
  nor_4  g0591(.A(new_n866), .B(new_n859), .Y(new_n867_1));
  nor_4  g0592(.A(new_n867_1), .B(new_n858_1), .Y(new_n868));
  nor_4  g0593(.A(new_n868), .B(new_n857), .Y(new_n869));
  not_3  g0594(.A(new_n869), .Y(new_n870_1));
  nand_4 g0595(.A(new_n870_1), .B(new_n856), .Y(new_n871));
  nand_4 g0596(.A(new_n871), .B(new_n855), .Y(new_n872));
  xnor_3 g0597(.A(new_n872), .B(new_n853), .Y(new_n873));
  nand_4 g0598(.A(new_n873), .B(new_n852), .Y(new_n874));
  not_3  g0599(.A(new_n874), .Y(new_n875));
  nor_4  g0600(.A(new_n873), .B(new_n852), .Y(new_n876));
  nor_4  g0601(.A(new_n876), .B(new_n875), .Y(new_n877));
  xnor_3 g0602(.A(new_n870_1), .B(new_n856), .Y(new_n878));
  nor_4  g0603(.A(new_n878), .B(new_n394), .Y(new_n879));
  not_3  g0604(.A(new_n878), .Y(new_n880));
  nor_4  g0605(.A(new_n880), .B(new_n395), .Y(new_n881));
  nor_4  g0606(.A(new_n881), .B(new_n879), .Y(new_n882_1));
  not_3  g0607(.A(new_n882_1), .Y(new_n883_1));
  nor_4  g0608(.A(new_n864), .B(new_n860), .Y(new_n884));
  not_3  g0609(.A(new_n866), .Y(new_n885));
  nor_4  g0610(.A(n1764), .B(n1145), .Y(new_n886));
  nor_4  g0611(.A(new_n886), .B(new_n861), .Y(new_n887));
  nand_4 g0612(.A(new_n887), .B(new_n407), .Y(new_n888_1));
  nand_4 g0613(.A(new_n888_1), .B(new_n885), .Y(new_n889));
  nor_4  g0614(.A(new_n889), .B(new_n884), .Y(new_n890));
  not_3  g0615(.A(new_n890), .Y(new_n891_1));
  not_3  g0616(.A(new_n415), .Y(new_n892_1));
  nor_4  g0617(.A(new_n888_1), .B(new_n865_1), .Y(new_n893));
  nor_4  g0618(.A(new_n893), .B(new_n890), .Y(new_n894));
  nand_4 g0619(.A(new_n894), .B(new_n892_1), .Y(new_n895));
  nand_4 g0620(.A(new_n895), .B(new_n891_1), .Y(new_n896));
  xnor_3 g0621(.A(new_n867_1), .B(new_n858_1), .Y(new_n897));
  not_3  g0622(.A(new_n897), .Y(new_n898));
  nor_4  g0623(.A(new_n898), .B(new_n896), .Y(new_n899));
  not_3  g0624(.A(new_n899), .Y(new_n900));
  not_3  g0625(.A(new_n424_1), .Y(new_n901));
  xnor_3 g0626(.A(new_n897), .B(new_n896), .Y(new_n902_1));
  nand_4 g0627(.A(new_n902_1), .B(new_n901), .Y(new_n903));
  nand_4 g0628(.A(new_n903), .B(new_n900), .Y(new_n904));
  nor_4  g0629(.A(new_n904), .B(new_n883_1), .Y(new_n905_1));
  nor_4  g0630(.A(new_n905_1), .B(new_n879), .Y(new_n906_1));
  xor_3  g0631(.A(new_n906_1), .B(new_n877), .Y(n74));
  not_3  g0632(.A(n171), .Y(new_n908));
  nor_4  g0633(.A(new_n480), .B(n1642), .Y(new_n909));
  xor_3  g0634(.A(new_n909), .B(new_n908), .Y(new_n910));
  nor_4  g0635(.A(new_n910), .B(new_n439), .Y(new_n911));
  xor_3  g0636(.A(new_n485), .B(new_n785), .Y(new_n912_1));
  not_3  g0637(.A(new_n912_1), .Y(new_n913));
  nor_4  g0638(.A(new_n913), .B(new_n436), .Y(new_n914));
  nor_4  g0639(.A(n402), .B(n171), .Y(new_n915));
  nor_4  g0640(.A(new_n915), .B(n1381), .Y(new_n916));
  not_3  g0641(.A(new_n916), .Y(new_n917));
  nor_4  g0642(.A(new_n917), .B(new_n914), .Y(new_n918));
  nor_4  g0643(.A(new_n918), .B(new_n911), .Y(new_n919));
  nor_4  g0644(.A(new_n919), .B(new_n560), .Y(new_n920));
  xor_3  g0645(.A(new_n788_1), .B(n1422), .Y(new_n921));
  not_3  g0646(.A(new_n921), .Y(new_n922));
  nor_4  g0647(.A(new_n922), .B(new_n436), .Y(new_n923));
  nor_4  g0648(.A(n557), .B(n402), .Y(new_n924));
  nor_4  g0649(.A(new_n924), .B(n1381), .Y(new_n925));
  not_3  g0650(.A(new_n925), .Y(new_n926));
  nor_4  g0651(.A(new_n926), .B(new_n923), .Y(new_n927_1));
  nand_4 g0652(.A(new_n909), .B(new_n908), .Y(new_n928));
  xor_3  g0653(.A(new_n928), .B(n557), .Y(new_n929));
  nor_4  g0654(.A(new_n929), .B(new_n439), .Y(new_n930));
  nor_4  g0655(.A(new_n930), .B(new_n927_1), .Y(new_n931_1));
  not_3  g0656(.A(new_n931_1), .Y(new_n932));
  nor_4  g0657(.A(new_n932), .B(new_n920), .Y(new_n933));
  nand_4 g0658(.A(new_n932), .B(new_n920), .Y(new_n934));
  not_3  g0659(.A(new_n934), .Y(new_n935_1));
  nor_4  g0660(.A(new_n935_1), .B(new_n933), .Y(n156));
  not_3  g0661(.A(new_n919), .Y(new_n937));
  nor_4  g0662(.A(new_n937), .B(new_n561), .Y(new_n938));
  nor_4  g0663(.A(new_n938), .B(new_n920), .Y(n1149));
  nand_4 g0664(.A(n1149), .B(new_n593), .Y(new_n940));
  not_3  g0665(.A(new_n940), .Y(new_n941));
  nor_4  g0666(.A(new_n941), .B(n156), .Y(new_n942_1));
  nor_4  g0667(.A(new_n940), .B(new_n931_1), .Y(new_n943));
  nor_4  g0668(.A(new_n943), .B(new_n942_1), .Y(n106));
  not_3  g0669(.A(new_n588_1), .Y(new_n945));
  xor_3  g0670(.A(new_n556), .B(new_n546), .Y(n1385));
  nor_4  g0671(.A(n1385), .B(new_n945), .Y(new_n947));
  nor_4  g0672(.A(new_n947), .B(new_n589), .Y(n126));
  xnor_3 g0673(.A(new_n765), .B(new_n725_1), .Y(n135));
  nor_4  g0674(.A(new_n641), .B(n1643), .Y(new_n950));
  xor_3  g0675(.A(new_n641), .B(n1643), .Y(new_n951));
  not_3  g0676(.A(new_n634), .Y(new_n952_1));
  nand_4 g0677(.A(new_n952_1), .B(new_n513), .Y(new_n953_1));
  not_3  g0678(.A(n353), .Y(new_n954));
  not_3  g0679(.A(new_n637), .Y(new_n955));
  nand_4 g0680(.A(new_n955), .B(new_n954), .Y(new_n956));
  xor_3  g0681(.A(new_n955), .B(new_n954), .Y(new_n957));
  not_3  g0682(.A(n952), .Y(new_n958));
  nand_4 g0683(.A(new_n674), .B(new_n958), .Y(new_n959));
  nand_4 g0684(.A(new_n729_1), .B(n1145), .Y(new_n960));
  xor_3  g0685(.A(new_n674), .B(new_n958), .Y(new_n961_1));
  nand_4 g0686(.A(new_n961_1), .B(new_n960), .Y(new_n962));
  nand_4 g0687(.A(new_n962), .B(new_n959), .Y(new_n963));
  nand_4 g0688(.A(new_n963), .B(new_n957), .Y(new_n964));
  nand_4 g0689(.A(new_n964), .B(new_n956), .Y(new_n965));
  xor_3  g0690(.A(new_n634), .B(n555), .Y(new_n966));
  nand_4 g0691(.A(new_n966), .B(new_n965), .Y(new_n967));
  nand_4 g0692(.A(new_n967), .B(new_n953_1), .Y(new_n968_1));
  nand_4 g0693(.A(new_n968_1), .B(new_n951), .Y(new_n969));
  not_3  g0694(.A(new_n969), .Y(new_n970));
  nor_4  g0695(.A(new_n970), .B(new_n950), .Y(new_n971));
  nand_4 g0696(.A(new_n971), .B(new_n630), .Y(new_n972));
  xor_3  g0697(.A(new_n972), .B(new_n649_1), .Y(n145));
  xor_3  g0698(.A(new_n404), .B(n347), .Y(n174));
  xnor_3 g0699(.A(new_n388), .B(new_n692), .Y(new_n975));
  not_3  g0700(.A(new_n975), .Y(new_n976));
  nand_4 g0701(.A(new_n391_1), .B(n682), .Y(new_n977));
  xnor_3 g0702(.A(new_n391_1), .B(new_n362), .Y(new_n978));
  nand_4 g0703(.A(new_n396), .B(n1435), .Y(new_n979_1));
  xnor_3 g0704(.A(new_n396), .B(new_n314), .Y(new_n980_1));
  nand_4 g0705(.A(new_n400), .B(n66), .Y(new_n981));
  not_3  g0706(.A(new_n981), .Y(new_n982));
  nor_4  g0707(.A(new_n400), .B(n66), .Y(new_n983));
  nor_4  g0708(.A(new_n983), .B(new_n982), .Y(new_n984));
  nor_4  g0709(.A(new_n410), .B(n968), .Y(new_n985));
  nor_4  g0710(.A(new_n465), .B(new_n350), .Y(new_n986));
  xnor_3 g0711(.A(new_n410), .B(n968), .Y(new_n987));
  nor_4  g0712(.A(new_n987), .B(new_n986), .Y(new_n988));
  nor_4  g0713(.A(new_n988), .B(new_n985), .Y(new_n989_1));
  nand_4 g0714(.A(new_n989_1), .B(new_n984), .Y(new_n990));
  nand_4 g0715(.A(new_n990), .B(new_n981), .Y(new_n991_1));
  nand_4 g0716(.A(new_n991_1), .B(new_n980_1), .Y(new_n992));
  nand_4 g0717(.A(new_n992), .B(new_n979_1), .Y(new_n993));
  nand_4 g0718(.A(new_n993), .B(new_n978), .Y(new_n994));
  nand_4 g0719(.A(new_n994), .B(new_n977), .Y(new_n995));
  xor_3  g0720(.A(new_n995), .B(new_n976), .Y(new_n996));
  xor_3  g0721(.A(new_n993), .B(new_n978), .Y(new_n997));
  not_3  g0722(.A(new_n997), .Y(new_n998));
  xor_3  g0723(.A(new_n989_1), .B(new_n984), .Y(n1426));
  xor_3  g0724(.A(new_n991_1), .B(new_n980_1), .Y(new_n1000_1));
  nor_4  g0725(.A(new_n1000_1), .B(n1426), .Y(new_n1001));
  nand_4 g0726(.A(new_n1001), .B(new_n998), .Y(new_n1002));
  xor_3  g0727(.A(new_n1002), .B(new_n996), .Y(n181));
  nor_4  g0728(.A(new_n421), .B(new_n419), .Y(new_n1004));
  xor_3  g0729(.A(new_n1004), .B(new_n901), .Y(n208));
  nor_4  g0730(.A(new_n637), .B(n213), .Y(new_n1006));
  not_3  g0731(.A(new_n1006), .Y(new_n1007));
  not_3  g0732(.A(n213), .Y(new_n1008));
  nor_4  g0733(.A(new_n955), .B(new_n1008), .Y(new_n1009));
  nor_4  g0734(.A(new_n1009), .B(new_n1006), .Y(new_n1010));
  nor_4  g0735(.A(new_n663), .B(n1743), .Y(new_n1011));
  not_3  g0736(.A(new_n1011), .Y(new_n1012_1));
  not_3  g0737(.A(n600), .Y(new_n1013));
  nor_4  g0738(.A(new_n669), .B(new_n1013), .Y(new_n1014));
  not_3  g0739(.A(new_n1014), .Y(new_n1015_1));
  not_3  g0740(.A(n1743), .Y(new_n1016_1));
  nor_4  g0741(.A(new_n674), .B(new_n1016_1), .Y(new_n1017));
  nor_4  g0742(.A(new_n1017), .B(new_n1011), .Y(new_n1018));
  nand_4 g0743(.A(new_n1018), .B(new_n1015_1), .Y(new_n1019));
  nand_4 g0744(.A(new_n1019), .B(new_n1012_1), .Y(new_n1020));
  nand_4 g0745(.A(new_n1020), .B(new_n1010), .Y(new_n1021));
  nand_4 g0746(.A(new_n1021), .B(new_n1007), .Y(new_n1022));
  nor_4  g0747(.A(new_n1022), .B(new_n952_1), .Y(new_n1023));
  nand_4 g0748(.A(new_n1023), .B(new_n641), .Y(new_n1024));
  xnor_3 g0749(.A(new_n1024), .B(new_n630), .Y(new_n1025_1));
  nor_4  g0750(.A(n1643), .B(n424), .Y(new_n1026));
  not_3  g0751(.A(new_n1026), .Y(new_n1027));
  xor_3  g0752(.A(n1643), .B(n424), .Y(new_n1028));
  nor_4  g0753(.A(n1363), .B(n555), .Y(new_n1029));
  not_3  g0754(.A(new_n1029), .Y(new_n1030_1));
  xor_3  g0755(.A(n1363), .B(n555), .Y(new_n1031));
  nor_4  g0756(.A(n498), .B(n353), .Y(new_n1032));
  not_3  g0757(.A(new_n1032), .Y(new_n1033));
  nand_4 g0758(.A(n498), .B(n353), .Y(new_n1034));
  not_3  g0759(.A(new_n1034), .Y(new_n1035));
  nor_4  g0760(.A(new_n1035), .B(new_n1032), .Y(new_n1036));
  nor_4  g0761(.A(n952), .B(n414), .Y(new_n1037));
  not_3  g0762(.A(new_n1037), .Y(new_n1038));
  nand_4 g0763(.A(n1145), .B(n183), .Y(new_n1039));
  nand_4 g0764(.A(n952), .B(n414), .Y(new_n1040));
  not_3  g0765(.A(new_n1040), .Y(new_n1041));
  nor_4  g0766(.A(new_n1041), .B(new_n1037), .Y(new_n1042));
  nand_4 g0767(.A(new_n1042), .B(new_n1039), .Y(new_n1043));
  nand_4 g0768(.A(new_n1043), .B(new_n1038), .Y(new_n1044));
  nand_4 g0769(.A(new_n1044), .B(new_n1036), .Y(new_n1045));
  nand_4 g0770(.A(new_n1045), .B(new_n1033), .Y(new_n1046));
  nand_4 g0771(.A(new_n1046), .B(new_n1031), .Y(new_n1047));
  nand_4 g0772(.A(new_n1047), .B(new_n1030_1), .Y(new_n1048));
  nand_4 g0773(.A(new_n1048), .B(new_n1028), .Y(new_n1049));
  nand_4 g0774(.A(new_n1049), .B(new_n1027), .Y(new_n1050));
  xnor_3 g0775(.A(new_n1050), .B(n17), .Y(new_n1051));
  xnor_3 g0776(.A(new_n1051), .B(new_n1025_1), .Y(new_n1052));
  not_3  g0777(.A(new_n1052), .Y(new_n1053));
  xnor_3 g0778(.A(new_n1023), .B(new_n642), .Y(new_n1054));
  xnor_3 g0779(.A(new_n1048), .B(new_n1028), .Y(new_n1055));
  nor_4  g0780(.A(new_n1055), .B(new_n1054), .Y(new_n1056));
  xnor_3 g0781(.A(new_n1022), .B(new_n952_1), .Y(new_n1057));
  xnor_3 g0782(.A(new_n1046), .B(new_n1031), .Y(new_n1058));
  not_3  g0783(.A(new_n1058), .Y(new_n1059));
  nand_4 g0784(.A(new_n1059), .B(new_n1057), .Y(new_n1060));
  xnor_3 g0785(.A(new_n1058), .B(new_n1057), .Y(new_n1061));
  xnor_3 g0786(.A(new_n1020), .B(new_n1010), .Y(new_n1062_1));
  not_3  g0787(.A(new_n1062_1), .Y(new_n1063));
  not_3  g0788(.A(new_n1045), .Y(new_n1064));
  nor_4  g0789(.A(new_n1044), .B(new_n1036), .Y(new_n1065));
  nor_4  g0790(.A(new_n1065), .B(new_n1064), .Y(new_n1066));
  nand_4 g0791(.A(new_n1066), .B(new_n1063), .Y(new_n1067_1));
  nor_4  g0792(.A(new_n1042), .B(new_n1039), .Y(new_n1068_1));
  not_3  g0793(.A(new_n1039), .Y(new_n1069));
  nor_4  g0794(.A(n1145), .B(n183), .Y(new_n1070));
  nor_4  g0795(.A(new_n1070), .B(new_n1069), .Y(new_n1071));
  nor_4  g0796(.A(new_n729_1), .B(n600), .Y(new_n1072));
  nor_4  g0797(.A(new_n1072), .B(new_n1014), .Y(new_n1073));
  nand_4 g0798(.A(new_n1073), .B(new_n1071), .Y(new_n1074));
  nand_4 g0799(.A(new_n1074), .B(new_n1043), .Y(new_n1075));
  nor_4  g0800(.A(new_n1075), .B(new_n1068_1), .Y(new_n1076));
  not_3  g0801(.A(new_n1076), .Y(new_n1077));
  xnor_3 g0802(.A(new_n1018), .B(new_n1014), .Y(new_n1078));
  not_3  g0803(.A(new_n1042), .Y(new_n1079));
  nor_4  g0804(.A(new_n1074), .B(new_n1079), .Y(new_n1080));
  nor_4  g0805(.A(new_n1080), .B(new_n1076), .Y(new_n1081));
  nand_4 g0806(.A(new_n1081), .B(new_n1078), .Y(new_n1082));
  nand_4 g0807(.A(new_n1082), .B(new_n1077), .Y(new_n1083));
  xnor_3 g0808(.A(new_n1066), .B(new_n1062_1), .Y(new_n1084));
  nand_4 g0809(.A(new_n1084), .B(new_n1083), .Y(new_n1085));
  nand_4 g0810(.A(new_n1085), .B(new_n1067_1), .Y(new_n1086));
  nand_4 g0811(.A(new_n1086), .B(new_n1061), .Y(new_n1087));
  nand_4 g0812(.A(new_n1087), .B(new_n1060), .Y(new_n1088));
  not_3  g0813(.A(new_n1054), .Y(new_n1089));
  not_3  g0814(.A(new_n1028), .Y(new_n1090));
  xnor_3 g0815(.A(new_n1048), .B(new_n1090), .Y(new_n1091));
  nor_4  g0816(.A(new_n1091), .B(new_n1089), .Y(new_n1092));
  nor_4  g0817(.A(new_n1092), .B(new_n1056), .Y(new_n1093));
  nand_4 g0818(.A(new_n1093), .B(new_n1088), .Y(new_n1094));
  not_3  g0819(.A(new_n1094), .Y(new_n1095));
  nor_4  g0820(.A(new_n1095), .B(new_n1056), .Y(new_n1096));
  xor_3  g0821(.A(new_n1096), .B(new_n1053), .Y(n216));
  not_3  g0822(.A(new_n1084), .Y(new_n1098));
  xor_3  g0823(.A(new_n1098), .B(new_n1083), .Y(n218));
  xnor_3 g0824(.A(new_n844), .B(new_n828), .Y(n231));
  not_3  g0825(.A(n1747), .Y(new_n1101));
  not_3  g0826(.A(n738), .Y(new_n1102));
  not_3  g0827(.A(n17), .Y(new_n1103_1));
  nor_4  g0828(.A(new_n1050), .B(new_n1103_1), .Y(new_n1104));
  nand_4 g0829(.A(new_n1104), .B(n961), .Y(new_n1105));
  nor_4  g0830(.A(new_n1105), .B(new_n1102), .Y(new_n1106));
  not_3  g0831(.A(new_n1106), .Y(new_n1107));
  xor_3  g0832(.A(new_n1107), .B(new_n1101), .Y(new_n1108));
  nor_4  g0833(.A(new_n1024), .B(new_n629), .Y(new_n1109));
  nand_4 g0834(.A(new_n1109), .B(new_n690), .Y(new_n1110));
  nor_4  g0835(.A(new_n1110), .B(new_n701), .Y(new_n1111));
  xnor_3 g0836(.A(new_n1111), .B(new_n780), .Y(new_n1112));
  xnor_3 g0837(.A(new_n1112), .B(new_n1108), .Y(new_n1113_1));
  xnor_3 g0838(.A(new_n1105), .B(n738), .Y(new_n1114));
  xnor_3 g0839(.A(new_n1110), .B(new_n700), .Y(new_n1115));
  nor_4  g0840(.A(new_n1115), .B(new_n1114), .Y(new_n1116));
  xnor_3 g0841(.A(new_n1115), .B(new_n1114), .Y(new_n1117));
  not_3  g0842(.A(n961), .Y(new_n1118));
  xnor_3 g0843(.A(new_n1104), .B(new_n1118), .Y(new_n1119_1));
  xnor_3 g0844(.A(new_n1109), .B(new_n649_1), .Y(new_n1120));
  nor_4  g0845(.A(new_n1120), .B(new_n1119_1), .Y(new_n1121));
  xnor_3 g0846(.A(new_n1120), .B(new_n1119_1), .Y(new_n1122));
  nor_4  g0847(.A(new_n1051), .B(new_n1025_1), .Y(new_n1123));
  nor_4  g0848(.A(new_n1096), .B(new_n1052), .Y(new_n1124));
  nor_4  g0849(.A(new_n1124), .B(new_n1123), .Y(new_n1125));
  nor_4  g0850(.A(new_n1125), .B(new_n1122), .Y(new_n1126));
  nor_4  g0851(.A(new_n1126), .B(new_n1121), .Y(new_n1127));
  nor_4  g0852(.A(new_n1127), .B(new_n1117), .Y(new_n1128));
  nor_4  g0853(.A(new_n1128), .B(new_n1116), .Y(new_n1129));
  xnor_3 g0854(.A(new_n1129), .B(new_n1113_1), .Y(n238));
  not_3  g0855(.A(n675), .Y(new_n1131));
  not_3  g0856(.A(n433), .Y(new_n1132));
  nor_4  g0857(.A(new_n302), .B(new_n1132), .Y(new_n1133));
  nand_4 g0858(.A(new_n1133), .B(n1537), .Y(new_n1134));
  nor_4  g0859(.A(new_n1134), .B(new_n1131), .Y(new_n1135_1));
  xor_3  g0860(.A(new_n1135_1), .B(n1263), .Y(new_n1136));
  not_3  g0861(.A(new_n1134), .Y(new_n1137));
  nor_4  g0862(.A(new_n1137), .B(n675), .Y(new_n1138_1));
  nor_4  g0863(.A(new_n1138_1), .B(new_n1135_1), .Y(new_n1139));
  not_3  g0864(.A(new_n1139), .Y(new_n1140_1));
  nor_4  g0865(.A(new_n1140_1), .B(new_n486), .Y(new_n1141));
  xnor_3 g0866(.A(new_n1139), .B(n379), .Y(new_n1142_1));
  xnor_3 g0867(.A(new_n1133), .B(n1537), .Y(new_n1143));
  nor_4  g0868(.A(new_n1143), .B(new_n483), .Y(new_n1144));
  xnor_3 g0869(.A(new_n1143), .B(n1527), .Y(new_n1145_1));
  nand_4 g0870(.A(new_n303_1), .B(n46), .Y(new_n1146));
  nand_4 g0871(.A(new_n388), .B(n1597), .Y(new_n1147));
  nand_4 g0872(.A(new_n995), .B(new_n975), .Y(new_n1148));
  nand_4 g0873(.A(new_n1148), .B(new_n1147), .Y(new_n1149_1));
  xnor_3 g0874(.A(new_n303_1), .B(new_n366), .Y(new_n1150));
  nand_4 g0875(.A(new_n1150), .B(new_n1149_1), .Y(new_n1151));
  nand_4 g0876(.A(new_n1151), .B(new_n1146), .Y(new_n1152));
  nand_4 g0877(.A(new_n1152), .B(new_n1145_1), .Y(new_n1153));
  not_3  g0878(.A(new_n1153), .Y(new_n1154));
  nor_4  g0879(.A(new_n1154), .B(new_n1144), .Y(new_n1155));
  nor_4  g0880(.A(new_n1155), .B(new_n1142_1), .Y(new_n1156));
  nor_4  g0881(.A(new_n1156), .B(new_n1141), .Y(new_n1157));
  nand_4 g0882(.A(new_n1157), .B(new_n1136), .Y(new_n1158));
  not_3  g0883(.A(new_n1158), .Y(new_n1159));
  nor_4  g0884(.A(new_n1157), .B(new_n1136), .Y(new_n1160));
  nor_4  g0885(.A(new_n1160), .B(new_n1159), .Y(new_n1161_1));
  not_3  g0886(.A(new_n1161_1), .Y(new_n1162_1));
  not_3  g0887(.A(new_n1142_1), .Y(new_n1163));
  xor_3  g0888(.A(new_n1155), .B(new_n1163), .Y(new_n1164));
  nor_4  g0889(.A(new_n1152), .B(new_n1145_1), .Y(new_n1165));
  nor_4  g0890(.A(new_n1165), .B(new_n1154), .Y(new_n1166));
  not_3  g0891(.A(new_n1166), .Y(new_n1167));
  nor_4  g0892(.A(new_n1000_1), .B(new_n997), .Y(new_n1168));
  nand_4 g0893(.A(new_n1168), .B(new_n996), .Y(new_n1169));
  xnor_3 g0894(.A(new_n1150), .B(new_n1149_1), .Y(new_n1170));
  not_3  g0895(.A(new_n1170), .Y(new_n1171));
  nor_4  g0896(.A(new_n1171), .B(new_n1169), .Y(new_n1172_1));
  nand_4 g0897(.A(new_n1172_1), .B(new_n1167), .Y(new_n1173));
  nor_4  g0898(.A(new_n1173), .B(n1426), .Y(new_n1174));
  nand_4 g0899(.A(new_n1174), .B(new_n1164), .Y(new_n1175_1));
  xnor_3 g0900(.A(new_n1175_1), .B(new_n1162_1), .Y(n270));
  xnor_3 g0901(.A(new_n721), .B(new_n391_1), .Y(new_n1177));
  not_3  g0902(.A(new_n1177), .Y(new_n1178));
  nor_4  g0903(.A(new_n736), .B(new_n397), .Y(new_n1179));
  nor_4  g0904(.A(new_n741), .B(new_n401_1), .Y(new_n1180));
  not_3  g0905(.A(new_n410), .Y(new_n1181));
  nand_4 g0906(.A(new_n749), .B(new_n404), .Y(new_n1182));
  nand_4 g0907(.A(new_n1182), .B(new_n1181), .Y(new_n1183_1));
  xnor_3 g0908(.A(new_n669), .B(new_n665_1), .Y(new_n1184));
  nor_4  g0909(.A(new_n1184), .B(new_n465), .Y(new_n1185));
  nor_4  g0910(.A(new_n1185), .B(new_n410), .Y(new_n1186));
  nor_4  g0911(.A(new_n1182), .B(new_n291), .Y(new_n1187));
  nor_4  g0912(.A(new_n1187), .B(new_n1186), .Y(new_n1188));
  nand_4 g0913(.A(new_n1188), .B(new_n754), .Y(new_n1189));
  nand_4 g0914(.A(new_n1189), .B(new_n1183_1), .Y(new_n1190));
  xnor_3 g0915(.A(new_n741), .B(new_n401_1), .Y(new_n1191_1));
  nor_4  g0916(.A(new_n1191_1), .B(new_n1190), .Y(new_n1192));
  nor_4  g0917(.A(new_n1192), .B(new_n1180), .Y(new_n1193));
  xnor_3 g0918(.A(new_n736), .B(new_n397), .Y(new_n1194_1));
  nor_4  g0919(.A(new_n1194_1), .B(new_n1193), .Y(new_n1195));
  nor_4  g0920(.A(new_n1195), .B(new_n1179), .Y(new_n1196));
  xor_3  g0921(.A(new_n1196), .B(new_n1178), .Y(n276));
  xor_3  g0922(.A(new_n887), .B(new_n407), .Y(n290));
  not_3  g0923(.A(new_n987), .Y(new_n1199_1));
  xor_3  g0924(.A(new_n1199_1), .B(new_n986), .Y(n292));
  not_3  g0925(.A(new_n809), .Y(new_n1201_1));
  nor_4  g0926(.A(new_n1201_1), .B(n266), .Y(new_n1202_1));
  not_3  g0927(.A(new_n1202_1), .Y(new_n1203));
  nand_4 g0928(.A(new_n1111), .B(new_n798), .Y(new_n1204));
  nor_4  g0929(.A(new_n1204), .B(new_n800), .Y(new_n1205));
  nand_4 g0930(.A(new_n1205), .B(new_n816), .Y(new_n1206));
  xor_3  g0931(.A(new_n1205), .B(new_n816), .Y(new_n1207));
  nor_4  g0932(.A(new_n1107), .B(new_n1101), .Y(new_n1208));
  xor_3  g0933(.A(new_n1204), .B(new_n800), .Y(new_n1209));
  nor_4  g0934(.A(new_n1209), .B(new_n1208), .Y(new_n1210));
  xnor_3 g0935(.A(new_n1209), .B(new_n1208), .Y(new_n1211));
  nor_4  g0936(.A(new_n1112), .B(new_n1108), .Y(new_n1212));
  nor_4  g0937(.A(new_n1129), .B(new_n1113_1), .Y(new_n1213));
  nor_4  g0938(.A(new_n1213), .B(new_n1212), .Y(new_n1214));
  nor_4  g0939(.A(new_n1214), .B(new_n1211), .Y(new_n1215));
  nor_4  g0940(.A(new_n1215), .B(new_n1210), .Y(new_n1216));
  nand_4 g0941(.A(new_n1216), .B(new_n1207), .Y(new_n1217));
  nand_4 g0942(.A(new_n1217), .B(new_n1206), .Y(new_n1218));
  nor_4  g0943(.A(new_n1218), .B(new_n1203), .Y(n299));
  nand_4 g0944(.A(new_n516), .B(n1341), .Y(new_n1220));
  xnor_3 g0945(.A(new_n517_1), .B(n1341), .Y(new_n1221));
  nand_4 g0946(.A(new_n442), .B(n69), .Y(new_n1222_1));
  nand_4 g0947(.A(new_n458), .B(new_n443), .Y(new_n1223));
  nand_4 g0948(.A(new_n1223), .B(new_n1222_1), .Y(new_n1224));
  nand_4 g0949(.A(new_n1224), .B(new_n1221), .Y(new_n1225));
  nand_4 g0950(.A(new_n1225), .B(new_n1220), .Y(new_n1226));
  nand_4 g0951(.A(new_n1226), .B(new_n509), .Y(new_n1227));
  not_3  g0952(.A(new_n1227), .Y(new_n1228));
  nand_4 g0953(.A(new_n1228), .B(new_n544), .Y(new_n1229));
  xnor_3 g0954(.A(new_n1229), .B(new_n556), .Y(new_n1230));
  not_3  g0955(.A(new_n1230), .Y(new_n1231));
  not_3  g0956(.A(n862), .Y(new_n1232));
  nor_4  g0957(.A(n1643), .B(n761), .Y(new_n1233));
  not_3  g0958(.A(new_n1233), .Y(new_n1234_1));
  xor_3  g0959(.A(n1643), .B(n761), .Y(new_n1235_1));
  nor_4  g0960(.A(n1172), .B(n555), .Y(new_n1236));
  not_3  g0961(.A(new_n1236), .Y(new_n1237_1));
  xor_3  g0962(.A(n1172), .B(n555), .Y(new_n1238));
  nor_4  g0963(.A(n695), .B(n353), .Y(new_n1239));
  nand_4 g0964(.A(n695), .B(n353), .Y(new_n1240));
  not_3  g0965(.A(new_n1240), .Y(new_n1241));
  nor_4  g0966(.A(new_n1241), .B(new_n1239), .Y(new_n1242));
  not_3  g0967(.A(new_n1242), .Y(new_n1243));
  nor_4  g0968(.A(n1296), .B(n952), .Y(new_n1244));
  nand_4 g0969(.A(n1145), .B(n1062), .Y(new_n1245));
  not_3  g0970(.A(new_n1245), .Y(new_n1246));
  not_3  g0971(.A(new_n1244), .Y(new_n1247));
  nand_4 g0972(.A(n1296), .B(n952), .Y(new_n1248));
  nand_4 g0973(.A(new_n1248), .B(new_n1247), .Y(new_n1249_1));
  nor_4  g0974(.A(new_n1249_1), .B(new_n1246), .Y(new_n1250));
  nor_4  g0975(.A(new_n1250), .B(new_n1244), .Y(new_n1251));
  nor_4  g0976(.A(new_n1251), .B(new_n1243), .Y(new_n1252));
  nor_4  g0977(.A(new_n1252), .B(new_n1239), .Y(new_n1253));
  not_3  g0978(.A(new_n1253), .Y(new_n1254));
  nand_4 g0979(.A(new_n1254), .B(new_n1238), .Y(new_n1255_1));
  nand_4 g0980(.A(new_n1255_1), .B(new_n1237_1), .Y(new_n1256));
  nand_4 g0981(.A(new_n1256), .B(new_n1235_1), .Y(new_n1257));
  nand_4 g0982(.A(new_n1257), .B(new_n1234_1), .Y(new_n1258));
  nor_4  g0983(.A(new_n1258), .B(new_n1232), .Y(new_n1259));
  nor_4  g0984(.A(new_n1259), .B(n1222), .Y(new_n1260_1));
  not_3  g0985(.A(n1222), .Y(new_n1261));
  not_3  g0986(.A(new_n1259), .Y(new_n1262));
  nor_4  g0987(.A(new_n1262), .B(new_n1261), .Y(new_n1263_1));
  nor_4  g0988(.A(new_n1263_1), .B(new_n1260_1), .Y(new_n1264));
  xnor_3 g0989(.A(new_n1264), .B(new_n1231), .Y(new_n1265));
  xnor_3 g0990(.A(new_n1227), .B(new_n545), .Y(new_n1266));
  xnor_3 g0991(.A(new_n1258), .B(new_n1232), .Y(new_n1267));
  nand_4 g0992(.A(new_n1267), .B(new_n1266), .Y(new_n1268));
  not_3  g0993(.A(new_n1268), .Y(new_n1269));
  xnor_3 g0994(.A(new_n1267), .B(new_n1266), .Y(new_n1270));
  xnor_3 g0995(.A(new_n1226), .B(new_n509), .Y(new_n1271));
  not_3  g0996(.A(new_n1271), .Y(new_n1272));
  xnor_3 g0997(.A(new_n1256), .B(new_n1235_1), .Y(new_n1273));
  nor_4  g0998(.A(new_n1273), .B(new_n1272), .Y(new_n1274));
  xnor_3 g0999(.A(new_n1273), .B(new_n1271), .Y(new_n1275));
  xnor_3 g1000(.A(new_n1224), .B(new_n1221), .Y(new_n1276));
  xnor_3 g1001(.A(new_n1253), .B(new_n1238), .Y(new_n1277_1));
  nand_4 g1002(.A(new_n1277_1), .B(new_n1276), .Y(new_n1278_1));
  not_3  g1003(.A(new_n1221), .Y(new_n1279));
  xnor_3 g1004(.A(new_n1224), .B(new_n1279), .Y(new_n1280));
  xnor_3 g1005(.A(new_n1277_1), .B(new_n1280), .Y(new_n1281));
  not_3  g1006(.A(new_n1251), .Y(new_n1282));
  nor_4  g1007(.A(new_n1282), .B(new_n1242), .Y(new_n1283_1));
  nor_4  g1008(.A(new_n1283_1), .B(new_n1252), .Y(new_n1284));
  nand_4 g1009(.A(new_n1284), .B(new_n461), .Y(new_n1285));
  xnor_3 g1010(.A(new_n1284), .B(new_n459), .Y(new_n1286));
  not_3  g1011(.A(new_n1249_1), .Y(new_n1287));
  nor_4  g1012(.A(new_n1287), .B(new_n1245), .Y(new_n1288));
  not_3  g1013(.A(new_n1250), .Y(new_n1289));
  nor_4  g1014(.A(n1145), .B(n1062), .Y(new_n1290));
  nor_4  g1015(.A(new_n1290), .B(new_n1246), .Y(new_n1291));
  nand_4 g1016(.A(new_n1291), .B(new_n466), .Y(new_n1292));
  nand_4 g1017(.A(new_n1292), .B(new_n1289), .Y(new_n1293));
  nor_4  g1018(.A(new_n1293), .B(new_n1288), .Y(new_n1294));
  not_3  g1019(.A(new_n1294), .Y(new_n1295));
  nor_4  g1020(.A(new_n1292), .B(new_n1249_1), .Y(new_n1296_1));
  nor_4  g1021(.A(new_n1296_1), .B(new_n1294), .Y(new_n1297));
  nand_4 g1022(.A(new_n1297), .B(new_n471), .Y(new_n1298));
  nand_4 g1023(.A(new_n1298), .B(new_n1295), .Y(new_n1299));
  nand_4 g1024(.A(new_n1299), .B(new_n1286), .Y(new_n1300));
  nand_4 g1025(.A(new_n1300), .B(new_n1285), .Y(new_n1301));
  nand_4 g1026(.A(new_n1301), .B(new_n1281), .Y(new_n1302));
  nand_4 g1027(.A(new_n1302), .B(new_n1278_1), .Y(new_n1303));
  nand_4 g1028(.A(new_n1303), .B(new_n1275), .Y(new_n1304));
  not_3  g1029(.A(new_n1304), .Y(new_n1305_1));
  nor_4  g1030(.A(new_n1305_1), .B(new_n1274), .Y(new_n1306));
  nor_4  g1031(.A(new_n1306), .B(new_n1270), .Y(new_n1307));
  nor_4  g1032(.A(new_n1307), .B(new_n1269), .Y(new_n1308));
  xor_3  g1033(.A(new_n1308), .B(new_n1265), .Y(n317));
  xor_3  g1034(.A(new_n1291), .B(new_n466), .Y(n372));
  xor_3  g1035(.A(new_n904), .B(new_n882_1), .Y(n378));
  not_3  g1036(.A(new_n816), .Y(new_n1312));
  nor_4  g1037(.A(new_n972), .B(new_n649_1), .Y(new_n1313));
  nand_4 g1038(.A(new_n1313), .B(new_n700), .Y(new_n1314));
  nor_4  g1039(.A(new_n1314), .B(new_n780), .Y(new_n1315_1));
  nand_4 g1040(.A(new_n1315_1), .B(new_n793), .Y(new_n1316));
  nor_4  g1041(.A(new_n1316), .B(new_n1312), .Y(new_n1317));
  xor_3  g1042(.A(new_n1317), .B(new_n1202_1), .Y(n1425));
  xor_3  g1043(.A(new_n1315_1), .B(new_n793), .Y(n1249));
  not_3  g1044(.A(n1249), .Y(new_n1320));
  xor_3  g1045(.A(new_n1313), .B(new_n700), .Y(n1119));
  not_3  g1046(.A(n1119), .Y(new_n1322));
  nand_4 g1047(.A(new_n669), .B(new_n524), .Y(new_n1323));
  and_4  g1048(.A(new_n1323), .B(new_n960), .Y(n647));
  not_3  g1049(.A(n647), .Y(n1255));
  xor_3  g1050(.A(new_n961_1), .B(new_n960), .Y(new_n1326));
  nand_4 g1051(.A(new_n1326), .B(n1255), .Y(new_n1327));
  xnor_3 g1052(.A(new_n963), .B(new_n957), .Y(n1016));
  nor_4  g1053(.A(n1016), .B(new_n1327), .Y(new_n1329));
  xnor_3 g1054(.A(new_n966), .B(new_n965), .Y(n1683));
  not_3  g1055(.A(n1683), .Y(new_n1331));
  nor_4  g1056(.A(new_n1331), .B(new_n1329), .Y(new_n1332_1));
  nor_4  g1057(.A(new_n968_1), .B(new_n951), .Y(new_n1333));
  nor_4  g1058(.A(new_n1333), .B(new_n970), .Y(new_n1334));
  not_3  g1059(.A(new_n1334), .Y(n569));
  nand_4 g1060(.A(n569), .B(new_n1332_1), .Y(new_n1336));
  xor_3  g1061(.A(new_n971), .B(new_n630), .Y(n773));
  not_3  g1062(.A(n773), .Y(new_n1338_1));
  nor_4  g1063(.A(new_n1338_1), .B(new_n1336), .Y(new_n1339));
  nand_4 g1064(.A(new_n1339), .B(new_n690), .Y(new_n1340_1));
  nor_4  g1065(.A(new_n1340_1), .B(new_n1322), .Y(new_n1341_1));
  nand_4 g1066(.A(new_n1341_1), .B(new_n798), .Y(new_n1342));
  nor_4  g1067(.A(new_n1342), .B(new_n1320), .Y(new_n1343));
  nand_4 g1068(.A(new_n1343), .B(new_n816), .Y(new_n1344));
  xnor_3 g1069(.A(new_n1344), .B(n1425), .Y(n387));
  nor_4  g1070(.A(new_n1229), .B(new_n567), .Y(new_n1346));
  nand_4 g1071(.A(new_n1346), .B(new_n563), .Y(new_n1347_1));
  not_3  g1072(.A(new_n1347_1), .Y(new_n1348_1));
  nor_4  g1073(.A(new_n1346), .B(new_n563), .Y(new_n1349_1));
  nor_4  g1074(.A(new_n1349_1), .B(new_n1348_1), .Y(new_n1350));
  xnor_3 g1075(.A(new_n1263_1), .B(n1757), .Y(new_n1351_1));
  not_3  g1076(.A(new_n1351_1), .Y(new_n1352));
  nor_4  g1077(.A(new_n1352), .B(new_n1350), .Y(new_n1353));
  not_3  g1078(.A(new_n1350), .Y(new_n1354));
  nor_4  g1079(.A(new_n1351_1), .B(new_n1354), .Y(new_n1355));
  nor_4  g1080(.A(new_n1355), .B(new_n1353), .Y(new_n1356));
  nor_4  g1081(.A(new_n1264), .B(new_n1230), .Y(new_n1357));
  not_3  g1082(.A(new_n1265), .Y(new_n1358));
  nor_4  g1083(.A(new_n1308), .B(new_n1358), .Y(new_n1359));
  nor_4  g1084(.A(new_n1359), .B(new_n1357), .Y(new_n1360));
  xor_3  g1085(.A(new_n1360), .B(new_n1356), .Y(n401));
  not_3  g1086(.A(new_n578), .Y(n416));
  xnor_3 g1087(.A(new_n898), .B(new_n896), .Y(new_n1363_1));
  xor_3  g1088(.A(new_n1363_1), .B(new_n424_1), .Y(n423));
  nor_4  g1089(.A(new_n1280), .B(new_n396), .Y(new_n1365));
  nor_4  g1090(.A(new_n1276), .B(new_n397), .Y(new_n1366));
  nor_4  g1091(.A(new_n1366), .B(new_n1365), .Y(new_n1367));
  not_3  g1092(.A(new_n1367), .Y(new_n1368));
  not_3  g1093(.A(new_n460_1), .Y(new_n1369_1));
  nand_4 g1094(.A(new_n476_1), .B(new_n463), .Y(new_n1370));
  nand_4 g1095(.A(new_n1370), .B(new_n1369_1), .Y(new_n1371));
  xor_3  g1096(.A(new_n1371), .B(new_n1368), .Y(n426));
  not_3  g1097(.A(new_n1344), .Y(new_n1373));
  xor_3  g1098(.A(new_n1316), .B(new_n1312), .Y(n493));
  nor_4  g1099(.A(n493), .B(new_n1343), .Y(new_n1375));
  nor_4  g1100(.A(new_n1375), .B(new_n1373), .Y(n429));
  xor_3  g1101(.A(new_n1338_1), .B(new_n1336), .Y(n432));
  xnor_3 g1102(.A(new_n1271), .B(new_n391_1), .Y(new_n1378));
  not_3  g1103(.A(new_n1378), .Y(new_n1379));
  not_3  g1104(.A(new_n1365), .Y(new_n1380));
  nand_4 g1105(.A(new_n1371), .B(new_n1367), .Y(new_n1381_1));
  nand_4 g1106(.A(new_n1381_1), .B(new_n1380), .Y(new_n1382));
  xor_3  g1107(.A(new_n1382), .B(new_n1379), .Y(n452));
  not_3  g1108(.A(new_n996), .Y(new_n1384));
  nor_4  g1109(.A(new_n1002), .B(new_n1384), .Y(new_n1385_1));
  xor_3  g1110(.A(new_n1171), .B(new_n1385_1), .Y(n457));
  xnor_3 g1111(.A(new_n1214), .B(new_n1211), .Y(n460));
  xor_3  g1112(.A(new_n749), .B(new_n747_1), .Y(n476));
  not_3  g1113(.A(new_n426_1), .Y(new_n1389));
  xor_3  g1114(.A(new_n1389), .B(new_n399), .Y(n482));
  nor_4  g1115(.A(new_n1347_1), .B(new_n496), .Y(new_n1391));
  xor_3  g1116(.A(new_n1391), .B(new_n937), .Y(new_n1392));
  xnor_3 g1117(.A(new_n1392), .B(new_n1135_1), .Y(new_n1393_1));
  xnor_3 g1118(.A(new_n1347_1), .B(new_n496), .Y(new_n1394));
  not_3  g1119(.A(new_n1394), .Y(new_n1395));
  nor_4  g1120(.A(new_n1395), .B(new_n1139), .Y(new_n1396));
  xnor_3 g1121(.A(new_n1394), .B(new_n1140_1), .Y(new_n1397));
  not_3  g1122(.A(new_n1143), .Y(new_n1398));
  nor_4  g1123(.A(new_n1350), .B(new_n1398), .Y(new_n1399_1));
  xnor_3 g1124(.A(new_n1350), .B(new_n1398), .Y(new_n1400));
  xnor_3 g1125(.A(new_n302), .B(new_n1132), .Y(new_n1401));
  nor_4  g1126(.A(new_n1231), .B(new_n1401), .Y(new_n1402));
  not_3  g1127(.A(new_n1402), .Y(new_n1403));
  not_3  g1128(.A(new_n1266), .Y(new_n1404));
  nor_4  g1129(.A(new_n1404), .B(new_n388), .Y(new_n1405));
  not_3  g1130(.A(new_n1405), .Y(new_n1406));
  nor_4  g1131(.A(new_n1266), .B(new_n385), .Y(new_n1407_1));
  nor_4  g1132(.A(new_n1407_1), .B(new_n1405), .Y(new_n1408));
  nand_4 g1133(.A(new_n1271), .B(new_n392), .Y(new_n1409));
  nand_4 g1134(.A(new_n1382), .B(new_n1378), .Y(new_n1410));
  nand_4 g1135(.A(new_n1410), .B(new_n1409), .Y(new_n1411));
  nand_4 g1136(.A(new_n1411), .B(new_n1408), .Y(new_n1412));
  nand_4 g1137(.A(new_n1412), .B(new_n1406), .Y(new_n1413));
  not_3  g1138(.A(new_n1413), .Y(new_n1414));
  nor_4  g1139(.A(new_n1230), .B(new_n303_1), .Y(new_n1415));
  nor_4  g1140(.A(new_n1415), .B(new_n1402), .Y(new_n1416));
  nand_4 g1141(.A(new_n1416), .B(new_n1414), .Y(new_n1417));
  nand_4 g1142(.A(new_n1417), .B(new_n1403), .Y(new_n1418));
  nor_4  g1143(.A(new_n1418), .B(new_n1400), .Y(new_n1419));
  nor_4  g1144(.A(new_n1419), .B(new_n1399_1), .Y(new_n1420));
  nor_4  g1145(.A(new_n1420), .B(new_n1397), .Y(new_n1421));
  nor_4  g1146(.A(new_n1421), .B(new_n1396), .Y(new_n1422_1));
  xnor_3 g1147(.A(new_n1422_1), .B(new_n1393_1), .Y(n510));
  xnor_3 g1148(.A(new_n1139), .B(new_n1112), .Y(new_n1424));
  nor_4  g1149(.A(new_n1398), .B(new_n1115), .Y(new_n1425_1));
  not_3  g1150(.A(new_n1425_1), .Y(new_n1426_1));
  not_3  g1151(.A(new_n1115), .Y(new_n1427));
  nor_4  g1152(.A(new_n1143), .B(new_n1427), .Y(new_n1428));
  nor_4  g1153(.A(new_n1428), .B(new_n1425_1), .Y(new_n1429));
  nor_4  g1154(.A(new_n1120), .B(new_n303_1), .Y(new_n1430));
  not_3  g1155(.A(new_n1430), .Y(new_n1431));
  not_3  g1156(.A(new_n1120), .Y(new_n1432));
  nor_4  g1157(.A(new_n1432), .B(new_n1401), .Y(new_n1433));
  nor_4  g1158(.A(new_n1433), .B(new_n1430), .Y(new_n1434));
  nor_4  g1159(.A(new_n1025_1), .B(new_n388), .Y(new_n1435_1));
  not_3  g1160(.A(new_n1435_1), .Y(new_n1436));
  not_3  g1161(.A(new_n1025_1), .Y(new_n1437));
  nor_4  g1162(.A(new_n1437), .B(new_n385), .Y(new_n1438));
  nor_4  g1163(.A(new_n1438), .B(new_n1435_1), .Y(new_n1439));
  nor_4  g1164(.A(new_n1089), .B(new_n392), .Y(new_n1440_1));
  nand_4 g1165(.A(new_n1057), .B(new_n397), .Y(new_n1441));
  xnor_3 g1166(.A(new_n1057), .B(new_n396), .Y(new_n1442));
  nor_4  g1167(.A(new_n1062_1), .B(new_n400), .Y(new_n1443));
  not_3  g1168(.A(new_n1443), .Y(new_n1444));
  nor_4  g1169(.A(new_n1063), .B(new_n401_1), .Y(new_n1445));
  nor_4  g1170(.A(new_n1445), .B(new_n1443), .Y(new_n1446));
  not_3  g1171(.A(new_n1073), .Y(new_n1447));
  nor_4  g1172(.A(new_n1447), .B(new_n465), .Y(new_n1448));
  nor_4  g1173(.A(new_n1448), .B(new_n410), .Y(new_n1449));
  not_3  g1174(.A(new_n1449), .Y(new_n1450));
  not_3  g1175(.A(new_n1448), .Y(new_n1451));
  nor_4  g1176(.A(new_n1451), .B(new_n291), .Y(new_n1452));
  nor_4  g1177(.A(new_n1452), .B(new_n1449), .Y(new_n1453_1));
  nand_4 g1178(.A(new_n1453_1), .B(new_n1078), .Y(new_n1454));
  nand_4 g1179(.A(new_n1454), .B(new_n1450), .Y(new_n1455));
  nand_4 g1180(.A(new_n1455), .B(new_n1446), .Y(new_n1456));
  nand_4 g1181(.A(new_n1456), .B(new_n1444), .Y(new_n1457_1));
  nand_4 g1182(.A(new_n1457_1), .B(new_n1442), .Y(new_n1458));
  nand_4 g1183(.A(new_n1458), .B(new_n1441), .Y(new_n1459));
  xnor_3 g1184(.A(new_n1054), .B(new_n391_1), .Y(new_n1460_1));
  nor_4  g1185(.A(new_n1460_1), .B(new_n1459), .Y(new_n1461_1));
  nor_4  g1186(.A(new_n1461_1), .B(new_n1440_1), .Y(new_n1462));
  nand_4 g1187(.A(new_n1462), .B(new_n1439), .Y(new_n1463_1));
  nand_4 g1188(.A(new_n1463_1), .B(new_n1436), .Y(new_n1464));
  nand_4 g1189(.A(new_n1464), .B(new_n1434), .Y(new_n1465));
  nand_4 g1190(.A(new_n1465), .B(new_n1431), .Y(new_n1466));
  nand_4 g1191(.A(new_n1466), .B(new_n1429), .Y(new_n1467));
  nand_4 g1192(.A(new_n1467), .B(new_n1426_1), .Y(new_n1468));
  xor_3  g1193(.A(new_n1468), .B(new_n1424), .Y(n517));
  xnor_3 g1194(.A(new_n1140_1), .B(new_n832), .Y(new_n1470_1));
  nand_4 g1195(.A(new_n1143), .B(new_n706), .Y(new_n1471));
  xnor_3 g1196(.A(new_n1143), .B(new_n838), .Y(new_n1472));
  nand_4 g1197(.A(new_n770_1), .B(new_n1401), .Y(new_n1473));
  nand_4 g1198(.A(new_n715_1), .B(new_n385), .Y(new_n1474));
  xnor_3 g1199(.A(new_n715_1), .B(new_n388), .Y(new_n1475));
  nand_4 g1200(.A(new_n721), .B(new_n392), .Y(new_n1476));
  nand_4 g1201(.A(new_n1196), .B(new_n1177), .Y(new_n1477));
  nand_4 g1202(.A(new_n1477), .B(new_n1476), .Y(new_n1478));
  nand_4 g1203(.A(new_n1478), .B(new_n1475), .Y(new_n1479));
  nand_4 g1204(.A(new_n1479), .B(new_n1474), .Y(new_n1480));
  xnor_3 g1205(.A(new_n712_1), .B(new_n1401), .Y(new_n1481_1));
  nand_4 g1206(.A(new_n1481_1), .B(new_n1480), .Y(new_n1482));
  nand_4 g1207(.A(new_n1482), .B(new_n1473), .Y(new_n1483));
  nand_4 g1208(.A(new_n1483), .B(new_n1472), .Y(new_n1484));
  nand_4 g1209(.A(new_n1484), .B(new_n1471), .Y(new_n1485));
  xnor_3 g1210(.A(new_n1485), .B(new_n1470_1), .Y(n522));
  xor_3  g1211(.A(new_n1155), .B(new_n1142_1), .Y(new_n1487));
  xnor_3 g1212(.A(new_n1173), .B(new_n1487), .Y(n532));
  not_3  g1213(.A(new_n318), .Y(new_n1489));
  nor_4  g1214(.A(new_n1201_1), .B(new_n1489), .Y(new_n1490));
  not_3  g1215(.A(new_n379_1), .Y(new_n1491));
  nor_4  g1216(.A(new_n1491), .B(new_n361), .Y(new_n1492));
  xor_3  g1217(.A(new_n373), .B(new_n478), .Y(new_n1493));
  nand_4 g1218(.A(new_n1493), .B(n1000), .Y(new_n1494));
  nor_4  g1219(.A(new_n693_1), .B(n682), .Y(new_n1495_1));
  nand_4 g1220(.A(new_n364), .B(n1527), .Y(new_n1496));
  not_3  g1221(.A(new_n1496), .Y(new_n1497));
  nor_4  g1222(.A(new_n1497), .B(new_n1495_1), .Y(new_n1498_1));
  nand_4 g1223(.A(new_n1498_1), .B(new_n305), .Y(new_n1499));
  nand_4 g1224(.A(new_n1499), .B(new_n1494), .Y(new_n1500));
  nand_4 g1225(.A(new_n1500), .B(new_n1492), .Y(new_n1501_1));
  xor_3  g1226(.A(new_n1495_1), .B(n379), .Y(new_n1502_1));
  nand_4 g1227(.A(new_n1502_1), .B(new_n305), .Y(new_n1503));
  nand_4 g1228(.A(new_n373), .B(n247), .Y(new_n1504));
  xor_3  g1229(.A(new_n1504), .B(new_n492), .Y(new_n1505));
  nand_4 g1230(.A(new_n1505), .B(n1000), .Y(new_n1506));
  nand_4 g1231(.A(new_n1506), .B(new_n1503), .Y(new_n1507_1));
  nor_4  g1232(.A(new_n1507_1), .B(new_n1501_1), .Y(new_n1508));
  nand_4 g1233(.A(new_n1495_1), .B(new_n486), .Y(new_n1509));
  nand_4 g1234(.A(new_n1509), .B(n1263), .Y(new_n1510));
  nor_4  g1235(.A(new_n810), .B(n682), .Y(new_n1511));
  nor_4  g1236(.A(new_n1511), .B(n1000), .Y(new_n1512));
  nand_4 g1237(.A(new_n1512), .B(new_n1510), .Y(new_n1513));
  nor_4  g1238(.A(new_n1504), .B(new_n492), .Y(new_n1514));
  xor_3  g1239(.A(new_n1514), .B(new_n908), .Y(new_n1515));
  nand_4 g1240(.A(new_n1515), .B(n1000), .Y(new_n1516));
  nand_4 g1241(.A(new_n1516), .B(new_n1513), .Y(new_n1517));
  nand_4 g1242(.A(new_n1517), .B(new_n1508), .Y(new_n1518));
  nand_4 g1243(.A(new_n1514), .B(n171), .Y(new_n1519));
  nand_4 g1244(.A(n1000), .B(n557), .Y(new_n1520));
  nor_4  g1245(.A(new_n1520), .B(new_n1519), .Y(new_n1521));
  nand_4 g1246(.A(new_n1512), .B(n1422), .Y(new_n1522));
  not_3  g1247(.A(new_n1520), .Y(new_n1523));
  nor_4  g1248(.A(new_n1519), .B(new_n305), .Y(new_n1524));
  nor_4  g1249(.A(new_n1524), .B(new_n1523), .Y(new_n1525_1));
  nand_4 g1250(.A(new_n1525_1), .B(new_n1522), .Y(new_n1526));
  nor_4  g1251(.A(new_n1526), .B(new_n1490), .Y(new_n1527_1));
  nor_4  g1252(.A(new_n1527_1), .B(new_n1521), .Y(new_n1528));
  nor_4  g1253(.A(new_n1528), .B(new_n1518), .Y(new_n1529));
  nor_4  g1254(.A(new_n1521), .B(new_n1490), .Y(new_n1530_1));
  and_4  g1255(.A(new_n1530_1), .B(new_n1529), .Y(new_n1531));
  nor_4  g1256(.A(new_n1531), .B(new_n1490), .Y(new_n1532));
  not_3  g1257(.A(new_n1518), .Y(new_n1533));
  xor_3  g1258(.A(new_n1528), .B(new_n1533), .Y(new_n1534));
  not_3  g1259(.A(new_n1534), .Y(new_n1535_1));
  not_3  g1260(.A(new_n322), .Y(new_n1536));
  xor_3  g1261(.A(n1597), .B(new_n362), .Y(new_n1537_1));
  nand_4 g1262(.A(new_n1537_1), .B(new_n305), .Y(new_n1538));
  not_3  g1263(.A(new_n326), .Y(new_n1539));
  nand_4 g1264(.A(new_n1539), .B(new_n1538), .Y(new_n1540));
  nor_4  g1265(.A(new_n1540), .B(new_n1536), .Y(new_n1541));
  nand_4 g1266(.A(new_n379_1), .B(new_n1541), .Y(new_n1542));
  xor_3  g1267(.A(new_n373), .B(n247), .Y(new_n1543));
  nor_4  g1268(.A(new_n1543), .B(new_n305), .Y(new_n1544_1));
  not_3  g1269(.A(new_n1499), .Y(new_n1545));
  nor_4  g1270(.A(new_n1545), .B(new_n1544_1), .Y(new_n1546));
  nor_4  g1271(.A(new_n1546), .B(new_n1542), .Y(new_n1547));
  xor_3  g1272(.A(new_n1495_1), .B(new_n486), .Y(new_n1548));
  nor_4  g1273(.A(new_n1548), .B(n1000), .Y(new_n1549));
  xor_3  g1274(.A(new_n1504), .B(n1642), .Y(new_n1550));
  nor_4  g1275(.A(new_n1550), .B(new_n305), .Y(new_n1551));
  nor_4  g1276(.A(new_n1551), .B(new_n1549), .Y(new_n1552));
  nor_4  g1277(.A(new_n1552), .B(new_n1547), .Y(new_n1553));
  nor_4  g1278(.A(new_n1553), .B(new_n1508), .Y(new_n1554));
  nor_4  g1279(.A(new_n380), .B(new_n360), .Y(new_n1555));
  xnor_3 g1280(.A(new_n1500), .B(new_n1492), .Y(new_n1556_1));
  nand_4 g1281(.A(new_n1556_1), .B(new_n1555), .Y(new_n1557));
  nor_4  g1282(.A(new_n1557), .B(new_n1554), .Y(new_n1558));
  xnor_3 g1283(.A(new_n1517), .B(new_n1508), .Y(new_n1559));
  nand_4 g1284(.A(new_n1559), .B(new_n1558), .Y(new_n1560));
  nor_4  g1285(.A(new_n1560), .B(new_n1535_1), .Y(new_n1561));
  nor_4  g1286(.A(new_n1561), .B(new_n1532), .Y(new_n1562));
  not_3  g1287(.A(new_n1562), .Y(new_n1563));
  xnor_3 g1288(.A(new_n1560), .B(new_n1534), .Y(new_n1564));
  not_3  g1289(.A(new_n1564), .Y(new_n1565));
  not_3  g1290(.A(n277), .Y(new_n1566));
  not_3  g1291(.A(n1622), .Y(new_n1567));
  not_3  g1292(.A(n49), .Y(new_n1568));
  nor_4  g1293(.A(n1643), .B(n469), .Y(new_n1569));
  not_3  g1294(.A(new_n1569), .Y(new_n1570));
  nand_4 g1295(.A(new_n872), .B(new_n853), .Y(new_n1571));
  nand_4 g1296(.A(new_n1571), .B(new_n1570), .Y(new_n1572));
  nor_4  g1297(.A(new_n1572), .B(new_n1568), .Y(new_n1573));
  not_3  g1298(.A(new_n1573), .Y(new_n1574));
  nor_4  g1299(.A(new_n1574), .B(new_n1567), .Y(new_n1575));
  nand_4 g1300(.A(new_n1575), .B(n906), .Y(new_n1576));
  nor_4  g1301(.A(new_n1576), .B(new_n1566), .Y(new_n1577));
  not_3  g1302(.A(new_n1560), .Y(new_n1578));
  nor_4  g1303(.A(new_n1559), .B(new_n1558), .Y(new_n1579));
  nor_4  g1304(.A(new_n1579), .B(new_n1578), .Y(new_n1580));
  nor_4  g1305(.A(new_n1580), .B(new_n1577), .Y(new_n1581));
  not_3  g1306(.A(new_n1581), .Y(new_n1582));
  not_3  g1307(.A(new_n1577), .Y(new_n1583));
  not_3  g1308(.A(new_n1580), .Y(new_n1584));
  nor_4  g1309(.A(new_n1584), .B(new_n1583), .Y(new_n1585));
  nor_4  g1310(.A(new_n1585), .B(new_n1581), .Y(new_n1586));
  not_3  g1311(.A(new_n1576), .Y(new_n1587));
  nor_4  g1312(.A(new_n1587), .B(n277), .Y(new_n1588));
  nor_4  g1313(.A(new_n1588), .B(new_n1577), .Y(new_n1589));
  xnor_3 g1314(.A(new_n1557), .B(new_n1554), .Y(new_n1590));
  not_3  g1315(.A(new_n1590), .Y(new_n1591));
  nor_4  g1316(.A(new_n1591), .B(new_n1589), .Y(new_n1592));
  not_3  g1317(.A(new_n1592), .Y(new_n1593));
  not_3  g1318(.A(new_n1589), .Y(new_n1594));
  nor_4  g1319(.A(new_n1590), .B(new_n1594), .Y(new_n1595_1));
  nor_4  g1320(.A(new_n1595_1), .B(new_n1592), .Y(new_n1596));
  nor_4  g1321(.A(new_n1575), .B(n906), .Y(new_n1597_1));
  nor_4  g1322(.A(new_n1597_1), .B(new_n1587), .Y(new_n1598));
  nor_4  g1323(.A(new_n1500), .B(new_n1492), .Y(new_n1599));
  nor_4  g1324(.A(new_n1599), .B(new_n1547), .Y(new_n1600_1));
  xnor_3 g1325(.A(new_n1600_1), .B(new_n1555), .Y(new_n1601_1));
  nor_4  g1326(.A(new_n1601_1), .B(new_n1598), .Y(new_n1602));
  not_3  g1327(.A(new_n1602), .Y(new_n1603));
  xnor_3 g1328(.A(new_n1601_1), .B(new_n1598), .Y(new_n1604));
  not_3  g1329(.A(new_n1604), .Y(new_n1605));
  not_3  g1330(.A(new_n381), .Y(new_n1606));
  nor_4  g1331(.A(new_n1573), .B(n1622), .Y(new_n1607));
  nor_4  g1332(.A(new_n1607), .B(new_n1575), .Y(new_n1608));
  nor_4  g1333(.A(new_n1608), .B(new_n1606), .Y(new_n1609));
  not_3  g1334(.A(new_n1609), .Y(new_n1610));
  xnor_3 g1335(.A(new_n1608), .B(new_n1606), .Y(new_n1611));
  not_3  g1336(.A(new_n1611), .Y(new_n1612));
  xnor_3 g1337(.A(new_n1572), .B(new_n1568), .Y(new_n1613_1));
  nor_4  g1338(.A(new_n1613_1), .B(new_n384), .Y(new_n1614));
  not_3  g1339(.A(new_n1614), .Y(new_n1615));
  xnor_3 g1340(.A(new_n1613_1), .B(new_n384), .Y(new_n1616));
  not_3  g1341(.A(new_n1616), .Y(new_n1617));
  nand_4 g1342(.A(new_n906_1), .B(new_n877), .Y(new_n1618));
  nand_4 g1343(.A(new_n1618), .B(new_n874), .Y(new_n1619));
  nand_4 g1344(.A(new_n1619), .B(new_n1617), .Y(new_n1620));
  nand_4 g1345(.A(new_n1620), .B(new_n1615), .Y(new_n1621));
  not_3  g1346(.A(new_n1621), .Y(new_n1622_1));
  nand_4 g1347(.A(new_n1622_1), .B(new_n1612), .Y(new_n1623));
  nand_4 g1348(.A(new_n1623), .B(new_n1610), .Y(new_n1624));
  nand_4 g1349(.A(new_n1624), .B(new_n1605), .Y(new_n1625));
  nand_4 g1350(.A(new_n1625), .B(new_n1603), .Y(new_n1626));
  nand_4 g1351(.A(new_n1626), .B(new_n1596), .Y(new_n1627));
  nand_4 g1352(.A(new_n1627), .B(new_n1593), .Y(new_n1628));
  nand_4 g1353(.A(new_n1628), .B(new_n1586), .Y(new_n1629_1));
  nand_4 g1354(.A(new_n1629_1), .B(new_n1582), .Y(new_n1630));
  nor_4  g1355(.A(new_n1630), .B(new_n1565), .Y(new_n1631));
  nor_4  g1356(.A(new_n1631), .B(new_n1563), .Y(n534));
  not_3  g1357(.A(new_n579), .Y(new_n1633_1));
  xor_3  g1358(.A(n1721), .B(new_n1633_1), .Y(n541));
  not_3  g1359(.A(n1426), .Y(n547));
  nor_4  g1360(.A(new_n1209), .B(new_n1135_1), .Y(new_n1636));
  xnor_3 g1361(.A(new_n1209), .B(new_n1135_1), .Y(new_n1637));
  nor_4  g1362(.A(new_n1139), .B(new_n1112), .Y(new_n1638));
  not_3  g1363(.A(new_n1468), .Y(new_n1639));
  nor_4  g1364(.A(new_n1639), .B(new_n1424), .Y(new_n1640));
  nor_4  g1365(.A(new_n1640), .B(new_n1638), .Y(new_n1641));
  nor_4  g1366(.A(new_n1641), .B(new_n1637), .Y(new_n1642_1));
  nor_4  g1367(.A(new_n1642_1), .B(new_n1636), .Y(new_n1643_1));
  nand_4 g1368(.A(new_n1643_1), .B(new_n1207), .Y(new_n1644));
  nand_4 g1369(.A(new_n1644), .B(new_n1206), .Y(new_n1645));
  nor_4  g1370(.A(new_n1645), .B(new_n1203), .Y(n549));
  xnor_3 g1371(.A(new_n1481_1), .B(new_n1480), .Y(n559));
  xor_3  g1372(.A(new_n1460_1), .B(new_n1459), .Y(n573));
  xnor_3 g1373(.A(new_n1641), .B(new_n1637), .Y(n588));
  not_3  g1374(.A(new_n575), .Y(new_n1650));
  xor_3  g1375(.A(new_n578), .B(new_n1650), .Y(n599));
  nor_4  g1376(.A(new_n1317), .B(new_n1203), .Y(n824));
  not_3  g1377(.A(n824), .Y(new_n1653));
  nor_4  g1378(.A(new_n1373), .B(new_n1653), .Y(n627));
  not_3  g1379(.A(new_n1207), .Y(new_n1655));
  xnor_3 g1380(.A(new_n1216), .B(new_n1655), .Y(n638));
  nor_4  g1381(.A(new_n928), .B(n557), .Y(new_n1657_1));
  nand_4 g1382(.A(new_n1657_1), .B(n1381), .Y(new_n1658));
  or_4   g1383(.A(new_n808), .B(new_n440), .Y(new_n1659));
  nand_4 g1384(.A(new_n1659), .B(new_n1658), .Y(new_n1660_1));
  nand_4 g1385(.A(new_n1660_1), .B(new_n934), .Y(new_n1661));
  not_3  g1386(.A(new_n1661), .Y(n643));
  not_3  g1387(.A(new_n960), .Y(new_n1663));
  xor_3  g1388(.A(new_n961_1), .B(new_n1663), .Y(n646));
  xor_3  g1389(.A(new_n1619), .B(new_n1617), .Y(n648));
  xnor_3 g1390(.A(new_n767), .B(new_n720), .Y(n665));
  xnor_3 g1391(.A(new_n1127), .B(new_n1117), .Y(n683));
  nor_4  g1392(.A(new_n1564), .B(new_n1135_1), .Y(new_n1668));
  not_3  g1393(.A(new_n1668), .Y(new_n1669));
  not_3  g1394(.A(new_n1135_1), .Y(new_n1670));
  xnor_3 g1395(.A(new_n1564), .B(new_n1670), .Y(new_n1671));
  nand_4 g1396(.A(new_n1584), .B(new_n1670), .Y(new_n1672));
  xnor_3 g1397(.A(new_n1580), .B(new_n1670), .Y(new_n1673));
  nand_4 g1398(.A(new_n1590), .B(new_n1140_1), .Y(new_n1674));
  xnor_3 g1399(.A(new_n1590), .B(new_n1139), .Y(new_n1675_1));
  xnor_3 g1400(.A(new_n1556_1), .B(new_n1555), .Y(new_n1676));
  nand_4 g1401(.A(new_n1676), .B(new_n1143), .Y(new_n1677_1));
  xnor_3 g1402(.A(new_n1601_1), .B(new_n1143), .Y(new_n1678_1));
  nand_4 g1403(.A(new_n381), .B(new_n1401), .Y(new_n1679));
  nand_4 g1404(.A(new_n433_1), .B(new_n382), .Y(new_n1680));
  nand_4 g1405(.A(new_n1680), .B(new_n1679), .Y(new_n1681));
  nand_4 g1406(.A(new_n1681), .B(new_n1678_1), .Y(new_n1682));
  nand_4 g1407(.A(new_n1682), .B(new_n1677_1), .Y(new_n1683_1));
  nand_4 g1408(.A(new_n1683_1), .B(new_n1675_1), .Y(new_n1684));
  nand_4 g1409(.A(new_n1684), .B(new_n1674), .Y(new_n1685));
  nand_4 g1410(.A(new_n1685), .B(new_n1673), .Y(new_n1686_1));
  nand_4 g1411(.A(new_n1686_1), .B(new_n1672), .Y(new_n1687));
  nand_4 g1412(.A(new_n1687), .B(new_n1671), .Y(new_n1688_1));
  nand_4 g1413(.A(new_n1688_1), .B(new_n1669), .Y(new_n1689));
  xor_3  g1414(.A(new_n1530_1), .B(new_n1529), .Y(new_n1690_1));
  xnor_3 g1415(.A(new_n1690_1), .B(new_n1561), .Y(new_n1691));
  nand_4 g1416(.A(new_n1691), .B(new_n1689), .Y(new_n1692));
  nor_4  g1417(.A(new_n1691), .B(new_n1135_1), .Y(new_n1693));
  not_3  g1418(.A(new_n1671), .Y(new_n1694));
  not_3  g1419(.A(new_n1687), .Y(new_n1695));
  nor_4  g1420(.A(new_n1695), .B(new_n1694), .Y(new_n1696));
  nor_4  g1421(.A(new_n1696), .B(new_n1670), .Y(new_n1697));
  nor_4  g1422(.A(new_n1697), .B(new_n1693), .Y(new_n1698));
  nand_4 g1423(.A(new_n1698), .B(new_n1692), .Y(new_n1699));
  xnor_3 g1424(.A(new_n1699), .B(new_n1562), .Y(n699));
  xor_3  g1425(.A(new_n894), .B(new_n415), .Y(n712));
  not_3  g1426(.A(new_n586), .Y(n715));
  not_3  g1427(.A(new_n1340_1), .Y(new_n1703));
  nor_4  g1428(.A(new_n1339), .B(n145), .Y(new_n1704));
  nor_4  g1429(.A(new_n1704), .B(new_n1703), .Y(n724));
  not_3  g1430(.A(n1016), .Y(new_n1706));
  xor_3  g1431(.A(new_n1706), .B(new_n1327), .Y(n725));
  xnor_3 g1432(.A(new_n1483), .B(new_n1472), .Y(n731));
  xnor_3 g1433(.A(new_n1681), .B(new_n1678_1), .Y(n748));
  xnor_3 g1434(.A(new_n1418), .B(new_n1400), .Y(n759));
  not_3  g1435(.A(new_n1173), .Y(new_n1711));
  nand_4 g1436(.A(new_n1711), .B(new_n1164), .Y(new_n1712));
  nor_4  g1437(.A(new_n1712), .B(new_n1162_1), .Y(new_n1713));
  nor_4  g1438(.A(new_n1135_1), .B(n1263), .Y(new_n1714));
  nor_4  g1439(.A(new_n1159), .B(new_n1714), .Y(new_n1715));
  nor_4  g1440(.A(new_n1715), .B(n1422), .Y(new_n1716));
  nand_4 g1441(.A(new_n1716), .B(new_n1713), .Y(new_n1717));
  not_3  g1442(.A(new_n1717), .Y(n770));
  not_3  g1443(.A(new_n1439), .Y(new_n1719));
  xor_3  g1444(.A(new_n1462), .B(new_n1719), .Y(n790));
  xor_3  g1445(.A(new_n1135_1), .B(new_n825), .Y(new_n1721_1));
  nor_4  g1446(.A(new_n1139), .B(new_n832), .Y(new_n1722));
  nand_4 g1447(.A(new_n1485), .B(new_n1470_1), .Y(new_n1723));
  not_3  g1448(.A(new_n1723), .Y(new_n1724));
  nor_4  g1449(.A(new_n1724), .B(new_n1722), .Y(new_n1725));
  xor_3  g1450(.A(new_n1725), .B(new_n1721_1), .Y(n792));
  not_3  g1451(.A(new_n1093), .Y(new_n1727_1));
  xor_3  g1452(.A(new_n1727_1), .B(new_n1088), .Y(n813));
  not_3  g1453(.A(new_n1286), .Y(new_n1729_1));
  xor_3  g1454(.A(new_n1299), .B(new_n1729_1), .Y(n823));
  not_3  g1455(.A(new_n471), .Y(new_n1731_1));
  xor_3  g1456(.A(new_n474), .B(new_n1731_1), .Y(n836));
  xnor_3 g1457(.A(new_n1683_1), .B(new_n1675_1), .Y(n846));
  not_3  g1458(.A(new_n1270), .Y(new_n1734));
  xor_3  g1459(.A(new_n1306), .B(new_n1734), .Y(n858));
  xor_3  g1460(.A(new_n1314), .B(new_n780), .Y(n865));
  not_3  g1461(.A(new_n1429), .Y(new_n1737_1));
  xor_3  g1462(.A(new_n1466), .B(new_n1737_1), .Y(n867));
  not_3  g1463(.A(new_n1391), .Y(new_n1739));
  nor_4  g1464(.A(new_n1739), .B(new_n919), .Y(new_n1740));
  not_3  g1465(.A(new_n1740), .Y(new_n1741));
  xor_3  g1466(.A(new_n1741), .B(new_n931_1), .Y(new_n1742));
  not_3  g1467(.A(new_n1742), .Y(new_n1743_1));
  nor_4  g1468(.A(new_n1392), .B(new_n1135_1), .Y(new_n1744));
  nor_4  g1469(.A(new_n1422_1), .B(new_n1393_1), .Y(new_n1745));
  nor_4  g1470(.A(new_n1745), .B(new_n1744), .Y(new_n1746_1));
  xnor_3 g1471(.A(new_n1746_1), .B(new_n1743_1), .Y(n883));
  not_3  g1472(.A(new_n771), .Y(new_n1748));
  xor_3  g1473(.A(new_n1748), .B(new_n769), .Y(n888));
  not_3  g1474(.A(new_n1392), .Y(new_n1750));
  not_3  g1475(.A(n839), .Y(new_n1751));
  nand_4 g1476(.A(new_n1263_1), .B(n1757), .Y(new_n1752));
  nor_4  g1477(.A(new_n1752), .B(new_n1751), .Y(new_n1753));
  not_3  g1478(.A(new_n1753), .Y(new_n1754));
  nand_4 g1479(.A(new_n1754), .B(new_n1750), .Y(new_n1755));
  not_3  g1480(.A(new_n1755), .Y(new_n1756));
  xnor_3 g1481(.A(new_n1753), .B(new_n1392), .Y(new_n1757_1));
  not_3  g1482(.A(new_n1752), .Y(new_n1758));
  nor_4  g1483(.A(new_n1758), .B(n839), .Y(new_n1759));
  nor_4  g1484(.A(new_n1759), .B(new_n1753), .Y(new_n1760));
  nor_4  g1485(.A(new_n1760), .B(new_n1395), .Y(new_n1761));
  not_3  g1486(.A(new_n1760), .Y(new_n1762));
  nor_4  g1487(.A(new_n1762), .B(new_n1394), .Y(new_n1763_1));
  nor_4  g1488(.A(new_n1763_1), .B(new_n1761), .Y(new_n1764_1));
  not_3  g1489(.A(new_n1764_1), .Y(new_n1765));
  not_3  g1490(.A(new_n1356), .Y(new_n1766));
  nor_4  g1491(.A(new_n1360), .B(new_n1766), .Y(new_n1767));
  nor_4  g1492(.A(new_n1767), .B(new_n1353), .Y(new_n1768));
  nor_4  g1493(.A(new_n1768), .B(new_n1765), .Y(new_n1769));
  nor_4  g1494(.A(new_n1769), .B(new_n1761), .Y(new_n1770));
  nor_4  g1495(.A(new_n1770), .B(new_n1757_1), .Y(new_n1771));
  nor_4  g1496(.A(new_n1771), .B(new_n1756), .Y(new_n1772));
  nand_4 g1497(.A(new_n1772), .B(new_n1742), .Y(new_n1773));
  not_3  g1498(.A(new_n1773), .Y(new_n1774));
  nor_4  g1499(.A(new_n1772), .B(new_n1742), .Y(new_n1775));
  nor_4  g1500(.A(new_n1775), .B(new_n1774), .Y(n891));
  not_3  g1501(.A(new_n1660_1), .Y(new_n1777));
  nor_4  g1502(.A(new_n1741), .B(new_n931_1), .Y(new_n1778));
  not_3  g1503(.A(new_n1778), .Y(new_n1779));
  nand_4 g1504(.A(new_n1773), .B(new_n1779), .Y(new_n1780));
  nor_4  g1505(.A(new_n1780), .B(new_n1777), .Y(n892));
  xor_3  g1506(.A(new_n1073), .B(new_n1071), .Y(n902));
  xor_3  g1507(.A(new_n1194_1), .B(new_n1193), .Y(n905));
  not_3  g1508(.A(new_n1174), .Y(new_n1784));
  nand_4 g1509(.A(new_n1170), .B(new_n1385_1), .Y(new_n1785));
  nand_4 g1510(.A(new_n1785), .B(new_n1166), .Y(new_n1786));
  nand_4 g1511(.A(new_n1786), .B(new_n1784), .Y(n912));
  nor_4  g1512(.A(n1149), .B(new_n593), .Y(new_n1788));
  nor_4  g1513(.A(new_n1788), .B(new_n941), .Y(n935));
  xor_3  g1514(.A(new_n1703), .B(n1119), .Y(n942));
  not_3  g1515(.A(new_n1122), .Y(new_n1791));
  xor_3  g1516(.A(new_n1125), .B(new_n1791), .Y(n944));
  nor_4  g1517(.A(new_n1175_1), .B(new_n1162_1), .Y(new_n1793));
  nand_4 g1518(.A(new_n1716), .B(new_n1793), .Y(new_n1794));
  not_3  g1519(.A(new_n1794), .Y(n974));
  not_3  g1520(.A(new_n389), .Y(new_n1796));
  xor_3  g1521(.A(new_n431), .B(new_n1796), .Y(n979));
  not_3  g1522(.A(new_n803), .Y(new_n1798));
  nor_4  g1523(.A(new_n817), .B(new_n1798), .Y(new_n1799));
  nor_4  g1524(.A(new_n816), .B(new_n804), .Y(new_n1800));
  nor_4  g1525(.A(new_n1202_1), .B(new_n1800), .Y(new_n1801));
  nor_4  g1526(.A(new_n1801), .B(new_n1799), .Y(new_n1802));
  not_3  g1527(.A(new_n1802), .Y(new_n1803));
  nor_4  g1528(.A(new_n1803), .B(new_n850), .Y(n980));
  not_3  g1529(.A(new_n1434), .Y(new_n1805));
  xor_3  g1530(.A(new_n1464), .B(new_n1805), .Y(n989));
  xor_3  g1531(.A(new_n1695), .B(new_n1671), .Y(n991));
  xor_3  g1532(.A(new_n1768), .B(new_n1764_1), .Y(n1005));
  xnor_3 g1533(.A(new_n1420), .B(new_n1397), .Y(n1012));
  xor_3  g1534(.A(new_n1168), .B(new_n1384), .Y(n1015));
  nand_4 g1535(.A(new_n1801), .B(new_n850), .Y(new_n1811));
  not_3  g1536(.A(new_n850), .Y(new_n1812));
  nand_4 g1537(.A(new_n1801), .B(new_n1799), .Y(new_n1813));
  and_4  g1538(.A(new_n1813), .B(new_n1803), .Y(new_n1814));
  not_3  g1539(.A(new_n1814), .Y(new_n1815));
  nand_4 g1540(.A(new_n1815), .B(new_n1812), .Y(new_n1816));
  nand_4 g1541(.A(new_n1816), .B(new_n1811), .Y(n1025));
  xnor_3 g1542(.A(new_n1770), .B(new_n1757_1), .Y(n1030));
  not_3  g1543(.A(new_n842), .Y(new_n1819));
  xor_3  g1544(.A(new_n1819), .B(new_n836_1), .Y(n1067));
  xnor_3 g1545(.A(new_n1780), .B(new_n1777), .Y(n1068));
  xor_3  g1546(.A(new_n586), .B(new_n583), .Y(n1103));
  xor_3  g1547(.A(new_n467), .B(new_n465), .Y(n1113));
  nor_4  g1548(.A(new_n1173), .B(new_n1487), .Y(new_n1824));
  nand_4 g1549(.A(new_n1824), .B(new_n1161_1), .Y(new_n1825));
  not_3  g1550(.A(new_n1715), .Y(new_n1826));
  nor_4  g1551(.A(new_n1826), .B(new_n806), .Y(new_n1827));
  nand_4 g1552(.A(new_n1827), .B(new_n1825), .Y(new_n1828));
  nand_4 g1553(.A(new_n1828), .B(new_n1717), .Y(n1135));
  nand_4 g1554(.A(new_n1690_1), .B(new_n1631), .Y(new_n1830));
  not_3  g1555(.A(new_n1631), .Y(new_n1831));
  nand_4 g1556(.A(new_n1691), .B(new_n1831), .Y(new_n1832));
  nand_4 g1557(.A(new_n1832), .B(new_n1830), .Y(n1142));
  not_3  g1558(.A(new_n1689), .Y(new_n1834));
  xnor_3 g1559(.A(new_n1691), .B(new_n1135_1), .Y(new_n1835));
  xnor_3 g1560(.A(new_n1835), .B(new_n1834), .Y(n1161));
  xor_3  g1561(.A(new_n1170), .B(new_n1169), .Y(n1162));
  not_3  g1562(.A(new_n1342), .Y(new_n1838));
  nor_4  g1563(.A(n865), .B(new_n1341_1), .Y(new_n1839));
  nor_4  g1564(.A(new_n1839), .B(new_n1838), .Y(n1175));
  nor_4  g1565(.A(new_n1135_1), .B(new_n819), .Y(new_n1841));
  nor_4  g1566(.A(new_n1135_1), .B(new_n824_1), .Y(new_n1842));
  and_4  g1567(.A(new_n1842), .B(new_n1725), .Y(new_n1843));
  not_3  g1568(.A(new_n1722), .Y(new_n1844));
  nand_4 g1569(.A(new_n1723), .B(new_n1844), .Y(new_n1845));
  nand_4 g1570(.A(new_n1845), .B(new_n1721_1), .Y(new_n1846));
  nor_4  g1571(.A(new_n1846), .B(new_n819), .Y(new_n1847));
  nor_4  g1572(.A(new_n1847), .B(new_n1843), .Y(new_n1848));
  nor_4  g1573(.A(new_n1848), .B(new_n1841), .Y(new_n1849));
  xnor_3 g1574(.A(new_n1849), .B(new_n1814), .Y(n1191));
  not_3  g1575(.A(new_n1172_1), .Y(new_n1851));
  xor_3  g1576(.A(new_n1851), .B(new_n1167), .Y(n1194));
  xor_3  g1577(.A(new_n429_1), .B(new_n428), .Y(n1199));
  not_3  g1578(.A(new_n1446), .Y(new_n1854));
  xor_3  g1579(.A(new_n1455), .B(new_n1854), .Y(n1201));
  not_3  g1580(.A(new_n962), .Y(new_n1856));
  nand_4 g1581(.A(new_n1323), .B(new_n1856), .Y(new_n1857));
  nand_4 g1582(.A(new_n1857), .B(new_n1327), .Y(n1202));
  xor_3  g1583(.A(n569), .B(new_n1332_1), .Y(n1234));
  xnor_3 g1584(.A(new_n1712), .B(new_n1162_1), .Y(n1235));
  not_3  g1585(.A(n1183), .Y(n1237));
  xnor_3 g1586(.A(new_n1218), .B(new_n1203), .Y(n1260));
  nor_4  g1587(.A(new_n1838), .B(n1249), .Y(new_n1863));
  nor_4  g1588(.A(new_n1863), .B(new_n1343), .Y(n1277));
  nand_4 g1589(.A(new_n1746_1), .B(new_n1742), .Y(new_n1865));
  nand_4 g1590(.A(new_n1865), .B(new_n1779), .Y(new_n1866));
  nor_4  g1591(.A(new_n1866), .B(new_n1777), .Y(n1278));
  nor_4  g1592(.A(new_n415), .B(new_n412), .Y(new_n1868));
  not_3  g1593(.A(new_n413), .Y(new_n1869));
  nor_4  g1594(.A(new_n892_1), .B(new_n1869), .Y(new_n1870));
  nor_4  g1595(.A(new_n1870), .B(new_n418), .Y(new_n1871));
  nor_4  g1596(.A(new_n1871), .B(new_n1868), .Y(n1283));
  nor_4  g1597(.A(new_n1784), .B(new_n1487), .Y(new_n1873));
  nand_4 g1598(.A(new_n1873), .B(new_n1161_1), .Y(new_n1874));
  nand_4 g1599(.A(new_n1827), .B(new_n1874), .Y(new_n1875));
  nand_4 g1600(.A(new_n1875), .B(new_n1794), .Y(n1305));
  xor_3  g1601(.A(new_n587), .B(n1727), .Y(n1315));
  not_3  g1602(.A(new_n1596), .Y(new_n1878));
  xor_3  g1603(.A(new_n1626), .B(new_n1878), .Y(n1330));
  not_3  g1604(.A(new_n1475), .Y(new_n1880));
  xor_3  g1605(.A(new_n1478), .B(new_n1880), .Y(n1338));
  not_3  g1606(.A(new_n754), .Y(new_n1882));
  xor_3  g1607(.A(new_n756), .B(new_n1882), .Y(n1340));
  not_3  g1608(.A(new_n1630), .Y(new_n1884));
  nor_4  g1609(.A(new_n1884), .B(new_n1564), .Y(new_n1885));
  nor_4  g1610(.A(new_n1885), .B(new_n1631), .Y(n1347));
  nor_4  g1611(.A(new_n1660_1), .B(new_n934), .Y(new_n1887));
  nor_4  g1612(.A(new_n1887), .B(n643), .Y(new_n1888));
  not_3  g1613(.A(new_n1888), .Y(n1348));
  not_3  g1614(.A(new_n1275), .Y(new_n1890));
  xor_3  g1615(.A(new_n1303), .B(new_n1890), .Y(n1349));
  nor_4  g1616(.A(new_n1827), .B(new_n1716), .Y(new_n1892));
  xnor_3 g1617(.A(new_n1892), .B(new_n1825), .Y(n1369));
  xnor_3 g1618(.A(new_n1892), .B(new_n1874), .Y(n1383));
  xor_3  g1619(.A(new_n1622_1), .B(new_n1611), .Y(n1393));
  not_3  g1620(.A(new_n1078), .Y(new_n1896));
  xor_3  g1621(.A(new_n1453_1), .B(new_n1896), .Y(n1399));
  xor_3  g1622(.A(new_n1191_1), .B(new_n1190), .Y(n1407));
  nor_4  g1623(.A(new_n1661), .B(new_n943), .Y(n1440));
  xor_3  g1624(.A(new_n1000_1), .B(new_n998), .Y(n1453));
  xor_3  g1625(.A(new_n1188), .B(new_n1882), .Y(n1460));
  not_3  g1626(.A(new_n1843), .Y(new_n1902));
  not_3  g1627(.A(new_n1846), .Y(new_n1903));
  nand_4 g1628(.A(new_n1903), .B(new_n1135_1), .Y(new_n1904));
  nand_4 g1629(.A(new_n1904), .B(new_n1902), .Y(new_n1905));
  xnor_3 g1630(.A(new_n1905), .B(new_n849), .Y(n1463));
  xnor_3 g1631(.A(new_n1784), .B(new_n1487), .Y(n1470));
  xor_3  g1632(.A(new_n1447), .B(new_n465), .Y(n1481));
  not_3  g1633(.A(new_n758), .Y(new_n1909));
  xor_3  g1634(.A(new_n761_1), .B(new_n1909), .Y(n1495));
  not_3  g1635(.A(new_n1061), .Y(new_n1911));
  xor_3  g1636(.A(new_n1086), .B(new_n1911), .Y(n1498));
  xor_3  g1637(.A(new_n1624), .B(new_n1604), .Y(n1502));
  not_3  g1638(.A(new_n1301), .Y(new_n1914));
  xor_3  g1639(.A(new_n1914), .B(new_n1281), .Y(n1507));
  xor_3  g1640(.A(new_n1331), .B(new_n1329), .Y(n1525));
  not_3  g1641(.A(new_n763), .Y(new_n1917));
  xor_3  g1642(.A(new_n1917), .B(new_n740), .Y(n1535));
  not_3  g1643(.A(new_n1000_1), .Y(n1601));
  xor_3  g1644(.A(n1601), .B(n1426), .Y(n1556));
  xnor_3 g1645(.A(new_n1888), .B(new_n943), .Y(n1595));
  xnor_3 g1646(.A(new_n1457_1), .B(new_n1442), .Y(n1600));
  not_3  g1647(.A(new_n528), .Y(new_n1923));
  and_4  g1648(.A(new_n573_1), .B(new_n1923), .Y(new_n1924));
  or_4   g1649(.A(new_n1924), .B(new_n575), .Y(n1613));
  xor_3  g1650(.A(new_n1297), .B(new_n1731_1), .Y(n1629));
  nor_4  g1651(.A(new_n1849), .B(new_n1802), .Y(new_n1927));
  nand_4 g1652(.A(new_n1843), .B(new_n819), .Y(new_n1928));
  nand_4 g1653(.A(new_n1928), .B(new_n1813), .Y(new_n1929));
  nor_4  g1654(.A(new_n1929), .B(new_n1927), .Y(n1633));
  xor_3  g1655(.A(new_n1001), .B(new_n997), .Y(n1635));
  xor_3  g1656(.A(new_n1416), .B(new_n1414), .Y(n1654));
  nor_4  g1657(.A(new_n589), .B(n1138), .Y(new_n1933));
  nor_4  g1658(.A(new_n1933), .B(new_n591), .Y(n1657));
  xnor_3 g1659(.A(new_n1866), .B(new_n1777), .Y(n1660));
  xor_3  g1660(.A(new_n1081), .B(new_n1896), .Y(n1675));
  xnor_3 g1661(.A(new_n1643_1), .B(new_n1655), .Y(n1686));
  xor_3  g1662(.A(new_n1184), .B(new_n465), .Y(n1688));
  xnor_3 g1663(.A(new_n1628), .B(new_n1586), .Y(n1690));
  xnor_3 g1664(.A(new_n1685), .B(new_n1673), .Y(n1729));
  xnor_3 g1665(.A(new_n1645), .B(new_n1203), .Y(n1737));
  not_3  g1666(.A(new_n1408), .Y(new_n1942));
  xor_3  g1667(.A(new_n1411), .B(new_n1942), .Y(n1746));
  xor_3  g1668(.A(new_n404), .B(n347), .Y(n488));
  xor_3  g1669(.A(new_n1199_1), .B(new_n986), .Y(n1677));
endmodule


