
module top_810222779_843330999_776144567_776418743_1234615 (n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82, n86, n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200, n219, n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273, n284, n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341, n344, n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420, n430, n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560, n561, n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609, n626, n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729, n734, n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831, n832, n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961, n969, n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061, n1071, n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164, n1172, n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246, n1250, n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305, n1345, n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411, n1415, n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470, n1474, n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536, n1566, n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627, n1644, n1647, n1656, n1750, n1753, n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181, n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362, n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501, n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669, n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918, n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063, n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285, n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368, n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588, n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752);
input n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82, n86, n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200, n219, n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273, n284, n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341, n344, n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420, n430, n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560, n561, n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609, n626, n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729, n734, n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831, n832, n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961, n969, n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061, n1071, n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164, n1172, n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246, n1250, n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305, n1345, n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411, n1415, n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470, n1474, n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536, n1566, n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627, n1644, n1647, n1656, n1750, n1753;
output n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181, n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362, n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501, n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669, n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918, n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063, n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285, n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368, n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588, n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752;
wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n12, n13, n14, n15, n16, n17, n18, n19, n20, n24, n25, n26, n28, n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42, n43, n44, n46, n47, n48, n49, n51, n53, n55, n57, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n78, n79, n80, n81, n83, n84, n88, n89, n90, n91, n92, n93, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n108, n109, n110, n111, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123, n124, n125, n127, n128, n129, n131, n132, n133, n134, n135, n136, n137, n139, n140, n141, n142, n144, n145, n146, n147, n148, n149, n150, n151, n152, n154, n157, n158, n160, n162, n163, n165, n166, n167, n168, n169, n170, n171, n172, n174, n175, n176, n177, n178, n179, n180, n182, n183, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n217, n218, n221, n224, n225, n226, n227, n228, n229, n231, n232, n234, n235, n236, n237, n238, n239, n240, n241, n242, n245, n248, n249, n250, n252, n253, n255, n256, n257, n258, n259, n260, n261, n263, n264, n265, n266, n267, n269, n270, n271, n272, n274, n276, n277, n278, n279, n280, n281, n282, n283, n285, n286, n287, n289, n290, n291, n294, n295, n296, n297, n298, n302, n303, n305, n306, n308, n309, n311, n313, n316, n317, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n342, n343, n345, n347, n348, n349, n350, n351, n353, n354, n355, n356, n357, n358, n359, n360, n361, n363, n365, n366, n367, n368, n369, n371, n372, n373, n375, n377, n379, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n393, n394, n395, n397, n398, n400, n401, n402, n403, n404, n405, n406, n407, n410, n411, n412, n413, n414, n415, n418, n419, n421, n422, n423, n424, n425, n426, n427, n429, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n454, n455, n456, n458, n459, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n479, n480, n481, n482, n483, n484, n485, n486, n488, n490, n491, n492, n493, n494, n495, n496, n499, n500, n503, n504, n505, n508, n511, n512, n513, n514, n515, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n546, n547, n548, n549, n550, n551, n552, n554, n555, n556, n557, n558, n562, n563, n564, n565, n566, n568, n569, n570, n571, n572, n573, n575, n576, n577, n578, n579, n580, n583, n584, n586, n587, n588, n590, n591, n592, n594, n596, n599, n601, n602, n603, n604, n605, n606, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n639, n642, n643, n644, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n664, n665, n666, n667, n668, n670, n672, n673, n674, n675, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n691, n692, n694, n696, n697, n698, n699, n700, n702, n703, n704, n705, n706, n707, n708, n709, n711, n712, n713, n715, n716, n717, n718, n720, n721, n722, n723, n724, n725, n728, n730, n731, n732, n733, n735, n736, n737, n738, n739, n740, n741, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n770, n771, n772, n774, n776, n777, n780, n781, n783, n784, n785, n786, n788, n789, n791, n792, n793, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n822, n824, n825, n826, n827, n828, n829, n830, n833, n834, n835, n836, n837, n838, n840, n841, n843, n844, n845, n846, n847, n848, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n880, n881, n883, n884, n886, n887, n888, n889, n890, n891, n892, n893, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n917, n919, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n948, n949, n950, n951, n954, n955, n956, n957, n958, n959, n960, n962, n963, n964, n965, n966, n967, n968, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n981, n982, n983, n985, n987, n988, n989, n991, n993, n994, n995, n996, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1018, n1019, n1020, n1021, n1022, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1041, n1043, n1045, n1046, n1047, n1048, n1049, n1052, n1053, n1055, n1056, n1057, n1059, n1062, n1064, n1066, n1067, n1068, n1069, n1070, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1115, n1116, n1117, n1118, n1119, n1120, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1153, n1155, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1173, n1174, n1176, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1188, n1189, n1190, n1192, n1194, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1206, n1207, n1208, n1210, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1226, n1228, n1229, n1230, n1232, n1233, n1235, n1236, n1237, n1238, n1240, n1241, n1242, n1243, n1244, n1245, n1247, n1248, n1249, n1251, n1252, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1279, n1280, n1282, n1284, n1287, n1290, n1291, n1293, n1294, n1295, n1297, n1298, n1300, n1303, n1304, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1321, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1347, n1348, n1349, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1360, n1362, n1363, n1364, n1365, n1366, n1367, n1369, n1370, n1371, n1372, n1373, n1374, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1388, n1390, n1392, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1412, n1413, n1414, n1416, n1417, n1419, n1422, n1423, n1424, n1425, n1426, n1429, n1430, n1431, n1432, n1433, n1434, n1436, n1437, n1439, n1440, n1441, n1442, n1444, n1445, n1447, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1464, n1465, n1466, n1467, n1468, n1469, n1471, n1472, n1473, n1475, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1501, n1503, n1504, n1505, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1517, n1518, n1519, n1522, n1524, n1525, n1526, n1528, n1529, n1530, n1531, n1532, n1533, n1535, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1567, n1568, n1570, n1571, n1572, n1573, n1574, n1575, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1587, n1589, n1590, n1591, n1593, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1610, n1611, n1612, n1614, n1615, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1628, n1629, n1630, n1631, n1633, n1634, n1635, n1636, n1637, n1638, n1640, n1641, n1642, n1643, n1646, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1751, n1754, n1755, n1756;
assign n426 = n422 | n1543;
assign n1664 = n889 | n1101;
assign n1637 = ~(n456 ^ n1142);
assign n1067 = ~(n1402 ^ n145);
assign n993 = ~(n780 ^ n1263);
assign n1517 = n206 ^ n1725;
assign n1735 = n1116 | n1429;
assign n1539 = n1683 & n1276;
assign n154 = ~n1002;
assign n1347 = ~(n142 | n1105);
assign n1537 = ~n1540;
assign n1608 = ~(n1573 ^ n866);
assign n960 = ~n1377;
assign n476 = n768 & n1126;
assign n805 = n1485 | n192;
assign n752 = ~(n88 ^ n540);
assign n1048 = ~n654;
assign n1698 = ~(n1343 | n109);
assign n1326 = ~(n289 | n1230);
assign n721 = ~n728;
assign n1555 = ~n886;
assign n1578 = n1194 | n25;
assign n1383 = n802 | n218;
assign n821 = n374;
assign n802 = ~n837;
assign n103 = n1706 | n1557;
assign n175 = n717 | n943;
assign n468 = ~n1419;
assign n38 = ~(n1207 ^ n557);
assign n1585 = n1115 | n238;
assign n1105 = n1416 | n467;
assign n1648 = n935 | n266;
assign n165 = ~n1664;
assign n212 = n1721 | n500;
assign n624 = n885 & n197;
assign n1218 = n986 & n0;
assign n1002 = n228 | n1551;
assign n256 = n1357 | n1533;
assign n102 = n1531 | n686;
assign n1617 = ~(n1373 ^ n1417);
assign n123 = ~(n1512 ^ n1355);
assign n272 = n1100 & n177;
assign n305 = n1481 | n272;
assign n104 = ~(n721 | n1401);
assign n973 = n1408 | n379;
assign n70 = ~n923;
assign n1365 = ~n1506;
assign n1316 = ~(n632 ^ n1595);
assign n1015 = n376 & n1168;
assign n1302 = ~(n837 ^ n933);
assign n1480 = n779 & n721;
assign n1719 = n251 & n1555;
assign n1188 = n1268 | n1458;
assign n148 = ~(n721 | n1138);
assign n436 = ~(n777 ^ n194);
assign n1247 = ~(n1037 ^ n72);
assign n747 = ~n1708;
assign n579 = ~n1293;
assign n1556 = ~(n723 ^ n518);
assign n471 = n1558 & n1312;
assign n327 = ~n843;
assign n846 = ~n324;
assign n1488 = ~(n623 ^ n1382);
assign n1237 = ~(n380 & n701);
assign n785 = n63 & n807;
assign n1370 = n559 & n491;
assign n388 = ~n1559;
assign n658 = n1696 | n835;
assign n914 = ~n1387;
assign n331 = ~(n1107 ^ n1707);
assign n1212 = ~(n999 ^ n24);
assign n1623 = ~n891;
assign n488 = ~(n1535 | n1628);
assign n681 = n1172 & n602;
assign n1017 = n1476;
assign n298 = ~n1521;
assign n923 = n1692 & n474;
assign n670 = ~n626;
assign n554 = n134 & n1400;
assign n1515 = ~n1008;
assign n1325 = n1579 | n423;
assign n1201 = n1623 | n1511;
assign n549 = ~(n63 | n32);
assign n1158 = n1241 | n1354;
assign n197 = ~n1314;
assign n861 = n64 | n1244;
assign n801 = ~(n1615 | n1336);
assign n151 = n312 & n1458;
assign n516 = n1187;
assign n1075 = n124 & n1482;
assign n946 = n568 | n999;
assign n1525 = ~(n1339 ^ n615);
assign n587 = ~(n1734 | n772);
assign n1179 = ~n545;
assign n686 = ~(n1178 | n175);
assign n1465 = n1254 | n1167;
assign n1477 = n89 & n495;
assign n1687 = n523 | n73;
assign n1538 = n1013 | n444;
assign n1355 = ~n188;
assign n1736 = n687 | n979;
assign n1119 = ~(n257 | n200);
assign n26 = ~n778;
assign n1714 = ~(n1445 ^ n1084);
assign n1658 = n1261 | n10;
assign n1596 = n1393 & n530;
assign n1673 = ~n993;
assign n1743 = n359 | n434;
assign n1335 = ~(n1686 | n1073);
assign n1612 = ~(n721 | n56);
assign n1458 = ~n808;
assign n182 = n1346 & n602;
assign n1468 = ~(n1597 ^ n980);
assign n195 = n1251 & n1598;
assign n1307 = ~(n1273 ^ n427);
assign n324 = ~(n1721 ^ n732);
assign n828 = n1752 | n493;
assign n958 = n1673 & n798;
assign n301 = n318;
assign n316 = ~n1201;
assign n174 = ~(n1597 ^ n923);
assign n119 = ~n567;
assign n124 = n395 & n1034;
assign n460 = n21;
assign n1496 = ~(n1049 ^ n630);
assign n1214 = ~n339;
assign n504 = ~(n49 ^ n1406);
assign n1107 = ~(n83 ^ n724);
assign n811 = ~n1475;
assign n1189 = n2 & n323;
assign n17 = ~n865;
assign n474 = n803 | n905;
assign n1084 = ~(n1648 ^ n1018);
assign n1287 = ~(n261 ^ n1727);
assign n252 = ~(n522 | n132);
assign n760 = n1230 & n873;
assign n1497 = n721 | n346;
assign n606 = ~(n1537 ^ n60);
assign n481 = n1182 | n1238;
assign n306 = n1577 | n1203;
assign n99 = ~(n1535 ^ n1442);
assign n35 = n636 | n1620;
assign n1394 = ~n1681;
assign n1099 = n1489 | n806;
assign n1306 = n1204 | n1619;
assign n302 = ~(n1173 ^ n608);
assign n1600 = ~(n32 ^ n1473);
assign n308 = ~n1239;
assign n611 = ~(n1166 ^ n1699);
assign n1058 = ~(n1667 ^ n810);
assign n687 = ~n1711;
assign n1430 = ~n307;
assign n414 = ~(n1470 | n910);
assign n1511 = ~n907;
assign n340 = n613 & n698;
assign n1621 = n934 & n1697;
assign n1532 = ~(n1667 | n840);
assign n1404 = n133 ^ n375;
assign n921 = n1644 & n1136;
assign n835 = ~n413;
assign n1395 = ~n738;
assign n1072 = ~(n899 ^ n938);
assign n492 = ~(n900 | n86);
assign n637 = n1672 & n1475;
assign n213 = n142 ^ n1083;
assign n1269 = ~(n999 | n703);
assign n999 = ~n1419;
assign n373 = ~(n740 ^ n407);
assign n1170 = n903 | n694;
assign n271 = n1750 & n238;
assign n177 = ~(n1230 | n1335);
assign n1689 = ~(n1200 ^ n707);
assign n1282 = n454 | n639;
assign n1235 = n1722 | n649;
assign n900 = ~n413;
assign n1747 = n1102 | n75;
assign n1148 = n798 | n1390;
assign n96 = n687 | n1139;
assign n140 = n651 & n248;
assign n1194 = ~(n1099 | n189);
assign n635 = n1668 | n197;
assign n137 = n1415 & n530;
assign n1018 = n479 & n840;
assign n530 = ~n808;
assign n1085 = n899 & n1264;
assign n1162 = n803 | n1191;
assign n357 = ~(n367 | n158);
assign n91 = n985 | n443;
assign n1083 = n1015 | n804;
assign n1091 = ~(n876 ^ n33);
assign n367 = n1360 & n575;
assign n1274 = n1698 | n1075;
assign n379 = n964 | n717;
assign n1229 = ~(n922 ^ n1651);
assign n1126 = ~n852;
assign n1197 = ~n179;
assign n962 = ~(n1686 ^ n1498);
assign n47 = n1083 & n1492;
assign n1113 = ~n1188;
assign n1457 = ~(n206 ^ n1343);
assign n1155 = n1405 | n567;
assign n866 = ~(n654 ^ n1629);
assign n1353 = n204 | n577;
assign n537 = n1291 | n1098;
assign n1618 = n761 | n465;
assign n1397 = n219 & n1168;
assign n758 = ~n565;
assign n1582 = ~(n1641 ^ n1476);
assign n1272 = ~(n146 | n481);
assign n592 = n760 | n1327;
assign n1226 = n1585 & n569;
assign n1642 = n1561 | n250;
assign n1380 = ~(n1573 ^ n1133);
assign n1132 = ~(n324 | n241);
assign n1135 = ~n888;
assign n746 = n1493 | n503;
assign n1320 = n1263;
assign n100 = ~(n354 | n1137);
assign n1009 = ~(n1340 ^ n1636);
assign n259 = ~n908;
assign n719 = n1361 | n1225;
assign n245 = ~(n803 | n769);
assign n486 = n614 | n1012;
assign n1604 = ~(n572 | n1682);
assign n525 = ~(n1673 ^ n1148);
assign n1056 = ~(n555 ^ n730);
assign n9 = ~n1284;
assign n1738 = n45;
assign n718 = n629 | n636;
assign n266 = n1552 | n1222;
assign n120 = n1288 | n1322;
assign n807 = n1136 | n1435;
assign n1565 = ~n1747;
assign n812 = n1623 ^ n907;
assign n874 = ~(n1535 | n1695);
assign n1190 = n695 | n653;
assign n646 = ~(n852 | n1436);
assign n1133 = n883 | n1048;
assign n229 = n793 | n59;
assign n383 = ~(n948 ^ n1148);
assign n1709 = n849 & n776;
assign n1358 = n1700 | n212;
assign n1215 = ~(n1601 | n998);
assign n348 = ~n1307;
assign n731 = ~n1694;
assign n1716 = n1304 | n333;
assign n798 = n249 & n1129;
assign n1381 = ~n1043;
assign n1493 = ~n225;
assign n180 = ~n1386;
assign n1399 = n930 & n655;
assign n1740 = n824 | n618;
assign n777 = n137 | n207;
assign n1315 = n1328 | n900;
assign n1513 = ~(n1405 | n823);
assign n199 = n915 | n257;
assign n1267 = n416 & n444;
assign n239 = ~n50;
assign n48 = ~(n613 ^ n405);
assign n800 = ~(n318 | n781);
assign n1033 = n514 | n989;
assign n738 = n682 | n668;
assign n536 = n790 & n240;
assign n551 = ~n1007;
assign n93 = ~(n899 ^ n960);
assign n639 = n1657 | n403;
assign n1037 = ~(n469 ^ n1055);
assign n511 = n637 & n1078;
assign n326 = n1333 | n1150;
assign n1297 = ~n1077;
assign n1741 = n1141 | n1731;
assign n80 = ~n938;
assign n1243 = n47 | n1022;
assign n1624 = n838 | n983;
assign n240 = ~n808;
assign n483 = n238 | n839;
assign n1718 = n5 | n1722;
assign n303 = n691 & n639;
assign n134 = ~n1261;
assign n1016 = n755 & n721;
assign n1150 = ~n668;
assign n422 = ~(n675 ^ n1398);
assign n817 = ~(n736 | n1422);
assign n88 = n20 | n864;
assign n1482 = n170 | n1545;
assign n1599 = ~n887;
assign n963 = n1461 | n444;
assign n1106 = n119 & n1002;
assign n230 = n831;
assign n1526 = ~(n630 | n1355);
assign n1570 = n1673 & n1390;
assign n1661 = ~(n99 ^ n129);
assign n242 = ~(n1637 ^ n606);
assign n1324 = ~n1396;
assign n1043 = n1724 | n386;
assign n509 = n769;
assign n1614 = n1298 | n1394;
assign n249 = ~n1116;
assign n1437 = n1542 | n875;
assign n378 = ~(n224 ^ n211);
assign n1087 = ~(n721 | n1502);
assign n1221 = ~(n1438 & n1536);
assign n437 = ~(n1220 ^ n394);
assign n1427 = n1407 | n1562;
assign n235 = n1377 | n1756;
assign n570 = ~(n708 ^ n948);
assign n1375 = n229 | n770;
assign n1455 = n1004 & n1044;
assign n90 = ~(n265 ^ n24);
assign n1486 = ~n1635;
assign n227 = n150 | n1290;
assign n1094 = n1319 & n205;
assign n1384 = n309 | n444;
assign n749 = ~n419;
assign n1417 = ~(n1303 ^ n1641);
assign n883 = ~n1629;
assign n1045 = ~(n43 ^ n33);
assign n387 = n217 | n877;
assign n820 = ~n203;
assign n1314 = ~n263;
assign n1144 = ~n212;
assign n466 = n441 | n636;
assign n950 = n1692 & n483;
assign n655 = n971 | n530;
assign n112 = ~(n42 ^ n907);
assign n794 = ~(n225 ^ n1208);
assign n167 = n238 | n222;
assign n1251 = n1293 | n708;
assign n1019 = n651 | n527;
assign n1396 = n100 & n1666;
assign n660 = n676 & n197;
assign n1078 = n248 & n527;
assign n135 = ~n1073;
assign n1051 = ~(n689 ^ n168);
assign n496 = n564 & n473;
assign n1339 = ~(n66 ^ n336);
assign n1629 = n2 | n684;
assign n1177 = n487;
assign n1639 = ~(n302 ^ n801);
assign n465 = n1152 & n491;
assign n433 = ~(n315 & n997);
assign n677 = n1648 | n1232;
assign n1011 = n1513 | n1426;
assign n740 = n1309 | n1742;
assign n1321 = ~n691;
assign n534 = ~(n248 ^ n472);
assign n515 = n579 | n706;
assign n386 = ~n1174;
assign n1459 = ~(n321 ^ n1507);
assign n490 = n1029 | n748;
assign n519 = n1682 & n994;
assign n1060 = n762 | n1702;
assign n850 = ~n1061;
assign n803 = ~n413;
assign n14 = ~n1279;
assign n1151 = n868 | n212;
assign n1501 = n1140 | n148;
assign n429 = ~n1629;
assign n1700 = ~n1582;
assign n231 = n565 & n1150;
assign n463 = n836 | n240;
assign n32 = n884 | n745;
assign n1527 = ~(n311 ^ n1706);
assign n768 = n214 & n981;
assign n1219 = ~n561;
assign n406 = n845 | n1070;
assign n662 = n282 | n496;
assign n943 = n1491 | n1722;
assign n1035 = n732 & n340;
assign n451 = n979 | n647;
assign n1454 = ~(n1742 | n1035);
assign n1349 = n1630 | n1405;
assign n228 = n268 & n1168;
assign n926 = n1413 | n356;
assign n991 = n1059 & n946;
assign n928 = ~(n1089 | n787);
assign n1216 = n1057 | n226;
assign n1597 = n1692 & n1509;
assign n1522 = n1103 & n491;
assign n292 = n408;
assign n1462 = ~(n1572 ^ n769);
assign n858 = ~(n490 | n1229);
assign n359 = n1216 | n932;
assign n419 = n591 | n530;
assign n221 = ~n605;
assign n867 = n1555 & n117;
assign n442 = ~(n1515 ^ n1487);
assign n765 = n774 | n982;
assign n533 = n1367 | n149;
assign n1142 = ~(n371 ^ n1665);
assign n784 = ~n1648;
assign n1020 = n906 & n1371;
assign n1607 = n679 | n389;
assign n41 = n721 | n223;
assign n1117 = ~(n408 | n704);
assign n1602 = n63 & n1374;
assign n1007 = n1349 & n1077;
assign n717 = ~(n1402 ^ n895);
assign n1086 = n1479 | n738;
assign n1228 = n84 & n777;
assign n289 = n811 | n1432;
assign n1708 = n529 | n1555;
assign n1715 = ~n1064;
assign n697 = n1493 | n677;
assign n121 = ~(n1623 ^ n739);
assign n1694 = ~(n841 ^ n1470);
assign n1080 = ~(n994 | n242);
assign n1467 = n1655 | n1119;
assign n69 = n1049 | n368;
assign n1655 = n589 & n835;
assign n989 = ~(n1399 | n452);
assign n1734 = ~(n1232 ^ n225);
assign n809 = ~(n1493 | n435);
assign n588 = ~(n18 | n1726);
assign n1076 = ~n1250;
assign n1169 = ~(n321 ^ n1336);
assign n1357 = ~n1432;
assign n1434 = ~(n1535 | n659);
assign n653 = n1528 & n1703;
assign n25 = ~(n144 | n306);
assign n956 = ~(n1364 | n901);
assign n930 = n238 | n1071;
assign n1323 = n40 & n257;
assign n364 = n1477 | n1508;
assign n1407 = n1212 & n1650;
assign n1279 = ~(n1530 ^ n138);
assign n183 = ~(n741 | n891);
assign n1484 = n467 | n363;
assign n1483 = ~(n1159 ^ n610);
assign n682 = n545 & n758;
assign n564 = ~n479;
assign n139 = ~n78;
assign n187 = ~(n38 ^ n1009);
assign n142 = n735 & n887;
assign n772 = ~(n859 ^ n825);
assign n661 = ~(n803 | n94);
assign n1028 = n921 | n1541;
assign n126 = n1449 | n566;
assign n12 = ~(n236 ^ n1496);
assign n869 = n1127 | n197;
assign n1543 = ~(n1659 ^ n111);
assign n1332 = n1379 | n578;
assign n1340 = ~(n874 ^ n1635);
assign n735 = n524 | n257;
assign n1173 = n1553 | n198;
assign n443 = ~(n1575 | n402);
assign n913 = n1106 | n1559;
assign n1727 = n949 ^ n857;
assign n896 = ~n1734;
assign n269 = ~n750;
assign n253 = ~(n1537 | n1307);
assign n1240 = n689 & n576;
assign n1545 = n169 | n1728;
assign n1196 = n1021 ^ n1301;
assign n659 = ~(n1405 | n1389);
assign n484 = ~n1202;
assign n250 = n1193 & n491;
assign n427 = ~(n470 ^ n157);
assign n819 = n159 & n835;
assign n390 = ~(n1026 | n340);
assign n190 = ~n1627;
assign n1253 = n1050;
assign n369 = ~(n66 ^ n172);
assign n1293 = n980 | n358;
assign n1166 = ~(n1249 ^ n957);
assign n683 = n1126 & n1204;
assign n333 = n1121 & n491;
assign n89 = ~(n249 ^ n327);
assign n1184 = n1672 & n1634;
assign n448 = n98 | n1383;
assign n505 = n976 | n1705;
assign n774 = ~(n205 | n1390);
assign n542 = ~(n654 ^ n1380);
assign n754 = ~(n752 ^ n851);
assign n602 = ~n413;
assign n1590 = n1483 | n1030;
assign n461 = ~n302;
assign n753 = ~(n543 ^ n1716);
assign n1414 = n446 & n476;
assign n0 = n627 | n1341;
assign n750 = n1210 | n747;
assign n1273 = ~(n1604 ^ n505);
assign n1392 = n1275 | n1046;
assign n1128 = ~(n896 | n783);
assign n211 = n1080 | n1621;
assign n815 = n1649 | n1088;
assign n1693 = ~(n1217 | n911);
assign n1571 = n879 & n900;
assign n573 = n1007 | n145;
assign n1717 = n1200 & n1664;
assign n1079 = ~n538;
assign n906 = ~n1733;
assign n181 = ~(n1468 ^ n1505);
assign n804 = n262 & n602;
assign n42 = ~n1743;
assign n512 = n369 | n1271;
assign n20 = n1419 & n237;
assign n1490 = n1518 | n1053;
assign n1171 = ~(n1260 ^ n1725);
assign n1070 = n409 & n1136;
assign n557 = ~(n1530 ^ n841);
assign n698 = n1324 | n61;
assign n377 = n1414 | n583;
assign n1507 = ~(n302 ^ n473);
assign n1622 = ~n941;
assign n1460 = ~(n811 | n1079);
assign n23 = n346;
assign n863 = n835 | n1500;
assign n957 = n653 ^ n972;
assign n97 = n1189 | n449;
assign n1534 = n920;
assign n616 = n687 | n979;
assign n418 = ~(n471 ^ n332);
assign n893 = ~(n1700 ^ n339);
assign n1676 = n1660 | n681;
assign n1568 = ~n1476;
assign n1050 = n1361 | n1237;
assign n771 = n1144 | n1579;
assign n651 = n287 & n1382;
assign n1352 = ~n972;
assign n129 = ~(n1434 ^ n488);
assign n432 = ~(n1135 | n265);
assign n618 = n87 & n602;
assign n709 = n110 | n377;
assign n908 = n1739 | n1116;
assign n813 = ~(n721 | n775);
assign n578 = ~n635;
assign n1236 = n531 | n1701;
assign n736 = n1190 | n1493;
assign n49 = n1180 & n163;
assign n1359 = ~(n654 ^ n901);
assign n1270 = n313 | n105;
assign n877 = n1276 & n757;
assign n1160 = ~(n570 | n1505);
assign n1318 = n668 & n754;
assign n363 = ~(n1416 ^ n142);
assign n1531 = ~(n573 | n759);
assign n1681 = n1560 & n1025;
assign n940 = ~(n579 ^ n756);
assign n886 = ~n728;
assign n1124 = ~(n257 | n1616);
assign n85 = n153;
assign n1207 = ~(n1317 ^ n1572);
assign n1542 = ~(n644 | n1484);
assign n1475 = ~(n1392 ^ n1592);
assign n619 = n107 & n1206;
assign n711 = ~(n1574 | n1650);
assign n1248 = n1321 | n1217;
assign n295 = n1396 & n326;
assign n766 = ~(n1019 ^ n203);
assign n53 = n1591 | n1478;
assign n173 = n823;
assign n384 = ~(n471 ^ n68);
assign n36 = n1681 & n1539;
assign n263 = ~n308;
assign n907 = ~(n750 ^ n293);
assign n297 = n345 | n384;
assign n558 = ~n977;
assign n844 = ~n1468;
assign n909 = n26 | n238;
assign n873 = n858 | n978;
assign n517 = n398 | n1198;
assign n751 = ~(n1021 ^ n725);
assign n453 = n1359;
assign n925 = ~n248;
assign n623 = n258 | n1113;
assign n1487 = n271 | n51;
assign n1029 = n1184 | n1153;
assign n208 = ~(n478 & n1095);
assign n672 = n468 & n322;
assign n767 = ~(n580 ^ n1043);
assign n1518 = n361 | n1272;
assign n1654 = n19 | n1098;
assign n1529 = n199 & n1451;
assign n72 = ~(n929 ^ n650);
assign n713 = n36 | n387;
assign n636 = ~(n133 ^ n857);
assign n464 = ~(n868 | n829);
assign n19 = ~(n353 ^ n1291);
assign n237 = ~(n722 ^ n222);
assign n1046 = ~n1310;
assign n351 = ~n613;
assign n825 = ~(n8 ^ n1262);
assign n1704 = n902 & n1650;
assign n68 = n909 & n1703;
assign n1595 = n1447 | n819;
assign n1588 = n956 | n1334;
assign n783 = ~n772;
assign n1453 = ~n441;
assign n786 = ~(n7 | n911);
assign n366 = n776 | n608;
assign n878 = n1041 & n899;
assign n1669 = n1713 & n1269;
assign n1294 = ~n1251;
assign n1062 = n900 | n727;
assign n1178 = n614 | n649;
assign n1258 = n1378 | n1348;
assign n1678 = n988 | n1743;
assign n945 = n508 | n1460;
assign n1304 = n1222 & n314;
assign n797 = ~n33;
assign n270 = n837 & n519;
assign n1697 = ~(n911 | n253);
assign n1587 = n1375 | n120;
assign n1112 = ~n945;
assign n583 = n446 & n646;
assign n44 = ~(n1583 ^ n856);
assign n1649 = ~(n721 | n399);
assign n1643 = ~(n636 | n1409);
assign n604 = n977 & n1756;
assign n995 = ~(n201 | n1395);
assign n8 = n784 | n321;
assign n792 = ~n1572;
assign n81 = n1120 | n994;
assign n1322 = n1590 | n426;
assign n446 = ~n28;
assign n205 = ~n993;
assign n428 = n1588;
assign n1755 = ~(n602 | n45);
assign n555 = n1331 | n1601;
assign n74 = ~n1226;
assign n1466 = n254 & n491;
assign n1561 = n1289 & n197;
assign n1632 = n1186;
assign n133 = n853 & n959;
assign n1254 = n673 & n1224;
assign n1422 = n461 | n1667;
assign n1611 = n1199 | n325;
assign n1424 = ~(n603 | n715);
assign n1111 = ~n489;
assign n854 = n1720 | n39;
assign n657 = n669 | n126;
assign n1042 = n1566;
assign n360 = n672 | n1395;
assign n493 = n1594 | n1587;
assign n540 = ~(n888 ^ n134);
assign n22 = n1027 | n1549;
assign n255 = ~(n1054 & n1040);
assign n322 = n568 & n703;
assign n1514 = n598 & n444;
assign n216 = ~(n1462 ^ n1746);
assign n708 = ~n706;
assign n757 = n462 | n1;
assign n902 = ~(n1311 ^ n991);
assign n725 = n660 | n1599;
assign n1089 = ~n1388;
assign n1598 = n515 & n495;
assign n1082 = ~(n611 ^ n1109);
assign n935 = ~n612;
assign n1729 = n138;
assign n1153 = n140 & n637;
assign n43 = n624 | n250;
assign n576 = n311 & n789;
assign n726 = n1296;
assign n903 = n1652 & n1708;
assign n1410 = ~(n613 ^ n968);
assign n1505 = ~n982;
assign n92 = ~(n513 ^ n90);
assign n1580 = ~(n587 | n1554);
assign n723 = n1579 ^ n1026;
assign n1285 = n1401;
assign n440 = ~(n846 | n1610);
assign n1102 = ~n984;
assign n884 = ~(n602 | n1656);
assign n1653 = ~(n1135 | n1125);
assign n585 = n553;
assign n281 = ~n295;
assign n319 = ~(n593 & n1286);
assign n445 = n1523 & n900;
assign n501 = n200;
assign n1257 = n1656 | n1486;
assign n450 = n1047 | n528;
assign n1665 = ~(n1694 ^ n1279);
assign n1141 = ~(n1196 | n342);
assign n356 = ~(n49 | n1718);
assign n528 = ~(n1248 | n320);
assign n186 = n19 | n1199;
assign n834 = n302 & n496;
assign n818 = n172 ^ n1456;
assign n330 = ~(n14 | n1284);
assign n122 = ~(n1640 | n718);
assign n791 = ~n998;
assign n28 = n1235 | n486;
assign n1450 = ~n742;
assign n597 = ~(n1179 ^ n321);
assign n1337 = n1138;
assign n402 = n1499 | n466;
assign n1031 = n34 | n1168;
assign n875 = ~(n974 | n1170);
assign n1010 = n303 | n160;
assign n656 = n190 | n1168;
assign n1110 = ~n323;
assign n495 = ~n982;
assign n1130 = ~(n79 ^ n535);
assign n1385 = n1596 | n1466;
assign n146 = n632 | n763;
assign n1198 = ~(n1072 | n42);
assign n1261 = ~(n154 ^ n567);
assign n1104 = ~n138;
assign n1485 = n1163 | n826;
assign n210 = n926 | n252;
assign n888 = ~(n1740 ^ n374);
assign n1619 = ~(n28 | n1754);
assign n898 = n68 ^ n406;
assign n796 = ~n243;
assign n1165 = ~n950;
assign n780 = ~n880;
assign n24 = ~n568;
assign n1147 = n1550 | n629;
assign n704 = ~n1303;
assign n1489 = n1535 | n928;
assign n1367 = ~(n769 | n792);
assign n497 = n1656;
assign n1351 = n1694 & n39;
assign n841 = n63 & n382;
assign n1402 = n1680 & n656;
assign n1711 = ~(n74 ^ n1344);
assign n904 = n558 & n960;
assign n584 = n471 | n647;
assign n1579 = n870 | n601;
assign n890 = ~n671;
assign n793 = ~(n1287 ^ n1661);
assign n168 = ~(n1228 | n576);
assign n538 = n140 | n1078;
assign n1266 = ~n1616;
assign n62 = ~n506;
assign n795 = ~(n385 ^ n92);
assign n688 = ~(n545 | n264);
assign n531 = n562 & n1356;
assign n277 = ~(n1577 ^ n815);
assign n629 = ~(n949 ^ n375);
assign n1328 = ~n1114;
assign n1115 = ~n392;
assign n1341 = ~n487;
assign n1720 = n1104 & n1530;
assign n304 = n420 & n832;
assign n543 = ~n1529;
assign n1131 = ~n1717;
assign n1309 = ~n500;
assign n164 = ~(n1672 ^ n482);
assign n739 = n37 & n1511;
assign n1161 = n1136 | n980;
assign n876 = n1093 & n1384;
assign n527 = n1228 & n689;
assign n264 = ~(n1714 ^ n954);
assign n1074 = ~n1283;
assign n901 = n639 | n1693;
assign n513 = n237 ^ n468;
assign n548 = n847 | n1222;
assign n983 = ~(n335 | n1663);
assign n523 = ~(n276 | n1134);
assign n762 = ~(n183 | n1678);
assign n467 = ~(n1083 ^ n1492);
assign n1635 = n1692 & n1372;
assign n565 = n1422 | n746;
assign n1343 = n658 & n869;
assign n1090 = ~(n1291 ^ n1165);
assign n191 = ~n604;
assign n703 = ~n237;
assign n149 = n586 & n1462;
assign n569 = n193 | n1222;
assign n613 = ~(n543 ^ n1401);
assign n401 = ~n589;
assign n675 = ~(n1546 ^ n1091);
assign n413 = ~n308;
assign n978 = n490 & n158;
assign n1097 = n1377 | n1201;
assign n345 = ~n101;
assign n415 = n958 & n490;
assign n1680 = n1089 | n153;
assign n1737 = ~(n785 ^ n1392);
assign n1030 = ~(n285 ^ n215);
assign n1731 = n899 & n499;
assign n1260 = n1605 | n618;
assign n918 = n657 | n828;
assign n700 = n1223 | n279;
assign n1159 = ~(n1404 ^ n1233);
assign n127 = ~(n1733 | n1000);
assign n518 = ~(n1742 ^ n893);
assign n939 = ~n1018;
assign n2 = ~n986;
assign n837 = ~(n1317 ^ n626);
assign n673 = ~n698;
assign n1388 = ~n1314;
assign n911 = ~n994;
assign n625 = ~(n1236 ^ n1465);
assign n1176 = n1260 & n1725;
assign n870 = n1631 & n580;
assign n16 = ~(n322 ^ n1270);
assign n508 = n296 | n1634;
assign n720 = ~(n996 | n1284);
assign n836 = ~n1156;
assign n605 = n291 | n530;
assign n1671 = ~(n1385 ^ n722);
assign n761 = ~(n257 | n408);
assign n521 = ~n1451;
assign n1329 = n979 | n647;
assign n816 = ~(n688 | n1580);
assign n354 = ~(n374 | n1646);
assign n1638 = n627 | n559;
assign n1705 = n533 | n9;
assign n196 = n835 | n1566;
assign n724 = n425 | n333;
assign n1503 = ~n347;
assign n1426 = n882 & n1405;
assign n472 = ~(n1019 | n1240);
assign n1232 = ~(n653 ^ n695);
assign n325 = n1118 | n404;
assign n381 = n267 | n705;
assign n1510 = ~n321;
assign n1577 = n1161 & n1538;
assign n1391 = ~(n14 ^ n833);
assign n696 = ~(n899 | n1264);
assign n398 = ~(n1085 | n830);
assign n1650 = ~n738;
assign n1100 = n1039 | n135;
assign n404 = ~n1593;
assign n1262 = n1677 | n939;
assign n666 = n607 & n1004;
assign n1723 = ~n502;
assign n782 = n222;
assign n630 = ~n1295;
assign n347 = n1614 | n295;
assign n830 = n696 | n1743;
assign n1003 = ~n227;
assign n1724 = n1576 & n1458;
assign n462 = n594 | n1741;
assign n1284 = n98 | n1064;
assign n294 = ~(n1263 | n780);
assign n648 = ~(n311 ^ n820);
assign n938 = n1584 | n1264;
assign n336 = ~n631;
assign n57 = n116 | n1405;
assign n1200 = n666 | n207;
assign n1362 = n1020 & n583;
assign n1421 = n695;
assign n892 = ~n507;
assign n1049 = n1535 | n661;
assign n1564 = ~n1385;
assign n612 = n1369 | n530;
assign n1 = ~(n1245 | n1444);
assign n759 = n1722 | n614;
assign n27 = n947;
assign n1001 = ~n622;
assign n1116 = ~(n278 ^ n346);
assign n83 = n1259 | n521;
assign n1423 = ~(n1145 | n1318);
assign n840 = n736 & n697;
assign n912 = n187 | n1130;
assign n1211 = n1241 | n897;
assign n342 = ~n904;
assign n61 = ~(n1333 | n1395);
assign n1535 = ~n1747;
assign n1651 = ~(n1123 ^ n940);
assign n1185 = ~(n721 | n1301);
assign n238 = ~n413;
assign n715 = ~(n680 | n622);
assign n1127 = ~n600;
assign n339 = ~(n1303 ^ n408);
assign n1601 = ~n266;
assign n37 = n293 | n269;
assign n827 = n127 | n1158;
assign n1575 = n629 | n1620;
assign n1280 = n1020 & n1414;
assign n1431 = n248 & n1240;
assign n355 = ~(n721 | n374);
assign n343 = n1453 | n1499;
assign n1620 = ~(n1494 ^ n664);
assign n5 = n57 & n605;
assign n634 = ~(n1581 | n1606);
assign n31 = n721 | n1592;
assign n714 = n1036 | n995;
assign n1055 = n1412 ^ n74;
assign n296 = n1342 & n1392;
assign n7 = n14 | n448;
assign n108 = ~n722;
assign n891 = ~(n1642 ^ n920);
assign n226 = ~(n1149 | n868);
assign n1412 = n1732 & n635;
assign n1390 = ~n756;
assign n352 = n1463;
assign n1630 = ~n77;
assign n1192 = ~(n547 | n942);
assign n417 = n399;
assign n1732 = n890 | n257;
assign n1242 = ~n601;
assign n1319 = n125 & n1602;
assign n942 = ~(n1181 | n599);
assign n494 = n1607 | n122;
assign n328 = ~(n900 | n831);
assign n603 = n680 & n274;
assign n915 = ~n82;
assign n1032 = n1376 | n238;
assign n965 = n1755 | n1709;
assign n321 = ~(n266 ^ n612);
assign n130 = n1592;
assign n553 = n450 | n1010;
assign n1498 = ~(n311 ^ n945);
assign n1068 = n1722 | n614;
assign n1296 = ~n992;
assign n1615 = n545 & n283;
assign n1583 = n1129 | n843;
assign n1667 = ~n473;
assign n1581 = n494 | n91;
assign n1252 = ~n1569;
assign n1540 = ~(n98 ^ n837);
assign n562 = ~(n698 | n1108);
assign n55 = ~(n628 | n1469);
assign n1186 = n1047 | n872;
assign n716 = n231 & n795;
assign n1101 = n969 & n1206;
assign n457 = n827 | n1452;
assign n1063 = ~(n613 ^ n136);
assign n1356 = n1444 | n1001;
assign n1331 = n1222 & n1411;
assign n1238 = n1171 | n1457;
assign n405 = n1353 | n290;
assign n756 = n141 & n1688;
assign n1069 = n257 | n220;
assign n1683 = n1669 & n682;
assign n1093 = n257 | n293;
assign n1004 = ~n1314;
assign n642 = n1450 | n530;
assign n217 = n550 | n415;
assign n160 = n485 | n563;
assign n1136 = ~n413;
assign n1373 = ~(n753 ^ n767);
assign n403 = n1351 | n720;
assign n763 = ~(n179 ^ n1595);
assign n1077 = n298 | n1458;
assign n730 = n1455 | n1348;
assign n1065 = ~(n592 ^ n305);
assign n1419 = ~(n1385 ^ n1463);
assign n678 = ~n1595;
assign n491 = ~n413;
assign n1000 = ~n1581;
assign n954 = ~(n896 ^ n1169);
assign n833 = n1705 | n480;
assign n198 = ~n569;
assign n776 = ~n1388;
assign n1657 = n414 | n329;
assign n162 = ~n1428;
assign n1471 = n316 | n191;
assign n951 = n19 | n1098;
assign n475 = ~n1149;
assign n1554 = n1179 | n1128;
assign n193 = ~n54;
assign n1330 = ~(n1165 | n970);
assign n110 = n1567 | n683;
assign n948 = n1293 & n844;
assign n1744 = ~(n55 | n911);
assign n1547 = n420;
assign n897 = ~(n1733 | n634);
assign n1405 = ~n728;
assign n1726 = ~(n1206 | n1205);
assign n712 = ~(n1041 | n904);
assign n1491 = ~n964;
assign n1377 = n725 ^ n1566;
assign n498 = n293;
assign n1672 = ~(n785 ^ n318);
assign n1433 = n95 | n332;
assign n1157 = n712 & n235;
assign n1591 = ~(n1512 | n69);
assign n1605 = n1753 & n1222;
assign n194 = n867 | n1522;
assign n1552 = ~n510;
assign n224 = n699 | n1744;
assign n407 = n1358 & n178;
assign n1473 = n182 | n328;
assign n649 = ~(n551 ^ n1011);
assign n1139 = n101 | n384;
assign n141 = ~(n1319 | n259);
assign n421 = ~(n652 ^ n1467);
assign n826 = n282 & n302;
assign n1464 = n784 | n1544;
assign n1574 = ~(n134 | n88);
assign n1610 = ~(n431 ^ n411);
assign n591 = ~n1647;
assign n1546 = ~(n1416 ^ n115);
assign n1551 = ~n869;
assign n1013 = ~n71;
assign n456 = n1705 ^ n572;
assign n1038 = ~(n283 | n1336);
assign n1181 = n1179 | n716;
assign n1682 = ~(n1635 ^ n1656);
assign n1066 = ~n1059;
assign n566 = ~(n1520 & n1613);
assign n1012 = n973 | n17;
assign n1557 = n367 & n1229;
assign n919 = n1658 & n711;
assign n852 = n1654 | n1611;
assign n1436 = ~n1490;
assign n974 = n876 | n1045;
assign n972 = n1397 | n1070;
assign n722 = n151 | n484;
assign n1369 = ~n1205;
assign n131 = n1117 | n106;
assign n934 = n1540 | n348;
assign n1451 = n850 | n1555;
assign n275 = n1296;
assign n917 = ~(n846 ^ n48);
assign n1118 = n232 | n67;
assign n444 = ~n808;
assign n1203 = n368 | n1014;
assign n479 = n45 | n1352;
assign n60 = ~(n1682 ^ n941);
assign n218 = ~n1682;
assign n459 = n300 & n835;
assign n1206 = ~n413;
assign n1298 = ~n1276;
assign n1005 = ~(n467 | n363);
assign n1544 = ~n571;
assign n1666 = ~(n338 | n1653);
assign n439 = ~(n814 ^ n256);
assign n215 = ~(n1439 ^ n1525);
assign n1008 = n104 | n15;
assign n1652 = n239 | n1405;
assign n1452 = n1280 | n1362;
assign n225 = ~(n972 ^ n45);
assign n449 = ~(n1638 ^ n986);
assign n1195 = n1704 | n919;
assign n764 = n1674 | n1143;
assign n368 = ~(n1295 ^ n188);
assign n499 = ~n235;
assign n526 = n294 | n1094;
assign n1685 = ~(n876 ^ n903);
assign n1413 = n1676 & n1618;
assign n982 = n490 | n937;
assign n1690 = n975 | n139;
assign n532 = ~n1573;
assign n1686 = ~n1039;
assign n1492 = n1185 | n1480;
assign n334 = ~(n405 | n855);
assign n6 = ~(n1489 ^ n806);
assign n106 = n204 & n339;
assign n931 = ~(n1123 ^ n383);
assign n105 = n913 | n554;
assign n773 = n980;
assign n1174 = n1074 | n1555;
assign n628 = ~(n1608 | n1282);
assign n1702 = ~(n121 | n42);
assign n814 = ~(n1228 | n311);
assign n1241 = n986 & n737;
assign n1567 = n1578 | n286;
assign n397 = ~n664;
assign n679 = n949 & n375;
assign n111 = ~(n438 ^ n410);
assign n353 = n31 & n1031;
assign n1308 = n1111 | n1555;
assign n1312 = n1723 | n444;
assign n1679 = ~(n962 ^ n860);
assign n317 = n834 | n817;
assign n247 = ~(n1700 ^ n1325);
assign n640 = n1345;
assign n1376 = ~n953;
assign n855 = ~(n1358 | n673);
assign n1027 = ~(n1570 | n765);
assign n1223 = ~(n993 | n908);
assign n349 = n1624 | n861;
assign n309 = ~n1448;
assign n985 = ~(n1147 | n1096);
assign n868 = n1214 | n1700;
assign n1026 = ~n267;
assign n617 = n685 | n336;
assign n535 = ~(n174 ^ n674);
assign n853 = n1206 | n138;
assign n971 = ~n341;
assign n1631 = ~n823;
assign n1208 = n78 & n435;
assign n370 = ~(n339 ^ n334);
assign n59 = ~(n546 ^ n12);
assign n851 = ~(n513 ^ n16);
assign n541 = n162 | n238;
assign n889 = ~(n257 | n1345);
assign n203 = ~(n811 ^ n1672);
assign n158 = ~(n44 ^ n931);
assign n748 = n1684 | n511;
assign n95 = ~n406;
assign n395 = ~(n1171 | n1457);
assign n201 = ~(n888 ^ n1270);
assign n937 = ~(n1360 | n1230);
assign n18 = n729 & n900;
assign n575 = ~n490;
assign n842 = n1205;
assign n1628 = ~(n257 | n246);
assign n144 = n1751 | n6;
assign n998 = n197 | n18;
assign n994 = n1503 | n713;
assign n529 = ~n641;
assign n1721 = ~n539;
assign n1562 = ~(n1748 | n360);
assign n741 = ~n37;
assign n1549 = ~(n525 | n495);
assign n3 = ~(n1206 | n487);
assign n684 = ~n1092;
assign n234 = ~(n93 ^ n1471);
assign n789 = n757 | n944;
assign n1429 = ~n1583;
assign n685 = n692 & n1188;
assign n371 = n586 | n1715;
assign n996 = n731 | n14;
assign n280 = n1418 & n257;
assign n241 = ~n1610;
assign n881 = ~(n166 ^ n520);
assign n1006 = ~(n237 ^ n1395);
assign n361 = ~(n702 | n147);
assign n1081 = n865 & n621;
assign n615 = ~(n165 ^ n1028);
assign n65 = ~(n368 | n1014);
assign n988 = ~n1756;
assign n622 = ~(n1441 ^ n234);
assign n860 = ~(n1256 ^ n766);
assign n1024 = ~(n812 ^ n1662);
assign n594 = n1603 | n878;
assign n632 = n167 & n1730;
assign n848 = n1516 & n1222;
assign n1096 = n924 | n35;
assign n455 = ~(n648 ^ n881);
assign n1508 = n1735 & n1710;
assign n101 = n266 | n791;
assign n922 = ~(n843 ^ n856);
assign n283 = n473 & n1677;
assign n236 = ~(n1489 ^ n1751);
assign n737 = n1638 | n1110;
assign n1379 = n310 & n240;
assign n172 = n541 & n419;
assign n1699 = ~(n1173 ^ n1332);
assign n707 = n400 | n1522;
assign n880 = n63 & n1069;
assign n1728 = ~(n451 | n96);
assign n1288 = n912 | n128;
assign n1047 = n1218 | n429;
assign n1703 = n1076 | n1004;
assign n788 = ~n1282;
assign n520 = n289 & n1112;
assign n1137 = n1106 & n888;
assign n976 = ~n448;
assign n1039 = ~(n689 ^ n925);
assign n1233 = ~(n924 ^ n1494);
assign n214 = n690 & n1711;
assign n1122 = n542 & n639;
assign n1593 = n65 & n365;
assign n643 = n637 & n1357;
assign n1408 = ~(n83 | n1008);
assign n1363 = ~(n1045 | n1685);
assign n1752 = n118 | n208;
assign n358 = ~n1597;
assign n1742 = n1472 | n1633;
assign n1371 = n590 & n1643;
assign n932 = n131 | n464;
assign n480 = n1462 & n270;
assign n680 = n1151 & n1444;
assign n424 = ~n1071;
assign n176 = ~(n1683 | n281);
assign n114 = n1533 | n1431;
assign n1053 = n1176 | n1274;
assign n1559 = n1066 & n1311;
assign n1589 = n154 ^ n1740;
assign n1528 = n1252 | n1136;
assign n702 = n1197 | n678;
assign n15 = n1227 & n602;
assign n169 = ~(n1433 | n616);
assign n1707 = n895 ^ n551;
assign n862 = ~n36;
assign n84 = ~n1345;
assign n1249 = ~(n871 ^ n1258);
assign n150 = ~n689;
assign n705 = ~n732;
assign n1603 = ~(n1301 | n1675);
assign n1670 = ~(n93 ^ n604);
assign n1245 = n1196 | n1097;
assign n610 = ~(n1600 ^ n421);
assign n1378 = n240 & n1281;
assign n857 = n1535 | n492;
assign n1368 = n420;
assign n1021 = n733 | n804;
assign n434 = ~(n1151 | n673);
assign n1445 = ~(n78 ^ n1507);
assign n1469 = ~(n542 | n788);
assign n454 = ~n1217;
assign n692 = n1749 | n835;
assign n824 = n645 & n1555;
assign n400 = n240 & n1023;
assign n1641 = n848 | n221;
assign n571 = n1179 | n1510;
assign n964 = n83 & n1008;
assign n1398 = ~(n504 ^ n1265);
assign n941 = n330 | n854;
assign n1572 = n63 & n393;
assign n952 = ~(n539 ^ n1454);
assign n1584 = ~n1097;
assign n1684 = n800 | n1425;
assign n627 = ~n156;
assign n1606 = n1371 & n709;
assign n1754 = ~(n768 | n1490);
assign n1333 = ~n1669;
assign n1696 = ~n288;
assign n291 = ~n710;
assign n39 = n1279 & n533;
assign n706 = ~(n923 ^ n399);
assign n1277 = ~(n1038 ^ n1690);
assign n968 = ~n893;
assign n157 = ~(n1519 ^ n1300);
assign n1550 = n1535 | n1087;
assign n411 = ~(n1410 ^ n373);
assign n147 = n1171 | n1457;
assign n621 = n210 | n102;
assign n1633 = ~n381;
assign n1725 = n355 | n1016;
assign n118 = ~(n581 & n743);
assign n1677 = ~n746;
assign n1220 = ~(n331 ^ n556);
assign n1271 = n1131 | n1098;
assign n1478 = n1593 & n349;
assign n1264 = ~n1157;
assign n1213 = ~(n249 | n1583);
assign n547 = ~(n545 | n1423);
assign n669 = n1221 | n433;
assign n1014 = ~(n1512 ^ n1049);
assign n1311 = ~n1261;
assign n375 = n1146 | n459;
assign n1553 = n1609 & n1555;
assign n966 = ~(n721 | n1263);
assign n577 = n870 & n1582;
assign n1634 = n987 & n1475;
assign n1640 = n397 | n260;
assign n620 = n153 | n1381;
assign n320 = ~n387;
assign n76 = n1136 | n626;
assign n1733 = n97;
assign n1134 = n1712 | n1743;
assign n163 = n180 | n1168;
assign n1342 = ~n1592;
assign n500 = n705 | n351;
assign n596 = ~(n667 ^ n751);
assign n595 = n1301;
assign n1303 = n1719 | n681;
assign n1143 = ~n124;
assign n665 = ~n829;
assign n1209 = n1071;
assign n394 = ~(n458 ^ n213);
assign n887 = n1625 | n1458;
assign n1057 = n339 & n577;
assign n125 = ~n346;
assign n66 = n1440 & n463;
assign n1509 = n835 | n1278;
assign n654 = ~(n1092 ^ n986);
assign n638 = n420;
assign n278 = ~n1602;
assign n539 = ~(n580 ^ n823);
assign n552 = ~n1739;
assign n674 = ~(n1602 ^ n880);
assign n843 = n552 | n1294;
assign n438 = ~(n1399 ^ n1344);
assign n745 = n663 & n1136;
assign n799 = ~(n436 ^ n1488);
assign n1123 = n708 ^ n1468;
assign n1125 = ~n554;
assign n644 = n1052 | n797;
assign n145 = ~n1011;
assign n1439 = ~(n353 ^ n970);
assign n1691 = ~n1173;
assign n599 = ~(n231 | n754);
assign n650 = n1343 ^ n1260;
assign n1292 = n1616;
assign n544 = n673 | n440;
assign n116 = ~n1586;
assign n550 = n526 | n700;
assign n1224 = ~(n917 ^ n1556);
assign n1230 = ~n789;
assign n1073 = ~(n439 ^ n455);
assign n1530 = n1692 & n863;
assign n894 = ~(n811 ^ n114);
assign n1745 = ~(n1617 ^ n596);
assign n1374 = n900 | n391;
assign n977 = n920 | n1504;
assign n1668 = ~n1175;
assign n452 = n1412 | n687;
assign n1425 = n296 & n1672;
assign n1268 = ~n1443;
assign n838 = ~(n617 | n1313);
assign n335 = n66 | n1199;
assign n1548 = n567;
assign n441 = n1535 | n209;
assign n847 = ~n936;
assign n51 = ~(n721 | n947);
assign n206 = n1155 & n548;
assign n189 = n368 | n1014;
assign n435 = n571 | n1232;
assign n232 = ~(n1200 | n1664);
assign n161 = n457;
assign n568 = n222 | n108;
assign n1265 = ~(n1067 ^ n442);
assign n425 = n1222 & n560;
assign n1499 = ~(n924 ^ n1550);
assign n469 = ~(n1056 ^ n898);
assign n1291 = n1032 & n1310;
assign n412 = ~(n941 | n786);
assign n276 = n960 & n191;
assign n1025 = ~n1151;
assign n113 = n892 | n1458;
assign n856 = ~(n205 ^ n249);
assign n808 = ~n263;
assign n1256 = n1228 ^ n1533;
assign n1701 = ~(n136 | n1424);
assign n1646 = ~n1740;
assign n689 = ~(n1382 ^ n1446);
assign n46 = ~n1566;
assign n152 = ~(n960 ^ n1471);
assign n1558 = n803 | n695;
assign n372 = ~(n353 | n537);
assign n1730 = n796 | n1168;
assign n1259 = n344 & n197;
assign n546 = ~(n1366 ^ n1090);
assign n1441 = ~(n812 ^ n13);
assign n1713 = ~(n1135 | n1261);
assign n128 = n1745 | n1082;
assign n1674 = n1215 | n297;
assign n423 = n539 & n1035;
assign n694 = n467 | n363;
assign n1533 = n987 | n538;
assign n1751 = n1535 | n350;
assign n1746 = ~(n371 | n270);
assign n179 = n1267 | n1466;
assign n927 = ~(n257 | n920);
assign n1041 = n46 & n725;
assign n652 = ~(n1370 | n3);
assign n899 = ~n1196;
assign n580 = n536 | n1297;
assign n389 = ~(n133 | n1495);
assign n1059 = n1463 | n1564;
assign n1659 = ~(n1517 ^ n1316);
assign n115 = ~n1492;
assign n949 = n63 & n41;
assign n458 = n903 ^ n43;
assign n274 = ~(n1670 ^ n1024);
assign n987 = n1266 & n623;
assign n967 = ~(n1577 ^ n1751);
assign n1145 = ~(n668 | n795);
assign n258 = n58 & n240;
assign n1354 = n1020 & n110;
assign n313 = n134 & n20;
assign n601 = n475 | n665;
assign n845 = n29 & n1004;
assign n1449 = ~(n284 & n574);
assign n1519 = n1403 | n371;
assign n1442 = ~(n1535 | n1612);
assign n1494 = n245 | n1571;
assign n1749 = ~n52;
assign n1199 = ~(n1456 ^ n631);
assign n279 = n205 & n1183;
assign n1406 = ~n1618;
assign n207 = n1246 & n491;
assign n1366 = ~(n1689 ^ n818);
assign n924 = n76 & n963;
assign n482 = ~(n945 | n1326);
assign n1400 = ~n946;
assign n13 = ~(n739 ^ n80);
assign n10 = ~n88;
assign n1036 = ~(n432 | n1086);
assign n1108 = ~(n359 | n274);
assign n1204 = n1437 | n1243;
assign n188 = n966 | n1323;
assign n1594 = n255 | n319;
assign n73 = ~(n152 | n42);
assign n1146 = ~(n1405 | n1470);
assign n1180 = n1405 | n1476;
assign n1710 = ~(n1213 | n495);
assign n1098 = ~(n950 ^ n633);
assign n1120 = n1608 & n744;
assign n1663 = n172 | n951;
assign n202 = ~(n1026 | n613);
assign n1688 = ~n1183;
assign n209 = ~n32;
assign n171 = n1458 & n961;
assign n136 = ~n698;
assign n975 = ~n503;
assign n396 = n195 | n1160;
assign n34 = ~n1305;
assign n1472 = ~n620;
assign n1244 = ~(n186 | n512);
assign n1625 = ~n1154;
assign n257 = ~n728;
assign n1348 = n299 & n491;
assign n781 = ~n785;
assign n944 = ~(n1394 | n176);
assign n4 = n1136 | n1299;
assign n1722 = ~(n1676 ^ n1618);
assign n1034 = ~(n763 | n185);
assign n1313 = n19 | n1098;
assign n1560 = ~n1245;
assign n1675 = ~n1021;
assign n431 = ~(n202 ^ n771);
assign n1310 = n1365 | n1458;
assign n871 = n171 | n1601;
assign n633 = n447 | n445;
assign n338 = ~(n1135 | n388);
assign n1222 = ~n886;
assign n285 = ~(n123 ^ n277);
assign n1129 = n706 & n1468;
assign n1255 = n62 | n1206;
assign n910 = ~n841;
assign n260 = ~n1494;
assign n1275 = n1474 & n1168;
assign n1512 = n1497 & n1308;
assign n1364 = ~(n1573 ^ n1629);
assign n1088 = n1164 & n257;
assign n859 = ~(n1459 ^ n1277);
assign n332 = ~n965;
assign n1416 = n196 & n113;
assign n572 = ~n1257;
assign n647 = ~(n406 ^ n965);
assign n916 = ~(n1682 ^ n911);
assign n1660 = n734 & n240;
assign n1563 = ~n200;
assign n524 = ~n273;
assign n556 = n5 ^ n1676;
assign n1756 = n37 | n1623;
assign n1327 = ~(n357 | n103);
assign n166 = n1003 | n1019;
assign n1168 = ~n1314;
assign n732 = ~(n1043 ^ n153);
assign n362 = n914 | n1361;
assign n1461 = ~n143;
assign n265 = ~n105;
assign n1432 = n925 | n227;
assign n282 = n424 & n1332;
assign n204 = n1568 & n1641;
assign n810 = n809 | n939;
assign n1440 = n1206 | n1446;
assign n1573 = ~(n0 ^ n986);
assign n970 = ~n633;
assign n929 = n1182 ^ n179;
assign n822 = ~(n584 | n1524);
assign n1456 = ~n685;
assign n1276 = n958 & n643;
assign n1092 = n627 | n1563;
assign n1479 = n1135 & n265;
assign n192 = ~(n1422 | n697);
assign n981 = ~(n1329 | n764);
assign n1210 = n244 & n197;
assign n614 = ~(n49 ^ n5);
assign n1217 = n996 | n448;
assign n329 = n1720 & n1694;
assign n959 = n1219 | n444;
assign n1334 = n1380 & n901;
assign n955 = ~(n588 ^ n1501);
assign n586 = n670 & n1317;
assign n770 = n437 | n1247;
assign n1662 = ~(n741 ^ n1157);
assign n79 = ~(n799 ^ n1737);
assign n1234 = n608;
assign n1692 = ~n1565;
assign n473 = ~(n1332 ^ n1071);
assign n1739 = n399 | n70;
assign n1338 = ~(n1535 | n813);
assign n590 = ~(n629 | n1620);
assign n184 = n420;
assign n1420 = ~(n1232 ^ n1464);
assign n1712 = ~(n960 | n191);
assign n1300 = n7 & n1622;
assign n311 = ~(n777 ^ n1345);
assign n979 = ~(n1399 ^ n1412);
assign n631 = n1124 | n280;
assign n1444 = ~n359;
assign n1706 = ~n789;
assign n1202 = n1430 | n240;
assign n1290 = ~n311;
assign n664 = n63 & n4;
assign n30 = n362;
assign n78 = n1190 & n677;
assign n287 = ~n1446;
assign n337 = n626;
assign n733 = n1350 & n530;
assign n323 = n156 & n401;
assign n1447 = ~(n1405 | n1463);
assign n1372 = n803 | n430;
assign n667 = ~(n1642 ^ n750);
assign n1524 = n68 | n1736;
assign n1064 = n1257 | n802;
assign n990 = ~(n1694 ^ n412);
assign n563 = ~(n1248 | n347);
assign n1403 = ~n1383;
assign n1295 = n1692 & n1062;
assign n267 = n1401 | n1529;
assign n1382 = n1514 | n749;
assign n895 = n1315 & n1174;
assign n1149 = n620 | n1721;
assign n261 = ~(n1550 ^ n397);
assign n1183 = n249 & n1294;
assign n1495 = n857 | n629;
assign n248 = ~(n623 ^ n1616);
assign n185 = ~(n632 ^ n1182);
assign n806 = ~n815;
assign n393 = n602 | n477;
assign n382 = n1206 | n582;
assign n447 = ~(n803 | n318);
assign n1636 = ~(n1535 ^ n1338);
assign n64 = n1330 | n372;
assign n1317 = n1692 & n1162;
assign n233 = ~(n1192 ^ n816);
assign n691 = n532 & n1048;
assign n1163 = ~(n608 | n1691);
assign n33 = n927 | n619;
assign n365 = ~(n6 | n967);
assign n744 = ~n639;
assign n286 = n1526 | n53;
assign n410 = ~(n418 ^ n955);
assign n1409 = n549 | n343;
assign n1748 = ~(n999 | n322);
assign n865 = n1005 & n1363;
assign n1344 = n366 & n642;
assign n1052 = ~n43;
assign n1481 = n1706 & n1679;
assign n470 = ~(n1682 ^ n1665);
assign n1182 = n1255 & n1202;
assign n290 = ~(n1700 | n1242);
assign n1504 = ~n1642;
assign n132 = n895 | n1068;
assign n350 = ~(n257 | n609);
assign n178 = ~n405;
assign n109 = n206 | n1171;
assign n1336 = n662 | n1532;
assign n98 = ~n1462;
assign n699 = ~(n1122 | n81);
assign n668 = n317 | n805;
assign n1109 = ~(n1671 ^ n1589);
assign n693 = ~(n732 ^ n390);
assign n385 = ~(n864 ^ n540);
assign n1645 = n1446;
assign n829 = n1721 | n381;
assign n75 = ~n11;
assign n170 = n1033 | n822;
assign n503 = n1510 | n1232;
assign n1140 = n155 & n803;
assign n1360 = ~n643;
assign n1231 = n1470;
assign n63 = ~n1565;
assign n728 = ~n308;
assign n864 = ~n991;
assign n1695 = ~(n257 | n1626);
assign n1167 = ~(n1132 | n544);
assign n522 = n1402 | n649;
assign n1022 = n1347 | n1081;
assign n485 = ~(n1248 | n862);
assign n67 = n1717 | n369;
assign n872 = n691 & n901;
assign n514 = ~(n1226 | n1344);
assign n933 = ~(n572 | n519);
assign n1541 = ~(n721 | n21);
endmodule
