// Benchmark "top_810222779_843330999_776144567_776418743_1234615" written by ABC on Fri Jun 14 22:41:39 2024

module top_810222779_843330999_776144567_776418743_1234615 ( 
    n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82, n86,
    n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200, n219,
    n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273, n284,
    n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341, n344,
    n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420, n430,
    n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560, n561,
    n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609, n626,
    n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729, n734,
    n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831, n832,
    n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961, n969,
    n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061, n1071,
    n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164, n1172,
    n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246, n1250,
    n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305, n1345,
    n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411, n1415,
    n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470, n1474,
    n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536, n1566,
    n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627, n1644,
    n1647, n1656, n1750, n1753,
    n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181,
    n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362,
    n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501,
    n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669,
    n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918,
    n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063,
    n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285,
    n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368,
    n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588,
    n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752  );
  input  n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82,
    n86, n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200,
    n219, n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273,
    n284, n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341,
    n344, n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420,
    n430, n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560,
    n561, n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609,
    n626, n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729,
    n734, n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831,
    n832, n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961,
    n969, n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061,
    n1071, n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164,
    n1172, n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246,
    n1250, n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305,
    n1345, n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411,
    n1415, n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470,
    n1474, n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536,
    n1566, n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627,
    n1644, n1647, n1656, n1750, n1753;
  output n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181,
    n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362,
    n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501,
    n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669,
    n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918,
    n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063,
    n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285,
    n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368,
    n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588,
    n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752;
  wire new_n316, new_n317, new_n318_1, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337_1, new_n338, new_n339, new_n340, new_n341_1,
    new_n342, new_n343, new_n344_1, new_n345, new_n346_1, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352_1, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362_1, new_n363, new_n364_1, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370_1, new_n371, new_n372, new_n373,
    new_n374_1, new_n375, new_n376_1, new_n377, new_n378_1, new_n379,
    new_n380_1, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391_1, new_n392_1,
    new_n393, new_n394, new_n395, new_n396_1, new_n397, new_n398,
    new_n399_1, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408_1, new_n409_1, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416_1, new_n417_1,
    new_n418, new_n419, new_n420_1, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428_1, new_n429, new_n430_1,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n443, new_n444,
    new_n445, new_n446, new_n447, new_n448, new_n449, new_n450, new_n451,
    new_n452, new_n453_1, new_n454, new_n455, new_n456, new_n457_1,
    new_n458, new_n459, new_n460_1, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477_1,
    new_n478_1, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487_1, new_n488, new_n489_1, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497_1,
    new_n498_1, new_n499, new_n500, new_n501_1, new_n502_1, new_n503,
    new_n504, new_n505, new_n506_1, new_n507_1, new_n508, new_n509_1,
    new_n510_1, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516_1, new_n517_1, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534_1, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545_1, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553_1, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559_1, new_n560_1, new_n561_1, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567_1, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574_1, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581_1, new_n582_1,
    new_n583, new_n584, new_n585_1, new_n586, new_n587, new_n588,
    new_n589_1, new_n590, new_n591, new_n592, new_n593_1, new_n594,
    new_n595_1, new_n596, new_n597_1, new_n598_1, new_n599, new_n600_1,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607_1,
    new_n608_1, new_n609_1, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625_1, new_n626_1,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638_1, new_n639,
    new_n640_1, new_n641_1, new_n642, new_n643, new_n644, new_n645_1,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n660, new_n661, new_n663_1,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669_1, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676_1,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690_1,
    new_n691, new_n692, new_n693_1, new_n694, new_n695_1, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701_1, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710_1,
    new_n711, new_n712, new_n713, new_n714_1, new_n715, new_n716, new_n717,
    new_n718, new_n719_1, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726_1, new_n727_1, new_n728, new_n729_1, new_n730,
    new_n731, new_n732, new_n733, new_n734_1, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742_1, new_n743_1,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755_1, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769_1, new_n770, new_n771,
    new_n772, new_n773_1, new_n774, new_n775_1, new_n776, new_n777,
    new_n778_1, new_n779_1, new_n780, new_n781, new_n782_1, new_n783,
    new_n784, new_n785, new_n786, new_n787_1, new_n788, new_n789,
    new_n790_1, new_n791, new_n792, new_n793, new_n794_1, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821_1, new_n822,
    new_n823_1, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831_1, new_n832_1, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839_1, new_n840, new_n841,
    new_n842_1, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849_1, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879_1, new_n880, new_n881, new_n882_1,
    new_n883, new_n884, new_n885_1, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894_1, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905_1, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916_1, new_n917,
    new_n918_1, new_n919, new_n920_1, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936_1, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947_1, new_n948, new_n949, new_n950, new_n951,
    new_n952_1, new_n953_1, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961_1, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969_1, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980_1, new_n981, new_n982, new_n983, new_n984_1,
    new_n985, new_n986_1, new_n987, new_n988, new_n989, new_n990_1,
    new_n991, new_n992_1, new_n993, new_n994, new_n995, new_n996,
    new_n997_1, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006_1, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017_1, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023_1, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040_1, new_n1041, new_n1042_1, new_n1043, new_n1044_1, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050_1, new_n1051_1,
    new_n1052, new_n1053, new_n1054_1, new_n1055, new_n1056, new_n1057,
    new_n1058_1, new_n1059, new_n1060_1, new_n1061_1, new_n1062,
    new_n1063_1, new_n1064, new_n1065_1, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071_1, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095_1,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103_1, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114_1,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121_1, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152_1, new_n1153, new_n1154_1, new_n1155, new_n1156_1,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164_1, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172_1, new_n1173, new_n1174, new_n1175_1,
    new_n1176, new_n1177_1, new_n1178, new_n1179, new_n1182, new_n1184,
    new_n1185, new_n1186_1, new_n1187_1, new_n1189, new_n1191_1, new_n1192,
    new_n1193_1, new_n1194, new_n1195_1, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205_1, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211_1, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225_1, new_n1226, new_n1227_1, new_n1228,
    new_n1229, new_n1230, new_n1231_1, new_n1232, new_n1233, new_n1234_1,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239_1, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246_1,
    new_n1247, new_n1248, new_n1249, new_n1250_1, new_n1251, new_n1252,
    new_n1253_1, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263_1, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278_1, new_n1279, new_n1280, new_n1281_1, new_n1282,
    new_n1283_1, new_n1284, new_n1285_1, new_n1286_1, new_n1287, new_n1290,
    new_n1291, new_n1292_1, new_n1293, new_n1294, new_n1295, new_n1296_1,
    new_n1297, new_n1298, new_n1299_1, new_n1300, new_n1301_1, new_n1303,
    new_n1305_1, new_n1306_1, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1318,
    new_n1319, new_n1320_1, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337_1, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345_1, new_n1346_1, new_n1347, new_n1348, new_n1349, new_n1350_1,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359_1, new_n1360, new_n1361_1, new_n1362,
    new_n1363, new_n1364, new_n1366, new_n1367, new_n1368_1, new_n1373,
    new_n1374, new_n1375_1, new_n1376, new_n1377, new_n1379, new_n1380,
    new_n1382, new_n1384, new_n1385, new_n1386_1, new_n1387_1, new_n1388,
    new_n1389_1, new_n1390, new_n1391_1, new_n1392, new_n1393_1, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401_1, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411_1, new_n1412,
    new_n1413, new_n1414, new_n1415_1, new_n1416, new_n1417, new_n1418_1,
    new_n1419, new_n1420_1, new_n1421_1, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427_1, new_n1428_1, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435_1, new_n1436,
    new_n1437, new_n1438_1, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443_1, new_n1444, new_n1445, new_n1446_1, new_n1447, new_n1448_1,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463_1, new_n1464, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1470_1, new_n1471, new_n1472, new_n1473,
    new_n1474_1, new_n1475, new_n1476_1, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500_1, new_n1501, new_n1502_1, new_n1503,
    new_n1504, new_n1505, new_n1506_1, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516_1, new_n1517, new_n1518, new_n1519, new_n1520_1, new_n1522,
    new_n1523_1, new_n1524, new_n1525, new_n1526, new_n1527_1, new_n1528,
    new_n1529, new_n1530, new_n1531, new_n1532, new_n1533, new_n1534_1,
    new_n1535, new_n1536_1, new_n1537, new_n1538, new_n1539, new_n1540,
    new_n1541, new_n1542, new_n1543, new_n1544, new_n1545, new_n1546,
    new_n1547_1, new_n1548_1, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1554, new_n1555, new_n1556, new_n1557, new_n1558,
    new_n1559, new_n1560, new_n1561, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1566_1, new_n1567, new_n1568, new_n1569_1, new_n1570,
    new_n1571, new_n1572, new_n1573, new_n1574, new_n1575, new_n1576_1,
    new_n1577, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1584, new_n1586_1, new_n1587, new_n1588_1, new_n1589,
    new_n1590, new_n1591, new_n1592_1, new_n1593, new_n1594_1, new_n1595,
    new_n1598, new_n1599, new_n1600, new_n1603, new_n1604, new_n1606,
    new_n1607, new_n1608, new_n1609_1, new_n1610, new_n1612, new_n1613_1,
    new_n1615, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626_1, new_n1627_1, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632_1, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639_1, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644_1, new_n1645_1, new_n1646,
    new_n1647_1, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656_1, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1671, new_n1675,
    new_n1676, new_n1677, new_n1681, new_n1683, new_n1684;
  not_3  g0000(.A(n1263), .Y(new_n316));
  nand_4 g0001(.A(n984), .B(n11), .Y(new_n317));
  not_3  g0002(.A(new_n317), .Y(new_n318_1));
  not_3  g0003(.A(n1239), .Y(new_n319));
  nor_4  g0004(.A(new_n319), .B(n220), .Y(new_n320));
  nor_4  g0005(.A(new_n320), .B(new_n318_1), .Y(new_n321));
  nand_4 g0006(.A(new_n321), .B(new_n316), .Y(new_n322));
  not_3  g0007(.A(new_n321), .Y(new_n323));
  nand_4 g0008(.A(new_n323), .B(n1263), .Y(new_n324));
  nand_4 g0009(.A(new_n324), .B(new_n322), .Y(new_n325));
  nor_4  g0010(.A(new_n319), .B(n391), .Y(new_n326));
  nor_4  g0011(.A(new_n326), .B(new_n318_1), .Y(new_n327));
  not_3  g0012(.A(new_n327), .Y(new_n328));
  nor_4  g0013(.A(new_n328), .B(n346), .Y(new_n329));
  not_3  g0014(.A(n346), .Y(new_n330));
  nor_4  g0015(.A(new_n327), .B(new_n330), .Y(new_n331));
  nor_4  g0016(.A(new_n319), .B(n905), .Y(new_n332));
  nor_4  g0017(.A(new_n332), .B(new_n318_1), .Y(new_n333));
  not_3  g0018(.A(new_n333), .Y(new_n334));
  nor_4  g0019(.A(new_n334), .B(n399), .Y(new_n335));
  not_3  g0020(.A(n399), .Y(new_n336));
  nor_4  g0021(.A(new_n333), .B(new_n336), .Y(new_n337_1));
  nor_4  g0022(.A(n1278), .B(new_n319), .Y(new_n338));
  nor_4  g0023(.A(new_n338), .B(new_n318_1), .Y(new_n339));
  not_3  g0024(.A(new_n339), .Y(new_n340));
  nor_4  g0025(.A(new_n340), .B(n980), .Y(new_n341_1));
  not_3  g0026(.A(new_n341_1), .Y(new_n342));
  nor_4  g0027(.A(new_n342), .B(new_n337_1), .Y(new_n343));
  nor_4  g0028(.A(new_n343), .B(new_n335), .Y(new_n344_1));
  nor_4  g0029(.A(new_n344_1), .B(new_n331), .Y(new_n345));
  nor_4  g0030(.A(new_n345), .B(new_n329), .Y(new_n346_1));
  not_3  g0031(.A(new_n346_1), .Y(new_n347));
  not_3  g0032(.A(n318), .Y(new_n348));
  nor_4  g0033(.A(n1435), .B(new_n319), .Y(new_n349));
  nor_4  g0034(.A(new_n349), .B(new_n318_1), .Y(new_n350));
  or_4   g0035(.A(new_n350), .B(new_n348), .Y(new_n351));
  nand_4 g0036(.A(new_n350), .B(new_n348), .Y(new_n352_1));
  nand_4 g0037(.A(n1415), .B(n1239), .Y(new_n353));
  not_3  g0038(.A(new_n353), .Y(new_n354));
  not_3  g0039(.A(n1246), .Y(new_n355));
  nor_4  g0040(.A(new_n355), .B(n1239), .Y(new_n356));
  nor_4  g0041(.A(new_n356), .B(new_n354), .Y(new_n357));
  nor_4  g0042(.A(new_n357), .B(n1345), .Y(new_n358));
  not_3  g0043(.A(n1345), .Y(new_n359));
  not_3  g0044(.A(new_n357), .Y(new_n360));
  nor_4  g0045(.A(new_n360), .B(new_n359), .Y(new_n361));
  nor_4  g0046(.A(new_n361), .B(new_n358), .Y(new_n362_1));
  not_3  g0047(.A(new_n362_1), .Y(new_n363));
  nand_4 g0048(.A(n1239), .B(n58), .Y(new_n364_1));
  not_3  g0049(.A(new_n364_1), .Y(new_n365));
  not_3  g0050(.A(n1443), .Y(new_n366));
  nor_4  g0051(.A(new_n366), .B(n1239), .Y(new_n367));
  nor_4  g0052(.A(new_n367), .B(new_n365), .Y(new_n368));
  xor_3  g0053(.A(new_n368), .B(n1616), .Y(new_n369));
  not_3  g0054(.A(new_n369), .Y(new_n370_1));
  not_3  g0055(.A(n1446), .Y(new_n371));
  nand_4 g0056(.A(n1239), .B(n598), .Y(new_n372));
  not_3  g0057(.A(new_n372), .Y(new_n373));
  not_3  g0058(.A(n1647), .Y(new_n374_1));
  nor_4  g0059(.A(new_n374_1), .B(n1239), .Y(new_n375));
  nor_4  g0060(.A(new_n375), .B(new_n373), .Y(new_n376_1));
  not_3  g0061(.A(new_n376_1), .Y(new_n377));
  nor_4  g0062(.A(new_n377), .B(new_n371), .Y(new_n378_1));
  nor_4  g0063(.A(new_n376_1), .B(n1446), .Y(new_n379));
  nor_4  g0064(.A(new_n379), .B(new_n378_1), .Y(new_n380_1));
  not_3  g0065(.A(new_n380_1), .Y(new_n381));
  nor_4  g0066(.A(new_n381), .B(new_n370_1), .Y(new_n382));
  not_3  g0067(.A(new_n382), .Y(new_n383));
  nor_4  g0068(.A(new_n383), .B(new_n363), .Y(new_n384));
  not_3  g0069(.A(new_n384), .Y(new_n385));
  nand_4 g0070(.A(n1474), .B(n1239), .Y(new_n386));
  not_3  g0071(.A(new_n386), .Y(new_n387));
  not_3  g0072(.A(n1506), .Y(new_n388));
  nor_4  g0073(.A(new_n388), .B(n1239), .Y(new_n389));
  nor_4  g0074(.A(new_n389), .B(new_n387), .Y(new_n390));
  and_4  g0075(.A(new_n390), .B(n1592), .Y(new_n391_1));
  nor_4  g0076(.A(new_n390), .B(n1592), .Y(new_n392_1));
  nor_4  g0077(.A(new_n392_1), .B(new_n391_1), .Y(new_n393));
  not_3  g0078(.A(new_n393), .Y(new_n394));
  nor_4  g0079(.A(new_n394), .B(new_n385), .Y(new_n395));
  not_3  g0080(.A(new_n395), .Y(new_n396_1));
  nand_4 g0081(.A(n1350), .B(n1239), .Y(new_n397));
  not_3  g0082(.A(new_n397), .Y(new_n398));
  not_3  g0083(.A(n262), .Y(new_n399_1));
  nor_4  g0084(.A(n1239), .B(new_n399_1), .Y(new_n400));
  nor_4  g0085(.A(new_n400), .B(new_n398), .Y(new_n401));
  nor_4  g0086(.A(new_n401), .B(n1301), .Y(new_n402));
  not_3  g0087(.A(n1301), .Y(new_n403));
  not_3  g0088(.A(new_n401), .Y(new_n404));
  nor_4  g0089(.A(new_n404), .B(new_n403), .Y(new_n405));
  nand_4 g0090(.A(n1239), .B(n676), .Y(new_n406));
  not_3  g0091(.A(new_n406), .Y(new_n407));
  not_3  g0092(.A(n1154), .Y(new_n408_1));
  nor_4  g0093(.A(n1239), .B(new_n408_1), .Y(new_n409_1));
  nor_4  g0094(.A(new_n409_1), .B(new_n407), .Y(new_n410));
  nor_4  g0095(.A(new_n410), .B(n1566), .Y(new_n411));
  not_3  g0096(.A(n1566), .Y(new_n412));
  not_3  g0097(.A(new_n410), .Y(new_n413));
  nor_4  g0098(.A(new_n413), .B(new_n412), .Y(new_n414));
  nand_4 g0099(.A(n1289), .B(n1239), .Y(new_n415));
  not_3  g0100(.A(new_n415), .Y(new_n416_1));
  not_3  g0101(.A(n1193), .Y(new_n417_1));
  nor_4  g0102(.A(n1239), .B(new_n417_1), .Y(new_n418));
  nor_4  g0103(.A(new_n418), .B(new_n416_1), .Y(new_n419));
  and_4  g0104(.A(new_n419), .B(n920), .Y(new_n420_1));
  nand_4 g0105(.A(n1239), .B(n244), .Y(new_n421));
  not_3  g0106(.A(new_n421), .Y(new_n422));
  not_3  g0107(.A(n641), .Y(new_n423));
  nor_4  g0108(.A(n1239), .B(new_n423), .Y(new_n424));
  nor_4  g0109(.A(new_n424), .B(new_n422), .Y(new_n425));
  nor_4  g0110(.A(new_n425), .B(n293), .Y(new_n426));
  nor_4  g0111(.A(new_n419), .B(n920), .Y(new_n427));
  nor_4  g0112(.A(new_n427), .B(new_n426), .Y(new_n428_1));
  nor_4  g0113(.A(new_n428_1), .B(new_n420_1), .Y(new_n429));
  not_3  g0114(.A(new_n429), .Y(new_n430_1));
  nor_4  g0115(.A(new_n430_1), .B(new_n414), .Y(new_n431));
  nor_4  g0116(.A(new_n431), .B(new_n411), .Y(new_n432));
  nor_4  g0117(.A(new_n432), .B(new_n405), .Y(new_n433));
  nor_4  g0118(.A(new_n433), .B(new_n402), .Y(new_n434));
  not_3  g0119(.A(new_n434), .Y(new_n435));
  not_3  g0120(.A(n293), .Y(new_n436));
  not_3  g0121(.A(new_n425), .Y(new_n437));
  nor_4  g0122(.A(new_n437), .B(new_n436), .Y(new_n438));
  nor_4  g0123(.A(new_n438), .B(new_n426), .Y(new_n439));
  nand_4 g0124(.A(n1239), .B(n251), .Y(new_n440));
  not_3  g0125(.A(new_n440), .Y(new_n441));
  not_3  g0126(.A(n1172), .Y(new_n442));
  nor_4  g0127(.A(n1239), .B(new_n442), .Y(new_n443));
  nor_4  g0128(.A(new_n443), .B(new_n441), .Y(new_n444));
  and_4  g0129(.A(new_n444), .B(n408), .Y(new_n445));
  nor_4  g0130(.A(new_n444), .B(n408), .Y(new_n446));
  not_3  g0131(.A(n1476), .Y(new_n447));
  nand_4 g0132(.A(n1516), .B(n1239), .Y(new_n448));
  not_3  g0133(.A(new_n448), .Y(new_n449));
  not_3  g0134(.A(n710), .Y(new_n450));
  nor_4  g0135(.A(n1239), .B(new_n450), .Y(new_n451));
  nor_4  g0136(.A(new_n451), .B(new_n449), .Y(new_n452));
  not_3  g0137(.A(new_n452), .Y(new_n453_1));
  nor_4  g0138(.A(new_n453_1), .B(new_n447), .Y(new_n454));
  nand_4 g0139(.A(n1239), .B(n82), .Y(new_n455));
  not_3  g0140(.A(new_n455), .Y(new_n456));
  not_3  g0141(.A(n1061), .Y(new_n457_1));
  nor_4  g0142(.A(n1239), .B(new_n457_1), .Y(new_n458));
  nor_4  g0143(.A(new_n458), .B(new_n456), .Y(new_n459));
  nor_4  g0144(.A(new_n459), .B(n1401), .Y(new_n460_1));
  not_3  g0145(.A(n1401), .Y(new_n461));
  not_3  g0146(.A(new_n459), .Y(new_n462));
  nor_4  g0147(.A(new_n462), .B(new_n461), .Y(new_n463));
  nor_4  g0148(.A(new_n463), .B(new_n460_1), .Y(new_n464));
  not_3  g0149(.A(new_n464), .Y(new_n465));
  nand_4 g0150(.A(n1239), .B(n790), .Y(new_n466));
  not_3  g0151(.A(new_n466), .Y(new_n467));
  not_3  g0152(.A(n1521), .Y(new_n468));
  nor_4  g0153(.A(new_n468), .B(n1239), .Y(new_n469));
  nor_4  g0154(.A(new_n469), .B(new_n467), .Y(new_n470));
  and_4  g0155(.A(new_n470), .B(n823), .Y(new_n471));
  nor_4  g0156(.A(new_n470), .B(n823), .Y(new_n472));
  nor_4  g0157(.A(new_n472), .B(new_n471), .Y(new_n473));
  not_3  g0158(.A(new_n473), .Y(new_n474));
  nand_4 g0159(.A(n1576), .B(n1239), .Y(new_n475));
  not_3  g0160(.A(new_n475), .Y(new_n476));
  not_3  g0161(.A(n1283), .Y(new_n477_1));
  nor_4  g0162(.A(new_n477_1), .B(n1239), .Y(new_n478_1));
  nor_4  g0163(.A(new_n478_1), .B(new_n476), .Y(new_n479));
  and_4  g0164(.A(new_n479), .B(n153), .Y(new_n480));
  nor_4  g0165(.A(new_n479), .B(n153), .Y(new_n481));
  nor_4  g0166(.A(new_n481), .B(new_n480), .Y(new_n482));
  not_3  g0167(.A(new_n482), .Y(new_n483));
  nor_4  g0168(.A(new_n483), .B(new_n474), .Y(new_n484));
  not_3  g0169(.A(new_n484), .Y(new_n485));
  nor_4  g0170(.A(new_n485), .B(new_n465), .Y(new_n486));
  not_3  g0171(.A(new_n486), .Y(new_n487_1));
  nor_4  g0172(.A(new_n487_1), .B(new_n454), .Y(new_n488));
  not_3  g0173(.A(n374), .Y(new_n489_1));
  nand_4 g0174(.A(n1239), .B(n645), .Y(new_n490));
  not_3  g0175(.A(new_n490), .Y(new_n491));
  not_3  g0176(.A(n87), .Y(new_n492));
  nor_4  g0177(.A(n1239), .B(new_n492), .Y(new_n493));
  nor_4  g0178(.A(new_n493), .B(new_n491), .Y(new_n494));
  not_3  g0179(.A(new_n494), .Y(new_n495));
  nor_4  g0180(.A(new_n495), .B(new_n489_1), .Y(new_n496));
  nand_4 g0181(.A(new_n495), .B(new_n489_1), .Y(new_n497_1));
  not_3  g0182(.A(n567), .Y(new_n498_1));
  nand_4 g0183(.A(n1239), .B(n268), .Y(new_n499));
  not_3  g0184(.A(new_n499), .Y(new_n500));
  not_3  g0185(.A(n600), .Y(new_n501_1));
  nor_4  g0186(.A(n1239), .B(new_n501_1), .Y(new_n502_1));
  nor_4  g0187(.A(new_n502_1), .B(new_n500), .Y(new_n503));
  not_3  g0188(.A(new_n503), .Y(new_n504));
  nor_4  g0189(.A(new_n504), .B(new_n498_1), .Y(new_n505));
  not_3  g0190(.A(new_n505), .Y(new_n506_1));
  nor_4  g0191(.A(new_n503), .B(n567), .Y(new_n507_1));
  not_3  g0192(.A(new_n507_1), .Y(new_n508));
  nand_4 g0193(.A(n1393), .B(n1239), .Y(new_n509_1));
  not_3  g0194(.A(new_n509_1), .Y(new_n510_1));
  not_3  g0195(.A(n254), .Y(new_n511));
  nor_4  g0196(.A(n1239), .B(new_n511), .Y(new_n512));
  nor_4  g0197(.A(new_n512), .B(new_n510_1), .Y(new_n513));
  nor_4  g0198(.A(new_n513), .B(n1463), .Y(new_n514));
  not_3  g0199(.A(n1463), .Y(new_n515));
  not_3  g0200(.A(new_n513), .Y(new_n516_1));
  nor_4  g0201(.A(new_n516_1), .B(new_n515), .Y(new_n517_1));
  nor_4  g0202(.A(new_n517_1), .B(new_n514), .Y(new_n518));
  nand_4 g0203(.A(n1239), .B(n312), .Y(new_n519));
  not_3  g0204(.A(new_n519), .Y(new_n520));
  not_3  g0205(.A(n307), .Y(new_n521));
  nor_4  g0206(.A(n1239), .B(new_n521), .Y(new_n522));
  nor_4  g0207(.A(new_n522), .B(new_n520), .Y(new_n523));
  nor_4  g0208(.A(new_n523), .B(n222), .Y(new_n524));
  not_3  g0209(.A(n222), .Y(new_n525));
  not_3  g0210(.A(new_n523), .Y(new_n526));
  nor_4  g0211(.A(new_n526), .B(new_n525), .Y(new_n527));
  nor_4  g0212(.A(new_n527), .B(new_n524), .Y(new_n528));
  nand_4 g0213(.A(new_n528), .B(new_n518), .Y(new_n529));
  not_3  g0214(.A(n608), .Y(new_n530));
  nand_4 g0215(.A(n1609), .B(n1239), .Y(new_n531));
  not_3  g0216(.A(new_n531), .Y(new_n532));
  not_3  g0217(.A(n54), .Y(new_n533));
  nor_4  g0218(.A(n1239), .B(new_n533), .Y(new_n534_1));
  nor_4  g0219(.A(new_n534_1), .B(new_n532), .Y(new_n535));
  not_3  g0220(.A(new_n535), .Y(new_n536));
  nor_4  g0221(.A(new_n536), .B(new_n530), .Y(new_n537));
  not_3  g0222(.A(new_n537), .Y(new_n538));
  nor_4  g0223(.A(new_n535), .B(n608), .Y(new_n539));
  not_3  g0224(.A(new_n539), .Y(new_n540));
  nand_4 g0225(.A(n1239), .B(n310), .Y(new_n541));
  not_3  g0226(.A(new_n541), .Y(new_n542));
  not_3  g0227(.A(n1175), .Y(new_n543));
  nor_4  g0228(.A(n1239), .B(new_n543), .Y(new_n544));
  nor_4  g0229(.A(new_n544), .B(new_n542), .Y(new_n545_1));
  nor_4  g0230(.A(new_n545_1), .B(n1071), .Y(new_n546));
  not_3  g0231(.A(new_n546), .Y(new_n547));
  not_3  g0232(.A(n1071), .Y(new_n548));
  not_3  g0233(.A(new_n545_1), .Y(new_n549));
  nor_4  g0234(.A(new_n549), .B(new_n548), .Y(new_n550));
  not_3  g0235(.A(new_n550), .Y(new_n551));
  nand_4 g0236(.A(n1239), .B(n219), .Y(new_n552));
  not_3  g0237(.A(new_n552), .Y(new_n553_1));
  not_3  g0238(.A(n409), .Y(new_n554));
  nor_4  g0239(.A(n1239), .B(new_n554), .Y(new_n555));
  nor_4  g0240(.A(new_n555), .B(new_n553_1), .Y(new_n556));
  nor_4  g0241(.A(new_n556), .B(n45), .Y(new_n557));
  not_3  g0242(.A(new_n557), .Y(new_n558));
  nand_4 g0243(.A(new_n556), .B(n45), .Y(new_n559_1));
  not_3  g0244(.A(n695), .Y(new_n560_1));
  nand_4 g0245(.A(n1569), .B(n1239), .Y(new_n561_1));
  not_3  g0246(.A(n1250), .Y(new_n562));
  nor_4  g0247(.A(new_n562), .B(n1239), .Y(new_n563));
  not_3  g0248(.A(new_n563), .Y(new_n564));
  nand_4 g0249(.A(new_n564), .B(new_n561_1), .Y(new_n565));
  nand_4 g0250(.A(new_n565), .B(new_n560_1), .Y(new_n566));
  not_3  g0251(.A(new_n561_1), .Y(new_n567_1));
  nor_4  g0252(.A(new_n563), .B(new_n567_1), .Y(new_n568));
  nand_4 g0253(.A(new_n568), .B(n695), .Y(new_n569));
  nand_4 g0254(.A(new_n319), .B(n510), .Y(new_n570));
  nor_4  g0255(.A(new_n570), .B(n1205), .Y(new_n571));
  nand_4 g0256(.A(new_n571), .B(new_n569), .Y(new_n572));
  nand_4 g0257(.A(new_n572), .B(new_n566), .Y(new_n573));
  nand_4 g0258(.A(new_n573), .B(new_n559_1), .Y(new_n574_1));
  nand_4 g0259(.A(new_n574_1), .B(new_n558), .Y(new_n575));
  nand_4 g0260(.A(new_n575), .B(new_n551), .Y(new_n576));
  nand_4 g0261(.A(new_n576), .B(new_n547), .Y(new_n577));
  not_3  g0262(.A(new_n559_1), .Y(new_n578));
  nor_4  g0263(.A(new_n578), .B(new_n557), .Y(new_n579));
  not_3  g0264(.A(new_n566), .Y(new_n580));
  not_3  g0265(.A(new_n569), .Y(new_n581_1));
  nor_4  g0266(.A(new_n581_1), .B(new_n580), .Y(new_n582_1));
  nand_4 g0267(.A(new_n582_1), .B(new_n579), .Y(new_n583));
  not_3  g0268(.A(n545), .Y(new_n584));
  not_3  g0269(.A(new_n571), .Y(new_n585_1));
  nor_4  g0270(.A(n1239), .B(n510), .Y(new_n586));
  nand_4 g0271(.A(new_n586), .B(n1205), .Y(new_n587));
  nand_4 g0272(.A(new_n587), .B(new_n585_1), .Y(new_n588));
  nor_4  g0273(.A(new_n588), .B(new_n584), .Y(new_n589_1));
  nor_4  g0274(.A(new_n550), .B(new_n546), .Y(new_n590));
  nand_4 g0275(.A(new_n590), .B(new_n589_1), .Y(new_n591));
  nor_4  g0276(.A(new_n591), .B(new_n583), .Y(new_n592));
  nor_4  g0277(.A(new_n592), .B(new_n577), .Y(new_n593_1));
  nand_4 g0278(.A(new_n593_1), .B(new_n540), .Y(new_n594));
  nand_4 g0279(.A(new_n594), .B(new_n538), .Y(new_n595_1));
  nor_4  g0280(.A(new_n595_1), .B(new_n529), .Y(new_n596));
  not_3  g0281(.A(new_n524), .Y(new_n597_1));
  nor_4  g0282(.A(new_n597_1), .B(new_n517_1), .Y(new_n598_1));
  nor_4  g0283(.A(new_n598_1), .B(new_n514), .Y(new_n599));
  not_3  g0284(.A(new_n599), .Y(new_n600_1));
  nor_4  g0285(.A(new_n600_1), .B(new_n596), .Y(new_n601));
  nand_4 g0286(.A(new_n601), .B(new_n508), .Y(new_n602));
  nand_4 g0287(.A(new_n602), .B(new_n506_1), .Y(new_n603));
  nand_4 g0288(.A(new_n603), .B(new_n497_1), .Y(new_n604));
  not_3  g0289(.A(new_n604), .Y(new_n605));
  nor_4  g0290(.A(new_n605), .B(new_n496), .Y(new_n606));
  nand_4 g0291(.A(new_n606), .B(new_n488), .Y(new_n607_1));
  nor_4  g0292(.A(new_n452), .B(n1476), .Y(new_n608_1));
  not_3  g0293(.A(new_n460_1), .Y(new_n609_1));
  nor_4  g0294(.A(new_n480), .B(new_n609_1), .Y(new_n610));
  nor_4  g0295(.A(new_n481), .B(new_n472), .Y(new_n611));
  not_3  g0296(.A(new_n611), .Y(new_n612));
  nor_4  g0297(.A(new_n612), .B(new_n610), .Y(new_n613));
  nor_4  g0298(.A(new_n613), .B(new_n471), .Y(new_n614));
  nor_4  g0299(.A(new_n614), .B(new_n608_1), .Y(new_n615));
  nor_4  g0300(.A(new_n615), .B(new_n454), .Y(new_n616));
  not_3  g0301(.A(new_n616), .Y(new_n617));
  nand_4 g0302(.A(new_n617), .B(new_n607_1), .Y(new_n618));
  nor_4  g0303(.A(new_n618), .B(new_n446), .Y(new_n619));
  nor_4  g0304(.A(new_n619), .B(new_n445), .Y(new_n620));
  nand_4 g0305(.A(new_n620), .B(new_n439), .Y(new_n621));
  nor_4  g0306(.A(new_n427), .B(new_n420_1), .Y(new_n622));
  not_3  g0307(.A(new_n622), .Y(new_n623));
  nor_4  g0308(.A(new_n405), .B(new_n402), .Y(new_n624));
  nor_4  g0309(.A(new_n414), .B(new_n411), .Y(new_n625_1));
  and_4  g0310(.A(new_n625_1), .B(new_n624), .Y(new_n626_1));
  not_3  g0311(.A(new_n626_1), .Y(new_n627));
  nor_4  g0312(.A(new_n627), .B(new_n623), .Y(new_n628));
  not_3  g0313(.A(new_n628), .Y(new_n629));
  nor_4  g0314(.A(new_n629), .B(new_n621), .Y(new_n630));
  nor_4  g0315(.A(new_n630), .B(new_n435), .Y(new_n631));
  nor_4  g0316(.A(new_n631), .B(new_n396_1), .Y(new_n632));
  not_3  g0317(.A(n1616), .Y(new_n633));
  not_3  g0318(.A(new_n368), .Y(new_n634));
  nand_4 g0319(.A(new_n634), .B(new_n633), .Y(new_n635));
  nor_4  g0320(.A(new_n379), .B(new_n358), .Y(new_n636));
  not_3  g0321(.A(new_n636), .Y(new_n637));
  nor_4  g0322(.A(new_n634), .B(new_n633), .Y(new_n638_1));
  nor_4  g0323(.A(new_n378_1), .B(new_n638_1), .Y(new_n639));
  nand_4 g0324(.A(new_n639), .B(new_n637), .Y(new_n640_1));
  nand_4 g0325(.A(new_n640_1), .B(new_n635), .Y(new_n641_1));
  nor_4  g0326(.A(new_n641_1), .B(new_n392_1), .Y(new_n642));
  nor_4  g0327(.A(new_n642), .B(new_n391_1), .Y(new_n643));
  nor_4  g0328(.A(new_n643), .B(new_n632), .Y(new_n644));
  nand_4 g0329(.A(new_n644), .B(new_n352_1), .Y(new_n645_1));
  nand_4 g0330(.A(new_n645_1), .B(new_n351), .Y(new_n646));
  nor_4  g0331(.A(new_n331), .B(new_n329), .Y(new_n647));
  nor_4  g0332(.A(new_n337_1), .B(new_n335), .Y(new_n648));
  not_3  g0333(.A(new_n648), .Y(new_n649));
  xor_3  g0334(.A(new_n340), .B(n980), .Y(new_n650));
  not_3  g0335(.A(new_n650), .Y(new_n651));
  nor_4  g0336(.A(new_n651), .B(new_n649), .Y(new_n652));
  nand_4 g0337(.A(new_n652), .B(new_n647), .Y(new_n653));
  nor_4  g0338(.A(new_n653), .B(new_n646), .Y(new_n654));
  nor_4  g0339(.A(new_n654), .B(new_n347), .Y(new_n655));
  xor_3  g0340(.A(new_n655), .B(new_n325), .Y(n22));
  not_3  g0341(.A(n1361), .Y(new_n657));
  nand_4 g0342(.A(n1387), .B(new_n657), .Y(n30));
  xor_3  g0343(.A(new_n620), .B(new_n439), .Y(n112));
  nand_4 g0344(.A(n1613), .B(n1520), .Y(new_n660));
  nand_4 g0345(.A(n574), .B(n284), .Y(new_n661));
  or_4   g0346(.A(new_n661), .B(new_n660), .Y(n126));
  nor_4  g0347(.A(new_n319), .B(n223), .Y(new_n663_1));
  nor_4  g0348(.A(new_n663_1), .B(new_n318_1), .Y(new_n664));
  not_3  g0349(.A(n300), .Y(new_n665));
  nor_4  g0350(.A(n1239), .B(new_n665), .Y(new_n666));
  nor_4  g0351(.A(n1470), .B(new_n319), .Y(new_n667));
  nor_4  g0352(.A(new_n667), .B(new_n666), .Y(new_n668));
  not_3  g0353(.A(new_n668), .Y(new_n669_1));
  nor_4  g0354(.A(new_n669_1), .B(new_n664), .Y(new_n670));
  nor_4  g0355(.A(new_n319), .B(n86), .Y(new_n671_1));
  nor_4  g0356(.A(new_n671_1), .B(new_n318_1), .Y(new_n672));
  not_3  g0357(.A(n561), .Y(new_n673));
  nor_4  g0358(.A(n1239), .B(new_n673), .Y(new_n674));
  nor_4  g0359(.A(new_n319), .B(n138), .Y(new_n675));
  or_4   g0360(.A(new_n675), .B(new_n674), .Y(new_n676_1));
  nor_4  g0361(.A(new_n676_1), .B(new_n672), .Y(new_n677));
  nor_4  g0362(.A(new_n677), .B(new_n670), .Y(new_n678));
  not_3  g0363(.A(new_n678), .Y(new_n679));
  nand_4 g0364(.A(new_n676_1), .B(new_n672), .Y(new_n680));
  nor_4  g0365(.A(n1299), .B(new_n319), .Y(new_n681));
  nor_4  g0366(.A(new_n681), .B(new_n318_1), .Y(new_n682));
  not_3  g0367(.A(n879), .Y(new_n683));
  nor_4  g0368(.A(n1239), .B(new_n683), .Y(new_n684));
  nor_4  g0369(.A(new_n319), .B(n769), .Y(new_n685));
  nor_4  g0370(.A(new_n685), .B(new_n684), .Y(new_n686));
  not_3  g0371(.A(new_n686), .Y(new_n687));
  nand_4 g0372(.A(new_n687), .B(new_n682), .Y(new_n688));
  nand_4 g0373(.A(new_n688), .B(new_n680), .Y(new_n689));
  nor_4  g0374(.A(n1502), .B(new_n319), .Y(new_n690_1));
  nor_4  g0375(.A(new_n690_1), .B(new_n318_1), .Y(new_n691));
  not_3  g0376(.A(n143), .Y(new_n692));
  nor_4  g0377(.A(n1239), .B(new_n692), .Y(new_n693_1));
  nor_4  g0378(.A(new_n319), .B(n626), .Y(new_n694));
  nor_4  g0379(.A(new_n694), .B(new_n693_1), .Y(new_n695_1));
  not_3  g0380(.A(new_n695_1), .Y(new_n696));
  nor_4  g0381(.A(new_n696), .B(new_n691), .Y(new_n697));
  nor_4  g0382(.A(new_n687), .B(new_n682), .Y(new_n698));
  nor_4  g0383(.A(new_n698), .B(new_n697), .Y(new_n699));
  not_3  g0384(.A(new_n699), .Y(new_n700));
  not_3  g0385(.A(n663), .Y(new_n701_1));
  nor_4  g0386(.A(n1239), .B(new_n701_1), .Y(new_n702));
  nor_4  g0387(.A(n1656), .B(new_n319), .Y(new_n703));
  nor_4  g0388(.A(new_n703), .B(new_n702), .Y(new_n704));
  nor_4  g0389(.A(new_n704), .B(new_n318_1), .Y(new_n705));
  not_3  g0390(.A(new_n691), .Y(new_n706));
  nor_4  g0391(.A(new_n695_1), .B(new_n706), .Y(new_n707));
  nor_4  g0392(.A(new_n707), .B(new_n705), .Y(new_n708));
  nor_4  g0393(.A(new_n708), .B(new_n700), .Y(new_n709));
  nor_4  g0394(.A(new_n709), .B(new_n689), .Y(new_n710_1));
  nor_4  g0395(.A(new_n710_1), .B(new_n679), .Y(new_n711));
  nor_4  g0396(.A(new_n319), .B(n787), .Y(new_n712));
  nor_4  g0397(.A(new_n712), .B(new_n318_1), .Y(new_n713));
  not_3  g0398(.A(n1164), .Y(new_n714_1));
  nor_4  g0399(.A(n1239), .B(new_n714_1), .Y(new_n715));
  nor_4  g0400(.A(new_n319), .B(n399), .Y(new_n716));
  nor_4  g0401(.A(new_n716), .B(new_n715), .Y(new_n717));
  not_3  g0402(.A(new_n717), .Y(new_n718));
  nor_4  g0403(.A(new_n718), .B(new_n713), .Y(new_n719_1));
  nor_4  g0404(.A(new_n319), .B(n727), .Y(new_n720));
  nor_4  g0405(.A(new_n720), .B(new_n318_1), .Y(new_n721));
  not_3  g0406(.A(n40), .Y(new_n722));
  nor_4  g0407(.A(n1239), .B(new_n722), .Y(new_n723));
  nor_4  g0408(.A(n1263), .B(new_n319), .Y(new_n724));
  nor_4  g0409(.A(new_n724), .B(new_n723), .Y(new_n725));
  not_3  g0410(.A(new_n725), .Y(new_n726_1));
  nor_4  g0411(.A(new_n726_1), .B(new_n721), .Y(new_n727_1));
  nor_4  g0412(.A(new_n319), .B(n94), .Y(new_n728));
  nor_4  g0413(.A(new_n728), .B(new_n318_1), .Y(new_n729_1));
  not_3  g0414(.A(n489), .Y(new_n730));
  nor_4  g0415(.A(n1239), .B(new_n730), .Y(new_n731));
  nor_4  g0416(.A(new_n319), .B(n346), .Y(new_n732));
  nor_4  g0417(.A(new_n732), .B(new_n731), .Y(new_n733));
  not_3  g0418(.A(new_n733), .Y(new_n734_1));
  nor_4  g0419(.A(new_n734_1), .B(new_n729_1), .Y(new_n735));
  nor_4  g0420(.A(new_n735), .B(new_n727_1), .Y(new_n736));
  not_3  g0421(.A(new_n736), .Y(new_n737));
  nor_4  g0422(.A(new_n737), .B(new_n719_1), .Y(new_n738));
  not_3  g0423(.A(new_n738), .Y(new_n739));
  not_3  g0424(.A(new_n713), .Y(new_n740));
  nor_4  g0425(.A(new_n717), .B(new_n740), .Y(new_n741));
  nor_4  g0426(.A(new_n319), .B(n609), .Y(new_n742_1));
  nor_4  g0427(.A(new_n742_1), .B(new_n318_1), .Y(new_n743_1));
  not_3  g0428(.A(new_n743_1), .Y(new_n744));
  not_3  g0429(.A(n71), .Y(new_n745));
  nor_4  g0430(.A(n1239), .B(new_n745), .Y(new_n746));
  nor_4  g0431(.A(new_n319), .B(n980), .Y(new_n747));
  nor_4  g0432(.A(new_n747), .B(new_n746), .Y(new_n748));
  nor_4  g0433(.A(new_n748), .B(new_n744), .Y(new_n749));
  nor_4  g0434(.A(new_n749), .B(new_n741), .Y(new_n750));
  nor_4  g0435(.A(new_n750), .B(new_n739), .Y(new_n751));
  not_3  g0436(.A(new_n721), .Y(new_n752));
  nor_4  g0437(.A(new_n725), .B(new_n752), .Y(new_n753));
  not_3  g0438(.A(new_n729_1), .Y(new_n754));
  nor_4  g0439(.A(new_n733), .B(new_n754), .Y(new_n755_1));
  nor_4  g0440(.A(new_n755_1), .B(new_n753), .Y(new_n756));
  nor_4  g0441(.A(new_n756), .B(new_n727_1), .Y(new_n757));
  nor_4  g0442(.A(new_n757), .B(new_n751), .Y(new_n758));
  nor_4  g0443(.A(new_n319), .B(n839), .Y(new_n759));
  nor_4  g0444(.A(new_n759), .B(new_n318_1), .Y(new_n760));
  not_3  g0445(.A(new_n760), .Y(new_n761));
  not_3  g0446(.A(n1523), .Y(new_n762));
  nor_4  g0447(.A(new_n762), .B(n1239), .Y(new_n763));
  nor_4  g0448(.A(new_n319), .B(n318), .Y(new_n764));
  nor_4  g0449(.A(new_n764), .B(new_n763), .Y(new_n765));
  nand_4 g0450(.A(new_n765), .B(new_n761), .Y(new_n766));
  not_3  g0451(.A(new_n750), .Y(new_n767));
  not_3  g0452(.A(new_n748), .Y(new_n768));
  nor_4  g0453(.A(new_n768), .B(new_n743_1), .Y(new_n769_1));
  nor_4  g0454(.A(new_n769_1), .B(new_n767), .Y(new_n770));
  nand_4 g0455(.A(new_n770), .B(new_n738), .Y(new_n771));
  nor_4  g0456(.A(new_n765), .B(new_n761), .Y(new_n772));
  nand_4 g0457(.A(n1239), .B(n953), .Y(new_n773_1));
  not_3  g0458(.A(new_n773_1), .Y(new_n774));
  nor_4  g0459(.A(new_n774), .B(new_n389), .Y(new_n775_1));
  not_3  g0460(.A(n1305), .Y(new_n776));
  nor_4  g0461(.A(new_n776), .B(n1239), .Y(new_n777));
  nor_4  g0462(.A(n1592), .B(new_n319), .Y(new_n778_1));
  nor_4  g0463(.A(new_n778_1), .B(new_n777), .Y(new_n779_1));
  nor_4  g0464(.A(new_n779_1), .B(new_n775_1), .Y(new_n780));
  nor_4  g0465(.A(new_n780), .B(new_n772), .Y(new_n781));
  and_4  g0466(.A(new_n779_1), .B(new_n775_1), .Y(new_n782_1));
  nand_4 g0467(.A(n1239), .B(n52), .Y(new_n783));
  not_3  g0468(.A(new_n783), .Y(new_n784));
  nor_4  g0469(.A(new_n784), .B(new_n367), .Y(new_n785));
  not_3  g0470(.A(n1418), .Y(new_n786));
  nor_4  g0471(.A(new_n786), .B(n1239), .Y(new_n787_1));
  nor_4  g0472(.A(n1616), .B(new_n319), .Y(new_n788));
  nor_4  g0473(.A(new_n788), .B(new_n787_1), .Y(new_n789));
  nor_4  g0474(.A(new_n789), .B(new_n785), .Y(new_n790_1));
  not_3  g0475(.A(new_n785), .Y(new_n791));
  not_3  g0476(.A(new_n789), .Y(new_n792));
  nor_4  g0477(.A(new_n792), .B(new_n791), .Y(new_n793));
  nand_4 g0478(.A(n1428), .B(n1239), .Y(new_n794_1));
  not_3  g0479(.A(new_n794_1), .Y(new_n795));
  nor_4  g0480(.A(new_n795), .B(new_n375), .Y(new_n796));
  not_3  g0481(.A(new_n796), .Y(new_n797));
  not_3  g0482(.A(n1156), .Y(new_n798));
  nor_4  g0483(.A(n1239), .B(new_n798), .Y(new_n799));
  nor_4  g0484(.A(n1446), .B(new_n319), .Y(new_n800));
  nor_4  g0485(.A(new_n800), .B(new_n799), .Y(new_n801));
  not_3  g0486(.A(new_n801), .Y(new_n802));
  nor_4  g0487(.A(new_n802), .B(new_n797), .Y(new_n803));
  nor_4  g0488(.A(new_n803), .B(new_n793), .Y(new_n804));
  nor_4  g0489(.A(new_n801), .B(new_n796), .Y(new_n805));
  nand_4 g0490(.A(n1239), .B(n607), .Y(new_n806));
  not_3  g0491(.A(new_n806), .Y(new_n807));
  nor_4  g0492(.A(new_n807), .B(new_n356), .Y(new_n808));
  not_3  g0493(.A(n969), .Y(new_n809));
  nor_4  g0494(.A(n1239), .B(new_n809), .Y(new_n810));
  nor_4  g0495(.A(n1345), .B(new_n319), .Y(new_n811));
  nor_4  g0496(.A(new_n811), .B(new_n810), .Y(new_n812));
  nor_4  g0497(.A(new_n812), .B(new_n808), .Y(new_n813));
  nor_4  g0498(.A(new_n813), .B(new_n805), .Y(new_n814));
  not_3  g0499(.A(new_n814), .Y(new_n815));
  and_4  g0500(.A(new_n815), .B(new_n804), .Y(new_n816));
  nor_4  g0501(.A(new_n816), .B(new_n790_1), .Y(new_n817));
  or_4   g0502(.A(new_n817), .B(new_n782_1), .Y(new_n818));
  nand_4 g0503(.A(new_n818), .B(new_n781), .Y(new_n819));
  nand_4 g0504(.A(n1239), .B(n376), .Y(new_n820));
  not_3  g0505(.A(new_n820), .Y(new_n821_1));
  nor_4  g0506(.A(new_n821_1), .B(new_n400), .Y(new_n822));
  not_3  g0507(.A(new_n822), .Y(new_n823_1));
  not_3  g0508(.A(n779), .Y(new_n824));
  nor_4  g0509(.A(n1239), .B(new_n824), .Y(new_n825));
  nor_4  g0510(.A(n1301), .B(new_n319), .Y(new_n826));
  nor_4  g0511(.A(new_n826), .B(new_n825), .Y(new_n827));
  not_3  g0512(.A(new_n827), .Y(new_n828));
  nor_4  g0513(.A(new_n828), .B(new_n823_1), .Y(new_n829));
  not_3  g0514(.A(new_n829), .Y(new_n830));
  nor_4  g0515(.A(new_n827), .B(new_n822), .Y(new_n831_1));
  nand_4 g0516(.A(n1239), .B(n273), .Y(new_n832_1));
  not_3  g0517(.A(new_n832_1), .Y(new_n833));
  nor_4  g0518(.A(new_n833), .B(new_n409_1), .Y(new_n834));
  not_3  g0519(.A(n507), .Y(new_n835));
  nor_4  g0520(.A(n1239), .B(new_n835), .Y(new_n836));
  nor_4  g0521(.A(n1566), .B(new_n319), .Y(new_n837));
  nor_4  g0522(.A(new_n837), .B(new_n836), .Y(new_n838));
  nor_4  g0523(.A(new_n838), .B(new_n834), .Y(new_n839_1));
  nor_4  g0524(.A(new_n839_1), .B(new_n831_1), .Y(new_n840));
  and_4  g0525(.A(new_n838), .B(new_n834), .Y(new_n841));
  nand_4 g0526(.A(n1239), .B(n885), .Y(new_n842_1));
  not_3  g0527(.A(new_n842_1), .Y(new_n843));
  nor_4  g0528(.A(new_n843), .B(new_n418), .Y(new_n844));
  not_3  g0529(.A(n107), .Y(new_n845));
  nor_4  g0530(.A(n1239), .B(new_n845), .Y(new_n846));
  nor_4  g0531(.A(new_n319), .B(n920), .Y(new_n847));
  nor_4  g0532(.A(new_n847), .B(new_n846), .Y(new_n848));
  and_4  g0533(.A(new_n848), .B(new_n844), .Y(new_n849_1));
  nor_4  g0534(.A(new_n849_1), .B(new_n841), .Y(new_n850));
  nor_4  g0535(.A(new_n848), .B(new_n844), .Y(new_n851));
  nand_4 g0536(.A(n1239), .B(n50), .Y(new_n852));
  not_3  g0537(.A(new_n852), .Y(new_n853));
  nor_4  g0538(.A(new_n853), .B(new_n424), .Y(new_n854));
  not_3  g0539(.A(n1448), .Y(new_n855));
  nor_4  g0540(.A(new_n855), .B(n1239), .Y(new_n856));
  nor_4  g0541(.A(new_n319), .B(n293), .Y(new_n857));
  nor_4  g0542(.A(new_n857), .B(new_n856), .Y(new_n858));
  nor_4  g0543(.A(new_n858), .B(new_n854), .Y(new_n859));
  nor_4  g0544(.A(new_n859), .B(new_n851), .Y(new_n860));
  nand_4 g0545(.A(n1239), .B(n734), .Y(new_n861));
  not_3  g0546(.A(new_n861), .Y(new_n862));
  nor_4  g0547(.A(new_n862), .B(new_n443), .Y(new_n863));
  not_3  g0548(.A(new_n863), .Y(new_n864));
  not_3  g0549(.A(n1152), .Y(new_n865));
  nor_4  g0550(.A(n1239), .B(new_n865), .Y(new_n866));
  nor_4  g0551(.A(new_n319), .B(n408), .Y(new_n867));
  nor_4  g0552(.A(new_n867), .B(new_n866), .Y(new_n868));
  not_3  g0553(.A(new_n868), .Y(new_n869));
  nor_4  g0554(.A(new_n869), .B(new_n864), .Y(new_n870));
  and_4  g0555(.A(new_n858), .B(new_n854), .Y(new_n871));
  nor_4  g0556(.A(new_n871), .B(new_n870), .Y(new_n872));
  nand_4 g0557(.A(n1586), .B(n1239), .Y(new_n873));
  not_3  g0558(.A(new_n873), .Y(new_n874));
  nor_4  g0559(.A(new_n874), .B(new_n451), .Y(new_n875));
  not_3  g0560(.A(n1386), .Y(new_n876));
  nor_4  g0561(.A(new_n876), .B(n1239), .Y(new_n877));
  nor_4  g0562(.A(n1476), .B(new_n319), .Y(new_n878));
  nor_4  g0563(.A(new_n878), .B(new_n877), .Y(new_n879_1));
  nor_4  g0564(.A(new_n879_1), .B(new_n875), .Y(new_n880));
  not_3  g0565(.A(new_n880), .Y(new_n881));
  nor_4  g0566(.A(new_n868), .B(new_n863), .Y(new_n882_1));
  nand_4 g0567(.A(n1239), .B(n1114), .Y(new_n883));
  not_3  g0568(.A(new_n883), .Y(new_n884));
  nor_4  g0569(.A(new_n884), .B(new_n478_1), .Y(new_n885_1));
  not_3  g0570(.A(n1627), .Y(new_n886));
  nor_4  g0571(.A(new_n886), .B(n1239), .Y(new_n887));
  nor_4  g0572(.A(new_n319), .B(n153), .Y(new_n888));
  nor_4  g0573(.A(new_n888), .B(new_n887), .Y(new_n889));
  nor_4  g0574(.A(new_n889), .B(new_n885_1), .Y(new_n890));
  nand_4 g0575(.A(n1239), .B(n77), .Y(new_n891));
  not_3  g0576(.A(new_n891), .Y(new_n892));
  nor_4  g0577(.A(new_n892), .B(new_n469), .Y(new_n893));
  not_3  g0578(.A(n882), .Y(new_n894_1));
  nor_4  g0579(.A(n1239), .B(new_n894_1), .Y(new_n895));
  nor_4  g0580(.A(new_n319), .B(n823), .Y(new_n896));
  nor_4  g0581(.A(new_n896), .B(new_n895), .Y(new_n897));
  nor_4  g0582(.A(new_n897), .B(new_n893), .Y(new_n898));
  nor_4  g0583(.A(new_n898), .B(new_n890), .Y(new_n899));
  not_3  g0584(.A(new_n899), .Y(new_n900));
  nand_4 g0585(.A(n1239), .B(n344), .Y(new_n901));
  not_3  g0586(.A(new_n901), .Y(new_n902));
  nor_4  g0587(.A(new_n902), .B(new_n458), .Y(new_n903));
  not_3  g0588(.A(n1227), .Y(new_n904));
  nor_4  g0589(.A(n1239), .B(new_n904), .Y(new_n905_1));
  nor_4  g0590(.A(n1401), .B(new_n319), .Y(new_n906));
  nor_4  g0591(.A(new_n906), .B(new_n905_1), .Y(new_n907));
  or_4   g0592(.A(new_n907), .B(new_n903), .Y(new_n908));
  not_3  g0593(.A(new_n885_1), .Y(new_n909));
  not_3  g0594(.A(new_n889), .Y(new_n910));
  nor_4  g0595(.A(new_n910), .B(new_n909), .Y(new_n911));
  nor_4  g0596(.A(new_n911), .B(new_n908), .Y(new_n912));
  nor_4  g0597(.A(new_n912), .B(new_n900), .Y(new_n913));
  and_4  g0598(.A(new_n897), .B(new_n893), .Y(new_n914));
  and_4  g0599(.A(new_n879_1), .B(new_n875), .Y(new_n915));
  or_4   g0600(.A(new_n915), .B(new_n914), .Y(new_n916_1));
  nor_4  g0601(.A(new_n916_1), .B(new_n913), .Y(new_n917));
  nor_4  g0602(.A(new_n917), .B(new_n882_1), .Y(new_n918_1));
  nand_4 g0603(.A(new_n918_1), .B(new_n881), .Y(new_n919));
  nand_4 g0604(.A(new_n919), .B(new_n872), .Y(new_n920_1));
  nand_4 g0605(.A(new_n920_1), .B(new_n860), .Y(new_n921));
  nand_4 g0606(.A(new_n921), .B(new_n850), .Y(new_n922));
  nand_4 g0607(.A(new_n922), .B(new_n840), .Y(new_n923));
  nand_4 g0608(.A(new_n923), .B(new_n830), .Y(new_n924));
  nand_4 g0609(.A(n1239), .B(n288), .Y(new_n925));
  not_3  g0610(.A(new_n925), .Y(new_n926));
  nor_4  g0611(.A(new_n926), .B(new_n502_1), .Y(new_n927));
  not_3  g0612(.A(new_n927), .Y(new_n928));
  not_3  g0613(.A(n936), .Y(new_n929));
  nor_4  g0614(.A(n1239), .B(new_n929), .Y(new_n930));
  nor_4  g0615(.A(new_n319), .B(n567), .Y(new_n931));
  nor_4  g0616(.A(new_n931), .B(new_n930), .Y(new_n932));
  not_3  g0617(.A(new_n932), .Y(new_n933));
  nand_4 g0618(.A(new_n933), .B(new_n928), .Y(new_n934));
  nor_4  g0619(.A(new_n933), .B(new_n928), .Y(new_n935));
  nand_4 g0620(.A(n1239), .B(n416), .Y(new_n936_1));
  not_3  g0621(.A(new_n936_1), .Y(new_n937));
  nor_4  g0622(.A(new_n937), .B(new_n512), .Y(new_n938));
  not_3  g0623(.A(n159), .Y(new_n939));
  nor_4  g0624(.A(n1239), .B(new_n939), .Y(new_n940));
  nor_4  g0625(.A(n1463), .B(new_n319), .Y(new_n941));
  nor_4  g0626(.A(new_n941), .B(new_n940), .Y(new_n942));
  or_4   g0627(.A(new_n942), .B(new_n938), .Y(new_n943));
  nand_4 g0628(.A(n1239), .B(n506), .Y(new_n944));
  not_3  g0629(.A(new_n944), .Y(new_n945));
  nor_4  g0630(.A(new_n945), .B(new_n522), .Y(new_n946));
  not_3  g0631(.A(n243), .Y(new_n947_1));
  nor_4  g0632(.A(n1239), .B(new_n947_1), .Y(new_n948));
  nor_4  g0633(.A(new_n319), .B(n222), .Y(new_n949));
  nor_4  g0634(.A(new_n949), .B(new_n948), .Y(new_n950));
  nand_4 g0635(.A(new_n950), .B(new_n946), .Y(new_n951));
  or_4   g0636(.A(new_n950), .B(new_n946), .Y(new_n952_1));
  nand_4 g0637(.A(n1239), .B(n671), .Y(new_n953_1));
  not_3  g0638(.A(new_n953_1), .Y(new_n954));
  nor_4  g0639(.A(new_n954), .B(new_n544), .Y(new_n955));
  not_3  g0640(.A(n341), .Y(new_n956));
  nor_4  g0641(.A(n1239), .B(new_n956), .Y(new_n957));
  nor_4  g0642(.A(new_n319), .B(n1071), .Y(new_n958));
  nor_4  g0643(.A(new_n958), .B(new_n957), .Y(new_n959));
  or_4   g0644(.A(new_n959), .B(new_n955), .Y(new_n960));
  nand_4 g0645(.A(n1239), .B(n392), .Y(new_n961_1));
  not_3  g0646(.A(new_n961_1), .Y(new_n962));
  nor_4  g0647(.A(new_n962), .B(new_n534_1), .Y(new_n963));
  not_3  g0648(.A(n742), .Y(new_n964));
  nor_4  g0649(.A(n1239), .B(new_n964), .Y(new_n965));
  nor_4  g0650(.A(new_n319), .B(n608), .Y(new_n966));
  nor_4  g0651(.A(new_n966), .B(new_n965), .Y(new_n967));
  nor_4  g0652(.A(new_n967), .B(new_n963), .Y(new_n968));
  nand_4 g0653(.A(n1239), .B(n29), .Y(new_n969_1));
  not_3  g0654(.A(new_n969_1), .Y(new_n970));
  nor_4  g0655(.A(new_n970), .B(new_n555), .Y(new_n971));
  not_3  g0656(.A(new_n971), .Y(new_n972));
  not_3  g0657(.A(n849), .Y(new_n973));
  nor_4  g0658(.A(n1239), .B(new_n973), .Y(new_n974));
  nor_4  g0659(.A(new_n319), .B(n45), .Y(new_n975));
  nor_4  g0660(.A(new_n975), .B(new_n974), .Y(new_n976));
  not_3  g0661(.A(new_n976), .Y(new_n977));
  nor_4  g0662(.A(new_n977), .B(new_n972), .Y(new_n978));
  nand_4 g0663(.A(n1239), .B(n778), .Y(new_n979));
  not_3  g0664(.A(new_n979), .Y(new_n980_1));
  nor_4  g0665(.A(new_n980_1), .B(new_n563), .Y(new_n981));
  not_3  g0666(.A(n502), .Y(new_n982));
  nor_4  g0667(.A(n1239), .B(new_n982), .Y(new_n983));
  nor_4  g0668(.A(new_n319), .B(n695), .Y(new_n984_1));
  nor_4  g0669(.A(new_n984_1), .B(new_n983), .Y(new_n985));
  nand_4 g0670(.A(new_n985), .B(new_n981), .Y(new_n986_1));
  not_3  g0671(.A(n690), .Y(new_n987));
  nor_4  g0672(.A(n1239), .B(n729), .Y(new_n988));
  or_4   g0673(.A(new_n988), .B(new_n987), .Y(new_n989));
  not_3  g0674(.A(new_n570), .Y(new_n990_1));
  or_4   g0675(.A(n729), .B(n690), .Y(new_n991));
  nand_4 g0676(.A(new_n991), .B(new_n990_1), .Y(new_n992_1));
  nand_4 g0677(.A(new_n992_1), .B(new_n989), .Y(new_n993));
  nand_4 g0678(.A(new_n993), .B(new_n986_1), .Y(new_n994));
  nor_4  g0679(.A(new_n976), .B(new_n971), .Y(new_n995));
  nor_4  g0680(.A(new_n985), .B(new_n981), .Y(new_n996));
  nor_4  g0681(.A(new_n996), .B(new_n995), .Y(new_n997_1));
  nand_4 g0682(.A(new_n997_1), .B(new_n994), .Y(new_n998));
  nand_4 g0683(.A(new_n959), .B(new_n955), .Y(new_n999));
  nand_4 g0684(.A(new_n999), .B(new_n998), .Y(new_n1000));
  nor_4  g0685(.A(new_n1000), .B(new_n978), .Y(new_n1001));
  nor_4  g0686(.A(new_n1001), .B(new_n968), .Y(new_n1002));
  nand_4 g0687(.A(new_n1002), .B(new_n960), .Y(new_n1003));
  nand_4 g0688(.A(new_n967), .B(new_n963), .Y(new_n1004));
  nand_4 g0689(.A(new_n1004), .B(new_n1003), .Y(new_n1005));
  nand_4 g0690(.A(new_n1005), .B(new_n952_1), .Y(new_n1006_1));
  nand_4 g0691(.A(new_n1006_1), .B(new_n951), .Y(new_n1007));
  nand_4 g0692(.A(new_n1007), .B(new_n943), .Y(new_n1008));
  nand_4 g0693(.A(new_n942), .B(new_n938), .Y(new_n1009));
  nand_4 g0694(.A(new_n1009), .B(new_n1008), .Y(new_n1010));
  nor_4  g0695(.A(new_n1010), .B(new_n935), .Y(new_n1011));
  nand_4 g0696(.A(n1753), .B(n1239), .Y(new_n1012));
  not_3  g0697(.A(new_n1012), .Y(new_n1013));
  nor_4  g0698(.A(new_n1013), .B(new_n493), .Y(new_n1014));
  not_3  g0699(.A(n755), .Y(new_n1015));
  nor_4  g0700(.A(n1239), .B(new_n1015), .Y(new_n1016));
  nor_4  g0701(.A(new_n319), .B(n374), .Y(new_n1017_1));
  nor_4  g0702(.A(new_n1017_1), .B(new_n1016), .Y(new_n1018));
  nor_4  g0703(.A(new_n1018), .B(new_n1014), .Y(new_n1019));
  nor_4  g0704(.A(new_n1019), .B(new_n1011), .Y(new_n1020));
  nand_4 g0705(.A(new_n1020), .B(new_n934), .Y(new_n1021));
  nand_4 g0706(.A(new_n1018), .B(new_n1014), .Y(new_n1022));
  nor_4  g0707(.A(new_n911), .B(new_n882_1), .Y(new_n1023_1));
  nand_4 g0708(.A(new_n1023_1), .B(new_n1022), .Y(new_n1024));
  nand_4 g0709(.A(new_n872), .B(new_n860), .Y(new_n1025));
  nor_4  g0710(.A(new_n1025), .B(new_n916_1), .Y(new_n1026));
  nor_4  g0711(.A(new_n880), .B(new_n829), .Y(new_n1027));
  nand_4 g0712(.A(new_n1027), .B(new_n840), .Y(new_n1028));
  and_4  g0713(.A(new_n899), .B(new_n850), .Y(new_n1029));
  xor_3  g0714(.A(new_n907), .B(new_n903), .Y(new_n1030));
  nand_4 g0715(.A(new_n1030), .B(new_n1029), .Y(new_n1031));
  nor_4  g0716(.A(new_n1031), .B(new_n1028), .Y(new_n1032));
  nand_4 g0717(.A(new_n1032), .B(new_n1026), .Y(new_n1033));
  nor_4  g0718(.A(new_n1033), .B(new_n1024), .Y(new_n1034));
  nand_4 g0719(.A(new_n1034), .B(new_n1021), .Y(new_n1035));
  nand_4 g0720(.A(new_n1035), .B(new_n924), .Y(n1306));
  nand_4 g0721(.A(new_n812), .B(new_n808), .Y(new_n1037));
  and_4  g0722(.A(new_n814), .B(new_n781), .Y(new_n1038));
  nand_4 g0723(.A(new_n1038), .B(new_n1037), .Y(new_n1039));
  nor_4  g0724(.A(new_n790_1), .B(new_n782_1), .Y(new_n1040_1));
  nand_4 g0725(.A(new_n1040_1), .B(new_n804), .Y(new_n1041));
  nor_4  g0726(.A(new_n1041), .B(new_n1039), .Y(new_n1042_1));
  nand_4 g0727(.A(new_n1042_1), .B(n1306), .Y(new_n1043));
  not_3  g0728(.A(new_n1043), .Y(new_n1044_1));
  nor_4  g0729(.A(new_n1044_1), .B(new_n819), .Y(new_n1045));
  nor_4  g0730(.A(new_n1045), .B(new_n771), .Y(new_n1046));
  nand_4 g0731(.A(new_n1046), .B(new_n766), .Y(new_n1047));
  nand_4 g0732(.A(new_n1047), .B(new_n758), .Y(new_n1048));
  nand_4 g0733(.A(new_n704), .B(new_n318_1), .Y(new_n1049));
  nand_4 g0734(.A(new_n1049), .B(new_n708), .Y(new_n1050_1));
  not_3  g0735(.A(new_n664), .Y(new_n1051_1));
  nor_4  g0736(.A(new_n668), .B(new_n1051_1), .Y(new_n1052));
  or_4   g0737(.A(new_n1052), .B(new_n700), .Y(new_n1053));
  nor_4  g0738(.A(new_n1053), .B(new_n689), .Y(new_n1054_1));
  nand_4 g0739(.A(new_n1054_1), .B(new_n678), .Y(new_n1055));
  nor_4  g0740(.A(new_n1055), .B(new_n1050_1), .Y(new_n1056));
  nand_4 g0741(.A(new_n1056), .B(new_n1048), .Y(new_n1057));
  not_3  g0742(.A(n986), .Y(new_n1058_1));
  nor_4  g0743(.A(n589), .B(n559), .Y(new_n1059));
  and_4  g0744(.A(new_n1059), .B(n156), .Y(new_n1060_1));
  or_4   g0745(.A(new_n1060_1), .B(new_n1058_1), .Y(new_n1061_1));
  not_3  g0746(.A(new_n1061_1), .Y(new_n1062));
  nor_4  g0747(.A(new_n1062), .B(new_n1052), .Y(new_n1063_1));
  nand_4 g0748(.A(new_n1063_1), .B(new_n1057), .Y(new_n1064));
  nor_4  g0749(.A(new_n1064), .B(new_n711), .Y(new_n1065_1));
  nand_4 g0750(.A(n589), .B(n559), .Y(new_n1066));
  nand_4 g0751(.A(new_n1066), .B(n156), .Y(new_n1067));
  nor_4  g0752(.A(new_n1067), .B(n986), .Y(new_n1068));
  nor_4  g0753(.A(new_n1068), .B(new_n1065_1), .Y(n161));
  xor_3  g0754(.A(new_n350), .B(new_n348), .Y(new_n1070));
  not_3  g0755(.A(new_n1070), .Y(new_n1071_1));
  xor_3  g0756(.A(new_n1071_1), .B(new_n644), .Y(n164));
  xor_3  g0757(.A(new_n651), .B(new_n646), .Y(n181));
  nor_4  g0758(.A(new_n319), .B(n477), .Y(new_n1074));
  nor_4  g0759(.A(new_n1074), .B(new_n318_1), .Y(new_n1075));
  not_3  g0760(.A(new_n1075), .Y(new_n1076));
  nor_4  g0761(.A(new_n1076), .B(n769), .Y(new_n1077));
  not_3  g0762(.A(n769), .Y(new_n1078));
  nor_4  g0763(.A(new_n1075), .B(new_n1078), .Y(new_n1079));
  nor_4  g0764(.A(new_n1079), .B(new_n1077), .Y(new_n1080));
  not_3  g0765(.A(n626), .Y(new_n1081));
  nor_4  g0766(.A(new_n319), .B(n1191), .Y(new_n1082));
  nor_4  g0767(.A(new_n1082), .B(new_n318_1), .Y(new_n1083));
  nand_4 g0768(.A(new_n1083), .B(new_n1081), .Y(new_n1084));
  not_3  g0769(.A(new_n1084), .Y(new_n1085));
  nor_4  g0770(.A(new_n319), .B(n430), .Y(new_n1086));
  nor_4  g0771(.A(new_n1086), .B(new_n318_1), .Y(new_n1087));
  not_3  g0772(.A(new_n1087), .Y(new_n1088));
  nor_4  g0773(.A(new_n1088), .B(n1656), .Y(new_n1089));
  nor_4  g0774(.A(new_n1089), .B(new_n1085), .Y(new_n1090));
  nand_4 g0775(.A(new_n655), .B(new_n322), .Y(new_n1091));
  nand_4 g0776(.A(new_n1091), .B(new_n324), .Y(new_n1092));
  nand_4 g0777(.A(new_n1092), .B(new_n1090), .Y(new_n1093));
  nor_4  g0778(.A(new_n1083), .B(new_n1081), .Y(new_n1094));
  not_3  g0779(.A(n1656), .Y(new_n1095_1));
  nor_4  g0780(.A(new_n1087), .B(new_n1095_1), .Y(new_n1096));
  nor_4  g0781(.A(new_n1096), .B(new_n1094), .Y(new_n1097));
  nor_4  g0782(.A(new_n1097), .B(new_n1085), .Y(new_n1098));
  not_3  g0783(.A(new_n1098), .Y(new_n1099));
  nand_4 g0784(.A(new_n1099), .B(new_n1093), .Y(new_n1100));
  xnor_3 g0785(.A(new_n1100), .B(new_n1080), .Y(n216));
  not_3  g0786(.A(new_n574_1), .Y(new_n1102));
  nor_4  g0787(.A(new_n573), .B(new_n557), .Y(new_n1103_1));
  nor_4  g0788(.A(new_n1103_1), .B(new_n1102), .Y(new_n1104));
  not_3  g0789(.A(new_n590), .Y(new_n1105));
  nor_4  g0790(.A(new_n539), .B(new_n537), .Y(new_n1106));
  xor_3  g0791(.A(new_n1106), .B(new_n1105), .Y(new_n1107));
  not_3  g0792(.A(new_n1107), .Y(new_n1108));
  xor_3  g0793(.A(new_n1108), .B(new_n588), .Y(new_n1109));
  nor_4  g0794(.A(new_n1109), .B(new_n571), .Y(new_n1110));
  nor_4  g0795(.A(new_n1108), .B(new_n585_1), .Y(new_n1111));
  nor_4  g0796(.A(new_n1111), .B(new_n1110), .Y(new_n1112));
  xor_3  g0797(.A(new_n1112), .B(new_n1104), .Y(new_n1113));
  not_3  g0798(.A(new_n577), .Y(new_n1114_1));
  xor_3  g0799(.A(new_n582_1), .B(new_n579), .Y(new_n1115));
  xor_3  g0800(.A(new_n1115), .B(new_n1114_1), .Y(new_n1116));
  nor_4  g0801(.A(new_n1116), .B(new_n1113), .Y(new_n1117));
  nand_4 g0802(.A(new_n1116), .B(new_n1113), .Y(new_n1118));
  nand_4 g0803(.A(new_n1118), .B(new_n584), .Y(new_n1119));
  nor_4  g0804(.A(new_n1119), .B(new_n1117), .Y(new_n1120));
  nor_4  g0805(.A(new_n587), .B(new_n580), .Y(new_n1121_1));
  nor_4  g0806(.A(new_n1121_1), .B(new_n581_1), .Y(new_n1122));
  xor_3  g0807(.A(new_n1122), .B(new_n1115), .Y(new_n1123));
  not_3  g0808(.A(new_n587), .Y(new_n1124));
  nand_4 g0809(.A(new_n1124), .B(new_n575), .Y(new_n1125));
  not_3  g0810(.A(new_n575), .Y(new_n1126));
  nor_4  g0811(.A(new_n588), .B(new_n583), .Y(new_n1127));
  nor_4  g0812(.A(new_n1127), .B(new_n1124), .Y(new_n1128));
  nand_4 g0813(.A(new_n1128), .B(new_n1126), .Y(new_n1129));
  nand_4 g0814(.A(new_n1129), .B(new_n1125), .Y(new_n1130));
  xor_3  g0815(.A(new_n1130), .B(new_n1123), .Y(new_n1131));
  not_3  g0816(.A(new_n1109), .Y(new_n1132));
  not_3  g0817(.A(new_n1127), .Y(new_n1133));
  nor_4  g0818(.A(new_n1133), .B(new_n550), .Y(new_n1134));
  nor_4  g0819(.A(new_n1134), .B(new_n577), .Y(new_n1135));
  xor_3  g0820(.A(new_n1135), .B(new_n1132), .Y(new_n1136));
  nor_4  g0821(.A(new_n1136), .B(new_n1131), .Y(new_n1137));
  nand_4 g0822(.A(new_n1136), .B(new_n1131), .Y(new_n1138_1));
  nand_4 g0823(.A(new_n1138_1), .B(n545), .Y(new_n1139));
  nor_4  g0824(.A(new_n1139), .B(new_n1137), .Y(new_n1140));
  nor_4  g0825(.A(new_n1140), .B(new_n1120), .Y(new_n1141));
  nor_4  g0826(.A(new_n599), .B(new_n507_1), .Y(new_n1142));
  nor_4  g0827(.A(new_n1142), .B(new_n505), .Y(new_n1143));
  not_3  g0828(.A(new_n529), .Y(new_n1144));
  not_3  g0829(.A(new_n527), .Y(new_n1145));
  nor_4  g0830(.A(new_n1145), .B(new_n517_1), .Y(new_n1146));
  nor_4  g0831(.A(new_n527), .B(new_n514), .Y(new_n1147));
  nor_4  g0832(.A(new_n1147), .B(new_n1146), .Y(new_n1148));
  nor_4  g0833(.A(new_n1148), .B(new_n1144), .Y(new_n1149));
  xor_3  g0834(.A(new_n494), .B(n374), .Y(new_n1150));
  not_3  g0835(.A(new_n1150), .Y(new_n1151));
  xor_3  g0836(.A(new_n1151), .B(new_n1149), .Y(new_n1152_1));
  xor_3  g0837(.A(new_n1152_1), .B(new_n1143), .Y(new_n1153));
  nand_4 g0838(.A(new_n1153), .B(new_n595_1), .Y(new_n1154_1));
  not_3  g0839(.A(new_n595_1), .Y(new_n1155));
  nor_4  g0840(.A(new_n600_1), .B(new_n1144), .Y(new_n1156_1));
  nor_4  g0841(.A(new_n1156_1), .B(new_n505), .Y(new_n1157));
  and_4  g0842(.A(new_n1156_1), .B(new_n508), .Y(new_n1158));
  nor_4  g0843(.A(new_n1158), .B(new_n1157), .Y(new_n1159));
  nor_4  g0844(.A(new_n524), .B(new_n518), .Y(new_n1160));
  not_3  g0845(.A(new_n598_1), .Y(new_n1161));
  nor_4  g0846(.A(new_n1161), .B(new_n514), .Y(new_n1162));
  nor_4  g0847(.A(new_n1162), .B(new_n1160), .Y(new_n1163));
  nor_4  g0848(.A(new_n507_1), .B(new_n505), .Y(new_n1164_1));
  not_3  g0849(.A(new_n1164_1), .Y(new_n1165));
  xor_3  g0850(.A(new_n1165), .B(new_n1151), .Y(new_n1166));
  xor_3  g0851(.A(new_n1166), .B(new_n1163), .Y(new_n1167));
  xor_3  g0852(.A(new_n1167), .B(new_n1159), .Y(new_n1168));
  nand_4 g0853(.A(new_n1168), .B(new_n1155), .Y(new_n1169));
  nand_4 g0854(.A(new_n1169), .B(new_n1154_1), .Y(new_n1170));
  xnor_3 g0855(.A(new_n1170), .B(new_n1141), .Y(n233));
  xor_3  g0856(.A(new_n452), .B(new_n447), .Y(new_n1172_1));
  not_3  g0857(.A(new_n606), .Y(new_n1173));
  nor_4  g0858(.A(new_n1173), .B(new_n465), .Y(new_n1174));
  nor_4  g0859(.A(new_n1174), .B(new_n460_1), .Y(new_n1175_1));
  nor_4  g0860(.A(new_n1175_1), .B(new_n483), .Y(new_n1176));
  nor_4  g0861(.A(new_n1176), .B(new_n481), .Y(new_n1177_1));
  nor_4  g0862(.A(new_n1177_1), .B(new_n474), .Y(new_n1178));
  nor_4  g0863(.A(new_n1178), .B(new_n472), .Y(new_n1179));
  xor_3  g0864(.A(new_n1179), .B(new_n1172_1), .Y(n247));
  not_3  g0865(.A(n992), .Y(n275));
  nand_4 g0866(.A(n832), .B(n420), .Y(new_n1182));
  not_3  g0867(.A(new_n1182), .Y(n304));
  nor_4  g0868(.A(new_n651), .B(new_n646), .Y(new_n1184));
  nor_4  g0869(.A(new_n1184), .B(new_n341_1), .Y(new_n1185));
  nor_4  g0870(.A(new_n1185), .B(new_n649), .Y(new_n1186_1));
  nor_4  g0871(.A(new_n1186_1), .B(new_n335), .Y(new_n1187_1));
  xnor_3 g0872(.A(new_n1187_1), .B(new_n647), .Y(n364));
  nor_4  g0873(.A(new_n446), .B(new_n445), .Y(new_n1189));
  xor_3  g0874(.A(new_n1189), .B(new_n618), .Y(n370));
  not_3  g0875(.A(new_n1092), .Y(new_n1191_1));
  not_3  g0876(.A(n138), .Y(new_n1192));
  nor_4  g0877(.A(n1500), .B(new_n319), .Y(new_n1193_1));
  nor_4  g0878(.A(new_n1193_1), .B(new_n318_1), .Y(new_n1194));
  nor_4  g0879(.A(new_n1194), .B(new_n1192), .Y(new_n1195_1));
  nor_4  g0880(.A(new_n1084), .B(new_n1079), .Y(new_n1196));
  nor_4  g0881(.A(new_n1196), .B(new_n1077), .Y(new_n1197));
  not_3  g0882(.A(new_n1197), .Y(new_n1198));
  nor_4  g0883(.A(new_n1198), .B(new_n1089), .Y(new_n1199));
  not_3  g0884(.A(new_n1080), .Y(new_n1200));
  nor_4  g0885(.A(new_n1094), .B(new_n1085), .Y(new_n1201));
  not_3  g0886(.A(new_n1201), .Y(new_n1202));
  nor_4  g0887(.A(new_n1202), .B(new_n1200), .Y(new_n1203));
  nor_4  g0888(.A(new_n1203), .B(new_n1198), .Y(new_n1204));
  nor_4  g0889(.A(new_n1204), .B(new_n1199), .Y(new_n1205_1));
  not_3  g0890(.A(new_n1194), .Y(new_n1206));
  nor_4  g0891(.A(new_n1206), .B(n138), .Y(new_n1207));
  nor_4  g0892(.A(new_n1207), .B(new_n1205_1), .Y(new_n1208));
  nor_4  g0893(.A(new_n1208), .B(new_n1195_1), .Y(new_n1209_1));
  not_3  g0894(.A(new_n1209_1), .Y(new_n1210));
  nor_4  g0895(.A(new_n1207), .B(new_n1195_1), .Y(new_n1211_1));
  nor_4  g0896(.A(new_n319), .B(n582), .Y(new_n1212));
  nor_4  g0897(.A(new_n1212), .B(new_n318_1), .Y(new_n1213));
  not_3  g0898(.A(new_n1213), .Y(new_n1214));
  nor_4  g0899(.A(new_n1214), .B(n1470), .Y(new_n1215));
  not_3  g0900(.A(n1470), .Y(new_n1216));
  nor_4  g0901(.A(new_n1213), .B(new_n1216), .Y(new_n1217));
  nor_4  g0902(.A(new_n1217), .B(new_n1215), .Y(new_n1218));
  xor_3  g0903(.A(new_n1218), .B(new_n1211_1), .Y(new_n1219));
  nor_4  g0904(.A(new_n1094), .B(new_n1090), .Y(new_n1220));
  xor_3  g0905(.A(new_n1220), .B(new_n1219), .Y(new_n1221));
  xor_3  g0906(.A(new_n1221), .B(new_n1210), .Y(new_n1222));
  not_3  g0907(.A(new_n1205_1), .Y(new_n1223));
  not_3  g0908(.A(new_n1211_1), .Y(new_n1224));
  not_3  g0909(.A(new_n1218), .Y(new_n1225_1));
  nor_4  g0910(.A(new_n1225_1), .B(new_n1224), .Y(new_n1226));
  not_3  g0911(.A(new_n1226), .Y(new_n1227_1));
  nor_4  g0912(.A(new_n1227_1), .B(new_n1223), .Y(new_n1228));
  not_3  g0913(.A(new_n1207), .Y(new_n1229));
  nor_4  g0914(.A(new_n1217), .B(new_n1229), .Y(new_n1230));
  nor_4  g0915(.A(new_n1230), .B(new_n1215), .Y(new_n1231_1));
  not_3  g0916(.A(new_n1231_1), .Y(new_n1232));
  nor_4  g0917(.A(new_n1232), .B(new_n1228), .Y(new_n1233));
  nand_4 g0918(.A(n487), .B(n156), .Y(new_n1234_1));
  nand_4 g0919(.A(n200), .B(n156), .Y(new_n1235));
  not_3  g0920(.A(new_n1235), .Y(new_n1236));
  nor_4  g0921(.A(new_n1236), .B(n986), .Y(new_n1237));
  xor_3  g0922(.A(new_n1237), .B(new_n1234_1), .Y(new_n1238));
  and_4  g0923(.A(new_n1238), .B(new_n1233), .Y(new_n1239_1));
  not_3  g0924(.A(new_n1234_1), .Y(new_n1240));
  nor_4  g0925(.A(new_n1240), .B(n986), .Y(new_n1241));
  nor_4  g0926(.A(new_n1235), .B(new_n1058_1), .Y(new_n1242));
  and_4  g0927(.A(new_n1242), .B(n487), .Y(new_n1243));
  nor_4  g0928(.A(new_n1243), .B(new_n1241), .Y(new_n1244));
  not_3  g0929(.A(new_n1244), .Y(new_n1245));
  nor_4  g0930(.A(new_n1236), .B(new_n1240), .Y(new_n1246_1));
  nor_4  g0931(.A(new_n1246_1), .B(new_n1245), .Y(new_n1247));
  not_3  g0932(.A(new_n1247), .Y(new_n1248));
  nor_4  g0933(.A(new_n1248), .B(new_n1233), .Y(new_n1249));
  nor_4  g0934(.A(new_n1249), .B(new_n1239_1), .Y(new_n1250_1));
  xnor_3 g0935(.A(new_n1250_1), .B(new_n1222), .Y(new_n1251));
  xor_3  g0936(.A(new_n1201), .B(new_n1200), .Y(new_n1252));
  nor_4  g0937(.A(new_n1096), .B(new_n1089), .Y(new_n1253_1));
  not_3  g0938(.A(new_n1089), .Y(new_n1254));
  nor_4  g0939(.A(new_n1204), .B(new_n1254), .Y(new_n1255));
  nor_4  g0940(.A(new_n1255), .B(new_n1199), .Y(new_n1256));
  nor_4  g0941(.A(new_n1256), .B(new_n1253_1), .Y(new_n1257));
  not_3  g0942(.A(new_n1253_1), .Y(new_n1258));
  nor_4  g0943(.A(new_n1258), .B(new_n1197), .Y(new_n1259));
  nor_4  g0944(.A(new_n1259), .B(new_n1257), .Y(new_n1260));
  xor_3  g0945(.A(new_n1260), .B(new_n1252), .Y(new_n1261));
  xnor_3 g0946(.A(new_n1261), .B(new_n1251), .Y(new_n1262));
  nor_4  g0947(.A(new_n1262), .B(new_n1191_1), .Y(new_n1263_1));
  not_3  g0948(.A(new_n1233), .Y(new_n1264));
  not_3  g0949(.A(new_n1203), .Y(new_n1265));
  nor_4  g0950(.A(new_n1258), .B(new_n1265), .Y(new_n1266));
  not_3  g0951(.A(new_n1266), .Y(new_n1267));
  nor_4  g0952(.A(new_n1267), .B(new_n1224), .Y(new_n1268));
  not_3  g0953(.A(new_n1268), .Y(new_n1269));
  nor_4  g0954(.A(new_n1269), .B(new_n1225_1), .Y(new_n1270));
  nor_4  g0955(.A(new_n1270), .B(new_n1264), .Y(new_n1271));
  and_4  g0956(.A(new_n1271), .B(new_n1238), .Y(new_n1272));
  nor_4  g0957(.A(new_n1271), .B(new_n1248), .Y(new_n1273));
  or_4   g0958(.A(new_n1273), .B(new_n1272), .Y(new_n1274));
  and_4  g0959(.A(new_n1256), .B(new_n1252), .Y(new_n1275));
  not_3  g0960(.A(new_n1256), .Y(new_n1276));
  nand_4 g0961(.A(new_n1267), .B(new_n1252), .Y(new_n1277));
  and_4  g0962(.A(new_n1277), .B(new_n1276), .Y(new_n1278_1));
  nor_4  g0963(.A(new_n1278_1), .B(new_n1275), .Y(new_n1279));
  xor_3  g0964(.A(new_n1279), .B(new_n1219), .Y(new_n1280));
  nor_4  g0965(.A(new_n1210), .B(new_n1099), .Y(new_n1281_1));
  nor_4  g0966(.A(new_n1268), .B(new_n1098), .Y(new_n1282));
  and_4  g0967(.A(new_n1282), .B(new_n1210), .Y(new_n1283_1));
  nor_4  g0968(.A(new_n1283_1), .B(new_n1281_1), .Y(new_n1284));
  xnor_3 g0969(.A(new_n1284), .B(new_n1280), .Y(new_n1285_1));
  xnor_3 g0970(.A(new_n1285_1), .B(new_n1274), .Y(new_n1286_1));
  nor_4  g0971(.A(new_n1286_1), .B(new_n1092), .Y(new_n1287));
  nor_4  g0972(.A(new_n1287), .B(new_n1263_1), .Y(n378));
  xor_3  g0973(.A(new_n1185), .B(new_n649), .Y(n396));
  nor_4  g0974(.A(new_n1258), .B(new_n1092), .Y(new_n1290));
  nand_4 g0975(.A(new_n1290), .B(new_n1203), .Y(new_n1291));
  nand_4 g0976(.A(new_n1291), .B(new_n1223), .Y(new_n1292_1));
  nand_4 g0977(.A(new_n1292_1), .B(new_n1226), .Y(new_n1293));
  nand_4 g0978(.A(new_n1293), .B(new_n1231_1), .Y(new_n1294));
  nand_4 g0979(.A(new_n1294), .B(new_n1238), .Y(new_n1295));
  nand_4 g0980(.A(new_n1253_1), .B(new_n1191_1), .Y(new_n1296_1));
  nor_4  g0981(.A(new_n1296_1), .B(new_n1265), .Y(new_n1297));
  nor_4  g0982(.A(new_n1297), .B(new_n1205_1), .Y(new_n1298));
  nor_4  g0983(.A(new_n1298), .B(new_n1227_1), .Y(new_n1299_1));
  nor_4  g0984(.A(new_n1299_1), .B(new_n1232), .Y(new_n1300));
  nand_4 g0985(.A(new_n1300), .B(new_n1248), .Y(new_n1301_1));
  nand_4 g0986(.A(new_n1301_1), .B(new_n1295), .Y(n428));
  nor_4  g0987(.A(new_n1242), .B(new_n1237), .Y(new_n1303));
  xnor_3 g0988(.A(new_n1303), .B(new_n1294), .Y(n453));
  or_4   g0989(.A(new_n429), .B(new_n411), .Y(new_n1305_1));
  nor_4  g0990(.A(new_n1305_1), .B(new_n620), .Y(new_n1306_1));
  not_3  g0991(.A(new_n432), .Y(new_n1307));
  not_3  g0992(.A(new_n439), .Y(new_n1308));
  nor_4  g0993(.A(new_n1308), .B(new_n414), .Y(new_n1309));
  and_4  g0994(.A(new_n1309), .B(new_n622), .Y(new_n1310));
  nor_4  g0995(.A(new_n1310), .B(new_n1307), .Y(new_n1311));
  nor_4  g0996(.A(new_n1311), .B(new_n1306_1), .Y(new_n1312));
  xor_3  g0997(.A(new_n1312), .B(new_n624), .Y(n517));
  nor_4  g0998(.A(new_n631), .B(new_n363), .Y(new_n1314));
  nor_4  g0999(.A(new_n1314), .B(new_n637), .Y(new_n1315));
  nor_4  g1000(.A(new_n1315), .B(new_n378_1), .Y(new_n1316));
  xor_3  g1001(.A(new_n1316), .B(new_n369), .Y(n534));
  nor_4  g1002(.A(new_n1294), .B(new_n1244), .Y(new_n1318));
  or_4   g1003(.A(new_n1246_1), .B(n986), .Y(new_n1319));
  not_3  g1004(.A(new_n1319), .Y(new_n1320_1));
  nor_4  g1005(.A(new_n1320_1), .B(new_n1318), .Y(n553));
  xor_3  g1006(.A(new_n588), .B(new_n584), .Y(n597));
  nor_4  g1007(.A(new_n481), .B(new_n460_1), .Y(new_n1323));
  nor_4  g1008(.A(new_n1323), .B(new_n610), .Y(new_n1324));
  xor_3  g1009(.A(new_n1324), .B(new_n614), .Y(new_n1325));
  xor_3  g1010(.A(new_n482), .B(new_n474), .Y(new_n1326));
  xor_3  g1011(.A(new_n1189), .B(new_n1172_1), .Y(new_n1327));
  xor_3  g1012(.A(new_n1327), .B(new_n1326), .Y(new_n1328));
  xor_3  g1013(.A(new_n617), .B(new_n464), .Y(new_n1329));
  not_3  g1014(.A(new_n1329), .Y(new_n1330));
  xnor_3 g1015(.A(new_n1330), .B(new_n1328), .Y(new_n1331));
  xnor_3 g1016(.A(new_n1331), .B(new_n1325), .Y(new_n1332));
  nand_4 g1017(.A(new_n1332), .B(new_n1173), .Y(new_n1333));
  nor_4  g1018(.A(new_n1329), .B(new_n488), .Y(new_n1334));
  xor_3  g1019(.A(new_n614), .B(new_n463), .Y(new_n1335));
  nor_4  g1020(.A(new_n1335), .B(new_n486), .Y(new_n1336));
  not_3  g1021(.A(new_n463), .Y(new_n1337_1));
  nor_4  g1022(.A(new_n481), .B(new_n1337_1), .Y(new_n1338));
  nor_4  g1023(.A(new_n1338), .B(new_n480), .Y(new_n1339));
  xnor_3 g1024(.A(new_n1339), .B(new_n1328), .Y(new_n1340));
  xnor_3 g1025(.A(new_n1340), .B(new_n1336), .Y(new_n1341));
  xnor_3 g1026(.A(new_n1341), .B(new_n1334), .Y(new_n1342));
  nand_4 g1027(.A(new_n1342), .B(new_n606), .Y(new_n1343));
  nand_4 g1028(.A(new_n1343), .B(new_n1333), .Y(new_n1344));
  xor_3  g1029(.A(new_n625_1), .B(new_n624), .Y(new_n1345_1));
  not_3  g1030(.A(new_n428_1), .Y(new_n1346_1));
  not_3  g1031(.A(new_n438), .Y(new_n1347));
  nor_4  g1032(.A(new_n1347), .B(new_n420_1), .Y(new_n1348));
  nor_4  g1033(.A(new_n1348), .B(new_n1346_1), .Y(new_n1349));
  not_3  g1034(.A(new_n426), .Y(new_n1350_1));
  not_3  g1035(.A(new_n427), .Y(new_n1351));
  nor_4  g1036(.A(new_n1351), .B(new_n1350_1), .Y(new_n1352));
  nor_4  g1037(.A(new_n1352), .B(new_n1349), .Y(new_n1353));
  xor_3  g1038(.A(new_n1353), .B(new_n1345_1), .Y(new_n1354));
  xor_3  g1039(.A(new_n1354), .B(new_n1311), .Y(new_n1355));
  nand_4 g1040(.A(new_n1355), .B(new_n620), .Y(new_n1356));
  not_3  g1041(.A(new_n620), .Y(new_n1357));
  xor_3  g1042(.A(new_n623), .B(new_n438), .Y(new_n1358));
  not_3  g1043(.A(new_n431), .Y(new_n1359_1));
  nand_4 g1044(.A(new_n1305_1), .B(new_n1359_1), .Y(new_n1360));
  xnor_3 g1045(.A(new_n1360), .B(new_n1345_1), .Y(new_n1361_1));
  xor_3  g1046(.A(new_n1361_1), .B(new_n1358), .Y(new_n1362));
  nand_4 g1047(.A(new_n1362), .B(new_n1357), .Y(new_n1363));
  nand_4 g1048(.A(new_n1363), .B(new_n1356), .Y(new_n1364));
  xnor_3 g1049(.A(new_n1364), .B(new_n1344), .Y(n625));
  nand_4 g1050(.A(n1536), .B(n1438), .Y(new_n1366));
  nand_4 g1051(.A(n997), .B(n315), .Y(new_n1367));
  nor_4  g1052(.A(new_n1367), .B(new_n1366), .Y(new_n1368_1));
  not_3  g1053(.A(new_n1368_1), .Y(n669));
  xor_3  g1054(.A(new_n1175_1), .B(new_n483), .Y(n693));
  xor_3  g1055(.A(new_n1151), .B(new_n603), .Y(n714));
  or_4   g1056(.A(n1361), .B(n1225), .Y(n719));
  not_3  g1057(.A(new_n579), .Y(new_n1373));
  not_3  g1058(.A(new_n582_1), .Y(new_n1374));
  nor_4  g1059(.A(new_n589_1), .B(new_n571), .Y(new_n1375_1));
  nor_4  g1060(.A(new_n1375_1), .B(new_n1374), .Y(new_n1376));
  nor_4  g1061(.A(new_n1376), .B(new_n580), .Y(new_n1377));
  xor_3  g1062(.A(new_n1377), .B(new_n1373), .Y(n794));
  nand_4 g1063(.A(new_n1316), .B(new_n369), .Y(new_n1379));
  nand_4 g1064(.A(new_n1379), .B(new_n635), .Y(new_n1380));
  xor_3  g1065(.A(new_n1380), .B(new_n393), .Y(n894));
  nor_4  g1066(.A(new_n1253_1), .B(new_n1191_1), .Y(new_n1382));
  nor_4  g1067(.A(new_n1382), .B(new_n1290), .Y(n916));
  nand_4 g1068(.A(n1411), .B(n1239), .Y(new_n1384));
  nand_4 g1069(.A(new_n1384), .B(new_n570), .Y(new_n1385));
  xor_3  g1070(.A(new_n1385), .B(new_n981), .Y(new_n1386_1));
  xor_3  g1071(.A(new_n971), .B(new_n938), .Y(new_n1387_1));
  xor_3  g1072(.A(new_n1387_1), .B(new_n1386_1), .Y(new_n1388));
  xor_3  g1073(.A(new_n1388), .B(new_n963), .Y(new_n1389_1));
  xor_3  g1074(.A(new_n955), .B(new_n946), .Y(new_n1390));
  not_3  g1075(.A(n299), .Y(new_n1391_1));
  nor_4  g1076(.A(n1239), .B(new_n1391_1), .Y(new_n1392));
  nand_4 g1077(.A(n1239), .B(n1044), .Y(new_n1393_1));
  not_3  g1078(.A(new_n1393_1), .Y(new_n1394));
  nor_4  g1079(.A(new_n1394), .B(new_n1392), .Y(new_n1395));
  xor_3  g1080(.A(new_n1014), .B(new_n927), .Y(new_n1396));
  xor_3  g1081(.A(new_n1396), .B(new_n1395), .Y(new_n1397));
  xor_3  g1082(.A(new_n1397), .B(new_n1390), .Y(new_n1398));
  nor_4  g1083(.A(new_n1398), .B(new_n1389_1), .Y(new_n1399));
  and_4  g1084(.A(new_n1398), .B(new_n1389_1), .Y(new_n1400));
  nor_4  g1085(.A(new_n1400), .B(new_n1399), .Y(new_n1401_1));
  nor_4  g1086(.A(new_n318_1), .B(new_n319), .Y(new_n1402));
  not_3  g1087(.A(n56), .Y(new_n1403));
  xor_3  g1088(.A(n1389), .B(n246), .Y(new_n1404));
  xor_3  g1089(.A(new_n1404), .B(new_n1403), .Y(new_n1405));
  and_4  g1090(.A(new_n1405), .B(new_n1402), .Y(new_n1406));
  and_4  g1091(.A(new_n690_1), .B(new_n682), .Y(new_n1407));
  not_3  g1092(.A(new_n681), .Y(new_n1408));
  nor_4  g1093(.A(new_n706), .B(new_n1408), .Y(new_n1409));
  nor_4  g1094(.A(new_n1409), .B(new_n1407), .Y(new_n1410));
  not_3  g1095(.A(new_n671_1), .Y(new_n1411_1));
  nor_4  g1096(.A(new_n1411_1), .B(new_n1051_1), .Y(new_n1412));
  and_4  g1097(.A(new_n672), .B(new_n663_1), .Y(new_n1413));
  nor_4  g1098(.A(new_n1413), .B(new_n1412), .Y(new_n1414));
  xor_3  g1099(.A(new_n1414), .B(new_n1410), .Y(new_n1415_1));
  xor_3  g1100(.A(new_n1415_1), .B(new_n1406), .Y(new_n1416));
  nor_4  g1101(.A(new_n1416), .B(new_n1401_1), .Y(new_n1417));
  not_3  g1102(.A(new_n712), .Y(new_n1418_1));
  nor_4  g1103(.A(new_n744), .B(new_n1418_1), .Y(new_n1419));
  not_3  g1104(.A(new_n742_1), .Y(new_n1420_1));
  nor_4  g1105(.A(new_n1420_1), .B(new_n740), .Y(new_n1421_1));
  nor_4  g1106(.A(new_n1421_1), .B(new_n1419), .Y(new_n1422));
  not_3  g1107(.A(n1103), .Y(new_n1423));
  nor_4  g1108(.A(n1239), .B(new_n1423), .Y(new_n1424));
  nand_4 g1109(.A(n1239), .B(n1023), .Y(new_n1425));
  not_3  g1110(.A(new_n1425), .Y(new_n1426));
  nor_4  g1111(.A(new_n1426), .B(new_n1424), .Y(new_n1427_1));
  xor_3  g1112(.A(new_n1427_1), .B(new_n808), .Y(new_n1428_1));
  xor_3  g1113(.A(new_n1428_1), .B(new_n1422), .Y(new_n1429));
  xor_3  g1114(.A(new_n797), .B(new_n785), .Y(new_n1430));
  not_3  g1115(.A(new_n728), .Y(new_n1431));
  nor_4  g1116(.A(new_n1431), .B(new_n752), .Y(new_n1432));
  not_3  g1117(.A(new_n720), .Y(new_n1433));
  nor_4  g1118(.A(new_n754), .B(new_n1433), .Y(new_n1434));
  nor_4  g1119(.A(new_n1434), .B(new_n1432), .Y(new_n1435_1));
  xor_3  g1120(.A(new_n775_1), .B(new_n760), .Y(new_n1436));
  xor_3  g1121(.A(new_n1436), .B(new_n1435_1), .Y(new_n1437));
  xor_3  g1122(.A(new_n1437), .B(new_n1430), .Y(new_n1438_1));
  xnor_3 g1123(.A(new_n1438_1), .B(new_n1429), .Y(new_n1439));
  xor_3  g1124(.A(new_n854), .B(new_n834), .Y(new_n1440));
  not_3  g1125(.A(n1121), .Y(new_n1441));
  nor_4  g1126(.A(n1239), .B(new_n1441), .Y(new_n1442));
  nand_4 g1127(.A(n1239), .B(n560), .Y(new_n1443_1));
  not_3  g1128(.A(new_n1443_1), .Y(new_n1444));
  nor_4  g1129(.A(new_n1444), .B(new_n1442), .Y(new_n1445));
  xor_3  g1130(.A(new_n1445), .B(new_n909), .Y(new_n1446_1));
  xor_3  g1131(.A(new_n1446_1), .B(new_n1440), .Y(new_n1447));
  xor_3  g1132(.A(new_n903), .B(new_n864), .Y(new_n1448_1));
  xor_3  g1133(.A(new_n1448_1), .B(new_n1447), .Y(new_n1449));
  not_3  g1134(.A(new_n893), .Y(new_n1450));
  xor_3  g1135(.A(new_n1450), .B(new_n844), .Y(new_n1451));
  xor_3  g1136(.A(new_n1451), .B(new_n875), .Y(new_n1452));
  xor_3  g1137(.A(new_n1452), .B(new_n823_1), .Y(new_n1453));
  xnor_3 g1138(.A(new_n1453), .B(new_n1449), .Y(new_n1454));
  nor_4  g1139(.A(new_n1454), .B(new_n1439), .Y(new_n1455));
  nand_4 g1140(.A(new_n1455), .B(new_n1417), .Y(n1375));
  xor_3  g1141(.A(new_n479), .B(new_n459), .Y(new_n1457));
  xor_3  g1142(.A(new_n444), .B(new_n413), .Y(new_n1458));
  xor_3  g1143(.A(new_n1458), .B(new_n1457), .Y(new_n1459));
  xor_3  g1144(.A(new_n1459), .B(new_n419), .Y(new_n1460));
  xor_3  g1145(.A(new_n452), .B(new_n401), .Y(new_n1461));
  nand_4 g1146(.A(n1239), .B(n314), .Y(new_n1462));
  not_3  g1147(.A(new_n1462), .Y(new_n1463_1));
  nor_4  g1148(.A(new_n1463_1), .B(new_n1442), .Y(new_n1464));
  xor_3  g1149(.A(new_n470), .B(new_n437), .Y(new_n1465));
  xor_3  g1150(.A(new_n1465), .B(new_n1464), .Y(new_n1466));
  xor_3  g1151(.A(new_n1466), .B(new_n1461), .Y(new_n1467));
  xnor_3 g1152(.A(new_n1467), .B(new_n1460), .Y(new_n1468));
  xor_3  g1153(.A(new_n503), .B(new_n495), .Y(new_n1469));
  xor_3  g1154(.A(new_n523), .B(new_n513), .Y(new_n1470_1));
  xor_3  g1155(.A(new_n1470_1), .B(new_n1469), .Y(new_n1471));
  nand_4 g1156(.A(n1281), .B(n1239), .Y(new_n1472));
  not_3  g1157(.A(new_n1472), .Y(new_n1473));
  nor_4  g1158(.A(new_n1473), .B(new_n1392), .Y(new_n1474_1));
  nand_4 g1159(.A(n1239), .B(n961), .Y(new_n1475));
  not_3  g1160(.A(new_n1475), .Y(new_n1476_1));
  nor_4  g1161(.A(new_n1476_1), .B(new_n990_1), .Y(new_n1477));
  xor_3  g1162(.A(new_n1477), .B(new_n1474_1), .Y(new_n1478));
  xor_3  g1163(.A(new_n556), .B(new_n549), .Y(new_n1479));
  xor_3  g1164(.A(new_n1479), .B(new_n1478), .Y(new_n1480));
  xor_3  g1165(.A(new_n568), .B(new_n535), .Y(new_n1481));
  xor_3  g1166(.A(new_n1481), .B(new_n1480), .Y(new_n1482));
  xnor_3 g1167(.A(new_n1482), .B(new_n1471), .Y(new_n1483));
  nor_4  g1168(.A(new_n1483), .B(new_n1468), .Y(new_n1484));
  not_3  g1169(.A(new_n320), .Y(new_n1485));
  nor_4  g1170(.A(new_n328), .B(new_n1485), .Y(new_n1486));
  not_3  g1171(.A(new_n326), .Y(new_n1487));
  nor_4  g1172(.A(new_n1487), .B(new_n323), .Y(new_n1488));
  nor_4  g1173(.A(new_n1488), .B(new_n1486), .Y(new_n1489));
  xor_3  g1174(.A(new_n634), .B(new_n350), .Y(new_n1490));
  xor_3  g1175(.A(new_n1490), .B(new_n1489), .Y(new_n1491));
  xor_3  g1176(.A(new_n390), .B(new_n376_1), .Y(new_n1492));
  not_3  g1177(.A(new_n332), .Y(new_n1493));
  nor_4  g1178(.A(new_n340), .B(new_n1493), .Y(new_n1494));
  not_3  g1179(.A(new_n338), .Y(new_n1495));
  nor_4  g1180(.A(new_n1495), .B(new_n334), .Y(new_n1496));
  nor_4  g1181(.A(new_n1496), .B(new_n1494), .Y(new_n1497));
  nand_4 g1182(.A(n1239), .B(n117), .Y(new_n1498));
  not_3  g1183(.A(new_n1498), .Y(new_n1499));
  nor_4  g1184(.A(new_n1499), .B(new_n1424), .Y(new_n1500_1));
  xor_3  g1185(.A(new_n1500_1), .B(new_n357), .Y(new_n1501));
  xor_3  g1186(.A(new_n1501), .B(new_n1497), .Y(new_n1502_1));
  xor_3  g1187(.A(new_n1502_1), .B(new_n1492), .Y(new_n1503));
  xnor_3 g1188(.A(new_n1503), .B(new_n1491), .Y(new_n1504));
  not_3  g1189(.A(n430), .Y(new_n1505));
  xor_3  g1190(.A(n1626), .B(n775), .Y(new_n1506_1));
  xor_3  g1191(.A(new_n1506_1), .B(new_n1505), .Y(new_n1507));
  and_4  g1192(.A(new_n1507), .B(new_n1402), .Y(new_n1508));
  not_3  g1193(.A(new_n1212), .Y(new_n1509));
  nor_4  g1194(.A(new_n1509), .B(new_n1206), .Y(new_n1510));
  not_3  g1195(.A(new_n1193_1), .Y(new_n1511));
  nor_4  g1196(.A(new_n1214), .B(new_n1511), .Y(new_n1512));
  nor_4  g1197(.A(new_n1512), .B(new_n1510), .Y(new_n1513));
  and_4  g1198(.A(new_n1083), .B(new_n1074), .Y(new_n1514));
  not_3  g1199(.A(new_n1082), .Y(new_n1515));
  nor_4  g1200(.A(new_n1515), .B(new_n1076), .Y(new_n1516_1));
  nor_4  g1201(.A(new_n1516_1), .B(new_n1514), .Y(new_n1517));
  xor_3  g1202(.A(new_n1517), .B(new_n1513), .Y(new_n1518));
  xor_3  g1203(.A(new_n1518), .B(new_n1508), .Y(new_n1519));
  nor_4  g1204(.A(new_n1519), .B(new_n1504), .Y(new_n1520_1));
  nand_4 g1205(.A(new_n1520_1), .B(new_n1484), .Y(n1288));
  nor_4  g1206(.A(n1288), .B(n1375), .Y(new_n1522));
  not_3  g1207(.A(n1346), .Y(new_n1523_1));
  nor_4  g1208(.A(new_n1523_1), .B(n1239), .Y(new_n1524));
  nor_4  g1209(.A(new_n319), .B(n831), .Y(new_n1525));
  nor_4  g1210(.A(new_n1525), .B(new_n1524), .Y(new_n1526));
  xor_3  g1211(.A(new_n695_1), .B(new_n686), .Y(new_n1527_1));
  xor_3  g1212(.A(new_n1527_1), .B(new_n1526), .Y(new_n1528));
  not_3  g1213(.A(new_n1066), .Y(new_n1529));
  nor_4  g1214(.A(new_n1529), .B(new_n1059), .Y(new_n1530));
  nor_4  g1215(.A(new_n1530), .B(n1239), .Y(new_n1531));
  xor_3  g1216(.A(n487), .B(n200), .Y(new_n1532));
  nor_4  g1217(.A(new_n1532), .B(new_n319), .Y(new_n1533));
  or_4   g1218(.A(new_n1533), .B(new_n1531), .Y(new_n1534_1));
  not_3  g1219(.A(new_n1534_1), .Y(new_n1535));
  xor_3  g1220(.A(new_n676_1), .B(new_n668), .Y(new_n1536_1));
  xor_3  g1221(.A(new_n1536_1), .B(new_n704), .Y(new_n1537));
  xnor_3 g1222(.A(new_n1537), .B(new_n1535), .Y(new_n1538));
  xnor_3 g1223(.A(new_n1538), .B(new_n1528), .Y(new_n1539));
  nand_4 g1224(.A(n1239), .B(n21), .Y(new_n1540));
  not_3  g1225(.A(new_n1540), .Y(new_n1541));
  nor_4  g1226(.A(n1644), .B(n1239), .Y(new_n1542));
  nor_4  g1227(.A(new_n1542), .B(new_n1541), .Y(new_n1543));
  xor_3  g1228(.A(new_n1543), .B(new_n779_1), .Y(new_n1544));
  xor_3  g1229(.A(new_n765), .B(new_n734_1), .Y(new_n1545));
  xor_3  g1230(.A(new_n1545), .B(new_n1544), .Y(new_n1546));
  xor_3  g1231(.A(new_n792), .B(new_n717), .Y(new_n1547_1));
  xor_3  g1232(.A(new_n812), .B(new_n801), .Y(new_n1548_1));
  xor_3  g1233(.A(new_n1548_1), .B(new_n1547_1), .Y(new_n1549));
  xor_3  g1234(.A(new_n748), .B(new_n726_1), .Y(new_n1550));
  xor_3  g1235(.A(new_n1550), .B(new_n1549), .Y(new_n1551));
  xnor_3 g1236(.A(new_n1551), .B(new_n1546), .Y(new_n1552));
  nor_4  g1237(.A(new_n1552), .B(new_n1539), .Y(new_n1553));
  nand_4 g1238(.A(n1239), .B(n947), .Y(new_n1554));
  not_3  g1239(.A(new_n1554), .Y(new_n1555));
  nor_4  g1240(.A(n1750), .B(n1239), .Y(new_n1556));
  nor_4  g1241(.A(new_n1556), .B(new_n1555), .Y(new_n1557));
  xor_3  g1242(.A(new_n1557), .B(new_n879_1), .Y(new_n1558));
  xor_3  g1243(.A(new_n897), .B(new_n869), .Y(new_n1559));
  xor_3  g1244(.A(new_n858), .B(new_n838), .Y(new_n1560));
  xor_3  g1245(.A(new_n1560), .B(new_n1559), .Y(new_n1561));
  xor_3  g1246(.A(new_n907), .B(new_n910), .Y(new_n1562));
  xor_3  g1247(.A(new_n848), .B(new_n827), .Y(new_n1563));
  xor_3  g1248(.A(new_n1563), .B(new_n1562), .Y(new_n1564));
  xnor_3 g1249(.A(new_n1564), .B(new_n1561), .Y(new_n1565));
  xnor_3 g1250(.A(new_n1565), .B(new_n1558), .Y(new_n1566_1));
  nand_4 g1251(.A(n1239), .B(n1205), .Y(new_n1567));
  not_3  g1252(.A(new_n1567), .Y(new_n1568));
  nor_4  g1253(.A(new_n1568), .B(new_n988), .Y(new_n1569_1));
  xor_3  g1254(.A(new_n1569_1), .B(new_n1018), .Y(new_n1570));
  not_3  g1255(.A(new_n942), .Y(new_n1571));
  nand_4 g1256(.A(n1239), .B(n1138), .Y(new_n1572));
  not_3  g1257(.A(new_n1572), .Y(new_n1573));
  nor_4  g1258(.A(n1239), .B(n155), .Y(new_n1574));
  nor_4  g1259(.A(new_n1574), .B(new_n1573), .Y(new_n1575));
  xor_3  g1260(.A(new_n1575), .B(new_n1571), .Y(new_n1576_1));
  xor_3  g1261(.A(new_n1576_1), .B(new_n1570), .Y(new_n1577));
  xor_3  g1262(.A(new_n985), .B(new_n977), .Y(new_n1578));
  xor_3  g1263(.A(new_n967), .B(new_n959), .Y(new_n1579));
  xor_3  g1264(.A(new_n1579), .B(new_n1578), .Y(new_n1580));
  xor_3  g1265(.A(new_n950), .B(new_n932), .Y(new_n1581));
  xor_3  g1266(.A(new_n1581), .B(new_n1580), .Y(new_n1582));
  xnor_3 g1267(.A(new_n1582), .B(new_n1577), .Y(new_n1583));
  nor_4  g1268(.A(new_n1583), .B(new_n1566_1), .Y(new_n1584));
  nand_4 g1269(.A(new_n1584), .B(new_n1553), .Y(n1322));
  nand_4 g1270(.A(n1095), .B(n743), .Y(new_n1586_1));
  nand_4 g1271(.A(n581), .B(n478), .Y(new_n1587));
  nor_4  g1272(.A(new_n1587), .B(new_n1586_1), .Y(new_n1588_1));
  nand_4 g1273(.A(n1286), .B(n1054), .Y(new_n1589));
  nand_4 g1274(.A(n1040), .B(n593), .Y(new_n1590));
  nor_4  g1275(.A(new_n1590), .B(new_n1589), .Y(new_n1591));
  nand_4 g1276(.A(new_n1591), .B(new_n1368_1), .Y(new_n1592_1));
  nor_4  g1277(.A(new_n1592_1), .B(n126), .Y(new_n1593));
  nand_4 g1278(.A(new_n1593), .B(new_n1588_1), .Y(new_n1594_1));
  nor_4  g1279(.A(new_n1594_1), .B(n1322), .Y(new_n1595));
  nand_4 g1280(.A(new_n1595), .B(new_n1522), .Y(n918));
  xor_3  g1281(.A(new_n1177_1), .B(new_n474), .Y(n952));
  not_3  g1282(.A(new_n1195_1), .Y(new_n1598));
  nand_4 g1283(.A(new_n1291), .B(new_n1208), .Y(new_n1599));
  nand_4 g1284(.A(new_n1599), .B(new_n1598), .Y(new_n1600));
  xnor_3 g1285(.A(new_n1600), .B(new_n1218), .Y(n990));
  xor_3  g1286(.A(new_n1155), .B(new_n528), .Y(n1006));
  not_3  g1287(.A(n380), .Y(new_n1603));
  nor_4  g1288(.A(n1361), .B(new_n1603), .Y(new_n1604));
  nand_4 g1289(.A(new_n1604), .B(n701), .Y(n1050));
  not_3  g1290(.A(new_n378_1), .Y(new_n1606));
  nand_4 g1291(.A(new_n1315), .B(new_n1606), .Y(new_n1607));
  nor_4  g1292(.A(new_n1314), .B(new_n358), .Y(new_n1608));
  nor_4  g1293(.A(new_n1608), .B(new_n380_1), .Y(new_n1609_1));
  not_3  g1294(.A(new_n1609_1), .Y(new_n1610));
  nand_4 g1295(.A(new_n1610), .B(new_n1607), .Y(n1051));
  nor_4  g1296(.A(new_n1377), .B(new_n1373), .Y(new_n1612));
  nor_4  g1297(.A(new_n1612), .B(new_n557), .Y(new_n1613_1));
  xor_3  g1298(.A(new_n1613_1), .B(new_n1105), .Y(n1058));
  nand_4 g1299(.A(new_n621), .B(new_n1350_1), .Y(new_n1615));
  xor_3  g1300(.A(new_n1615), .B(new_n622), .Y(n1060));
  xor_3  g1301(.A(new_n606), .B(new_n464), .Y(n1063));
  not_3  g1302(.A(new_n631), .Y(new_n1618));
  xor_3  g1303(.A(new_n380_1), .B(new_n370_1), .Y(new_n1619));
  xor_3  g1304(.A(new_n1071_1), .B(new_n393), .Y(new_n1620));
  xor_3  g1305(.A(new_n1620), .B(new_n1619), .Y(new_n1621));
  not_3  g1306(.A(new_n1621), .Y(new_n1622));
  not_3  g1307(.A(new_n358), .Y(new_n1623));
  nor_4  g1308(.A(new_n378_1), .B(new_n1623), .Y(new_n1624));
  nor_4  g1309(.A(new_n1624), .B(new_n636), .Y(new_n1625));
  xor_3  g1310(.A(new_n1625), .B(new_n641_1), .Y(new_n1626_1));
  xor_3  g1311(.A(new_n1626_1), .B(new_n1622), .Y(new_n1627_1));
  xor_3  g1312(.A(new_n643), .B(new_n363), .Y(new_n1628));
  xor_3  g1313(.A(new_n1628), .B(new_n1627_1), .Y(new_n1629));
  nor_4  g1314(.A(new_n1629), .B(new_n1618), .Y(new_n1630));
  xor_3  g1315(.A(new_n641_1), .B(new_n361), .Y(new_n1631));
  nor_4  g1316(.A(new_n1631), .B(new_n384), .Y(new_n1632_1));
  nand_4 g1317(.A(new_n1632_1), .B(new_n1628), .Y(new_n1633));
  not_3  g1318(.A(new_n1628), .Y(new_n1634));
  nor_4  g1319(.A(new_n1632_1), .B(new_n395), .Y(new_n1635));
  nand_4 g1320(.A(new_n1635), .B(new_n1634), .Y(new_n1636));
  nand_4 g1321(.A(new_n1636), .B(new_n1633), .Y(new_n1637));
  not_3  g1322(.A(new_n361), .Y(new_n1638));
  nor_4  g1323(.A(new_n379), .B(new_n1638), .Y(new_n1639_1));
  nor_4  g1324(.A(new_n1639_1), .B(new_n378_1), .Y(new_n1640));
  xor_3  g1325(.A(new_n1640), .B(new_n1622), .Y(new_n1641));
  xor_3  g1326(.A(new_n1641), .B(new_n1637), .Y(new_n1642));
  nor_4  g1327(.A(new_n1642), .B(new_n631), .Y(new_n1643));
  nor_4  g1328(.A(new_n1643), .B(new_n1630), .Y(new_n1644_1));
  not_3  g1329(.A(new_n335), .Y(new_n1645_1));
  nor_4  g1330(.A(new_n650), .B(new_n1645_1), .Y(new_n1646));
  not_3  g1331(.A(new_n344_1), .Y(new_n1647_1));
  nor_4  g1332(.A(new_n652), .B(new_n1647_1), .Y(new_n1648));
  not_3  g1333(.A(new_n1648), .Y(new_n1649));
  and_4  g1334(.A(new_n651), .B(new_n337_1), .Y(new_n1650));
  nor_4  g1335(.A(new_n1650), .B(new_n1649), .Y(new_n1651));
  nor_4  g1336(.A(new_n1651), .B(new_n1646), .Y(new_n1652));
  xor_3  g1337(.A(new_n647), .B(new_n325), .Y(new_n1653));
  xor_3  g1338(.A(new_n1653), .B(new_n342), .Y(new_n1654));
  not_3  g1339(.A(new_n1654), .Y(new_n1655));
  xor_3  g1340(.A(new_n1655), .B(new_n1652), .Y(new_n1656_1));
  xor_3  g1341(.A(new_n1656_1), .B(new_n347), .Y(new_n1657));
  nand_4 g1342(.A(new_n1657), .B(new_n646), .Y(new_n1658));
  not_3  g1343(.A(new_n329), .Y(new_n1659));
  nor_4  g1344(.A(new_n1649), .B(new_n1659), .Y(new_n1660));
  not_3  g1345(.A(new_n331), .Y(new_n1661));
  nor_4  g1346(.A(new_n1648), .B(new_n1661), .Y(new_n1662));
  nor_4  g1347(.A(new_n1662), .B(new_n1660), .Y(new_n1663));
  xor_3  g1348(.A(new_n1663), .B(new_n1655), .Y(new_n1664));
  xor_3  g1349(.A(new_n1664), .B(new_n648), .Y(new_n1665));
  nor_4  g1350(.A(new_n1665), .B(new_n646), .Y(new_n1666));
  not_3  g1351(.A(new_n1666), .Y(new_n1667));
  nand_4 g1352(.A(new_n1667), .B(new_n1658), .Y(new_n1668));
  xnor_3 g1353(.A(new_n1668), .B(new_n1644_1), .Y(n1065));
  xor_3  g1354(.A(new_n1165), .B(new_n601), .Y(n1195));
  nor_4  g1355(.A(new_n1290), .B(new_n1089), .Y(new_n1671));
  xnor_3 g1356(.A(new_n1671), .B(new_n1201), .Y(n1302));
  xnor_3 g1357(.A(new_n1292_1), .B(new_n1224), .Y(n1391));
  xor_3  g1358(.A(new_n1375_1), .B(new_n1374), .Y(n1420));
  nand_4 g1359(.A(new_n1155), .B(new_n528), .Y(new_n1675));
  and_4  g1360(.A(new_n1675), .B(new_n1160), .Y(new_n1676));
  or_4   g1361(.A(new_n1676), .B(new_n596), .Y(new_n1677));
  nor_4  g1362(.A(new_n1677), .B(new_n1162), .Y(n1427));
  xor_3  g1363(.A(new_n631), .B(new_n363), .Y(n1527));
  not_3  g1364(.A(new_n1591), .Y(n1594));
  not_3  g1365(.A(new_n593_1), .Y(new_n1681));
  xor_3  g1366(.A(new_n1106), .B(new_n1681), .Y(n1639));
  nor_4  g1367(.A(new_n1615), .B(new_n623), .Y(new_n1683));
  nor_4  g1368(.A(new_n1683), .B(new_n420_1), .Y(new_n1684));
  xor_3  g1369(.A(new_n1684), .B(new_n625_1), .Y(n1687));
  not_3  g1370(.A(new_n1588_1), .Y(n1752));
  buf_2  g1371(.A(n346), .Y(n23));
  buf_2  g1372(.A(n947), .Y(n27));
  buf_2  g1373(.A(n153), .Y(n85));
  buf_2  g1374(.A(n1592), .Y(n130));
  buf_2  g1375(.A(n823), .Y(n173));
  buf_2  g1376(.A(n420), .Y(n184));
  buf_2  g1377(.A(n831), .Y(n230));
  buf_2  g1378(.A(n408), .Y(n292));
  buf_2  g1379(.A(n318), .Y(n301));
  buf_2  g1380(.A(n626), .Y(n337));
  buf_2  g1381(.A(n1463), .Y(n352));
  nand_4 g1382(.A(n1387), .B(new_n657), .Y(n362));
  buf_2  g1383(.A(n399), .Y(n417));
  nor_4  g1384(.A(new_n1068), .B(new_n1065_1), .Y(n457));
  buf_2  g1385(.A(n21), .Y(n460));
  buf_2  g1386(.A(n1656), .Y(n497));
  buf_2  g1387(.A(n293), .Y(n498));
  buf_2  g1388(.A(n200), .Y(n501));
  buf_2  g1389(.A(n769), .Y(n509));
  buf_2  g1390(.A(n1187), .Y(n516));
  nor_4  g1391(.A(new_n1320_1), .B(new_n1318), .Y(n585));
  buf_2  g1392(.A(n1301), .Y(n595));
  buf_2  g1393(.A(n420), .Y(n638));
  buf_2  g1394(.A(n1345), .Y(n640));
  not_3  g1395(.A(n992), .Y(n726));
  buf_2  g1396(.A(n980), .Y(n773));
  buf_2  g1397(.A(n222), .Y(n782));
  buf_2  g1398(.A(n374), .Y(n821));
  buf_2  g1399(.A(n1205), .Y(n842));
  buf_2  g1400(.A(n1476), .Y(n1017));
  buf_2  g1401(.A(n1566), .Y(n1042));
  buf_2  g1402(.A(n487), .Y(n1177));
  nor_4  g1403(.A(new_n1320_1), .B(new_n1318), .Y(n1186));
  buf_2  g1404(.A(n1071), .Y(n1209));
  nor_4  g1405(.A(new_n1068), .B(new_n1065_1), .Y(n1211));
  buf_2  g1406(.A(n1470), .Y(n1231));
  buf_2  g1407(.A(n608), .Y(n1234));
  nand_4 g1408(.A(new_n1604), .B(n701), .Y(n1253));
  buf_2  g1409(.A(n1401), .Y(n1285));
  buf_2  g1410(.A(n1616), .Y(n1292));
  not_3  g1411(.A(n992), .Y(n1296));
  buf_2  g1412(.A(n1263), .Y(n1320));
  buf_2  g1413(.A(n1138), .Y(n1337));
  xnor_3 g1414(.A(new_n1303), .B(new_n1294), .Y(n1359));
  buf_2  g1415(.A(n420), .Y(n1368));
  buf_2  g1416(.A(n695), .Y(n1421));
  buf_2  g1417(.A(n920), .Y(n1534));
  buf_2  g1418(.A(n420), .Y(n1547));
  buf_2  g1419(.A(n567), .Y(n1548));
  nand_4 g1420(.A(new_n1301_1), .B(new_n1295), .Y(n1588));
  nor_4  g1421(.A(new_n1320_1), .B(new_n1318), .Y(n1632));
  buf_2  g1422(.A(n1446), .Y(n1645));
  buf_2  g1423(.A(n138), .Y(n1729));
  buf_2  g1424(.A(n45), .Y(n1738));
endmodule


