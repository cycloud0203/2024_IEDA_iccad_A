// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Fri Jun 14 22:43:13 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1,
    new_n993, new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067_1, new_n1068, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094_1, new_n1095, new_n1096,
    new_n1097_1, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136_1, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1199_1, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269_1, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333_1, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355, new_n1356,
    new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471_1, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1, new_n2432,
    new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498_1,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1, new_n2510,
    new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522_1,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558_1,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564_1,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1, new_n2582,
    new_n2583, new_n2584, new_n2585_1, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172_1, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214_1, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230_1,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272_1,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3282, new_n3283, new_n3284, new_n3285,
    new_n3286, new_n3287_1, new_n3288, new_n3289, new_n3290, new_n3291,
    new_n3292, new_n3293, new_n3294, new_n3295, new_n3296, new_n3297,
    new_n3298, new_n3299, new_n3300, new_n3301, new_n3302, new_n3303,
    new_n3304, new_n3305, new_n3306, new_n3307, new_n3308, new_n3309,
    new_n3310, new_n3311, new_n3312, new_n3313, new_n3314, new_n3315,
    new_n3316, new_n3317, new_n3318, new_n3319, new_n3320, new_n3321,
    new_n3322, new_n3323, new_n3324, new_n3325, new_n3326, new_n3327,
    new_n3328, new_n3329, new_n3330, new_n3331, new_n3332, new_n3333,
    new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339_1,
    new_n3340, new_n3341, new_n3342_1, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357,
    new_n3358, new_n3359, new_n3360, new_n3361, new_n3362, new_n3363,
    new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369,
    new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627_1,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719_1, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754_1, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849_1,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865_1, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986_1, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005_1, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086_1, new_n4087, new_n4088_1, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094_1, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141_1, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155_1, new_n4156,
    new_n4157, new_n4158, new_n4159_1, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187_1, new_n4188, new_n4189_1, new_n4190_1, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203_1, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226_1, new_n4227, new_n4228, new_n4229,
    new_n4230_1, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300_1, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312_1, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326_1, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333_1, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370_1, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378_1, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397_1,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436_1, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499_1,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516_1, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553_1,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4575, new_n4577, new_n4579, new_n4580, new_n4581,
    new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587,
    new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593,
    new_n4594, new_n4595, new_n4596, new_n4597, new_n4598, new_n4599,
    new_n4600, new_n4601, new_n4602, new_n4603, new_n4604, new_n4605,
    new_n4606, new_n4607, new_n4608, new_n4609, new_n4610, new_n4611,
    new_n4612, new_n4613, new_n4614, new_n4615, new_n4616, new_n4617,
    new_n4618, new_n4619, new_n4620, new_n4621, new_n4622, new_n4623,
    new_n4624, new_n4625, new_n4626, new_n4627, new_n4628, new_n4629,
    new_n4630, new_n4631, new_n4632, new_n4633, new_n4634_1, new_n4635,
    new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641,
    new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686_1, new_n4687, new_n4688, new_n4689_1,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733_1, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757_1, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805_1, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817_1, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826_1, new_n4827,
    new_n4828_1, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903_1, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921_1, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928_1, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1, new_n4971_1,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1, new_n5031,
    new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069_1, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094_1, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105_1, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132_1, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153_1, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191_1, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198_1, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212_1, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314_1, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1,
    new_n5320_1, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579_1, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641_1, new_n5642, new_n5643, new_n5644,
    new_n5645_1, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670_1, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693_1, new_n5694_1, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760_1, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767_1, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798_1, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814_1, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857_1, new_n5858, new_n5859, new_n5860_1,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934_1, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016_1, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038_1, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089_1,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126_1, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192_1, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254_1, new_n6255, new_n6256, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271, new_n6272, new_n6273_1, new_n6274, new_n6275,
    new_n6276, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281,
    new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294_1,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358_1, new_n6359_1, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429_1, new_n6430, new_n6431_1, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441_1, new_n6442, new_n6443, new_n6444,
    new_n6445_1, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504,
    new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559,
    new_n6560, new_n6561, new_n6564, new_n6565, new_n6566, new_n6567,
    new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573,
    new_n6574, new_n6575, new_n6576, new_n6577, new_n6578_1, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604_1, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611_1, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645_1,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687_1,
    new_n6688, new_n6689_1, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703_1, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742_1, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770_1, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776_1, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797_1, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806_1, new_n6807,
    new_n6808, new_n6809_1, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822_1, new_n6823, new_n6824, new_n6825,
    new_n6826_1, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860_1, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877_1, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986_1, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159_1, new_n7160_1, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193_1,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236_1, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265_1,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270_1, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294_1, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320_1, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331,
    new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354_1, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388_1, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436_1, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456_1, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500_1, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523_1,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546_1, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568_1, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646_1, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7712, new_n7714, new_n7715, new_n7718, new_n7720,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946_1, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965_1, new_n7966_1, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981_1, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997,
    new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003,
    new_n8004, new_n8005, new_n8006, new_n8007, new_n8008, new_n8009,
    new_n8010, new_n8011, new_n8012, new_n8013, new_n8014, new_n8015,
    new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021,
    new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027,
    new_n8028_1, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033,
    new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039,
    new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045,
    new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051,
    new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057,
    new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063,
    new_n8064, new_n8065_1, new_n8066, new_n8067, new_n8068, new_n8069,
    new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075,
    new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081,
    new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087,
    new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093,
    new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099,
    new_n8100_1, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105,
    new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129,
    new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135,
    new_n8136, new_n8137, new_n8138_1, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202_1, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236_1, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255,
    new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8261,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303_1, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336_1, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384_1, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398_1, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8427,
    new_n8428, new_n8429, new_n8430, new_n8431, new_n8432, new_n8433_1,
    new_n8434, new_n8435, new_n8436, new_n8438, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476_1, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550, new_n8551, new_n8552, new_n8554, new_n8555, new_n8557,
    new_n8558, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595_1, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665_1, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717_1, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759_1, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804,
    new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819_1, new_n8820, new_n8821, new_n8822,
    new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834,
    new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840,
    new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846,
    new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852,
    new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858,
    new_n8859, new_n8860, new_n8861, new_n8862, new_n8863, new_n8864,
    new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870,
    new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876,
    new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882,
    new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888,
    new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894,
    new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900,
    new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906,
    new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912,
    new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918,
    new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924,
    new_n8925, new_n8926, new_n8927, new_n8928, new_n8929, new_n8930,
    new_n8931, new_n8932, new_n8933, new_n8934, new_n8935, new_n8936,
    new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942,
    new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948,
    new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954,
    new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080_1,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111_1, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137_1, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189_1, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195_1, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241_1, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260,
    new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272,
    new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278,
    new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284,
    new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290,
    new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296,
    new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302,
    new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308,
    new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314,
    new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320,
    new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326,
    new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332,
    new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9338,
    new_n9339, new_n9340, new_n9341, new_n9342, new_n9343, new_n9346,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387_1, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400_1, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457_1, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571_1, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578_1, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583_1, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637_1, new_n9638, new_n9639, new_n9640_1, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706_1, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725_1,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756_1, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820_1, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920_1, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938_1, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956_1, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022_1, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066,
    new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072,
    new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078,
    new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090,
    new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102,
    new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108,
    new_n10109, new_n10110, new_n10111, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150,
    new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156,
    new_n10157, new_n10158, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174_1, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202,
    new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208,
    new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214,
    new_n10215, new_n10216, new_n10217_1, new_n10218, new_n10219,
    new_n10220, new_n10221, new_n10222, new_n10223_1, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278_1, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285,
    new_n10286, new_n10287, new_n10288, new_n10289, new_n10290, new_n10291,
    new_n10292, new_n10293, new_n10294, new_n10295, new_n10296, new_n10297,
    new_n10298, new_n10299, new_n10300, new_n10301, new_n10302, new_n10303,
    new_n10304, new_n10305, new_n10306, new_n10307, new_n10308, new_n10309,
    new_n10310, new_n10311, new_n10312, new_n10313, new_n10314, new_n10315,
    new_n10316, new_n10317, new_n10318, new_n10319, new_n10320, new_n10321,
    new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327_1, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361,
    new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367,
    new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385,
    new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391_1, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439_1, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451_1, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476_1,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510_1, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545_1, new_n10546,
    new_n10547_1, new_n10548, new_n10549, new_n10550, new_n10551,
    new_n10552, new_n10553, new_n10554, new_n10555, new_n10556, new_n10557,
    new_n10558, new_n10559, new_n10560, new_n10562, new_n10566, new_n10567,
    new_n10570, new_n10571, new_n10572, new_n10573, new_n10574, new_n10575,
    new_n10576, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588, new_n10589_1, new_n10590, new_n10591, new_n10592,
    new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611, new_n10612, new_n10613, new_n10614, new_n10615, new_n10616,
    new_n10617, new_n10618, new_n10619, new_n10620, new_n10621, new_n10622,
    new_n10623, new_n10624, new_n10625, new_n10626, new_n10627, new_n10628,
    new_n10629, new_n10630, new_n10631, new_n10632, new_n10633, new_n10634,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644_1, new_n10645,
    new_n10646, new_n10647, new_n10648, new_n10649, new_n10650, new_n10651,
    new_n10652, new_n10653, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678_1, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685_1,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695_1, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789_1, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839,
    new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845,
    new_n10846, new_n10847, new_n10848_1, new_n10849, new_n10850,
    new_n10851_1, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898_1, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913_1,
    new_n10914, new_n10915, new_n10916, new_n10917, new_n10918, new_n10919,
    new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925,
    new_n10926, new_n10927, new_n10928_1, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949_1, new_n10950, new_n10951, new_n10952, new_n10953,
    new_n10954, new_n10955, new_n10956, new_n10957, new_n10958, new_n10959,
    new_n10960, new_n10961, new_n10962, new_n10963, new_n10964,
    new_n10965_1, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975,
    new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981,
    new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987,
    new_n10988, new_n10989, new_n10990_1, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023_1, new_n11024, new_n11025, new_n11026, new_n11027,
    new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033,
    new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039,
    new_n11040, new_n11041, new_n11042, new_n11043, new_n11044, new_n11045,
    new_n11046, new_n11047, new_n11048, new_n11049, new_n11050, new_n11051,
    new_n11052, new_n11053, new_n11054, new_n11055, new_n11056, new_n11057,
    new_n11058, new_n11059, new_n11060, new_n11061, new_n11062, new_n11063,
    new_n11064, new_n11065, new_n11066, new_n11067, new_n11068, new_n11069,
    new_n11070, new_n11071, new_n11072, new_n11073, new_n11074, new_n11075,
    new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094, new_n11096, new_n11098, new_n11100, new_n11101, new_n11102,
    new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114,
    new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120,
    new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153_1, new_n11154, new_n11155,
    new_n11156, new_n11157, new_n11158, new_n11159, new_n11160, new_n11161,
    new_n11162, new_n11163, new_n11164, new_n11165, new_n11166, new_n11167,
    new_n11168, new_n11169, new_n11170, new_n11171, new_n11172, new_n11173,
    new_n11174, new_n11175, new_n11176, new_n11177, new_n11178, new_n11179,
    new_n11180, new_n11181, new_n11182, new_n11183, new_n11184, new_n11185,
    new_n11186, new_n11187, new_n11188, new_n11189, new_n11190, new_n11191,
    new_n11192, new_n11193, new_n11194, new_n11195, new_n11196, new_n11197,
    new_n11198, new_n11199, new_n11200, new_n11201, new_n11202, new_n11203,
    new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209,
    new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215,
    new_n11216_1, new_n11217, new_n11218, new_n11219, new_n11220,
    new_n11221, new_n11222_1, new_n11223, new_n11224, new_n11225,
    new_n11226, new_n11227, new_n11228, new_n11229, new_n11230, new_n11231,
    new_n11232, new_n11233, new_n11234, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245, new_n11246, new_n11247, new_n11248, new_n11249,
    new_n11250, new_n11251, new_n11252, new_n11253, new_n11254, new_n11256,
    new_n11257_1, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296_1,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311_1, new_n11312, new_n11313,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325,
    new_n11326_1, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407_1,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419,
    new_n11420, new_n11421, new_n11422, new_n11423_1, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478_1, new_n11479, new_n11480, new_n11481, new_n11482,
    new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488,
    new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494,
    new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536_1, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607, new_n11608, new_n11609, new_n11610, new_n11611, new_n11612,
    new_n11613, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618,
    new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624,
    new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662_1, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667, new_n11668, new_n11669, new_n11670, new_n11671,
    new_n11672, new_n11673, new_n11674, new_n11675, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707_1, new_n11708, new_n11709, new_n11710, new_n11711,
    new_n11712, new_n11713, new_n11714, new_n11715, new_n11716, new_n11717,
    new_n11718, new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724, new_n11725, new_n11726, new_n11727, new_n11728_1,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755_1, new_n11756, new_n11757_1,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780_1,
    new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786,
    new_n11787, new_n11788, new_n11789, new_n11790, new_n11791_1,
    new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821_1, new_n11822, new_n11823, new_n11824, new_n11825,
    new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831,
    new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837,
    new_n11838, new_n11839, new_n11840, new_n11841, new_n11842, new_n11843,
    new_n11844, new_n11845, new_n11846, new_n11847, new_n11848, new_n11849,
    new_n11850, new_n11851, new_n11852, new_n11853, new_n11854, new_n11855,
    new_n11856, new_n11857, new_n11858, new_n11859, new_n11860, new_n11861,
    new_n11862, new_n11863, new_n11864, new_n11865, new_n11866, new_n11867,
    new_n11868, new_n11869, new_n11870, new_n11871, new_n11872, new_n11873,
    new_n11874, new_n11875, new_n11876_1, new_n11877_1, new_n11878,
    new_n11879, new_n11880, new_n11881, new_n11882, new_n11883, new_n11884,
    new_n11885, new_n11886, new_n11887, new_n11888, new_n11889, new_n11890,
    new_n11891, new_n11892_1, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917_1, new_n11918,
    new_n11919_1, new_n11920, new_n11921, new_n11922_1, new_n11923,
    new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965,
    new_n11966, new_n11967_1, new_n11968, new_n11969, new_n11970,
    new_n11971, new_n11972, new_n11973, new_n11974, new_n11975, new_n11976,
    new_n11977, new_n11978, new_n11979, new_n11980, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11998, new_n11999_1,
    new_n12000_1, new_n12001, new_n12002, new_n12003, new_n12004,
    new_n12005_1, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011, new_n12012, new_n12013, new_n12014_1,
    new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020_1, new_n12021, new_n12022, new_n12023, new_n12024,
    new_n12025_1, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044_1, new_n12045, new_n12046,
    new_n12047, new_n12048, new_n12049, new_n12050, new_n12051, new_n12052,
    new_n12053, new_n12054, new_n12055, new_n12056, new_n12057, new_n12058,
    new_n12059, new_n12060, new_n12061, new_n12062, new_n12063, new_n12064,
    new_n12065, new_n12066, new_n12067, new_n12068, new_n12069_1,
    new_n12070, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075,
    new_n12076_1, new_n12077, new_n12078, new_n12079, new_n12080,
    new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086,
    new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092,
    new_n12093, new_n12094, new_n12095, new_n12096, new_n12097, new_n12098,
    new_n12099, new_n12100, new_n12101, new_n12102, new_n12103, new_n12104,
    new_n12105, new_n12106, new_n12107, new_n12108, new_n12109, new_n12110,
    new_n12111_1, new_n12112, new_n12113, new_n12114, new_n12115,
    new_n12116, new_n12117, new_n12118, new_n12119, new_n12120, new_n12121,
    new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127,
    new_n12128, new_n12129, new_n12130, new_n12131, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145_1, new_n12146, new_n12147, new_n12148, new_n12149,
    new_n12150, new_n12151, new_n12152, new_n12153, new_n12154, new_n12155,
    new_n12156, new_n12157, new_n12158, new_n12159, new_n12160, new_n12161,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12177, new_n12178,
    new_n12181, new_n12184, new_n12186, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221_1, new_n12222, new_n12223, new_n12224, new_n12225,
    new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247_1, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299_1, new_n12300, new_n12301,
    new_n12302, new_n12303, new_n12304, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315, new_n12316, new_n12317, new_n12318, new_n12319,
    new_n12320, new_n12321, new_n12322, new_n12323, new_n12324, new_n12325,
    new_n12326, new_n12327, new_n12328, new_n12329, new_n12330, new_n12331,
    new_n12332, new_n12333, new_n12334, new_n12335, new_n12336, new_n12337,
    new_n12338, new_n12339, new_n12340, new_n12341, new_n12342, new_n12343,
    new_n12344, new_n12345, new_n12346, new_n12347, new_n12348, new_n12349,
    new_n12350, new_n12351, new_n12352, new_n12353, new_n12354, new_n12355,
    new_n12356, new_n12357, new_n12358, new_n12359, new_n12360, new_n12361,
    new_n12362, new_n12363, new_n12364, new_n12365, new_n12366, new_n12367,
    new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373,
    new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380, new_n12381, new_n12382, new_n12383, new_n12384, new_n12385,
    new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391_1, new_n12392, new_n12393, new_n12394, new_n12395,
    new_n12396, new_n12397, new_n12398, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408, new_n12409, new_n12410, new_n12411, new_n12412, new_n12413,
    new_n12414, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419,
    new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425,
    new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444_1, new_n12445, new_n12446, new_n12447, new_n12448,
    new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454,
    new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460,
    new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489_1,
    new_n12490, new_n12491, new_n12492, new_n12493, new_n12494, new_n12495,
    new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501,
    new_n12502, new_n12503, new_n12504, new_n12505, new_n12506, new_n12507,
    new_n12508, new_n12509, new_n12510, new_n12511_1, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538,
    new_n12539, new_n12540, new_n12541, new_n12542, new_n12543, new_n12544,
    new_n12545, new_n12546, new_n12547, new_n12548, new_n12549, new_n12550,
    new_n12551, new_n12552, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561, new_n12562,
    new_n12563, new_n12564, new_n12565, new_n12566, new_n12567, new_n12568,
    new_n12569, new_n12570, new_n12571, new_n12572, new_n12573, new_n12574,
    new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580,
    new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587, new_n12588, new_n12589, new_n12590, new_n12591_1,
    new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597,
    new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603,
    new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615,
    new_n12616, new_n12617, new_n12618, new_n12619, new_n12620, new_n12621,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626, new_n12627,
    new_n12628, new_n12629, new_n12630, new_n12631, new_n12632, new_n12633,
    new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639,
    new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648_1, new_n12649, new_n12650,
    new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656,
    new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662,
    new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12699, new_n12700, new_n12701, new_n12702, new_n12703,
    new_n12704_1, new_n12705_1, new_n12706_1, new_n12707, new_n12708,
    new_n12709_1, new_n12710, new_n12711, new_n12712, new_n12713,
    new_n12714, new_n12715, new_n12716, new_n12717, new_n12718, new_n12719,
    new_n12720_1, new_n12721, new_n12722, new_n12723, new_n12724,
    new_n12725, new_n12726, new_n12727, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12741, new_n12745, new_n12747,
    new_n12749, new_n12751, new_n12753_1, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777_1, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807_1,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826_1, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925_1,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947_1, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13129, new_n13131, new_n13134,
    new_n13136, new_n13138, new_n13140, new_n13142, new_n13144, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263, new_n13264, new_n13265, new_n13266,
    new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272,
    new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284,
    new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290,
    new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296,
    new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302,
    new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308,
    new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320,
    new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326,
    new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332,
    new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13347, new_n13348, new_n13350, new_n13351, new_n13352,
    new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358,
    new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364,
    new_n13365, new_n13366, new_n13367, new_n13368, new_n13369, new_n13370,
    new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13376,
    new_n13377, new_n13378, new_n13379, new_n13380, new_n13381, new_n13382,
    new_n13383, new_n13384, new_n13385, new_n13386, new_n13387, new_n13388,
    new_n13389, new_n13390, new_n13391, new_n13392, new_n13393, new_n13394,
    new_n13395, new_n13396, new_n13397, new_n13398, new_n13399, new_n13400,
    new_n13401, new_n13402, new_n13403, new_n13404, new_n13405, new_n13406,
    new_n13407, new_n13408, new_n13409, new_n13410, new_n13411, new_n13412,
    new_n13413, new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419, new_n13420, new_n13421, new_n13422, new_n13423, new_n13424,
    new_n13425, new_n13426, new_n13427, new_n13428, new_n13429, new_n13430,
    new_n13431, new_n13432, new_n13433, new_n13434, new_n13435, new_n13436,
    new_n13437, new_n13438, new_n13439, new_n13440, new_n13441, new_n13442,
    new_n13443, new_n13444, new_n13445, new_n13446, new_n13447, new_n13448,
    new_n13449, new_n13450, new_n13451, new_n13452, new_n13453, new_n13454,
    new_n13455, new_n13456, new_n13457, new_n13458, new_n13459, new_n13460,
    new_n13461, new_n13462, new_n13463, new_n13464, new_n13465, new_n13466,
    new_n13467, new_n13468, new_n13469, new_n13470, new_n13471, new_n13472,
    new_n13473, new_n13474, new_n13475, new_n13476, new_n13477, new_n13478,
    new_n13479, new_n13480, new_n13481, new_n13482, new_n13483, new_n13484,
    new_n13485, new_n13486, new_n13487, new_n13488, new_n13489, new_n13490,
    new_n13491, new_n13492, new_n13493, new_n13494, new_n13495, new_n13496,
    new_n13497, new_n13498, new_n13499, new_n13500, new_n13501, new_n13502,
    new_n13503, new_n13504, new_n13505, new_n13506, new_n13507, new_n13508,
    new_n13509, new_n13510, new_n13511, new_n13512, new_n13513, new_n13514,
    new_n13515, new_n13516, new_n13517, new_n13518, new_n13519, new_n13520,
    new_n13521, new_n13522, new_n13523, new_n13524, new_n13525, new_n13526,
    new_n13527, new_n13528, new_n13529, new_n13530, new_n13531, new_n13532,
    new_n13533, new_n13534, new_n13535, new_n13536, new_n13537, new_n13538,
    new_n13539, new_n13540, new_n13541, new_n13542, new_n13543, new_n13544,
    new_n13545, new_n13547, new_n13549, new_n13552, new_n13554, new_n13556,
    new_n13558, new_n13560, new_n13563, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591,
    new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597,
    new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603,
    new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609,
    new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615,
    new_n13616, new_n13617, new_n13618, new_n13619, new_n13620, new_n13621,
    new_n13622, new_n13623, new_n13624, new_n13625, new_n13626, new_n13627,
    new_n13628, new_n13629, new_n13630, new_n13631, new_n13632, new_n13633,
    new_n13634, new_n13635, new_n13636, new_n13637, new_n13638, new_n13639,
    new_n13640, new_n13641, new_n13642, new_n13643, new_n13644, new_n13645,
    new_n13646, new_n13647, new_n13648, new_n13649, new_n13650, new_n13651,
    new_n13652, new_n13653, new_n13654, new_n13655, new_n13656, new_n13657,
    new_n13658, new_n13659, new_n13660, new_n13661, new_n13662, new_n13663,
    new_n13664, new_n13665, new_n13666, new_n13667, new_n13668, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677, new_n13678, new_n13679, new_n13680, new_n13681,
    new_n13682, new_n13683, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708, new_n13709, new_n13710, new_n13711,
    new_n13712, new_n13713, new_n13714, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719, new_n13720, new_n13721, new_n13722, new_n13723,
    new_n13724, new_n13725, new_n13726, new_n13727, new_n13728, new_n13729,
    new_n13730, new_n13731, new_n13732, new_n13733, new_n13734, new_n13735,
    new_n13736, new_n13737, new_n13738, new_n13739, new_n13740, new_n13741,
    new_n13742, new_n13743, new_n13744, new_n13745, new_n13746, new_n13747,
    new_n13748, new_n13749, new_n13750, new_n13751, new_n13752, new_n13753,
    new_n13754, new_n13755, new_n13756, new_n13757, new_n13758, new_n13759,
    new_n13760, new_n13761, new_n13762, new_n13764, new_n13766, new_n13770,
    new_n13772, new_n13773, new_n13776, new_n13781, new_n13782, new_n13783,
    new_n13784, new_n13785, new_n13786, new_n13787, new_n13788, new_n13789,
    new_n13790, new_n13791, new_n13792, new_n13793, new_n13794, new_n13795,
    new_n13796, new_n13797, new_n13798, new_n13799, new_n13800, new_n13801,
    new_n13802, new_n13803, new_n13804, new_n13805, new_n13806, new_n13807,
    new_n13808, new_n13809, new_n13810, new_n13811, new_n13812, new_n13813,
    new_n13814, new_n13815, new_n13816, new_n13817, new_n13818, new_n13819,
    new_n13820, new_n13821, new_n13822, new_n13823, new_n13824, new_n13825,
    new_n13826, new_n13827, new_n13828, new_n13829, new_n13830, new_n13831,
    new_n13832, new_n13833, new_n13834, new_n13835, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843,
    new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850, new_n13851, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13981, new_n13984,
    new_n13988, new_n13990, new_n13994;
  nand_4 g00000(.A(n6687), .B(n6038), .Y(new_n377));
  not_3  g00001(.A(new_n377), .Y(new_n378));
  nand_4 g00002(.A(n8336), .B(n7354), .Y(new_n379));
  not_3  g00003(.A(new_n379), .Y(new_n380));
  nand_4 g00004(.A(n11222), .B(n8028), .Y(new_n381_1));
  nand_4 g00005(.A(n12069), .B(n1564), .Y(new_n382));
  not_3  g00006(.A(new_n382), .Y(new_n383));
  xor_3  g00007(.A(new_n383), .B(new_n381_1), .Y(new_n384));
  not_3  g00008(.A(new_n384), .Y(new_n385));
  xor_3  g00009(.A(new_n385), .B(new_n380), .Y(new_n386));
  xor_3  g00010(.A(new_n386), .B(new_n378), .Y(n112));
  nand_4 g00011(.A(n7436), .B(n1209), .Y(new_n388));
  nand_4 g00012(.A(n8276), .B(n7500), .Y(new_n389));
  nand_4 g00013(.A(n9241), .B(n7354), .Y(new_n390));
  xnor_3 g00014(.A(new_n390), .B(new_n389), .Y(new_n391));
  nor_4  g00015(.A(new_n391), .B(new_n388), .Y(new_n392));
  not_3  g00016(.A(new_n388), .Y(new_n393));
  not_3  g00017(.A(new_n391), .Y(new_n394));
  nor_4  g00018(.A(new_n394), .B(new_n393), .Y(new_n395));
  nor_4  g00019(.A(new_n395), .B(new_n392), .Y(new_n396));
  nand_4 g00020(.A(n8276), .B(n7354), .Y(new_n397_1));
  not_3  g00021(.A(new_n397_1), .Y(new_n398));
  nand_4 g00022(.A(n12299), .B(n1209), .Y(new_n399));
  not_3  g00023(.A(new_n399), .Y(new_n400));
  nor_4  g00024(.A(new_n400), .B(new_n398), .Y(new_n401));
  nand_4 g00025(.A(n7500), .B(n7436), .Y(new_n402));
  not_3  g00026(.A(new_n402), .Y(new_n403));
  xnor_3 g00027(.A(new_n399), .B(new_n397_1), .Y(new_n404));
  nor_4  g00028(.A(new_n404), .B(new_n403), .Y(new_n405_1));
  nor_4  g00029(.A(new_n405_1), .B(new_n401), .Y(new_n406));
  xnor_3 g00030(.A(new_n406), .B(new_n396), .Y(new_n407));
  nand_4 g00031(.A(n6776), .B(n4141), .Y(new_n408));
  nand_4 g00032(.A(n12299), .B(n5105), .Y(new_n409));
  xor_3  g00033(.A(new_n409), .B(new_n408), .Y(new_n410));
  xnor_3 g00034(.A(new_n410), .B(new_n407), .Y(new_n411));
  nand_4 g00035(.A(n6776), .B(n5105), .Y(new_n412));
  not_3  g00036(.A(new_n412), .Y(new_n413));
  nand_4 g00037(.A(n7436), .B(n7354), .Y(new_n414));
  not_3  g00038(.A(new_n414), .Y(new_n415));
  nand_4 g00039(.A(n6776), .B(n1209), .Y(new_n416));
  not_3  g00040(.A(new_n416), .Y(new_n417));
  nor_4  g00041(.A(new_n417), .B(new_n415), .Y(new_n418));
  nand_4 g00042(.A(n12299), .B(n7500), .Y(new_n419));
  not_3  g00043(.A(new_n419), .Y(new_n420));
  xnor_3 g00044(.A(new_n416), .B(new_n414), .Y(new_n421));
  nor_4  g00045(.A(new_n421), .B(new_n420), .Y(new_n422));
  nor_4  g00046(.A(new_n422), .B(new_n418), .Y(new_n423));
  nand_4 g00047(.A(new_n423), .B(new_n413), .Y(new_n424));
  xnor_3 g00048(.A(new_n423), .B(new_n413), .Y(new_n425));
  not_3  g00049(.A(new_n425), .Y(new_n426));
  xnor_3 g00050(.A(new_n404), .B(new_n402), .Y(new_n427));
  not_3  g00051(.A(new_n427), .Y(new_n428));
  nand_4 g00052(.A(new_n428), .B(new_n426), .Y(new_n429));
  nand_4 g00053(.A(new_n429), .B(new_n424), .Y(new_n430));
  xnor_3 g00054(.A(new_n430), .B(new_n411), .Y(new_n431));
  not_3  g00055(.A(new_n431), .Y(new_n432));
  nand_4 g00056(.A(n8759), .B(n4141), .Y(new_n433));
  not_3  g00057(.A(new_n433), .Y(new_n434));
  xnor_3 g00058(.A(new_n427), .B(new_n425), .Y(new_n435));
  not_3  g00059(.A(new_n435), .Y(new_n436));
  nand_4 g00060(.A(new_n436), .B(new_n434), .Y(new_n437));
  not_3  g00061(.A(new_n437), .Y(new_n438));
  nor_4  g00062(.A(new_n436), .B(new_n434), .Y(new_n439));
  nor_4  g00063(.A(new_n439), .B(new_n438), .Y(new_n440));
  nand_4 g00064(.A(n8759), .B(n5105), .Y(new_n441));
  not_3  g00065(.A(new_n441), .Y(new_n442));
  nand_4 g00066(.A(n12299), .B(n7354), .Y(new_n443));
  nand_4 g00067(.A(n8759), .B(n1209), .Y(new_n444));
  nand_4 g00068(.A(new_n444), .B(new_n443), .Y(new_n445));
  not_3  g00069(.A(new_n445), .Y(new_n446));
  nor_4  g00070(.A(new_n444), .B(new_n443), .Y(new_n447_1));
  nand_4 g00071(.A(n7500), .B(n6776), .Y(new_n448));
  not_3  g00072(.A(new_n448), .Y(new_n449));
  nor_4  g00073(.A(new_n449), .B(new_n447_1), .Y(new_n450));
  nor_4  g00074(.A(new_n450), .B(new_n446), .Y(new_n451));
  nand_4 g00075(.A(new_n451), .B(new_n442), .Y(new_n452));
  not_3  g00076(.A(new_n452), .Y(new_n453));
  xnor_3 g00077(.A(new_n451), .B(new_n442), .Y(new_n454));
  xnor_3 g00078(.A(new_n421), .B(new_n419), .Y(new_n455));
  nor_4  g00079(.A(new_n455), .B(new_n454), .Y(new_n456));
  nor_4  g00080(.A(new_n456), .B(new_n453), .Y(new_n457));
  not_3  g00081(.A(new_n457), .Y(new_n458));
  nand_4 g00082(.A(new_n458), .B(new_n440), .Y(new_n459));
  nand_4 g00083(.A(new_n459), .B(new_n437), .Y(new_n460));
  nand_4 g00084(.A(new_n460), .B(new_n432), .Y(new_n461));
  nand_4 g00085(.A(new_n406), .B(new_n396), .Y(new_n462));
  not_3  g00086(.A(new_n462), .Y(new_n463));
  nor_4  g00087(.A(new_n463), .B(new_n392), .Y(new_n464));
  not_3  g00088(.A(new_n464), .Y(new_n465));
  nand_4 g00089(.A(n6776), .B(n4928), .Y(new_n466));
  nand_4 g00090(.A(n12299), .B(n4141), .Y(new_n467));
  nand_4 g00091(.A(n8759), .B(n8236), .Y(new_n468));
  not_3  g00092(.A(new_n468), .Y(new_n469));
  xor_3  g00093(.A(new_n469), .B(new_n467), .Y(new_n470));
  xnor_3 g00094(.A(new_n470), .B(new_n466), .Y(new_n471));
  xnor_3 g00095(.A(new_n471), .B(new_n465), .Y(new_n472));
  nor_4  g00096(.A(new_n390), .B(new_n389), .Y(new_n473));
  not_3  g00097(.A(new_n473), .Y(new_n474));
  nand_4 g00098(.A(n7436), .B(n5105), .Y(new_n475));
  xor_3  g00099(.A(new_n475), .B(new_n474), .Y(new_n476));
  nand_4 g00100(.A(n9241), .B(n7500), .Y(new_n477));
  not_3  g00101(.A(new_n477), .Y(new_n478));
  nand_4 g00102(.A(n8276), .B(n1209), .Y(new_n479));
  nand_4 g00103(.A(n10510), .B(n7354), .Y(new_n480));
  xor_3  g00104(.A(new_n480), .B(new_n479), .Y(new_n481));
  xnor_3 g00105(.A(new_n481), .B(new_n478), .Y(new_n482));
  xnor_3 g00106(.A(new_n482), .B(new_n476), .Y(new_n483));
  xnor_3 g00107(.A(new_n483), .B(new_n472), .Y(new_n484));
  not_3  g00108(.A(new_n407), .Y(new_n485));
  nand_4 g00109(.A(new_n410), .B(new_n485), .Y(new_n486));
  nor_4  g00110(.A(new_n409), .B(new_n408), .Y(new_n487));
  not_3  g00111(.A(new_n487), .Y(new_n488));
  nand_4 g00112(.A(new_n430), .B(new_n411), .Y(new_n489));
  xnor_3 g00113(.A(new_n489), .B(new_n488), .Y(new_n490));
  nand_4 g00114(.A(new_n490), .B(new_n486), .Y(new_n491));
  xnor_3 g00115(.A(new_n491), .B(new_n484), .Y(new_n492));
  xnor_3 g00116(.A(new_n492), .B(new_n461), .Y(new_n493));
  nand_4 g00117(.A(n8759), .B(n4928), .Y(new_n494));
  not_3  g00118(.A(new_n494), .Y(new_n495));
  xnor_3 g00119(.A(new_n460), .B(new_n431), .Y(new_n496));
  nand_4 g00120(.A(new_n496), .B(new_n495), .Y(new_n497));
  xnor_3 g00121(.A(new_n455), .B(new_n454), .Y(new_n498));
  nand_4 g00122(.A(n8759), .B(n7354), .Y(new_n499));
  not_3  g00123(.A(new_n499), .Y(new_n500));
  nor_4  g00124(.A(new_n500), .B(new_n448), .Y(new_n501));
  nor_4  g00125(.A(new_n501), .B(new_n445), .Y(new_n502));
  nor_4  g00126(.A(new_n502), .B(new_n447_1), .Y(new_n503_1));
  nor_4  g00127(.A(new_n503_1), .B(new_n448), .Y(new_n504));
  not_3  g00128(.A(new_n504), .Y(new_n505));
  nor_4  g00129(.A(new_n505), .B(new_n498), .Y(new_n506));
  not_3  g00130(.A(new_n506), .Y(new_n507));
  xnor_3 g00131(.A(new_n458), .B(new_n440), .Y(new_n508));
  nor_4  g00132(.A(new_n508), .B(new_n507), .Y(new_n509));
  xnor_3 g00133(.A(new_n496), .B(new_n494), .Y(new_n510));
  nand_4 g00134(.A(new_n510), .B(new_n509), .Y(new_n511));
  nand_4 g00135(.A(new_n511), .B(new_n497), .Y(new_n512));
  xnor_3 g00136(.A(new_n512), .B(new_n493), .Y(new_n513));
  nand_4 g00137(.A(n12648), .B(n533), .Y(new_n514));
  nand_4 g00138(.A(n10545), .B(n1512), .Y(new_n515));
  nand_4 g00139(.A(n7690), .B(n1564), .Y(new_n516));
  xnor_3 g00140(.A(new_n516), .B(new_n515), .Y(new_n517));
  nor_4  g00141(.A(new_n517), .B(new_n514), .Y(new_n518));
  not_3  g00142(.A(new_n514), .Y(new_n519));
  not_3  g00143(.A(new_n517), .Y(new_n520));
  nor_4  g00144(.A(new_n520), .B(new_n519), .Y(new_n521_1));
  nor_4  g00145(.A(new_n521_1), .B(new_n518), .Y(new_n522));
  nand_4 g00146(.A(n10545), .B(n1564), .Y(new_n523));
  not_3  g00147(.A(new_n523), .Y(new_n524));
  nand_4 g00148(.A(n2530), .B(n533), .Y(new_n525));
  not_3  g00149(.A(new_n525), .Y(new_n526));
  nor_4  g00150(.A(new_n526), .B(new_n524), .Y(new_n527));
  nand_4 g00151(.A(n12648), .B(n1512), .Y(new_n528));
  not_3  g00152(.A(new_n528), .Y(new_n529));
  xnor_3 g00153(.A(new_n525), .B(new_n523), .Y(new_n530));
  nor_4  g00154(.A(new_n530), .B(new_n529), .Y(new_n531));
  nor_4  g00155(.A(new_n531), .B(new_n527), .Y(new_n532));
  xnor_3 g00156(.A(new_n532), .B(new_n522), .Y(new_n533_1));
  nand_4 g00157(.A(n8476), .B(n6806), .Y(new_n534));
  nand_4 g00158(.A(n2802), .B(n2530), .Y(new_n535));
  xor_3  g00159(.A(new_n535), .B(new_n534), .Y(new_n536));
  xnor_3 g00160(.A(new_n536), .B(new_n533_1), .Y(new_n537));
  nand_4 g00161(.A(n8476), .B(n2802), .Y(new_n538));
  not_3  g00162(.A(new_n538), .Y(new_n539));
  nand_4 g00163(.A(n12648), .B(n1564), .Y(new_n540));
  not_3  g00164(.A(new_n540), .Y(new_n541));
  nand_4 g00165(.A(n8476), .B(n533), .Y(new_n542));
  not_3  g00166(.A(new_n542), .Y(new_n543));
  nor_4  g00167(.A(new_n543), .B(new_n541), .Y(new_n544));
  nand_4 g00168(.A(n2530), .B(n1512), .Y(new_n545));
  not_3  g00169(.A(new_n545), .Y(new_n546));
  xnor_3 g00170(.A(new_n542), .B(new_n540), .Y(new_n547));
  nor_4  g00171(.A(new_n547), .B(new_n546), .Y(new_n548));
  nor_4  g00172(.A(new_n548), .B(new_n544), .Y(new_n549));
  nand_4 g00173(.A(new_n549), .B(new_n539), .Y(new_n550));
  not_3  g00174(.A(new_n550), .Y(new_n551));
  nor_4  g00175(.A(new_n549), .B(new_n539), .Y(new_n552));
  nor_4  g00176(.A(new_n552), .B(new_n551), .Y(new_n553));
  xnor_3 g00177(.A(new_n530), .B(new_n528), .Y(new_n554));
  not_3  g00178(.A(new_n554), .Y(new_n555));
  nand_4 g00179(.A(new_n555), .B(new_n553), .Y(new_n556));
  nand_4 g00180(.A(new_n556), .B(new_n550), .Y(new_n557));
  xnor_3 g00181(.A(new_n557), .B(new_n537), .Y(new_n558));
  nand_4 g00182(.A(n6806), .B(n5331), .Y(new_n559));
  not_3  g00183(.A(new_n559), .Y(new_n560));
  xnor_3 g00184(.A(new_n555), .B(new_n553), .Y(new_n561));
  not_3  g00185(.A(new_n561), .Y(new_n562));
  nand_4 g00186(.A(new_n562), .B(new_n560), .Y(new_n563));
  xnor_3 g00187(.A(new_n561), .B(new_n560), .Y(new_n564));
  nand_4 g00188(.A(n5331), .B(n2802), .Y(new_n565));
  not_3  g00189(.A(new_n565), .Y(new_n566));
  nand_4 g00190(.A(n2530), .B(n1564), .Y(new_n567));
  nand_4 g00191(.A(n5331), .B(n533), .Y(new_n568));
  nand_4 g00192(.A(new_n568), .B(new_n567), .Y(new_n569));
  not_3  g00193(.A(new_n569), .Y(new_n570));
  nor_4  g00194(.A(new_n568), .B(new_n567), .Y(new_n571));
  nand_4 g00195(.A(n8476), .B(n1512), .Y(new_n572));
  not_3  g00196(.A(new_n572), .Y(new_n573));
  nor_4  g00197(.A(new_n573), .B(new_n571), .Y(new_n574));
  nor_4  g00198(.A(new_n574), .B(new_n570), .Y(new_n575));
  nand_4 g00199(.A(new_n575), .B(new_n566), .Y(new_n576));
  not_3  g00200(.A(new_n576), .Y(new_n577));
  xnor_3 g00201(.A(new_n575), .B(new_n566), .Y(new_n578));
  xnor_3 g00202(.A(new_n547), .B(new_n545), .Y(new_n579));
  nor_4  g00203(.A(new_n579), .B(new_n578), .Y(new_n580));
  nor_4  g00204(.A(new_n580), .B(new_n577), .Y(new_n581));
  not_3  g00205(.A(new_n581), .Y(new_n582));
  nand_4 g00206(.A(new_n582), .B(new_n564), .Y(new_n583));
  nand_4 g00207(.A(new_n583), .B(new_n563), .Y(new_n584));
  not_3  g00208(.A(new_n584), .Y(new_n585));
  nor_4  g00209(.A(new_n585), .B(new_n558), .Y(new_n586));
  not_3  g00210(.A(new_n586), .Y(new_n587));
  nand_4 g00211(.A(new_n532), .B(new_n522), .Y(new_n588));
  not_3  g00212(.A(new_n588), .Y(new_n589));
  nor_4  g00213(.A(new_n589), .B(new_n518), .Y(new_n590));
  not_3  g00214(.A(new_n590), .Y(new_n591));
  nand_4 g00215(.A(n8476), .B(n5069), .Y(new_n592));
  nand_4 g00216(.A(n6806), .B(n2530), .Y(new_n593));
  nand_4 g00217(.A(n12044), .B(n5331), .Y(new_n594));
  not_3  g00218(.A(new_n594), .Y(new_n595));
  xor_3  g00219(.A(new_n595), .B(new_n593), .Y(new_n596));
  xnor_3 g00220(.A(new_n596), .B(new_n592), .Y(new_n597));
  xnor_3 g00221(.A(new_n597), .B(new_n591), .Y(new_n598));
  nor_4  g00222(.A(new_n516), .B(new_n515), .Y(new_n599));
  nand_4 g00223(.A(n12648), .B(n2802), .Y(new_n600));
  not_3  g00224(.A(new_n600), .Y(new_n601));
  xor_3  g00225(.A(new_n601), .B(new_n599), .Y(new_n602));
  not_3  g00226(.A(new_n602), .Y(new_n603));
  nand_4 g00227(.A(n7690), .B(n1512), .Y(new_n604));
  not_3  g00228(.A(new_n604), .Y(new_n605));
  nand_4 g00229(.A(n10545), .B(n533), .Y(new_n606));
  nand_4 g00230(.A(n3616), .B(n1564), .Y(new_n607));
  not_3  g00231(.A(new_n607), .Y(new_n608));
  xor_3  g00232(.A(new_n608), .B(new_n606), .Y(new_n609));
  xnor_3 g00233(.A(new_n609), .B(new_n605), .Y(new_n610));
  xnor_3 g00234(.A(new_n610), .B(new_n603), .Y(new_n611));
  xnor_3 g00235(.A(new_n611), .B(new_n598), .Y(new_n612));
  not_3  g00236(.A(new_n533_1), .Y(new_n613));
  nand_4 g00237(.A(new_n536), .B(new_n613), .Y(new_n614));
  nor_4  g00238(.A(new_n535), .B(new_n534), .Y(new_n615_1));
  nand_4 g00239(.A(new_n557), .B(new_n537), .Y(new_n616));
  not_3  g00240(.A(new_n616), .Y(new_n617));
  xnor_3 g00241(.A(new_n617), .B(new_n615_1), .Y(new_n618));
  nand_4 g00242(.A(new_n618), .B(new_n614), .Y(new_n619));
  xnor_3 g00243(.A(new_n619), .B(new_n612), .Y(new_n620));
  xnor_3 g00244(.A(new_n620), .B(new_n587), .Y(new_n621));
  nand_4 g00245(.A(n5331), .B(n5069), .Y(new_n622));
  xnor_3 g00246(.A(new_n585), .B(new_n558), .Y(new_n623));
  nand_4 g00247(.A(new_n623), .B(new_n622), .Y(new_n624));
  xnor_3 g00248(.A(new_n579), .B(new_n578), .Y(new_n625));
  nand_4 g00249(.A(n5331), .B(n1564), .Y(new_n626));
  not_3  g00250(.A(new_n626), .Y(new_n627));
  nor_4  g00251(.A(new_n627), .B(new_n572), .Y(new_n628));
  not_3  g00252(.A(new_n628), .Y(new_n629));
  xnor_3 g00253(.A(new_n568), .B(new_n567), .Y(new_n630));
  nand_4 g00254(.A(new_n630), .B(new_n629), .Y(new_n631));
  nor_4  g00255(.A(new_n631), .B(new_n572), .Y(new_n632));
  not_3  g00256(.A(new_n632), .Y(new_n633));
  nor_4  g00257(.A(new_n633), .B(new_n625), .Y(new_n634));
  not_3  g00258(.A(new_n634), .Y(new_n635));
  xnor_3 g00259(.A(new_n582), .B(new_n564), .Y(new_n636));
  nor_4  g00260(.A(new_n636), .B(new_n635), .Y(new_n637));
  not_3  g00261(.A(new_n637), .Y(new_n638));
  xnor_3 g00262(.A(new_n623), .B(new_n622), .Y(new_n639));
  not_3  g00263(.A(new_n639), .Y(new_n640));
  nand_4 g00264(.A(new_n640), .B(new_n638), .Y(new_n641));
  nand_4 g00265(.A(new_n641), .B(new_n624), .Y(new_n642));
  xnor_3 g00266(.A(new_n642), .B(new_n621), .Y(new_n643));
  nand_4 g00267(.A(n2393), .B(n1980), .Y(new_n644));
  nand_4 g00268(.A(n8028), .B(n3986), .Y(new_n645));
  nand_4 g00269(.A(n10848), .B(n5860), .Y(new_n646));
  xnor_3 g00270(.A(new_n646), .B(new_n645), .Y(new_n647));
  nor_4  g00271(.A(new_n647), .B(new_n644), .Y(new_n648));
  not_3  g00272(.A(new_n644), .Y(new_n649));
  not_3  g00273(.A(new_n647), .Y(new_n650));
  nor_4  g00274(.A(new_n650), .B(new_n649), .Y(new_n651));
  nor_4  g00275(.A(new_n651), .B(new_n648), .Y(new_n652));
  nand_4 g00276(.A(n8028), .B(n5860), .Y(new_n653));
  not_3  g00277(.A(new_n653), .Y(new_n654));
  nand_4 g00278(.A(n11892), .B(n1980), .Y(new_n655));
  not_3  g00279(.A(new_n655), .Y(new_n656));
  nor_4  g00280(.A(new_n656), .B(new_n654), .Y(new_n657));
  nor_4  g00281(.A(new_n655), .B(new_n653), .Y(new_n658_1));
  nand_4 g00282(.A(n10848), .B(n2393), .Y(new_n659));
  not_3  g00283(.A(new_n659), .Y(new_n660));
  nor_4  g00284(.A(new_n660), .B(new_n658_1), .Y(new_n661));
  nor_4  g00285(.A(new_n661), .B(new_n657), .Y(new_n662));
  xnor_3 g00286(.A(new_n662), .B(new_n652), .Y(new_n663));
  nand_4 g00287(.A(n12704), .B(n7388), .Y(new_n664));
  nand_4 g00288(.A(n11892), .B(n7294), .Y(new_n665));
  not_3  g00289(.A(new_n665), .Y(new_n666));
  xor_3  g00290(.A(new_n666), .B(new_n664), .Y(new_n667));
  xnor_3 g00291(.A(new_n667), .B(new_n663), .Y(new_n668));
  nand_4 g00292(.A(n7388), .B(n7294), .Y(new_n669));
  not_3  g00293(.A(new_n669), .Y(new_n670));
  nand_4 g00294(.A(n7388), .B(n1980), .Y(new_n671_1));
  not_3  g00295(.A(new_n671_1), .Y(new_n672));
  nand_4 g00296(.A(n8028), .B(n2393), .Y(new_n673));
  not_3  g00297(.A(new_n673), .Y(new_n674));
  nor_4  g00298(.A(new_n674), .B(new_n672), .Y(new_n675));
  nor_4  g00299(.A(new_n673), .B(new_n671_1), .Y(new_n676));
  nand_4 g00300(.A(n11892), .B(n10848), .Y(new_n677));
  not_3  g00301(.A(new_n677), .Y(new_n678));
  nor_4  g00302(.A(new_n678), .B(new_n676), .Y(new_n679));
  nor_4  g00303(.A(new_n679), .B(new_n675), .Y(new_n680));
  and_4  g00304(.A(new_n680), .B(new_n670), .Y(new_n681));
  xnor_3 g00305(.A(new_n680), .B(new_n670), .Y(new_n682));
  nor_4  g00306(.A(new_n658_1), .B(new_n657), .Y(new_n683));
  xnor_3 g00307(.A(new_n683), .B(new_n660), .Y(new_n684));
  nor_4  g00308(.A(new_n684), .B(new_n682), .Y(new_n685));
  nor_4  g00309(.A(new_n685), .B(new_n681), .Y(new_n686));
  xnor_3 g00310(.A(new_n686), .B(new_n668), .Y(new_n687));
  nand_4 g00311(.A(n12704), .B(n7965), .Y(new_n688));
  xnor_3 g00312(.A(new_n684), .B(new_n682), .Y(new_n689));
  nor_4  g00313(.A(new_n689), .B(new_n688), .Y(new_n690));
  not_3  g00314(.A(new_n690), .Y(new_n691));
  not_3  g00315(.A(new_n688), .Y(new_n692));
  not_3  g00316(.A(new_n689), .Y(new_n693));
  nor_4  g00317(.A(new_n693), .B(new_n692), .Y(new_n694));
  nor_4  g00318(.A(new_n694), .B(new_n690), .Y(new_n695));
  nand_4 g00319(.A(n7965), .B(n7294), .Y(new_n696));
  not_3  g00320(.A(new_n696), .Y(new_n697));
  nand_4 g00321(.A(n11892), .B(n8028), .Y(new_n698));
  not_3  g00322(.A(new_n698), .Y(new_n699));
  nand_4 g00323(.A(n7965), .B(n1980), .Y(new_n700));
  not_3  g00324(.A(new_n700), .Y(new_n701));
  nor_4  g00325(.A(new_n701), .B(new_n699), .Y(new_n702));
  nor_4  g00326(.A(new_n700), .B(new_n698), .Y(new_n703));
  nand_4 g00327(.A(n10848), .B(n7388), .Y(new_n704));
  not_3  g00328(.A(new_n704), .Y(new_n705));
  nor_4  g00329(.A(new_n705), .B(new_n703), .Y(new_n706));
  nor_4  g00330(.A(new_n706), .B(new_n702), .Y(new_n707));
  nand_4 g00331(.A(new_n707), .B(new_n697), .Y(new_n708));
  xnor_3 g00332(.A(new_n707), .B(new_n697), .Y(new_n709));
  not_3  g00333(.A(new_n709), .Y(new_n710));
  xnor_3 g00334(.A(new_n673), .B(new_n671_1), .Y(new_n711));
  xnor_3 g00335(.A(new_n711), .B(new_n677), .Y(new_n712));
  not_3  g00336(.A(new_n712), .Y(new_n713));
  nand_4 g00337(.A(new_n713), .B(new_n710), .Y(new_n714));
  nand_4 g00338(.A(new_n714), .B(new_n708), .Y(new_n715));
  nand_4 g00339(.A(new_n715), .B(new_n695), .Y(new_n716));
  nand_4 g00340(.A(new_n716), .B(new_n691), .Y(new_n717));
  not_3  g00341(.A(new_n717), .Y(new_n718));
  nor_4  g00342(.A(new_n718), .B(new_n687), .Y(new_n719));
  not_3  g00343(.A(new_n648), .Y(new_n720));
  nand_4 g00344(.A(new_n662), .B(new_n652), .Y(new_n721));
  nand_4 g00345(.A(new_n721), .B(new_n720), .Y(new_n722));
  nand_4 g00346(.A(n7388), .B(n5814), .Y(new_n723));
  nand_4 g00347(.A(n12704), .B(n11892), .Y(new_n724));
  nand_4 g00348(.A(n7965), .B(n4903), .Y(new_n725));
  not_3  g00349(.A(new_n725), .Y(new_n726));
  xor_3  g00350(.A(new_n726), .B(new_n724), .Y(new_n727));
  xnor_3 g00351(.A(new_n727), .B(new_n723), .Y(new_n728));
  not_3  g00352(.A(new_n728), .Y(new_n729));
  and_4  g00353(.A(new_n729), .B(new_n722), .Y(new_n730));
  nor_4  g00354(.A(new_n729), .B(new_n722), .Y(new_n731));
  nor_4  g00355(.A(new_n731), .B(new_n730), .Y(new_n732));
  nor_4  g00356(.A(new_n646), .B(new_n645), .Y(new_n733));
  not_3  g00357(.A(new_n733), .Y(new_n734));
  nand_4 g00358(.A(n7294), .B(n2393), .Y(new_n735));
  xor_3  g00359(.A(new_n735), .B(new_n734), .Y(new_n736));
  nand_4 g00360(.A(n10848), .B(n3986), .Y(new_n737));
  nand_4 g00361(.A(n5860), .B(n1980), .Y(new_n738));
  nand_4 g00362(.A(n8028), .B(n5857), .Y(new_n739));
  not_3  g00363(.A(new_n739), .Y(new_n740));
  xor_3  g00364(.A(new_n740), .B(new_n738), .Y(new_n741));
  xnor_3 g00365(.A(new_n741), .B(new_n737), .Y(new_n742));
  xnor_3 g00366(.A(new_n742), .B(new_n736), .Y(new_n743));
  xnor_3 g00367(.A(new_n743), .B(new_n732), .Y(new_n744));
  nor_4  g00368(.A(new_n667), .B(new_n663), .Y(new_n745));
  not_3  g00369(.A(new_n745), .Y(new_n746));
  nor_4  g00370(.A(new_n665), .B(new_n664), .Y(new_n747));
  nor_4  g00371(.A(new_n686), .B(new_n668), .Y(new_n748));
  xnor_3 g00372(.A(new_n748), .B(new_n747), .Y(new_n749));
  nand_4 g00373(.A(new_n749), .B(new_n746), .Y(new_n750));
  xnor_3 g00374(.A(new_n750), .B(new_n744), .Y(new_n751));
  xnor_3 g00375(.A(new_n751), .B(new_n719), .Y(new_n752));
  nand_4 g00376(.A(n7965), .B(n5814), .Y(new_n753_1));
  not_3  g00377(.A(new_n753_1), .Y(new_n754));
  xnor_3 g00378(.A(new_n717), .B(new_n687), .Y(new_n755));
  nand_4 g00379(.A(new_n755), .B(new_n754), .Y(new_n756));
  not_3  g00380(.A(new_n755), .Y(new_n757));
  nand_4 g00381(.A(new_n757), .B(new_n753_1), .Y(new_n758));
  xnor_3 g00382(.A(new_n712), .B(new_n709), .Y(new_n759));
  not_3  g00383(.A(new_n703), .Y(new_n760));
  nand_4 g00384(.A(n8028), .B(n7965), .Y(new_n761));
  nand_4 g00385(.A(new_n761), .B(new_n705), .Y(new_n762));
  nand_4 g00386(.A(new_n762), .B(new_n702), .Y(new_n763));
  nand_4 g00387(.A(new_n763), .B(new_n760), .Y(new_n764));
  not_3  g00388(.A(new_n764), .Y(new_n765));
  nor_4  g00389(.A(new_n765), .B(new_n704), .Y(new_n766));
  not_3  g00390(.A(new_n766), .Y(new_n767));
  nor_4  g00391(.A(new_n767), .B(new_n759), .Y(new_n768));
  not_3  g00392(.A(new_n768), .Y(new_n769));
  xnor_3 g00393(.A(new_n715), .B(new_n695), .Y(new_n770));
  nor_4  g00394(.A(new_n770), .B(new_n769), .Y(new_n771));
  nand_4 g00395(.A(new_n771), .B(new_n758), .Y(new_n772));
  nand_4 g00396(.A(new_n772), .B(new_n756), .Y(new_n773));
  xnor_3 g00397(.A(new_n773), .B(new_n752), .Y(new_n774));
  xnor_3 g00398(.A(new_n774), .B(new_n643), .Y(new_n775));
  xnor_3 g00399(.A(new_n636), .B(new_n635), .Y(new_n776));
  not_3  g00400(.A(new_n625), .Y(new_n777));
  nor_4  g00401(.A(new_n632), .B(new_n777), .Y(new_n778));
  nor_4  g00402(.A(new_n778), .B(new_n634), .Y(new_n779));
  not_3  g00403(.A(new_n759), .Y(new_n780));
  nor_4  g00404(.A(new_n766), .B(new_n780), .Y(new_n781));
  nor_4  g00405(.A(new_n781), .B(new_n768), .Y(new_n782));
  nor_4  g00406(.A(new_n782), .B(new_n779), .Y(new_n783_1));
  not_3  g00407(.A(new_n783_1), .Y(new_n784));
  not_3  g00408(.A(new_n782), .Y(new_n785));
  xnor_3 g00409(.A(new_n785), .B(new_n779), .Y(new_n786));
  nor_4  g00410(.A(new_n762), .B(new_n702), .Y(new_n787));
  nor_4  g00411(.A(new_n787), .B(new_n764), .Y(new_n788));
  nand_4 g00412(.A(new_n628), .B(new_n569), .Y(new_n789));
  nand_4 g00413(.A(new_n789), .B(new_n631), .Y(new_n790));
  not_3  g00414(.A(new_n790), .Y(new_n791));
  nand_4 g00415(.A(new_n791), .B(new_n788), .Y(new_n792));
  not_3  g00416(.A(new_n792), .Y(new_n793));
  xnor_3 g00417(.A(new_n791), .B(new_n788), .Y(new_n794));
  not_3  g00418(.A(new_n761), .Y(new_n795));
  nand_4 g00419(.A(new_n795), .B(new_n627), .Y(new_n796));
  nand_4 g00420(.A(n5331), .B(n1512), .Y(new_n797));
  nand_4 g00421(.A(n8476), .B(n1564), .Y(new_n798));
  xnor_3 g00422(.A(new_n798), .B(new_n797), .Y(new_n799));
  nor_4  g00423(.A(new_n799), .B(new_n796), .Y(new_n800));
  xnor_3 g00424(.A(new_n799), .B(new_n796), .Y(new_n801));
  nand_4 g00425(.A(n8028), .B(n7388), .Y(new_n802));
  nand_4 g00426(.A(n10848), .B(n7965), .Y(new_n803));
  xnor_3 g00427(.A(new_n803), .B(new_n802), .Y(new_n804));
  nor_4  g00428(.A(new_n804), .B(new_n801), .Y(new_n805));
  nor_4  g00429(.A(new_n805), .B(new_n800), .Y(new_n806_1));
  nor_4  g00430(.A(new_n806_1), .B(new_n794), .Y(new_n807));
  nor_4  g00431(.A(new_n807), .B(new_n793), .Y(new_n808));
  nand_4 g00432(.A(new_n808), .B(new_n786), .Y(new_n809));
  nand_4 g00433(.A(new_n809), .B(new_n784), .Y(new_n810));
  nand_4 g00434(.A(new_n810), .B(new_n776), .Y(new_n811));
  not_3  g00435(.A(new_n811), .Y(new_n812));
  not_3  g00436(.A(new_n770), .Y(new_n813));
  nor_4  g00437(.A(new_n813), .B(new_n768), .Y(new_n814));
  nor_4  g00438(.A(new_n814), .B(new_n771), .Y(new_n815));
  xnor_3 g00439(.A(new_n810), .B(new_n776), .Y(new_n816));
  nor_4  g00440(.A(new_n816), .B(new_n815), .Y(new_n817));
  nor_4  g00441(.A(new_n817), .B(new_n812), .Y(new_n818));
  xnor_3 g00442(.A(new_n639), .B(new_n638), .Y(new_n819));
  not_3  g00443(.A(new_n819), .Y(new_n820));
  nand_4 g00444(.A(new_n820), .B(new_n818), .Y(new_n821));
  xnor_3 g00445(.A(new_n819), .B(new_n818), .Y(new_n822));
  nand_4 g00446(.A(new_n758), .B(new_n756), .Y(new_n823));
  xnor_3 g00447(.A(new_n823), .B(new_n771), .Y(new_n824));
  nand_4 g00448(.A(new_n824), .B(new_n822), .Y(new_n825));
  nand_4 g00449(.A(new_n825), .B(new_n821), .Y(new_n826));
  xnor_3 g00450(.A(new_n826), .B(new_n775), .Y(new_n827));
  xnor_3 g00451(.A(new_n827), .B(new_n513), .Y(new_n828));
  not_3  g00452(.A(new_n510), .Y(new_n829));
  xnor_3 g00453(.A(new_n829), .B(new_n509), .Y(new_n830));
  xnor_3 g00454(.A(new_n508), .B(new_n507), .Y(new_n831));
  not_3  g00455(.A(new_n498), .Y(new_n832));
  nor_4  g00456(.A(new_n504), .B(new_n832), .Y(new_n833));
  nor_4  g00457(.A(new_n833), .B(new_n506), .Y(new_n834));
  not_3  g00458(.A(new_n834), .Y(new_n835));
  xnor_3 g00459(.A(new_n761), .B(new_n626), .Y(new_n836));
  nor_4  g00460(.A(new_n836), .B(new_n499), .Y(new_n837_1));
  not_3  g00461(.A(new_n837_1), .Y(new_n838));
  nand_4 g00462(.A(n7354), .B(n6776), .Y(new_n839));
  nand_4 g00463(.A(n8759), .B(n7500), .Y(new_n840));
  xnor_3 g00464(.A(new_n840), .B(new_n839), .Y(new_n841));
  nand_4 g00465(.A(new_n841), .B(new_n838), .Y(new_n842));
  xnor_3 g00466(.A(new_n804), .B(new_n801), .Y(new_n843));
  xnor_3 g00467(.A(new_n841), .B(new_n837_1), .Y(new_n844_1));
  nand_4 g00468(.A(new_n844_1), .B(new_n843), .Y(new_n845));
  nand_4 g00469(.A(new_n845), .B(new_n842), .Y(new_n846));
  not_3  g00470(.A(new_n503_1), .Y(new_n847));
  not_3  g00471(.A(new_n501), .Y(new_n848));
  nor_4  g00472(.A(new_n848), .B(new_n446), .Y(new_n849));
  nor_4  g00473(.A(new_n849), .B(new_n847), .Y(new_n850));
  not_3  g00474(.A(new_n850), .Y(new_n851));
  nand_4 g00475(.A(new_n851), .B(new_n846), .Y(new_n852));
  xnor_3 g00476(.A(new_n806_1), .B(new_n794), .Y(new_n853));
  xnor_3 g00477(.A(new_n850), .B(new_n846), .Y(new_n854));
  nand_4 g00478(.A(new_n854), .B(new_n853), .Y(new_n855));
  nand_4 g00479(.A(new_n855), .B(new_n852), .Y(new_n856));
  nand_4 g00480(.A(new_n856), .B(new_n835), .Y(new_n857));
  not_3  g00481(.A(new_n808), .Y(new_n858));
  xnor_3 g00482(.A(new_n858), .B(new_n786), .Y(new_n859));
  xnor_3 g00483(.A(new_n856), .B(new_n834), .Y(new_n860));
  nand_4 g00484(.A(new_n860), .B(new_n859), .Y(new_n861));
  nand_4 g00485(.A(new_n861), .B(new_n857), .Y(new_n862));
  nand_4 g00486(.A(new_n862), .B(new_n831), .Y(new_n863));
  not_3  g00487(.A(new_n815), .Y(new_n864));
  xnor_3 g00488(.A(new_n816), .B(new_n864), .Y(new_n865));
  not_3  g00489(.A(new_n863), .Y(new_n866));
  nor_4  g00490(.A(new_n862), .B(new_n831), .Y(new_n867));
  nor_4  g00491(.A(new_n867), .B(new_n866), .Y(new_n868));
  nand_4 g00492(.A(new_n868), .B(new_n865), .Y(new_n869));
  nand_4 g00493(.A(new_n869), .B(new_n863), .Y(new_n870));
  not_3  g00494(.A(new_n870), .Y(new_n871));
  nor_4  g00495(.A(new_n871), .B(new_n830), .Y(new_n872));
  xnor_3 g00496(.A(new_n870), .B(new_n830), .Y(new_n873));
  not_3  g00497(.A(new_n873), .Y(new_n874));
  xnor_3 g00498(.A(new_n820), .B(new_n818), .Y(new_n875));
  xnor_3 g00499(.A(new_n824), .B(new_n875), .Y(new_n876));
  nor_4  g00500(.A(new_n876), .B(new_n874), .Y(new_n877));
  nor_4  g00501(.A(new_n877), .B(new_n872), .Y(new_n878));
  xnor_3 g00502(.A(new_n878), .B(new_n828), .Y(new_n879));
  nand_4 g00503(.A(n12720), .B(n4312), .Y(new_n880));
  not_3  g00504(.A(new_n880), .Y(new_n881));
  nand_4 g00505(.A(n12025), .B(n6038), .Y(new_n882));
  nand_4 g00506(.A(n12705), .B(n2509), .Y(new_n883));
  not_3  g00507(.A(new_n883), .Y(new_n884));
  xor_3  g00508(.A(new_n884), .B(new_n882), .Y(new_n885));
  not_3  g00509(.A(new_n885), .Y(new_n886));
  xor_3  g00510(.A(new_n886), .B(new_n881), .Y(new_n887));
  nand_4 g00511(.A(n12705), .B(n6038), .Y(new_n888));
  not_3  g00512(.A(new_n888), .Y(new_n889));
  nand_4 g00513(.A(n12720), .B(n1097), .Y(new_n890));
  not_3  g00514(.A(new_n890), .Y(new_n891));
  nor_4  g00515(.A(new_n891), .B(new_n889), .Y(new_n892));
  nand_4 g00516(.A(n4312), .B(n2509), .Y(new_n893));
  not_3  g00517(.A(new_n893), .Y(new_n894));
  xor_3  g00518(.A(new_n891), .B(new_n888), .Y(new_n895));
  nor_4  g00519(.A(new_n895), .B(new_n894), .Y(new_n896));
  nor_4  g00520(.A(new_n896), .B(new_n892), .Y(new_n897));
  xnor_3 g00521(.A(new_n897), .B(new_n887), .Y(new_n898));
  nand_4 g00522(.A(n2508), .B(n1097), .Y(new_n899));
  nand_4 g00523(.A(n5964), .B(n2585), .Y(new_n900));
  xor_3  g00524(.A(new_n900), .B(new_n899), .Y(new_n901));
  not_3  g00525(.A(new_n901), .Y(new_n902));
  nor_4  g00526(.A(new_n902), .B(new_n898), .Y(new_n903));
  not_3  g00527(.A(new_n898), .Y(new_n904));
  nor_4  g00528(.A(new_n901), .B(new_n904), .Y(new_n905));
  nor_4  g00529(.A(new_n905), .B(new_n903), .Y(new_n906));
  nand_4 g00530(.A(n5964), .B(n2508), .Y(new_n907));
  not_3  g00531(.A(new_n907), .Y(new_n908));
  xnor_3 g00532(.A(new_n895), .B(new_n893), .Y(new_n909));
  not_3  g00533(.A(new_n909), .Y(new_n910));
  nor_4  g00534(.A(new_n910), .B(new_n908), .Y(new_n911_1));
  xor_3  g00535(.A(new_n910), .B(new_n907), .Y(new_n912));
  nand_4 g00536(.A(n6038), .B(n4312), .Y(new_n913));
  not_3  g00537(.A(new_n913), .Y(new_n914));
  nand_4 g00538(.A(n12720), .B(n5964), .Y(new_n915));
  not_3  g00539(.A(new_n915), .Y(new_n916));
  nor_4  g00540(.A(new_n916), .B(new_n914), .Y(new_n917));
  nor_4  g00541(.A(new_n915), .B(new_n913), .Y(new_n918));
  nand_4 g00542(.A(n2509), .B(n1097), .Y(new_n919));
  not_3  g00543(.A(new_n919), .Y(new_n920));
  nor_4  g00544(.A(new_n920), .B(new_n918), .Y(new_n921));
  nor_4  g00545(.A(new_n921), .B(new_n917), .Y(new_n922));
  nor_4  g00546(.A(new_n922), .B(new_n912), .Y(new_n923));
  nor_4  g00547(.A(new_n923), .B(new_n911_1), .Y(new_n924));
  not_3  g00548(.A(new_n924), .Y(new_n925));
  xnor_3 g00549(.A(new_n925), .B(new_n906), .Y(new_n926));
  nand_4 g00550(.A(n5305), .B(n2585), .Y(new_n927));
  not_3  g00551(.A(new_n922), .Y(new_n928));
  xnor_3 g00552(.A(new_n928), .B(new_n912), .Y(new_n929));
  nand_4 g00553(.A(new_n929), .B(new_n927), .Y(new_n930));
  not_3  g00554(.A(new_n930), .Y(new_n931));
  nor_4  g00555(.A(new_n929), .B(new_n927), .Y(new_n932));
  nor_4  g00556(.A(new_n932), .B(new_n931), .Y(new_n933));
  nand_4 g00557(.A(n5305), .B(n2508), .Y(new_n934));
  nand_4 g00558(.A(n6038), .B(n1097), .Y(new_n935));
  not_3  g00559(.A(new_n935), .Y(new_n936));
  nand_4 g00560(.A(n12720), .B(n5305), .Y(new_n937));
  not_3  g00561(.A(new_n937), .Y(new_n938));
  nand_4 g00562(.A(new_n938), .B(new_n936), .Y(new_n939));
  nand_4 g00563(.A(new_n937), .B(new_n935), .Y(new_n940));
  nand_4 g00564(.A(n5964), .B(n2509), .Y(new_n941));
  not_3  g00565(.A(new_n941), .Y(new_n942));
  nand_4 g00566(.A(new_n942), .B(new_n940), .Y(new_n943));
  nand_4 g00567(.A(new_n943), .B(new_n939), .Y(new_n944));
  not_3  g00568(.A(new_n944), .Y(new_n945));
  nor_4  g00569(.A(new_n945), .B(new_n934), .Y(new_n946));
  xor_3  g00570(.A(new_n944), .B(new_n934), .Y(new_n947));
  nor_4  g00571(.A(new_n918), .B(new_n917), .Y(new_n948));
  xor_3  g00572(.A(new_n948), .B(new_n919), .Y(new_n949));
  nor_4  g00573(.A(new_n949), .B(new_n947), .Y(new_n950));
  nor_4  g00574(.A(new_n950), .B(new_n946), .Y(new_n951));
  nand_4 g00575(.A(new_n951), .B(new_n933), .Y(new_n952));
  nand_4 g00576(.A(new_n952), .B(new_n930), .Y(new_n953));
  not_3  g00577(.A(new_n953), .Y(new_n954));
  nand_4 g00578(.A(new_n954), .B(new_n926), .Y(new_n955));
  nor_4  g00579(.A(new_n885), .B(new_n880), .Y(new_n956));
  nand_4 g00580(.A(new_n897), .B(new_n887), .Y(new_n957));
  not_3  g00581(.A(new_n957), .Y(new_n958));
  nor_4  g00582(.A(new_n958), .B(new_n956), .Y(new_n959));
  not_3  g00583(.A(new_n959), .Y(new_n960));
  nand_4 g00584(.A(n5964), .B(n4005), .Y(new_n961));
  nand_4 g00585(.A(n2585), .B(n1097), .Y(new_n962));
  nand_4 g00586(.A(n12706), .B(n5305), .Y(new_n963));
  nand_4 g00587(.A(new_n963), .B(new_n962), .Y(new_n964));
  not_3  g00588(.A(new_n962), .Y(new_n965));
  not_3  g00589(.A(new_n963), .Y(new_n966));
  nand_4 g00590(.A(new_n966), .B(new_n965), .Y(new_n967));
  and_4  g00591(.A(new_n967), .B(new_n964), .Y(new_n968));
  xor_3  g00592(.A(new_n968), .B(new_n961), .Y(new_n969));
  xnor_3 g00593(.A(new_n969), .B(new_n960), .Y(new_n970));
  nor_4  g00594(.A(new_n883), .B(new_n882), .Y(new_n971));
  nand_4 g00595(.A(n4312), .B(n2508), .Y(new_n972));
  not_3  g00596(.A(new_n972), .Y(new_n973));
  xor_3  g00597(.A(new_n973), .B(new_n971), .Y(new_n974));
  nand_4 g00598(.A(n12025), .B(n2509), .Y(new_n975));
  not_3  g00599(.A(new_n975), .Y(new_n976));
  nand_4 g00600(.A(n12720), .B(n12705), .Y(new_n977));
  nand_4 g00601(.A(n11257), .B(n6038), .Y(new_n978));
  not_3  g00602(.A(new_n978), .Y(new_n979));
  xor_3  g00603(.A(new_n979), .B(new_n977), .Y(new_n980));
  xnor_3 g00604(.A(new_n980), .B(new_n976), .Y(new_n981));
  xnor_3 g00605(.A(new_n981), .B(new_n974), .Y(new_n982));
  not_3  g00606(.A(new_n982), .Y(new_n983));
  xnor_3 g00607(.A(new_n983), .B(new_n970), .Y(new_n984));
  nor_4  g00608(.A(new_n900), .B(new_n899), .Y(new_n985));
  nand_4 g00609(.A(new_n924), .B(new_n906), .Y(new_n986));
  xnor_3 g00610(.A(new_n986), .B(new_n985), .Y(new_n987));
  nor_4  g00611(.A(new_n987), .B(new_n903), .Y(new_n988));
  xnor_3 g00612(.A(new_n988), .B(new_n984), .Y(new_n989));
  xnor_3 g00613(.A(new_n989), .B(new_n955), .Y(new_n990));
  nand_4 g00614(.A(n5305), .B(n4005), .Y(new_n991));
  not_3  g00615(.A(new_n926), .Y(new_n992_1));
  xnor_3 g00616(.A(new_n953), .B(new_n992_1), .Y(new_n993));
  nor_4  g00617(.A(new_n993), .B(new_n991), .Y(new_n994));
  not_3  g00618(.A(new_n994), .Y(new_n995));
  nand_4 g00619(.A(new_n993), .B(new_n991), .Y(new_n996_1));
  and_4  g00620(.A(new_n940), .B(new_n939), .Y(new_n997));
  nand_4 g00621(.A(n6038), .B(n5964), .Y(new_n998));
  nand_4 g00622(.A(n5305), .B(n2509), .Y(new_n999));
  nor_4  g00623(.A(new_n999), .B(new_n998), .Y(new_n1000));
  not_3  g00624(.A(new_n1000), .Y(new_n1001));
  nor_4  g00625(.A(new_n1001), .B(new_n997), .Y(new_n1002));
  not_3  g00626(.A(new_n1002), .Y(new_n1003));
  xnor_3 g00627(.A(new_n949), .B(new_n947), .Y(new_n1004));
  nor_4  g00628(.A(new_n1004), .B(new_n1003), .Y(new_n1005));
  xnor_3 g00629(.A(new_n951), .B(new_n933), .Y(new_n1006));
  nand_4 g00630(.A(new_n1006), .B(new_n1005), .Y(new_n1007));
  not_3  g00631(.A(new_n1007), .Y(new_n1008));
  nand_4 g00632(.A(new_n1008), .B(new_n996_1), .Y(new_n1009));
  nand_4 g00633(.A(new_n1009), .B(new_n995), .Y(new_n1010));
  xnor_3 g00634(.A(new_n1010), .B(new_n990), .Y(new_n1011));
  xnor_3 g00635(.A(new_n876), .B(new_n874), .Y(new_n1012));
  xnor_3 g00636(.A(new_n993), .B(new_n991), .Y(new_n1013));
  xnor_3 g00637(.A(new_n1013), .B(new_n1008), .Y(new_n1014));
  nor_4  g00638(.A(new_n1014), .B(new_n1012), .Y(new_n1015));
  xnor_3 g00639(.A(new_n876), .B(new_n873), .Y(new_n1016));
  xnor_3 g00640(.A(new_n1013), .B(new_n1007), .Y(new_n1017));
  nor_4  g00641(.A(new_n1017), .B(new_n1016), .Y(new_n1018));
  xnor_3 g00642(.A(new_n1006), .B(new_n1005), .Y(new_n1019));
  xnor_3 g00643(.A(new_n868), .B(new_n865), .Y(new_n1020_1));
  not_3  g00644(.A(new_n1020_1), .Y(new_n1021));
  nor_4  g00645(.A(new_n1021), .B(new_n1019), .Y(new_n1022));
  not_3  g00646(.A(new_n1022), .Y(new_n1023));
  xnor_3 g00647(.A(new_n1020_1), .B(new_n1019), .Y(new_n1024));
  not_3  g00648(.A(new_n1004), .Y(new_n1025));
  xor_3  g00649(.A(new_n1025), .B(new_n1003), .Y(new_n1026));
  xnor_3 g00650(.A(new_n860), .B(new_n859), .Y(new_n1027));
  not_3  g00651(.A(new_n1027), .Y(new_n1028));
  nor_4  g00652(.A(new_n1028), .B(new_n1026), .Y(new_n1029));
  not_3  g00653(.A(new_n1029), .Y(new_n1030));
  not_3  g00654(.A(new_n853), .Y(new_n1031));
  xor_3  g00655(.A(new_n854), .B(new_n1031), .Y(new_n1032));
  nand_4 g00656(.A(n6038), .B(n5305), .Y(new_n1033));
  not_3  g00657(.A(new_n1033), .Y(new_n1034));
  nor_4  g00658(.A(new_n1034), .B(new_n941), .Y(new_n1035));
  nor_4  g00659(.A(new_n1035), .B(new_n997), .Y(new_n1036));
  nor_4  g00660(.A(new_n1034), .B(new_n943), .Y(new_n1037));
  nor_4  g00661(.A(new_n1037), .B(new_n1036), .Y(new_n1038));
  nor_4  g00662(.A(new_n1038), .B(new_n1032), .Y(new_n1039));
  not_3  g00663(.A(new_n1032), .Y(new_n1040));
  xor_3  g00664(.A(new_n1038), .B(new_n1040), .Y(new_n1041));
  xor_3  g00665(.A(new_n836), .B(new_n499), .Y(new_n1042));
  not_3  g00666(.A(new_n1042), .Y(new_n1043));
  nor_4  g00667(.A(new_n1043), .B(new_n1033), .Y(new_n1044));
  not_3  g00668(.A(new_n1044), .Y(new_n1045));
  xor_3  g00669(.A(new_n999), .B(new_n998), .Y(new_n1046));
  not_3  g00670(.A(new_n1046), .Y(new_n1047));
  nor_4  g00671(.A(new_n1047), .B(new_n1045), .Y(new_n1048));
  xor_3  g00672(.A(new_n844_1), .B(new_n843), .Y(new_n1049));
  xor_3  g00673(.A(new_n1047), .B(new_n1044), .Y(new_n1050));
  nor_4  g00674(.A(new_n1050), .B(new_n1049), .Y(new_n1051));
  nor_4  g00675(.A(new_n1051), .B(new_n1048), .Y(new_n1052));
  not_3  g00676(.A(new_n1052), .Y(new_n1053));
  nor_4  g00677(.A(new_n1053), .B(new_n1041), .Y(new_n1054));
  nor_4  g00678(.A(new_n1054), .B(new_n1039), .Y(new_n1055));
  not_3  g00679(.A(new_n1026), .Y(new_n1056));
  nor_4  g00680(.A(new_n1027), .B(new_n1056), .Y(new_n1057));
  nor_4  g00681(.A(new_n1057), .B(new_n1029), .Y(new_n1058));
  nand_4 g00682(.A(new_n1058), .B(new_n1055), .Y(new_n1059));
  nand_4 g00683(.A(new_n1059), .B(new_n1030), .Y(new_n1060));
  nand_4 g00684(.A(new_n1060), .B(new_n1024), .Y(new_n1061));
  nand_4 g00685(.A(new_n1061), .B(new_n1023), .Y(new_n1062));
  nor_4  g00686(.A(new_n1062), .B(new_n1018), .Y(new_n1063));
  nor_4  g00687(.A(new_n1063), .B(new_n1015), .Y(new_n1064));
  nor_4  g00688(.A(new_n1064), .B(new_n1011), .Y(new_n1065));
  nand_4 g00689(.A(new_n1064), .B(new_n1011), .Y(new_n1066));
  not_3  g00690(.A(new_n1066), .Y(new_n1067_1));
  nor_4  g00691(.A(new_n1067_1), .B(new_n1065), .Y(new_n1068));
  xnor_3 g00692(.A(new_n1068), .B(new_n879), .Y(n226));
  nand_4 g00693(.A(n5305), .B(n4634), .Y(new_n1070));
  not_3  g00694(.A(new_n1070), .Y(new_n1071));
  nand_4 g00695(.A(n10223), .B(n5305), .Y(new_n1072));
  not_3  g00696(.A(new_n1072), .Y(new_n1073));
  nand_4 g00697(.A(n7265), .B(n1097), .Y(new_n1074));
  not_3  g00698(.A(new_n1074), .Y(new_n1075));
  nor_4  g00699(.A(new_n1075), .B(new_n1073), .Y(new_n1076));
  nor_4  g00700(.A(new_n1074), .B(new_n1072), .Y(new_n1077));
  nand_4 g00701(.A(n5964), .B(n2879), .Y(new_n1078));
  not_3  g00702(.A(new_n1078), .Y(new_n1079));
  nor_4  g00703(.A(new_n1079), .B(new_n1077), .Y(new_n1080));
  nor_4  g00704(.A(new_n1080), .B(new_n1076), .Y(new_n1081));
  nand_4 g00705(.A(new_n1081), .B(new_n1071), .Y(new_n1082));
  not_3  g00706(.A(new_n1082), .Y(new_n1083));
  nor_4  g00707(.A(new_n1081), .B(new_n1071), .Y(new_n1084));
  nor_4  g00708(.A(new_n1084), .B(new_n1083), .Y(new_n1085));
  nand_4 g00709(.A(n2879), .B(n1097), .Y(new_n1086));
  not_3  g00710(.A(new_n1086), .Y(new_n1087));
  nand_4 g00711(.A(n10223), .B(n5964), .Y(new_n1088));
  nand_4 g00712(.A(n7265), .B(n4312), .Y(new_n1089));
  xnor_3 g00713(.A(new_n1089), .B(new_n1088), .Y(new_n1090));
  xnor_3 g00714(.A(new_n1090), .B(new_n1087), .Y(new_n1091));
  xor_3  g00715(.A(new_n1091), .B(new_n1085), .Y(new_n1092));
  not_3  g00716(.A(new_n1092), .Y(new_n1093));
  nand_4 g00717(.A(n7265), .B(n5305), .Y(new_n1094_1));
  not_3  g00718(.A(new_n1094_1), .Y(new_n1095));
  nor_4  g00719(.A(new_n1095), .B(new_n1078), .Y(new_n1096));
  nor_4  g00720(.A(new_n1077), .B(new_n1076), .Y(new_n1097_1));
  nor_4  g00721(.A(new_n1097_1), .B(new_n1096), .Y(new_n1098));
  not_3  g00722(.A(new_n1098), .Y(new_n1099));
  nor_4  g00723(.A(new_n1099), .B(new_n1078), .Y(new_n1100));
  not_3  g00724(.A(new_n1100), .Y(new_n1101));
  xor_3  g00725(.A(new_n1101), .B(new_n1093), .Y(new_n1102));
  nand_4 g00726(.A(n8759), .B(n7946), .Y(new_n1103));
  nand_4 g00727(.A(n5331), .B(n2558), .Y(new_n1104));
  nand_4 g00728(.A(n9763), .B(n7965), .Y(new_n1105));
  xnor_3 g00729(.A(new_n1105), .B(new_n1104), .Y(new_n1106));
  nor_4  g00730(.A(new_n1106), .B(new_n1103), .Y(new_n1107));
  not_3  g00731(.A(new_n1107), .Y(new_n1108));
  nand_4 g00732(.A(n7946), .B(n6776), .Y(new_n1109));
  nand_4 g00733(.A(n8759), .B(n2024), .Y(new_n1110));
  xnor_3 g00734(.A(new_n1110), .B(new_n1109), .Y(new_n1111));
  nor_4  g00735(.A(new_n1111), .B(new_n1108), .Y(new_n1112));
  not_3  g00736(.A(new_n1112), .Y(new_n1113));
  nor_4  g00737(.A(new_n1105), .B(new_n1104), .Y(new_n1114));
  nand_4 g00738(.A(n9111), .B(n7965), .Y(new_n1115));
  nand_4 g00739(.A(n9763), .B(n7388), .Y(new_n1116));
  xnor_3 g00740(.A(new_n1116), .B(new_n1115), .Y(new_n1117));
  not_3  g00741(.A(new_n1117), .Y(new_n1118));
  xnor_3 g00742(.A(new_n1118), .B(new_n1114), .Y(new_n1119));
  nand_4 g00743(.A(n5331), .B(n2498), .Y(new_n1120));
  nand_4 g00744(.A(n8476), .B(n2558), .Y(new_n1121));
  and_4  g00745(.A(new_n1121), .B(new_n1120), .Y(new_n1122));
  nor_4  g00746(.A(new_n1121), .B(new_n1120), .Y(new_n1123));
  nor_4  g00747(.A(new_n1123), .B(new_n1122), .Y(new_n1124));
  xnor_3 g00748(.A(new_n1124), .B(new_n1119), .Y(new_n1125));
  not_3  g00749(.A(new_n1111), .Y(new_n1126));
  nor_4  g00750(.A(new_n1126), .B(new_n1107), .Y(new_n1127));
  nor_4  g00751(.A(new_n1127), .B(new_n1112), .Y(new_n1128));
  nand_4 g00752(.A(new_n1128), .B(new_n1125), .Y(new_n1129));
  nand_4 g00753(.A(new_n1129), .B(new_n1113), .Y(new_n1130));
  not_3  g00754(.A(new_n1130), .Y(new_n1131));
  not_3  g00755(.A(new_n1103), .Y(new_n1132));
  nand_4 g00756(.A(n6776), .B(n2024), .Y(new_n1133));
  nor_4  g00757(.A(new_n1133), .B(new_n1132), .Y(new_n1134));
  nand_4 g00758(.A(n12299), .B(n7946), .Y(new_n1135));
  not_3  g00759(.A(new_n1135), .Y(new_n1136_1));
  nand_4 g00760(.A(n9189), .B(n8759), .Y(new_n1137));
  not_3  g00761(.A(new_n1137), .Y(new_n1138_1));
  nand_4 g00762(.A(new_n1138_1), .B(new_n1136_1), .Y(new_n1139));
  nand_4 g00763(.A(new_n1137), .B(new_n1135), .Y(new_n1140));
  nand_4 g00764(.A(new_n1140), .B(new_n1139), .Y(new_n1141));
  not_3  g00765(.A(new_n1141), .Y(new_n1142));
  nor_4  g00766(.A(new_n1142), .B(new_n1134), .Y(new_n1143));
  not_3  g00767(.A(new_n1133), .Y(new_n1144));
  nand_4 g00768(.A(new_n1140), .B(new_n1144), .Y(new_n1145));
  nor_4  g00769(.A(new_n1145), .B(new_n1132), .Y(new_n1146));
  nor_4  g00770(.A(new_n1146), .B(new_n1143), .Y(new_n1147));
  not_3  g00771(.A(new_n1147), .Y(new_n1148));
  nor_4  g00772(.A(new_n1148), .B(new_n1131), .Y(new_n1149));
  nor_4  g00773(.A(new_n1147), .B(new_n1130), .Y(new_n1150));
  nor_4  g00774(.A(new_n1150), .B(new_n1149), .Y(new_n1151));
  nor_4  g00775(.A(new_n1118), .B(new_n1114), .Y(new_n1152));
  nor_4  g00776(.A(new_n1124), .B(new_n1119), .Y(new_n1153));
  nor_4  g00777(.A(new_n1153), .B(new_n1152), .Y(new_n1154));
  not_3  g00778(.A(new_n1105), .Y(new_n1155));
  nand_4 g00779(.A(n9111), .B(n7388), .Y(new_n1156));
  nor_4  g00780(.A(new_n1156), .B(new_n1155), .Y(new_n1157));
  nand_4 g00781(.A(n11892), .B(n9763), .Y(new_n1158));
  nand_4 g00782(.A(n7965), .B(n3342), .Y(new_n1159));
  nand_4 g00783(.A(new_n1159), .B(new_n1158), .Y(new_n1160));
  nor_4  g00784(.A(new_n1159), .B(new_n1158), .Y(new_n1161));
  not_3  g00785(.A(new_n1161), .Y(new_n1162));
  nand_4 g00786(.A(new_n1162), .B(new_n1160), .Y(new_n1163));
  not_3  g00787(.A(new_n1163), .Y(new_n1164));
  nor_4  g00788(.A(new_n1164), .B(new_n1157), .Y(new_n1165));
  not_3  g00789(.A(new_n1156), .Y(new_n1166));
  nand_4 g00790(.A(new_n1160), .B(new_n1166), .Y(new_n1167));
  nor_4  g00791(.A(new_n1167), .B(new_n1155), .Y(new_n1168));
  nor_4  g00792(.A(new_n1168), .B(new_n1165), .Y(new_n1169));
  xnor_3 g00793(.A(new_n1169), .B(new_n1154), .Y(new_n1170));
  not_3  g00794(.A(new_n1104), .Y(new_n1171));
  nand_4 g00795(.A(n8476), .B(n2498), .Y(new_n1172));
  nor_4  g00796(.A(new_n1172), .B(new_n1171), .Y(new_n1173));
  not_3  g00797(.A(new_n1173), .Y(new_n1174));
  nand_4 g00798(.A(n2558), .B(n2530), .Y(new_n1175));
  nand_4 g00799(.A(n5579), .B(n5331), .Y(new_n1176));
  nand_4 g00800(.A(new_n1176), .B(new_n1175), .Y(new_n1177));
  nor_4  g00801(.A(new_n1177), .B(new_n1174), .Y(new_n1178));
  not_3  g00802(.A(new_n1177), .Y(new_n1179));
  nor_4  g00803(.A(new_n1176), .B(new_n1175), .Y(new_n1180));
  nor_4  g00804(.A(new_n1180), .B(new_n1179), .Y(new_n1181));
  not_3  g00805(.A(new_n1181), .Y(new_n1182));
  nor_4  g00806(.A(new_n1182), .B(new_n1173), .Y(new_n1183));
  nor_4  g00807(.A(new_n1183), .B(new_n1178), .Y(new_n1184));
  not_3  g00808(.A(new_n1184), .Y(new_n1185));
  nor_4  g00809(.A(new_n1185), .B(new_n1170), .Y(new_n1186));
  not_3  g00810(.A(new_n1170), .Y(new_n1187));
  nor_4  g00811(.A(new_n1184), .B(new_n1187), .Y(new_n1188));
  nor_4  g00812(.A(new_n1188), .B(new_n1186), .Y(new_n1189));
  xnor_3 g00813(.A(new_n1189), .B(new_n1151), .Y(new_n1190));
  not_3  g00814(.A(new_n1190), .Y(new_n1191));
  not_3  g00815(.A(new_n1076), .Y(new_n1192));
  nand_4 g00816(.A(new_n1096), .B(new_n1192), .Y(new_n1193));
  nand_4 g00817(.A(new_n1193), .B(new_n1099), .Y(new_n1194));
  nor_4  g00818(.A(new_n1194), .B(new_n1191), .Y(new_n1195));
  not_3  g00819(.A(new_n1195), .Y(new_n1196));
  xor_3  g00820(.A(new_n1106), .B(new_n1103), .Y(new_n1197));
  nand_4 g00821(.A(new_n1197), .B(new_n1095), .Y(new_n1198_1));
  nand_4 g00822(.A(n7265), .B(n5964), .Y(new_n1199_1));
  nand_4 g00823(.A(n5305), .B(n2879), .Y(new_n1200));
  not_3  g00824(.A(new_n1200), .Y(new_n1201));
  xor_3  g00825(.A(new_n1201), .B(new_n1199_1), .Y(new_n1202));
  nand_4 g00826(.A(new_n1202), .B(new_n1198_1), .Y(new_n1203));
  not_3  g00827(.A(new_n1203), .Y(new_n1204));
  xor_3  g00828(.A(new_n1128), .B(new_n1125), .Y(new_n1205));
  not_3  g00829(.A(new_n1198_1), .Y(new_n1206));
  xor_3  g00830(.A(new_n1202), .B(new_n1206), .Y(new_n1207));
  nor_4  g00831(.A(new_n1207), .B(new_n1205), .Y(new_n1208));
  nor_4  g00832(.A(new_n1208), .B(new_n1204), .Y(new_n1209_1));
  not_3  g00833(.A(new_n1194), .Y(new_n1210));
  nor_4  g00834(.A(new_n1210), .B(new_n1190), .Y(new_n1211));
  nor_4  g00835(.A(new_n1211), .B(new_n1195), .Y(new_n1212));
  nand_4 g00836(.A(new_n1212), .B(new_n1209_1), .Y(new_n1213));
  nand_4 g00837(.A(new_n1213), .B(new_n1196), .Y(new_n1214));
  xnor_3 g00838(.A(new_n1214), .B(new_n1102), .Y(new_n1215));
  nand_4 g00839(.A(n8759), .B(n2522), .Y(new_n1216));
  nand_4 g00840(.A(new_n1145), .B(new_n1139), .Y(new_n1217));
  xnor_3 g00841(.A(new_n1217), .B(new_n1216), .Y(new_n1218));
  not_3  g00842(.A(new_n1218), .Y(new_n1219));
  nand_4 g00843(.A(n12299), .B(n2024), .Y(new_n1220));
  not_3  g00844(.A(new_n1220), .Y(new_n1221));
  nand_4 g00845(.A(n7946), .B(n7436), .Y(new_n1222));
  nand_4 g00846(.A(n9189), .B(n6776), .Y(new_n1223));
  xnor_3 g00847(.A(new_n1223), .B(new_n1222), .Y(new_n1224));
  xnor_3 g00848(.A(new_n1224), .B(new_n1221), .Y(new_n1225));
  xor_3  g00849(.A(new_n1225), .B(new_n1219), .Y(new_n1226));
  not_3  g00850(.A(new_n1143), .Y(new_n1227));
  nor_4  g00851(.A(new_n1227), .B(new_n1133), .Y(new_n1228));
  not_3  g00852(.A(new_n1228), .Y(new_n1229));
  xnor_3 g00853(.A(new_n1229), .B(new_n1226), .Y(new_n1230));
  not_3  g00854(.A(new_n1150), .Y(new_n1231));
  nand_4 g00855(.A(new_n1189), .B(new_n1151), .Y(new_n1232));
  nand_4 g00856(.A(new_n1232), .B(new_n1231), .Y(new_n1233));
  xnor_3 g00857(.A(new_n1233), .B(new_n1230), .Y(new_n1234));
  nand_4 g00858(.A(n5331), .B(n521), .Y(new_n1235));
  not_3  g00859(.A(new_n1172), .Y(new_n1236));
  nand_4 g00860(.A(new_n1177), .B(new_n1236), .Y(new_n1237));
  not_3  g00861(.A(new_n1237), .Y(new_n1238));
  nor_4  g00862(.A(new_n1238), .B(new_n1180), .Y(new_n1239));
  xnor_3 g00863(.A(new_n1239), .B(new_n1235), .Y(new_n1240));
  nand_4 g00864(.A(n12648), .B(n2558), .Y(new_n1241));
  nand_4 g00865(.A(n8476), .B(n5579), .Y(new_n1242));
  not_3  g00866(.A(new_n1242), .Y(new_n1243));
  nand_4 g00867(.A(n2530), .B(n2498), .Y(new_n1244));
  not_3  g00868(.A(new_n1244), .Y(new_n1245));
  nor_4  g00869(.A(new_n1245), .B(new_n1243), .Y(new_n1246));
  nor_4  g00870(.A(new_n1244), .B(new_n1242), .Y(new_n1247));
  nor_4  g00871(.A(new_n1247), .B(new_n1246), .Y(new_n1248));
  xnor_3 g00872(.A(new_n1248), .B(new_n1241), .Y(new_n1249));
  not_3  g00873(.A(new_n1249), .Y(new_n1250));
  xnor_3 g00874(.A(new_n1250), .B(new_n1240), .Y(new_n1251));
  not_3  g00875(.A(new_n1123), .Y(new_n1252));
  nor_4  g00876(.A(new_n1181), .B(new_n1252), .Y(new_n1253));
  not_3  g00877(.A(new_n1253), .Y(new_n1254));
  nor_4  g00878(.A(new_n1254), .B(new_n1251), .Y(new_n1255));
  not_3  g00879(.A(new_n1251), .Y(new_n1256));
  nor_4  g00880(.A(new_n1253), .B(new_n1256), .Y(new_n1257));
  nor_4  g00881(.A(new_n1257), .B(new_n1255), .Y(new_n1258));
  nand_4 g00882(.A(n7965), .B(n806), .Y(new_n1259));
  not_3  g00883(.A(new_n1167), .Y(new_n1260));
  nor_4  g00884(.A(new_n1260), .B(new_n1161), .Y(new_n1261));
  xnor_3 g00885(.A(new_n1261), .B(new_n1259), .Y(new_n1262));
  nand_4 g00886(.A(n9763), .B(n2393), .Y(new_n1263));
  nand_4 g00887(.A(n7388), .B(n3342), .Y(new_n1264));
  not_3  g00888(.A(new_n1264), .Y(new_n1265));
  nand_4 g00889(.A(n11892), .B(n9111), .Y(new_n1266));
  not_3  g00890(.A(new_n1266), .Y(new_n1267));
  nor_4  g00891(.A(new_n1267), .B(new_n1265), .Y(new_n1268));
  nor_4  g00892(.A(new_n1266), .B(new_n1264), .Y(new_n1269_1));
  nor_4  g00893(.A(new_n1269_1), .B(new_n1268), .Y(new_n1270));
  xnor_3 g00894(.A(new_n1270), .B(new_n1263), .Y(new_n1271));
  not_3  g00895(.A(new_n1271), .Y(new_n1272));
  xnor_3 g00896(.A(new_n1272), .B(new_n1262), .Y(new_n1273));
  not_3  g00897(.A(new_n1165), .Y(new_n1274));
  nor_4  g00898(.A(new_n1274), .B(new_n1156), .Y(new_n1275));
  not_3  g00899(.A(new_n1275), .Y(new_n1276));
  nor_4  g00900(.A(new_n1276), .B(new_n1273), .Y(new_n1277));
  not_3  g00901(.A(new_n1273), .Y(new_n1278));
  nor_4  g00902(.A(new_n1275), .B(new_n1278), .Y(new_n1279));
  nor_4  g00903(.A(new_n1279), .B(new_n1277), .Y(new_n1280));
  xnor_3 g00904(.A(new_n1280), .B(new_n1258), .Y(new_n1281));
  not_3  g00905(.A(new_n1281), .Y(new_n1282));
  nor_4  g00906(.A(new_n1169), .B(new_n1154), .Y(new_n1283));
  nor_4  g00907(.A(new_n1186), .B(new_n1283), .Y(new_n1284));
  not_3  g00908(.A(new_n1284), .Y(new_n1285));
  nor_4  g00909(.A(new_n1285), .B(new_n1282), .Y(new_n1286));
  nor_4  g00910(.A(new_n1284), .B(new_n1281), .Y(new_n1287));
  nor_4  g00911(.A(new_n1287), .B(new_n1286), .Y(new_n1288));
  xnor_3 g00912(.A(new_n1288), .B(new_n1234), .Y(new_n1289));
  xor_3  g00913(.A(new_n1289), .B(new_n1215), .Y(n381));
  nand_4 g00914(.A(n7862), .B(n6038), .Y(new_n1291));
  nand_4 g00915(.A(n7354), .B(n6877), .Y(new_n1292));
  nand_4 g00916(.A(n4805), .B(n1564), .Y(new_n1293));
  nand_4 g00917(.A(n8028), .B(n7236), .Y(new_n1294));
  not_3  g00918(.A(new_n1294), .Y(new_n1295));
  xor_3  g00919(.A(new_n1295), .B(new_n1293), .Y(new_n1296));
  xor_3  g00920(.A(new_n1296), .B(new_n1292), .Y(new_n1297));
  not_3  g00921(.A(new_n1297), .Y(new_n1298));
  xor_3  g00922(.A(new_n1298), .B(new_n1291), .Y(n397));
  nand_4 g00923(.A(n6687), .B(n4370), .Y(new_n1300));
  nand_4 g00924(.A(n11407), .B(n4189), .Y(new_n1301));
  nand_4 g00925(.A(n11877), .B(n6687), .Y(new_n1302));
  nand_4 g00926(.A(new_n1302), .B(new_n1301), .Y(new_n1303));
  not_3  g00927(.A(new_n1303), .Y(new_n1304));
  nor_4  g00928(.A(new_n1302), .B(new_n1301), .Y(new_n1305));
  nand_4 g00929(.A(n5212), .B(n2564), .Y(new_n1306));
  not_3  g00930(.A(new_n1306), .Y(new_n1307));
  nor_4  g00931(.A(new_n1307), .B(new_n1305), .Y(new_n1308));
  nor_4  g00932(.A(new_n1308), .B(new_n1304), .Y(new_n1309));
  xor_3  g00933(.A(new_n1309), .B(new_n1300), .Y(new_n1310));
  nand_4 g00934(.A(n5212), .B(n4189), .Y(new_n1311));
  not_3  g00935(.A(new_n1311), .Y(new_n1312));
  nand_4 g00936(.A(n11407), .B(n6770), .Y(new_n1313));
  nand_4 g00937(.A(n11877), .B(n2564), .Y(new_n1314));
  xnor_3 g00938(.A(new_n1314), .B(new_n1313), .Y(new_n1315));
  xor_3  g00939(.A(new_n1315), .B(new_n1312), .Y(new_n1316));
  xnor_3 g00940(.A(new_n1316), .B(new_n1310), .Y(new_n1317));
  not_3  g00941(.A(new_n1317), .Y(new_n1318));
  nand_4 g00942(.A(n11407), .B(n6687), .Y(new_n1319));
  not_3  g00943(.A(new_n1319), .Y(new_n1320));
  nor_4  g00944(.A(new_n1320), .B(new_n1306), .Y(new_n1321));
  nor_4  g00945(.A(new_n1321), .B(new_n1303), .Y(new_n1322));
  nor_4  g00946(.A(new_n1322), .B(new_n1305), .Y(new_n1323));
  nor_4  g00947(.A(new_n1323), .B(new_n1306), .Y(new_n1324));
  xor_3  g00948(.A(new_n1324), .B(new_n1318), .Y(new_n1325));
  not_3  g00949(.A(new_n1325), .Y(new_n1326));
  nand_4 g00950(.A(n12709), .B(n8336), .Y(new_n1327));
  nand_4 g00951(.A(n11222), .B(n10990), .Y(new_n1328));
  nand_4 g00952(.A(n12489), .B(n12069), .Y(new_n1329));
  xnor_3 g00953(.A(new_n1329), .B(new_n1328), .Y(new_n1330));
  nor_4  g00954(.A(new_n1330), .B(new_n1327), .Y(new_n1331));
  not_3  g00955(.A(new_n1331), .Y(new_n1332));
  nand_4 g00956(.A(n11728), .B(n8336), .Y(new_n1333_1));
  nand_4 g00957(.A(n12709), .B(n10928), .Y(new_n1334));
  not_3  g00958(.A(new_n1334), .Y(new_n1335));
  xor_3  g00959(.A(new_n1335), .B(new_n1333_1), .Y(new_n1336));
  nand_4 g00960(.A(new_n1336), .B(new_n1332), .Y(new_n1337));
  nor_4  g00961(.A(new_n1329), .B(new_n1328), .Y(new_n1338));
  not_3  g00962(.A(new_n1338), .Y(new_n1339));
  nand_4 g00963(.A(n11222), .B(n5760), .Y(new_n1340));
  nand_4 g00964(.A(n11153), .B(n10990), .Y(new_n1341));
  xnor_3 g00965(.A(new_n1341), .B(new_n1340), .Y(new_n1342));
  xnor_3 g00966(.A(new_n1342), .B(new_n1339), .Y(new_n1343));
  nand_4 g00967(.A(n12069), .B(n7159), .Y(new_n1344));
  nand_4 g00968(.A(n12489), .B(n12391), .Y(new_n1345));
  xor_3  g00969(.A(new_n1345), .B(new_n1344), .Y(new_n1346));
  not_3  g00970(.A(new_n1346), .Y(new_n1347));
  xnor_3 g00971(.A(new_n1347), .B(new_n1343), .Y(new_n1348));
  not_3  g00972(.A(new_n1337), .Y(new_n1349));
  nor_4  g00973(.A(new_n1336), .B(new_n1332), .Y(new_n1350));
  nor_4  g00974(.A(new_n1350), .B(new_n1349), .Y(new_n1351));
  nand_4 g00975(.A(new_n1351), .B(new_n1348), .Y(new_n1352));
  nand_4 g00976(.A(new_n1352), .B(new_n1337), .Y(new_n1353_1));
  not_3  g00977(.A(new_n1327), .Y(new_n1354));
  nand_4 g00978(.A(n11728), .B(n10928), .Y(new_n1355));
  nor_4  g00979(.A(new_n1355), .B(new_n1354), .Y(new_n1356));
  nand_4 g00980(.A(n12709), .B(n6986), .Y(new_n1357_1));
  not_3  g00981(.A(new_n1357_1), .Y(new_n1358));
  nand_4 g00982(.A(n8336), .B(n6429), .Y(new_n1359));
  not_3  g00983(.A(new_n1359), .Y(new_n1360));
  nor_4  g00984(.A(new_n1360), .B(new_n1358), .Y(new_n1361));
  nor_4  g00985(.A(new_n1359), .B(new_n1357_1), .Y(new_n1362));
  nor_4  g00986(.A(new_n1362), .B(new_n1361), .Y(new_n1363));
  nor_4  g00987(.A(new_n1363), .B(new_n1356), .Y(new_n1364));
  not_3  g00988(.A(new_n1364), .Y(new_n1365));
  not_3  g00989(.A(new_n1361), .Y(new_n1366));
  nand_4 g00990(.A(new_n1366), .B(new_n1356), .Y(new_n1367));
  nand_4 g00991(.A(new_n1367), .B(new_n1365), .Y(new_n1368));
  xnor_3 g00992(.A(new_n1368), .B(new_n1353_1), .Y(new_n1369));
  not_3  g00993(.A(new_n1329), .Y(new_n1370));
  nand_4 g00994(.A(n12391), .B(n7159), .Y(new_n1371));
  nor_4  g00995(.A(new_n1371), .B(new_n1370), .Y(new_n1372));
  nand_4 g00996(.A(n12489), .B(n7891), .Y(new_n1373));
  nand_4 g00997(.A(n12777), .B(n12069), .Y(new_n1374));
  nand_4 g00998(.A(new_n1374), .B(new_n1373), .Y(new_n1375));
  nor_4  g00999(.A(new_n1375), .B(new_n1372), .Y(new_n1376));
  nor_4  g01000(.A(new_n1374), .B(new_n1373), .Y(new_n1377));
  nor_4  g01001(.A(new_n1377), .B(new_n1376), .Y(new_n1378));
  nand_4 g01002(.A(new_n1375), .B(new_n1372), .Y(new_n1379));
  nand_4 g01003(.A(new_n1379), .B(new_n1378), .Y(new_n1380));
  nand_4 g01004(.A(n11153), .B(n5760), .Y(new_n1381));
  not_3  g01005(.A(new_n1381), .Y(new_n1382));
  nand_4 g01006(.A(new_n1382), .B(new_n1328), .Y(new_n1383));
  nand_4 g01007(.A(n10990), .B(n5314), .Y(new_n1384));
  not_3  g01008(.A(new_n1384), .Y(new_n1385));
  nand_4 g01009(.A(n11222), .B(n1478), .Y(new_n1386));
  not_3  g01010(.A(new_n1386), .Y(new_n1387));
  nand_4 g01011(.A(new_n1387), .B(new_n1385), .Y(new_n1388));
  nand_4 g01012(.A(new_n1386), .B(new_n1384), .Y(new_n1389));
  nand_4 g01013(.A(new_n1389), .B(new_n1388), .Y(new_n1390));
  nand_4 g01014(.A(new_n1390), .B(new_n1383), .Y(new_n1391));
  nand_4 g01015(.A(new_n1389), .B(new_n1382), .Y(new_n1392));
  not_3  g01016(.A(new_n1392), .Y(new_n1393));
  nand_4 g01017(.A(new_n1393), .B(new_n1328), .Y(new_n1394));
  nand_4 g01018(.A(new_n1394), .B(new_n1391), .Y(new_n1395));
  xnor_3 g01019(.A(new_n1395), .B(new_n1380), .Y(new_n1396));
  nor_4  g01020(.A(new_n1342), .B(new_n1339), .Y(new_n1397));
  nor_4  g01021(.A(new_n1347), .B(new_n1343), .Y(new_n1398));
  nor_4  g01022(.A(new_n1398), .B(new_n1397), .Y(new_n1399));
  nor_4  g01023(.A(new_n1399), .B(new_n1396), .Y(new_n1400));
  and_4  g01024(.A(new_n1399), .B(new_n1396), .Y(new_n1401));
  nor_4  g01025(.A(new_n1401), .B(new_n1400), .Y(new_n1402));
  xnor_3 g01026(.A(new_n1402), .B(new_n1369), .Y(new_n1403));
  not_3  g01027(.A(new_n1403), .Y(new_n1404));
  not_3  g01028(.A(new_n1323), .Y(new_n1405));
  not_3  g01029(.A(new_n1321), .Y(new_n1406));
  nor_4  g01030(.A(new_n1406), .B(new_n1304), .Y(new_n1407));
  nor_4  g01031(.A(new_n1407), .B(new_n1405), .Y(new_n1408));
  not_3  g01032(.A(new_n1408), .Y(new_n1409));
  nand_4 g01033(.A(new_n1409), .B(new_n1404), .Y(new_n1410));
  xnor_3 g01034(.A(new_n1409), .B(new_n1403), .Y(new_n1411));
  xor_3  g01035(.A(new_n1330), .B(new_n1327), .Y(new_n1412));
  nand_4 g01036(.A(new_n1412), .B(new_n1320), .Y(new_n1413));
  not_3  g01037(.A(new_n1413), .Y(new_n1414));
  nand_4 g01038(.A(n11407), .B(n2564), .Y(new_n1415));
  nand_4 g01039(.A(n6687), .B(n5212), .Y(new_n1416));
  xor_3  g01040(.A(new_n1416), .B(new_n1415), .Y(new_n1417));
  nor_4  g01041(.A(new_n1417), .B(new_n1414), .Y(new_n1418));
  not_3  g01042(.A(new_n1418), .Y(new_n1419));
  not_3  g01043(.A(new_n1348), .Y(new_n1420));
  xnor_3 g01044(.A(new_n1351), .B(new_n1420), .Y(new_n1421));
  xor_3  g01045(.A(new_n1417), .B(new_n1414), .Y(new_n1422));
  nand_4 g01046(.A(new_n1422), .B(new_n1421), .Y(new_n1423));
  nand_4 g01047(.A(new_n1423), .B(new_n1419), .Y(new_n1424));
  nand_4 g01048(.A(new_n1424), .B(new_n1411), .Y(new_n1425));
  nand_4 g01049(.A(new_n1425), .B(new_n1410), .Y(new_n1426));
  nor_4  g01050(.A(new_n1426), .B(new_n1326), .Y(new_n1427));
  not_3  g01051(.A(new_n1426), .Y(new_n1428));
  nor_4  g01052(.A(new_n1428), .B(new_n1325), .Y(new_n1429));
  nor_4  g01053(.A(new_n1429), .B(new_n1427), .Y(new_n1430));
  nand_4 g01054(.A(n8819), .B(n8336), .Y(new_n1431));
  nand_4 g01055(.A(n11728), .B(n6986), .Y(new_n1432));
  not_3  g01056(.A(new_n1432), .Y(new_n1433));
  nand_4 g01057(.A(n10928), .B(n6429), .Y(new_n1434));
  nand_4 g01058(.A(n12709), .B(n2226), .Y(new_n1435));
  xnor_3 g01059(.A(new_n1435), .B(new_n1434), .Y(new_n1436));
  xnor_3 g01060(.A(new_n1436), .B(new_n1433), .Y(new_n1437));
  not_3  g01061(.A(new_n1437), .Y(new_n1438));
  xor_3  g01062(.A(new_n1438), .B(new_n1431), .Y(new_n1439));
  not_3  g01063(.A(new_n1355), .Y(new_n1440));
  nor_4  g01064(.A(new_n1362), .B(new_n1440), .Y(new_n1441));
  nor_4  g01065(.A(new_n1441), .B(new_n1361), .Y(new_n1442));
  xnor_3 g01066(.A(new_n1442), .B(new_n1439), .Y(new_n1443));
  nor_4  g01067(.A(new_n1365), .B(new_n1355), .Y(new_n1444));
  xnor_3 g01068(.A(new_n1444), .B(new_n1443), .Y(new_n1445));
  nand_4 g01069(.A(n12069), .B(n6254), .Y(new_n1446));
  not_3  g01070(.A(new_n1446), .Y(new_n1447));
  not_3  g01071(.A(new_n1375), .Y(new_n1448));
  not_3  g01072(.A(new_n1371), .Y(new_n1449));
  nor_4  g01073(.A(new_n1377), .B(new_n1449), .Y(new_n1450));
  nor_4  g01074(.A(new_n1450), .B(new_n1448), .Y(new_n1451));
  xnor_3 g01075(.A(new_n1451), .B(new_n1447), .Y(new_n1452));
  nand_4 g01076(.A(n12489), .B(n7160), .Y(new_n1453));
  nand_4 g01077(.A(n12777), .B(n12391), .Y(new_n1454));
  not_3  g01078(.A(new_n1454), .Y(new_n1455));
  nand_4 g01079(.A(n7891), .B(n7159), .Y(new_n1456));
  not_3  g01080(.A(new_n1456), .Y(new_n1457));
  nor_4  g01081(.A(new_n1457), .B(new_n1455), .Y(new_n1458));
  nor_4  g01082(.A(new_n1456), .B(new_n1454), .Y(new_n1459));
  nor_4  g01083(.A(new_n1459), .B(new_n1458), .Y(new_n1460));
  xnor_3 g01084(.A(new_n1460), .B(new_n1453), .Y(new_n1461));
  not_3  g01085(.A(new_n1461), .Y(new_n1462));
  xnor_3 g01086(.A(new_n1462), .B(new_n1452), .Y(new_n1463));
  nor_4  g01087(.A(new_n1378), .B(new_n1371), .Y(new_n1464));
  not_3  g01088(.A(new_n1464), .Y(new_n1465));
  nor_4  g01089(.A(new_n1465), .B(new_n1463), .Y(new_n1466));
  not_3  g01090(.A(new_n1463), .Y(new_n1467));
  nor_4  g01091(.A(new_n1464), .B(new_n1467), .Y(new_n1468));
  nor_4  g01092(.A(new_n1468), .B(new_n1466), .Y(new_n1469));
  nand_4 g01093(.A(n11791), .B(n11222), .Y(new_n1470));
  nand_4 g01094(.A(new_n1392), .B(new_n1388), .Y(new_n1471_1));
  not_3  g01095(.A(new_n1471_1), .Y(new_n1472));
  xnor_3 g01096(.A(new_n1472), .B(new_n1470), .Y(new_n1473));
  nand_4 g01097(.A(n5760), .B(n5314), .Y(new_n1474));
  nand_4 g01098(.A(n10990), .B(n996), .Y(new_n1475));
  nand_4 g01099(.A(n11153), .B(n1478), .Y(new_n1476));
  xnor_3 g01100(.A(new_n1476), .B(new_n1475), .Y(new_n1477));
  xnor_3 g01101(.A(new_n1477), .B(new_n1474), .Y(new_n1478_1));
  xnor_3 g01102(.A(new_n1478_1), .B(new_n1473), .Y(new_n1479));
  nor_4  g01103(.A(new_n1391), .B(new_n1381), .Y(new_n1480));
  not_3  g01104(.A(new_n1480), .Y(new_n1481));
  nor_4  g01105(.A(new_n1481), .B(new_n1479), .Y(new_n1482));
  not_3  g01106(.A(new_n1479), .Y(new_n1483));
  nor_4  g01107(.A(new_n1480), .B(new_n1483), .Y(new_n1484));
  nor_4  g01108(.A(new_n1484), .B(new_n1482), .Y(new_n1485));
  xnor_3 g01109(.A(new_n1485), .B(new_n1469), .Y(new_n1486));
  nor_4  g01110(.A(new_n1395), .B(new_n1380), .Y(new_n1487));
  not_3  g01111(.A(new_n1487), .Y(new_n1488));
  not_3  g01112(.A(new_n1400), .Y(new_n1489));
  nand_4 g01113(.A(new_n1489), .B(new_n1488), .Y(new_n1490));
  xnor_3 g01114(.A(new_n1490), .B(new_n1486), .Y(new_n1491));
  xnor_3 g01115(.A(new_n1491), .B(new_n1445), .Y(new_n1492));
  nand_4 g01116(.A(new_n1368), .B(new_n1353_1), .Y(new_n1493));
  not_3  g01117(.A(new_n1493), .Y(new_n1494));
  nor_4  g01118(.A(new_n1402), .B(new_n1369), .Y(new_n1495));
  nor_4  g01119(.A(new_n1495), .B(new_n1494), .Y(new_n1496));
  not_3  g01120(.A(new_n1496), .Y(new_n1497));
  nor_4  g01121(.A(new_n1497), .B(new_n1492), .Y(new_n1498));
  not_3  g01122(.A(new_n1492), .Y(new_n1499));
  nor_4  g01123(.A(new_n1496), .B(new_n1499), .Y(new_n1500));
  nor_4  g01124(.A(new_n1500), .B(new_n1498), .Y(new_n1501));
  xor_3  g01125(.A(new_n1501), .B(new_n1430), .Y(n658));
  nand_4 g01126(.A(n7862), .B(n2585), .Y(new_n1503));
  not_3  g01127(.A(new_n1503), .Y(new_n1504));
  nand_4 g01128(.A(n2508), .B(n1333), .Y(new_n1505));
  not_3  g01129(.A(new_n1505), .Y(new_n1506));
  nand_4 g01130(.A(n11757), .B(n6038), .Y(new_n1507));
  not_3  g01131(.A(new_n1507), .Y(new_n1508));
  nand_4 g01132(.A(n12720), .B(n1333), .Y(new_n1509));
  not_3  g01133(.A(new_n1509), .Y(new_n1510_1));
  nor_4  g01134(.A(new_n1510_1), .B(new_n1508), .Y(new_n1511));
  nor_4  g01135(.A(new_n1509), .B(new_n1507), .Y(new_n1512_1));
  nand_4 g01136(.A(n3172), .B(n2509), .Y(new_n1513));
  not_3  g01137(.A(new_n1513), .Y(new_n1514));
  nor_4  g01138(.A(new_n1514), .B(new_n1512_1), .Y(new_n1515));
  nor_4  g01139(.A(new_n1515), .B(new_n1511), .Y(new_n1516));
  xnor_3 g01140(.A(new_n1516), .B(new_n1506), .Y(new_n1517));
  nand_4 g01141(.A(n11757), .B(n2509), .Y(new_n1518));
  nand_4 g01142(.A(n6038), .B(n5240), .Y(new_n1519));
  nand_4 g01143(.A(n12720), .B(n3172), .Y(new_n1520));
  xnor_3 g01144(.A(new_n1520), .B(new_n1519), .Y(new_n1521));
  xnor_3 g01145(.A(new_n1521), .B(new_n1518), .Y(new_n1522));
  xnor_3 g01146(.A(new_n1522), .B(new_n1517), .Y(new_n1523_1));
  not_3  g01147(.A(new_n1523_1), .Y(new_n1524));
  nor_4  g01148(.A(new_n1524), .B(new_n1504), .Y(new_n1525));
  not_3  g01149(.A(new_n1525), .Y(new_n1526));
  nor_4  g01150(.A(new_n1523_1), .B(new_n1503), .Y(new_n1527));
  nor_4  g01151(.A(new_n1527), .B(new_n1525), .Y(new_n1528));
  nand_4 g01152(.A(n7862), .B(n2508), .Y(new_n1529));
  nand_4 g01153(.A(n2509), .B(n1333), .Y(new_n1530));
  not_3  g01154(.A(new_n1530), .Y(new_n1531));
  nand_4 g01155(.A(n6038), .B(n3172), .Y(new_n1532));
  nand_4 g01156(.A(n12720), .B(n7862), .Y(new_n1533));
  nand_4 g01157(.A(new_n1533), .B(new_n1532), .Y(new_n1534));
  nand_4 g01158(.A(new_n1534), .B(new_n1531), .Y(new_n1535));
  not_3  g01159(.A(new_n1532), .Y(new_n1536));
  not_3  g01160(.A(new_n1533), .Y(new_n1537));
  nand_4 g01161(.A(new_n1537), .B(new_n1536), .Y(new_n1538));
  nand_4 g01162(.A(new_n1538), .B(new_n1535), .Y(new_n1539));
  not_3  g01163(.A(new_n1539), .Y(new_n1540));
  nor_4  g01164(.A(new_n1540), .B(new_n1529), .Y(new_n1541));
  xor_3  g01165(.A(new_n1539), .B(new_n1529), .Y(new_n1542));
  nor_4  g01166(.A(new_n1512_1), .B(new_n1511), .Y(new_n1543));
  xor_3  g01167(.A(new_n1543), .B(new_n1513), .Y(new_n1544));
  nor_4  g01168(.A(new_n1544), .B(new_n1542), .Y(new_n1545));
  nor_4  g01169(.A(new_n1545), .B(new_n1541), .Y(new_n1546));
  nand_4 g01170(.A(new_n1546), .B(new_n1528), .Y(new_n1547));
  nand_4 g01171(.A(new_n1547), .B(new_n1526), .Y(new_n1548));
  not_3  g01172(.A(new_n1548), .Y(new_n1549));
  nand_4 g01173(.A(n12720), .B(n11757), .Y(new_n1550));
  nand_4 g01174(.A(n5240), .B(n2509), .Y(new_n1551));
  nand_4 g01175(.A(n11821), .B(n6038), .Y(new_n1552));
  xnor_3 g01176(.A(new_n1552), .B(new_n1551), .Y(new_n1553));
  nor_4  g01177(.A(new_n1553), .B(new_n1550), .Y(new_n1554));
  not_3  g01178(.A(new_n1550), .Y(new_n1555));
  not_3  g01179(.A(new_n1553), .Y(new_n1556));
  nor_4  g01180(.A(new_n1556), .B(new_n1555), .Y(new_n1557));
  nor_4  g01181(.A(new_n1557), .B(new_n1554), .Y(new_n1558));
  not_3  g01182(.A(new_n1519), .Y(new_n1559));
  not_3  g01183(.A(new_n1520), .Y(new_n1560));
  nor_4  g01184(.A(new_n1560), .B(new_n1559), .Y(new_n1561));
  not_3  g01185(.A(new_n1518), .Y(new_n1562));
  nor_4  g01186(.A(new_n1521), .B(new_n1562), .Y(new_n1563));
  nor_4  g01187(.A(new_n1563), .B(new_n1561), .Y(new_n1564_1));
  xnor_3 g01188(.A(new_n1564_1), .B(new_n1558), .Y(new_n1565));
  not_3  g01189(.A(new_n1565), .Y(new_n1566));
  nand_4 g01190(.A(new_n1516), .B(new_n1506), .Y(new_n1567));
  not_3  g01191(.A(new_n1567), .Y(new_n1568));
  nor_4  g01192(.A(new_n1522), .B(new_n1517), .Y(new_n1569));
  nor_4  g01193(.A(new_n1569), .B(new_n1568), .Y(new_n1570));
  not_3  g01194(.A(new_n1570), .Y(new_n1571));
  nand_4 g01195(.A(n2585), .B(n1333), .Y(new_n1572));
  nand_4 g01196(.A(n3172), .B(n2508), .Y(new_n1573));
  xor_3  g01197(.A(new_n1573), .B(new_n1572), .Y(new_n1574));
  nor_4  g01198(.A(new_n1574), .B(new_n1571), .Y(new_n1575));
  not_3  g01199(.A(new_n1574), .Y(new_n1576_1));
  nor_4  g01200(.A(new_n1576_1), .B(new_n1570), .Y(new_n1577));
  nor_4  g01201(.A(new_n1577), .B(new_n1575), .Y(new_n1578));
  xnor_3 g01202(.A(new_n1578), .B(new_n1566), .Y(new_n1579));
  not_3  g01203(.A(new_n1579), .Y(new_n1580));
  nand_4 g01204(.A(new_n1580), .B(new_n1549), .Y(new_n1581));
  not_3  g01205(.A(new_n1577), .Y(new_n1582));
  nor_4  g01206(.A(new_n1573), .B(new_n1572), .Y(new_n1583));
  nor_4  g01207(.A(new_n1575), .B(new_n1565), .Y(new_n1584));
  xnor_3 g01208(.A(new_n1584), .B(new_n1583), .Y(new_n1585));
  nand_4 g01209(.A(new_n1585), .B(new_n1582), .Y(new_n1586));
  nor_4  g01210(.A(new_n1552), .B(new_n1551), .Y(new_n1587));
  nand_4 g01211(.A(n11757), .B(n2508), .Y(new_n1588));
  not_3  g01212(.A(new_n1588), .Y(new_n1589));
  xor_3  g01213(.A(new_n1589), .B(new_n1587), .Y(new_n1590));
  nand_4 g01214(.A(n11821), .B(n2509), .Y(new_n1591));
  not_3  g01215(.A(new_n1591), .Y(new_n1592));
  nand_4 g01216(.A(n12720), .B(n5240), .Y(new_n1593));
  nand_4 g01217(.A(n9080), .B(n6038), .Y(new_n1594));
  xnor_3 g01218(.A(new_n1594), .B(new_n1593), .Y(new_n1595));
  xnor_3 g01219(.A(new_n1595), .B(new_n1592), .Y(new_n1596));
  not_3  g01220(.A(new_n1596), .Y(new_n1597));
  xnor_3 g01221(.A(new_n1597), .B(new_n1590), .Y(new_n1598));
  not_3  g01222(.A(new_n1554), .Y(new_n1599));
  nand_4 g01223(.A(new_n1564_1), .B(new_n1558), .Y(new_n1600));
  nand_4 g01224(.A(new_n1600), .B(new_n1599), .Y(new_n1601));
  nand_4 g01225(.A(n4005), .B(n1333), .Y(new_n1602));
  nand_4 g01226(.A(n3172), .B(n2585), .Y(new_n1603));
  nand_4 g01227(.A(n12706), .B(n7862), .Y(new_n1604));
  nand_4 g01228(.A(new_n1604), .B(new_n1603), .Y(new_n1605));
  not_3  g01229(.A(new_n1603), .Y(new_n1606));
  not_3  g01230(.A(new_n1604), .Y(new_n1607));
  nand_4 g01231(.A(new_n1607), .B(new_n1606), .Y(new_n1608));
  nand_4 g01232(.A(new_n1608), .B(new_n1605), .Y(new_n1609));
  xor_3  g01233(.A(new_n1609), .B(new_n1602), .Y(new_n1610));
  xnor_3 g01234(.A(new_n1610), .B(new_n1601), .Y(new_n1611));
  xnor_3 g01235(.A(new_n1611), .B(new_n1598), .Y(new_n1612));
  not_3  g01236(.A(new_n1612), .Y(new_n1613));
  xnor_3 g01237(.A(new_n1613), .B(new_n1586), .Y(new_n1614));
  xnor_3 g01238(.A(new_n1614), .B(new_n1581), .Y(new_n1615));
  nand_4 g01239(.A(n7862), .B(n4005), .Y(new_n1616));
  not_3  g01240(.A(new_n1616), .Y(new_n1617));
  xnor_3 g01241(.A(new_n1579), .B(new_n1548), .Y(new_n1618));
  not_3  g01242(.A(new_n1618), .Y(new_n1619));
  nand_4 g01243(.A(new_n1619), .B(new_n1617), .Y(new_n1620));
  and_4  g01244(.A(new_n1538), .B(new_n1534), .Y(new_n1621));
  nand_4 g01245(.A(n6038), .B(n1333), .Y(new_n1622));
  nand_4 g01246(.A(n7862), .B(n2509), .Y(new_n1623));
  nor_4  g01247(.A(new_n1623), .B(new_n1622), .Y(new_n1624));
  not_3  g01248(.A(new_n1624), .Y(new_n1625));
  nor_4  g01249(.A(new_n1625), .B(new_n1621), .Y(new_n1626));
  not_3  g01250(.A(new_n1542), .Y(new_n1627));
  not_3  g01251(.A(new_n1544), .Y(new_n1628));
  xor_3  g01252(.A(new_n1628), .B(new_n1627), .Y(new_n1629));
  nand_4 g01253(.A(new_n1629), .B(new_n1626), .Y(new_n1630));
  not_3  g01254(.A(new_n1547), .Y(new_n1631));
  nor_4  g01255(.A(new_n1546), .B(new_n1528), .Y(new_n1632));
  nor_4  g01256(.A(new_n1632), .B(new_n1631), .Y(new_n1633));
  nor_4  g01257(.A(new_n1633), .B(new_n1630), .Y(new_n1634));
  nor_4  g01258(.A(new_n1618), .B(new_n1616), .Y(new_n1635));
  nor_4  g01259(.A(new_n1619), .B(new_n1617), .Y(new_n1636));
  nor_4  g01260(.A(new_n1636), .B(new_n1635), .Y(new_n1637));
  nand_4 g01261(.A(new_n1637), .B(new_n1634), .Y(new_n1638));
  nand_4 g01262(.A(new_n1638), .B(new_n1620), .Y(new_n1639));
  xnor_3 g01263(.A(new_n1639), .B(new_n1615), .Y(new_n1640));
  not_3  g01264(.A(new_n1640), .Y(new_n1641));
  nand_4 g01265(.A(n2464), .B(n1209), .Y(new_n1642));
  nor_4  g01266(.A(new_n1642), .B(new_n1292), .Y(new_n1643));
  nand_4 g01267(.A(n7354), .B(n2464), .Y(new_n1644));
  nand_4 g01268(.A(n6877), .B(n1209), .Y(new_n1645));
  nand_4 g01269(.A(new_n1645), .B(new_n1644), .Y(new_n1646));
  not_3  g01270(.A(new_n1646), .Y(new_n1647));
  nor_4  g01271(.A(new_n1647), .B(new_n1643), .Y(new_n1648));
  nand_4 g01272(.A(n9400), .B(n7354), .Y(new_n1649));
  nand_4 g01273(.A(n7500), .B(n6877), .Y(new_n1650));
  nor_4  g01274(.A(new_n1650), .B(new_n1649), .Y(new_n1651));
  not_3  g01275(.A(new_n1651), .Y(new_n1652));
  nor_4  g01276(.A(new_n1652), .B(new_n1648), .Y(new_n1653));
  not_3  g01277(.A(new_n1653), .Y(new_n1654));
  nand_4 g01278(.A(n6877), .B(n5105), .Y(new_n1655));
  not_3  g01279(.A(new_n1655), .Y(new_n1656));
  not_3  g01280(.A(new_n1643), .Y(new_n1657));
  nand_4 g01281(.A(n9400), .B(n7500), .Y(new_n1658_1));
  not_3  g01282(.A(new_n1658_1), .Y(new_n1659));
  nand_4 g01283(.A(new_n1659), .B(new_n1646), .Y(new_n1660));
  nand_4 g01284(.A(new_n1660), .B(new_n1657), .Y(new_n1661));
  nand_4 g01285(.A(new_n1661), .B(new_n1656), .Y(new_n1662));
  not_3  g01286(.A(new_n1662), .Y(new_n1663));
  nor_4  g01287(.A(new_n1661), .B(new_n1656), .Y(new_n1664));
  nor_4  g01288(.A(new_n1664), .B(new_n1663), .Y(new_n1665));
  nand_4 g01289(.A(n7500), .B(n2464), .Y(new_n1666));
  nand_4 g01290(.A(n9400), .B(n1209), .Y(new_n1667));
  not_3  g01291(.A(new_n1667), .Y(new_n1668));
  nand_4 g01292(.A(n11311), .B(n7354), .Y(new_n1669));
  not_3  g01293(.A(new_n1669), .Y(new_n1670));
  nor_4  g01294(.A(new_n1670), .B(new_n1668), .Y(new_n1671));
  nor_4  g01295(.A(new_n1669), .B(new_n1667), .Y(new_n1672));
  nor_4  g01296(.A(new_n1672), .B(new_n1671), .Y(new_n1673));
  xnor_3 g01297(.A(new_n1673), .B(new_n1666), .Y(new_n1674));
  xor_3  g01298(.A(new_n1674), .B(new_n1665), .Y(new_n1675));
  not_3  g01299(.A(new_n1675), .Y(new_n1676));
  nor_4  g01300(.A(new_n1676), .B(new_n1654), .Y(new_n1677));
  not_3  g01301(.A(new_n1677), .Y(new_n1678));
  nand_4 g01302(.A(n11311), .B(n7500), .Y(new_n1679));
  not_3  g01303(.A(new_n1679), .Y(new_n1680));
  nand_4 g01304(.A(n7354), .B(n4187), .Y(new_n1681));
  xnor_3 g01305(.A(new_n1681), .B(new_n1642), .Y(new_n1682));
  xnor_3 g01306(.A(new_n1682), .B(new_n1680), .Y(new_n1683));
  not_3  g01307(.A(new_n1683), .Y(new_n1684));
  nand_4 g01308(.A(n9400), .B(n5105), .Y(new_n1685));
  not_3  g01309(.A(new_n1666), .Y(new_n1686));
  nor_4  g01310(.A(new_n1672), .B(new_n1686), .Y(new_n1687));
  nor_4  g01311(.A(new_n1687), .B(new_n1671), .Y(new_n1688));
  xnor_3 g01312(.A(new_n1688), .B(new_n1685), .Y(new_n1689));
  xnor_3 g01313(.A(new_n1689), .B(new_n1684), .Y(new_n1690));
  nand_4 g01314(.A(n6877), .B(n4141), .Y(new_n1691));
  not_3  g01315(.A(new_n1691), .Y(new_n1692));
  nand_4 g01316(.A(new_n1674), .B(new_n1665), .Y(new_n1693));
  nand_4 g01317(.A(new_n1693), .B(new_n1662), .Y(new_n1694));
  xnor_3 g01318(.A(new_n1694), .B(new_n1692), .Y(new_n1695));
  xor_3  g01319(.A(new_n1695), .B(new_n1690), .Y(new_n1696));
  nor_4  g01320(.A(new_n1696), .B(new_n1678), .Y(new_n1697));
  not_3  g01321(.A(new_n1697), .Y(new_n1698));
  nand_4 g01322(.A(n6877), .B(n4928), .Y(new_n1699));
  nor_4  g01323(.A(new_n1694), .B(new_n1692), .Y(new_n1700));
  nor_4  g01324(.A(new_n1695), .B(new_n1690), .Y(new_n1701));
  nor_4  g01325(.A(new_n1701), .B(new_n1700), .Y(new_n1702));
  not_3  g01326(.A(new_n1702), .Y(new_n1703));
  nand_4 g01327(.A(n11311), .B(n1209), .Y(new_n1704));
  nand_4 g01328(.A(n7500), .B(n4187), .Y(new_n1705));
  nand_4 g01329(.A(n7354), .B(n4203), .Y(new_n1706));
  xnor_3 g01330(.A(new_n1706), .B(new_n1705), .Y(new_n1707));
  nor_4  g01331(.A(new_n1707), .B(new_n1704), .Y(new_n1708));
  not_3  g01332(.A(new_n1704), .Y(new_n1709));
  not_3  g01333(.A(new_n1707), .Y(new_n1710));
  nor_4  g01334(.A(new_n1710), .B(new_n1709), .Y(new_n1711));
  nor_4  g01335(.A(new_n1711), .B(new_n1708), .Y(new_n1712));
  and_4  g01336(.A(new_n1681), .B(new_n1642), .Y(new_n1713));
  nor_4  g01337(.A(new_n1682), .B(new_n1680), .Y(new_n1714));
  nor_4  g01338(.A(new_n1714), .B(new_n1713), .Y(new_n1715));
  xnor_3 g01339(.A(new_n1715), .B(new_n1712), .Y(new_n1716));
  not_3  g01340(.A(new_n1685), .Y(new_n1717));
  nand_4 g01341(.A(new_n1688), .B(new_n1717), .Y(new_n1718));
  nand_4 g01342(.A(new_n1689), .B(new_n1683), .Y(new_n1719));
  nand_4 g01343(.A(new_n1719), .B(new_n1718), .Y(new_n1720));
  nand_4 g01344(.A(n9400), .B(n4141), .Y(new_n1721));
  nand_4 g01345(.A(n5105), .B(n2464), .Y(new_n1722));
  xor_3  g01346(.A(new_n1722), .B(new_n1721), .Y(new_n1723));
  xnor_3 g01347(.A(new_n1723), .B(new_n1720), .Y(new_n1724));
  xnor_3 g01348(.A(new_n1724), .B(new_n1716), .Y(new_n1725));
  nor_4  g01349(.A(new_n1725), .B(new_n1703), .Y(new_n1726));
  not_3  g01350(.A(new_n1725), .Y(new_n1727));
  nor_4  g01351(.A(new_n1727), .B(new_n1702), .Y(new_n1728));
  nor_4  g01352(.A(new_n1728), .B(new_n1726), .Y(new_n1729));
  xnor_3 g01353(.A(new_n1729), .B(new_n1699), .Y(new_n1730));
  xnor_3 g01354(.A(new_n1730), .B(new_n1698), .Y(new_n1731));
  not_3  g01355(.A(new_n1731), .Y(new_n1732));
  nand_4 g01356(.A(n7294), .B(n7236), .Y(new_n1733));
  not_3  g01357(.A(new_n1733), .Y(new_n1734));
  nand_4 g01358(.A(n10848), .B(n3992), .Y(new_n1735));
  not_3  g01359(.A(new_n1735), .Y(new_n1736));
  nand_4 g01360(.A(n8384), .B(n8028), .Y(new_n1737));
  nand_4 g01361(.A(n7236), .B(n1980), .Y(new_n1738));
  nand_4 g01362(.A(new_n1738), .B(new_n1737), .Y(new_n1739));
  nand_4 g01363(.A(new_n1739), .B(new_n1736), .Y(new_n1740));
  not_3  g01364(.A(new_n1737), .Y(new_n1741));
  not_3  g01365(.A(new_n1738), .Y(new_n1742));
  nand_4 g01366(.A(new_n1742), .B(new_n1741), .Y(new_n1743));
  nand_4 g01367(.A(new_n1743), .B(new_n1740), .Y(new_n1744));
  nand_4 g01368(.A(new_n1744), .B(new_n1734), .Y(new_n1745));
  not_3  g01369(.A(new_n1745), .Y(new_n1746));
  nor_4  g01370(.A(new_n1744), .B(new_n1734), .Y(new_n1747));
  nor_4  g01371(.A(new_n1747), .B(new_n1746), .Y(new_n1748));
  nand_4 g01372(.A(n8028), .B(n6358), .Y(new_n1749));
  nand_4 g01373(.A(n3992), .B(n1980), .Y(new_n1750));
  nand_4 g01374(.A(n10848), .B(n8384), .Y(new_n1751));
  xnor_3 g01375(.A(new_n1751), .B(new_n1750), .Y(new_n1752));
  xnor_3 g01376(.A(new_n1752), .B(new_n1749), .Y(new_n1753));
  not_3  g01377(.A(new_n1753), .Y(new_n1754));
  xnor_3 g01378(.A(new_n1754), .B(new_n1748), .Y(new_n1755));
  nand_4 g01379(.A(new_n1743), .B(new_n1739), .Y(new_n1756));
  not_3  g01380(.A(new_n1756), .Y(new_n1757));
  nand_4 g01381(.A(n10848), .B(n7236), .Y(new_n1758));
  nand_4 g01382(.A(n8028), .B(n3992), .Y(new_n1759));
  nor_4  g01383(.A(new_n1759), .B(new_n1758), .Y(new_n1760));
  not_3  g01384(.A(new_n1760), .Y(new_n1761));
  nor_4  g01385(.A(new_n1761), .B(new_n1757), .Y(new_n1762));
  not_3  g01386(.A(new_n1762), .Y(new_n1763));
  nor_4  g01387(.A(new_n1763), .B(new_n1755), .Y(new_n1764));
  nand_4 g01388(.A(n10848), .B(n6358), .Y(new_n1765));
  not_3  g01389(.A(new_n1765), .Y(new_n1766));
  nand_4 g01390(.A(n8384), .B(n1980), .Y(new_n1767));
  nand_4 g01391(.A(n8028), .B(n5198), .Y(new_n1768));
  xnor_3 g01392(.A(new_n1768), .B(new_n1767), .Y(new_n1769));
  nor_4  g01393(.A(new_n1769), .B(new_n1766), .Y(new_n1770));
  not_3  g01394(.A(new_n1769), .Y(new_n1771));
  nor_4  g01395(.A(new_n1771), .B(new_n1765), .Y(new_n1772));
  nor_4  g01396(.A(new_n1772), .B(new_n1770), .Y(new_n1773));
  nand_4 g01397(.A(n7294), .B(n3992), .Y(new_n1774));
  not_3  g01398(.A(new_n1750), .Y(new_n1775));
  not_3  g01399(.A(new_n1751), .Y(new_n1776));
  nor_4  g01400(.A(new_n1776), .B(new_n1775), .Y(new_n1777));
  not_3  g01401(.A(new_n1749), .Y(new_n1778));
  nor_4  g01402(.A(new_n1752), .B(new_n1778), .Y(new_n1779));
  nor_4  g01403(.A(new_n1779), .B(new_n1777), .Y(new_n1780));
  xnor_3 g01404(.A(new_n1780), .B(new_n1774), .Y(new_n1781));
  xnor_3 g01405(.A(new_n1781), .B(new_n1773), .Y(new_n1782));
  nand_4 g01406(.A(n12704), .B(n7236), .Y(new_n1783));
  not_3  g01407(.A(new_n1783), .Y(new_n1784));
  nand_4 g01408(.A(new_n1754), .B(new_n1748), .Y(new_n1785));
  nand_4 g01409(.A(new_n1785), .B(new_n1745), .Y(new_n1786));
  xnor_3 g01410(.A(new_n1786), .B(new_n1784), .Y(new_n1787));
  xnor_3 g01411(.A(new_n1787), .B(new_n1782), .Y(new_n1788));
  nand_4 g01412(.A(new_n1788), .B(new_n1764), .Y(new_n1789));
  nand_4 g01413(.A(n7236), .B(n5814), .Y(new_n1790));
  not_3  g01414(.A(new_n1790), .Y(new_n1791));
  not_3  g01415(.A(new_n1774), .Y(new_n1792));
  nand_4 g01416(.A(new_n1780), .B(new_n1792), .Y(new_n1793));
  not_3  g01417(.A(new_n1773), .Y(new_n1794));
  nand_4 g01418(.A(new_n1781), .B(new_n1794), .Y(new_n1795));
  nand_4 g01419(.A(new_n1795), .B(new_n1793), .Y(new_n1796));
  nand_4 g01420(.A(n8384), .B(n7294), .Y(new_n1797));
  nand_4 g01421(.A(n12704), .B(n3992), .Y(new_n1798_1));
  xor_3  g01422(.A(new_n1798_1), .B(new_n1797), .Y(new_n1799));
  xnor_3 g01423(.A(new_n1799), .B(new_n1796), .Y(new_n1800));
  nand_4 g01424(.A(n6358), .B(n1980), .Y(new_n1801));
  not_3  g01425(.A(new_n1767), .Y(new_n1802));
  not_3  g01426(.A(new_n1768), .Y(new_n1803));
  nor_4  g01427(.A(new_n1803), .B(new_n1802), .Y(new_n1804));
  nor_4  g01428(.A(new_n1770), .B(new_n1804), .Y(new_n1805));
  xnor_3 g01429(.A(new_n1805), .B(new_n1801), .Y(new_n1806));
  nand_4 g01430(.A(n10848), .B(n5198), .Y(new_n1807));
  nand_4 g01431(.A(n8028), .B(n1471), .Y(new_n1808));
  xor_3  g01432(.A(new_n1808), .B(new_n1807), .Y(new_n1809));
  xnor_3 g01433(.A(new_n1809), .B(new_n1806), .Y(new_n1810));
  xnor_3 g01434(.A(new_n1810), .B(new_n1800), .Y(new_n1811));
  nor_4  g01435(.A(new_n1786), .B(new_n1784), .Y(new_n1812));
  nor_4  g01436(.A(new_n1787), .B(new_n1782), .Y(new_n1813));
  nor_4  g01437(.A(new_n1813), .B(new_n1812), .Y(new_n1814));
  xnor_3 g01438(.A(new_n1814), .B(new_n1811), .Y(new_n1815));
  xnor_3 g01439(.A(new_n1815), .B(new_n1791), .Y(new_n1816));
  nor_4  g01440(.A(new_n1816), .B(new_n1789), .Y(new_n1817));
  not_3  g01441(.A(new_n1789), .Y(new_n1818));
  not_3  g01442(.A(new_n1816), .Y(new_n1819));
  nor_4  g01443(.A(new_n1819), .B(new_n1818), .Y(new_n1820));
  nor_4  g01444(.A(new_n1820), .B(new_n1817), .Y(new_n1821));
  nand_4 g01445(.A(n4805), .B(n533), .Y(new_n1822));
  nand_4 g01446(.A(n5283), .B(n1564), .Y(new_n1823));
  nand_4 g01447(.A(new_n1823), .B(new_n1822), .Y(new_n1824));
  nor_4  g01448(.A(new_n1823), .B(new_n1822), .Y(new_n1825));
  not_3  g01449(.A(new_n1825), .Y(new_n1826));
  nand_4 g01450(.A(new_n1826), .B(new_n1824), .Y(new_n1827));
  not_3  g01451(.A(new_n1827), .Y(new_n1828));
  nand_4 g01452(.A(n11478), .B(n1564), .Y(new_n1829));
  nand_4 g01453(.A(n4805), .B(n1512), .Y(new_n1830));
  nor_4  g01454(.A(new_n1830), .B(new_n1829), .Y(new_n1831));
  not_3  g01455(.A(new_n1831), .Y(new_n1832));
  nor_4  g01456(.A(new_n1832), .B(new_n1828), .Y(new_n1833));
  not_3  g01457(.A(new_n1833), .Y(new_n1834));
  nand_4 g01458(.A(n4805), .B(n2802), .Y(new_n1835_1));
  nand_4 g01459(.A(n11478), .B(n1512), .Y(new_n1836));
  not_3  g01460(.A(new_n1836), .Y(new_n1837));
  nand_4 g01461(.A(new_n1837), .B(new_n1824), .Y(new_n1838));
  nand_4 g01462(.A(new_n1838), .B(new_n1826), .Y(new_n1839));
  not_3  g01463(.A(new_n1839), .Y(new_n1840));
  xnor_3 g01464(.A(new_n1840), .B(new_n1835_1), .Y(new_n1841));
  nand_4 g01465(.A(n1564), .B(n137), .Y(new_n1842));
  nand_4 g01466(.A(n5283), .B(n1512), .Y(new_n1843));
  nand_4 g01467(.A(n11478), .B(n533), .Y(new_n1844));
  xnor_3 g01468(.A(new_n1844), .B(new_n1843), .Y(new_n1845));
  xnor_3 g01469(.A(new_n1845), .B(new_n1842), .Y(new_n1846));
  xnor_3 g01470(.A(new_n1846), .B(new_n1841), .Y(new_n1847_1));
  nor_4  g01471(.A(new_n1847_1), .B(new_n1834), .Y(new_n1848));
  not_3  g01472(.A(new_n1848), .Y(new_n1849));
  nand_4 g01473(.A(n6806), .B(n4805), .Y(new_n1850));
  nand_4 g01474(.A(n11478), .B(n2802), .Y(new_n1851));
  not_3  g01475(.A(new_n1851), .Y(new_n1852));
  not_3  g01476(.A(new_n1843), .Y(new_n1853));
  not_3  g01477(.A(new_n1844), .Y(new_n1854));
  nor_4  g01478(.A(new_n1854), .B(new_n1853), .Y(new_n1855));
  not_3  g01479(.A(new_n1842), .Y(new_n1856));
  nor_4  g01480(.A(new_n1845), .B(new_n1856), .Y(new_n1857));
  nor_4  g01481(.A(new_n1857), .B(new_n1855), .Y(new_n1858));
  xnor_3 g01482(.A(new_n1858), .B(new_n1852), .Y(new_n1859));
  nand_4 g01483(.A(n1512), .B(n137), .Y(new_n1860));
  nand_4 g01484(.A(n5283), .B(n533), .Y(new_n1861));
  nand_4 g01485(.A(n6294), .B(n1564), .Y(new_n1862));
  xnor_3 g01486(.A(new_n1862), .B(new_n1861), .Y(new_n1863));
  xnor_3 g01487(.A(new_n1863), .B(new_n1860), .Y(new_n1864));
  xnor_3 g01488(.A(new_n1864), .B(new_n1859), .Y(new_n1865));
  nand_4 g01489(.A(new_n1865), .B(new_n1850), .Y(new_n1866));
  not_3  g01490(.A(new_n1866), .Y(new_n1867));
  nor_4  g01491(.A(new_n1865), .B(new_n1850), .Y(new_n1868));
  nor_4  g01492(.A(new_n1868), .B(new_n1867), .Y(new_n1869));
  nor_4  g01493(.A(new_n1840), .B(new_n1835_1), .Y(new_n1870));
  nor_4  g01494(.A(new_n1846), .B(new_n1841), .Y(new_n1871));
  nor_4  g01495(.A(new_n1871), .B(new_n1870), .Y(new_n1872));
  nand_4 g01496(.A(new_n1872), .B(new_n1869), .Y(new_n1873));
  not_3  g01497(.A(new_n1873), .Y(new_n1874));
  nor_4  g01498(.A(new_n1872), .B(new_n1869), .Y(new_n1875));
  nor_4  g01499(.A(new_n1875), .B(new_n1874), .Y(new_n1876));
  nor_4  g01500(.A(new_n1876), .B(new_n1849), .Y(new_n1877));
  nand_4 g01501(.A(n5069), .B(n4805), .Y(new_n1878));
  nand_4 g01502(.A(n533), .B(n137), .Y(new_n1879));
  nand_4 g01503(.A(n6294), .B(n1512), .Y(new_n1880));
  nand_4 g01504(.A(n6797), .B(n1564), .Y(new_n1881));
  xnor_3 g01505(.A(new_n1881), .B(new_n1880), .Y(new_n1882));
  nor_4  g01506(.A(new_n1882), .B(new_n1879), .Y(new_n1883));
  not_3  g01507(.A(new_n1879), .Y(new_n1884));
  not_3  g01508(.A(new_n1882), .Y(new_n1885));
  nor_4  g01509(.A(new_n1885), .B(new_n1884), .Y(new_n1886));
  nor_4  g01510(.A(new_n1886), .B(new_n1883), .Y(new_n1887));
  and_4  g01511(.A(new_n1862), .B(new_n1861), .Y(new_n1888));
  not_3  g01512(.A(new_n1860), .Y(new_n1889));
  nor_4  g01513(.A(new_n1863), .B(new_n1889), .Y(new_n1890));
  nor_4  g01514(.A(new_n1890), .B(new_n1888), .Y(new_n1891));
  xnor_3 g01515(.A(new_n1891), .B(new_n1887), .Y(new_n1892));
  not_3  g01516(.A(new_n1892), .Y(new_n1893));
  nand_4 g01517(.A(n11478), .B(n6806), .Y(new_n1894));
  nand_4 g01518(.A(n5283), .B(n2802), .Y(new_n1895));
  xor_3  g01519(.A(new_n1895), .B(new_n1894), .Y(new_n1896));
  xnor_3 g01520(.A(new_n1896), .B(new_n1893), .Y(new_n1897));
  nand_4 g01521(.A(new_n1858), .B(new_n1852), .Y(new_n1898));
  not_3  g01522(.A(new_n1898), .Y(new_n1899));
  nor_4  g01523(.A(new_n1864), .B(new_n1859), .Y(new_n1900));
  nor_4  g01524(.A(new_n1900), .B(new_n1899), .Y(new_n1901));
  xnor_3 g01525(.A(new_n1901), .B(new_n1897), .Y(new_n1902));
  nand_4 g01526(.A(new_n1873), .B(new_n1866), .Y(new_n1903));
  xnor_3 g01527(.A(new_n1903), .B(new_n1902), .Y(new_n1904));
  nor_4  g01528(.A(new_n1904), .B(new_n1878), .Y(new_n1905));
  not_3  g01529(.A(new_n1878), .Y(new_n1906_1));
  not_3  g01530(.A(new_n1904), .Y(new_n1907));
  nor_4  g01531(.A(new_n1907), .B(new_n1906_1), .Y(new_n1908));
  nor_4  g01532(.A(new_n1908), .B(new_n1905), .Y(new_n1909));
  xnor_3 g01533(.A(new_n1909), .B(new_n1877), .Y(new_n1910));
  xnor_3 g01534(.A(new_n1910), .B(new_n1821), .Y(new_n1911));
  nor_4  g01535(.A(new_n1788), .B(new_n1764), .Y(new_n1912));
  nor_4  g01536(.A(new_n1912), .B(new_n1818), .Y(new_n1913));
  xnor_3 g01537(.A(new_n1847_1), .B(new_n1834), .Y(new_n1914));
  not_3  g01538(.A(new_n1914), .Y(new_n1915));
  not_3  g01539(.A(new_n1755), .Y(new_n1916));
  nor_4  g01540(.A(new_n1762), .B(new_n1916), .Y(new_n1917));
  nor_4  g01541(.A(new_n1917), .B(new_n1764), .Y(new_n1918));
  nor_4  g01542(.A(new_n1918), .B(new_n1915), .Y(new_n1919));
  nor_4  g01543(.A(new_n1294), .B(new_n1293), .Y(new_n1920));
  xnor_3 g01544(.A(new_n1830), .B(new_n1829), .Y(new_n1921));
  not_3  g01545(.A(new_n1921), .Y(new_n1922));
  nor_4  g01546(.A(new_n1922), .B(new_n1920), .Y(new_n1923));
  not_3  g01547(.A(new_n1923), .Y(new_n1924));
  not_3  g01548(.A(new_n1920), .Y(new_n1925));
  nor_4  g01549(.A(new_n1921), .B(new_n1925), .Y(new_n1926));
  nor_4  g01550(.A(new_n1926), .B(new_n1923), .Y(new_n1927));
  not_3  g01551(.A(new_n1759), .Y(new_n1928));
  xor_3  g01552(.A(new_n1928), .B(new_n1758), .Y(new_n1929));
  nand_4 g01553(.A(new_n1929), .B(new_n1927), .Y(new_n1930));
  nand_4 g01554(.A(new_n1930), .B(new_n1924), .Y(new_n1931));
  not_3  g01555(.A(new_n1293), .Y(new_n1932));
  nor_4  g01556(.A(new_n1836), .B(new_n1932), .Y(new_n1933));
  nor_4  g01557(.A(new_n1933), .B(new_n1828), .Y(new_n1934));
  nor_4  g01558(.A(new_n1838), .B(new_n1932), .Y(new_n1935));
  nor_4  g01559(.A(new_n1935), .B(new_n1934), .Y(new_n1936));
  not_3  g01560(.A(new_n1936), .Y(new_n1937));
  nand_4 g01561(.A(new_n1937), .B(new_n1931), .Y(new_n1938));
  not_3  g01562(.A(new_n1938), .Y(new_n1939));
  xnor_3 g01563(.A(new_n1937), .B(new_n1931), .Y(new_n1940));
  nor_4  g01564(.A(new_n1735), .B(new_n1295), .Y(new_n1941));
  nor_4  g01565(.A(new_n1941), .B(new_n1757), .Y(new_n1942));
  nor_4  g01566(.A(new_n1740), .B(new_n1295), .Y(new_n1943));
  nor_4  g01567(.A(new_n1943), .B(new_n1942), .Y(new_n1944));
  nor_4  g01568(.A(new_n1944), .B(new_n1940), .Y(new_n1945));
  nor_4  g01569(.A(new_n1945), .B(new_n1939), .Y(new_n1946));
  not_3  g01570(.A(new_n1918), .Y(new_n1947));
  nor_4  g01571(.A(new_n1947), .B(new_n1914), .Y(new_n1948));
  nor_4  g01572(.A(new_n1948), .B(new_n1919), .Y(new_n1949));
  not_3  g01573(.A(new_n1949), .Y(new_n1950));
  nor_4  g01574(.A(new_n1950), .B(new_n1946), .Y(new_n1951));
  nor_4  g01575(.A(new_n1951), .B(new_n1919), .Y(new_n1952));
  nor_4  g01576(.A(new_n1952), .B(new_n1913), .Y(new_n1953));
  not_3  g01577(.A(new_n1876), .Y(new_n1954));
  nor_4  g01578(.A(new_n1954), .B(new_n1848), .Y(new_n1955));
  nor_4  g01579(.A(new_n1955), .B(new_n1877), .Y(new_n1956));
  not_3  g01580(.A(new_n1913), .Y(new_n1957));
  not_3  g01581(.A(new_n1919), .Y(new_n1958));
  nor_4  g01582(.A(new_n1937), .B(new_n1931), .Y(new_n1959));
  nor_4  g01583(.A(new_n1959), .B(new_n1939), .Y(new_n1960));
  not_3  g01584(.A(new_n1944), .Y(new_n1961));
  nand_4 g01585(.A(new_n1961), .B(new_n1960), .Y(new_n1962));
  nand_4 g01586(.A(new_n1962), .B(new_n1938), .Y(new_n1963));
  nand_4 g01587(.A(new_n1949), .B(new_n1963), .Y(new_n1964));
  nand_4 g01588(.A(new_n1964), .B(new_n1958), .Y(new_n1965));
  xnor_3 g01589(.A(new_n1965), .B(new_n1957), .Y(new_n1966));
  nor_4  g01590(.A(new_n1966), .B(new_n1956), .Y(new_n1967));
  nor_4  g01591(.A(new_n1967), .B(new_n1953), .Y(new_n1968));
  xnor_3 g01592(.A(new_n1968), .B(new_n1911), .Y(new_n1969));
  nand_4 g01593(.A(new_n1969), .B(new_n1732), .Y(new_n1970));
  xnor_3 g01594(.A(new_n1969), .B(new_n1731), .Y(new_n1971));
  not_3  g01595(.A(new_n1696), .Y(new_n1972));
  nor_4  g01596(.A(new_n1972), .B(new_n1677), .Y(new_n1973));
  nor_4  g01597(.A(new_n1973), .B(new_n1697), .Y(new_n1974));
  not_3  g01598(.A(new_n1974), .Y(new_n1975));
  not_3  g01599(.A(new_n1956), .Y(new_n1976));
  xnor_3 g01600(.A(new_n1966), .B(new_n1976), .Y(new_n1977));
  nor_4  g01601(.A(new_n1977), .B(new_n1975), .Y(new_n1978));
  xnor_3 g01602(.A(new_n1966), .B(new_n1956), .Y(new_n1979));
  xnor_3 g01603(.A(new_n1979), .B(new_n1974), .Y(new_n1980_1));
  xor_3  g01604(.A(new_n1676), .B(new_n1654), .Y(new_n1981));
  not_3  g01605(.A(new_n1981), .Y(new_n1982));
  nor_4  g01606(.A(new_n1949), .B(new_n1963), .Y(new_n1983));
  nor_4  g01607(.A(new_n1983), .B(new_n1951), .Y(new_n1984));
  nor_4  g01608(.A(new_n1984), .B(new_n1982), .Y(new_n1985));
  xnor_3 g01609(.A(new_n1984), .B(new_n1982), .Y(new_n1986));
  xnor_3 g01610(.A(new_n1944), .B(new_n1940), .Y(new_n1987));
  not_3  g01611(.A(new_n1987), .Y(new_n1988));
  not_3  g01612(.A(new_n1292), .Y(new_n1989));
  nor_4  g01613(.A(new_n1658_1), .B(new_n1989), .Y(new_n1990));
  nor_4  g01614(.A(new_n1990), .B(new_n1648), .Y(new_n1991));
  nor_4  g01615(.A(new_n1660), .B(new_n1989), .Y(new_n1992));
  nor_4  g01616(.A(new_n1992), .B(new_n1991), .Y(new_n1993));
  not_3  g01617(.A(new_n1993), .Y(new_n1994));
  nor_4  g01618(.A(new_n1994), .B(new_n1988), .Y(new_n1995));
  xor_3  g01619(.A(new_n1994), .B(new_n1988), .Y(new_n1996));
  not_3  g01620(.A(new_n1996), .Y(new_n1997));
  xnor_3 g01621(.A(new_n1929), .B(new_n1927), .Y(new_n1998));
  not_3  g01622(.A(new_n1998), .Y(new_n1999));
  xor_3  g01623(.A(new_n1650), .B(new_n1649), .Y(new_n2000));
  not_3  g01624(.A(new_n2000), .Y(new_n2001));
  nor_4  g01625(.A(new_n2001), .B(new_n1999), .Y(new_n2002));
  nor_4  g01626(.A(new_n1296), .B(new_n1292), .Y(new_n2003));
  not_3  g01627(.A(new_n2003), .Y(new_n2004));
  xor_3  g01628(.A(new_n2000), .B(new_n1999), .Y(new_n2005));
  nor_4  g01629(.A(new_n2005), .B(new_n2004), .Y(new_n2006));
  nor_4  g01630(.A(new_n2006), .B(new_n2002), .Y(new_n2007));
  nor_4  g01631(.A(new_n2007), .B(new_n1997), .Y(new_n2008));
  nor_4  g01632(.A(new_n2008), .B(new_n1995), .Y(new_n2009));
  nor_4  g01633(.A(new_n2009), .B(new_n1986), .Y(new_n2010));
  nor_4  g01634(.A(new_n2010), .B(new_n1985), .Y(new_n2011));
  nor_4  g01635(.A(new_n2011), .B(new_n1980_1), .Y(new_n2012));
  nor_4  g01636(.A(new_n2012), .B(new_n1978), .Y(new_n2013));
  nand_4 g01637(.A(new_n2013), .B(new_n1971), .Y(new_n2014));
  nand_4 g01638(.A(new_n2014), .B(new_n1970), .Y(new_n2015));
  not_3  g01639(.A(new_n1726), .Y(new_n2016));
  nand_4 g01640(.A(new_n1715), .B(new_n1712), .Y(new_n2017));
  not_3  g01641(.A(new_n2017), .Y(new_n2018));
  nor_4  g01642(.A(new_n2018), .B(new_n1708), .Y(new_n2019));
  not_3  g01643(.A(new_n2019), .Y(new_n2020));
  nand_4 g01644(.A(n9400), .B(n4928), .Y(new_n2021));
  not_3  g01645(.A(new_n2021), .Y(new_n2022));
  nand_4 g01646(.A(n4141), .B(n2464), .Y(new_n2023));
  nand_4 g01647(.A(n8236), .B(n6877), .Y(new_n2024_1));
  nand_4 g01648(.A(new_n2024_1), .B(new_n2023), .Y(new_n2025));
  not_3  g01649(.A(new_n2023), .Y(new_n2026));
  not_3  g01650(.A(new_n2024_1), .Y(new_n2027));
  nand_4 g01651(.A(new_n2027), .B(new_n2026), .Y(new_n2028));
  nand_4 g01652(.A(new_n2028), .B(new_n2025), .Y(new_n2029));
  xor_3  g01653(.A(new_n2029), .B(new_n2022), .Y(new_n2030));
  xnor_3 g01654(.A(new_n2030), .B(new_n2020), .Y(new_n2031));
  nor_4  g01655(.A(new_n1706), .B(new_n1705), .Y(new_n2032));
  nand_4 g01656(.A(n11311), .B(n5105), .Y(new_n2033));
  xnor_3 g01657(.A(new_n2033), .B(new_n2032), .Y(new_n2034));
  nand_4 g01658(.A(n7500), .B(n4203), .Y(new_n2035));
  not_3  g01659(.A(new_n2035), .Y(new_n2036));
  nand_4 g01660(.A(n4187), .B(n1209), .Y(new_n2037));
  nand_4 g01661(.A(n12753), .B(n7354), .Y(new_n2038));
  xnor_3 g01662(.A(new_n2038), .B(new_n2037), .Y(new_n2039));
  xnor_3 g01663(.A(new_n2039), .B(new_n2036), .Y(new_n2040));
  not_3  g01664(.A(new_n2040), .Y(new_n2041));
  xor_3  g01665(.A(new_n2041), .B(new_n2034), .Y(new_n2042));
  xnor_3 g01666(.A(new_n2042), .B(new_n2031), .Y(new_n2043));
  not_3  g01667(.A(new_n2043), .Y(new_n2044));
  nand_4 g01668(.A(new_n1723), .B(new_n1720), .Y(new_n2045));
  nor_4  g01669(.A(new_n1722), .B(new_n1721), .Y(new_n2046));
  nor_4  g01670(.A(new_n1723), .B(new_n1720), .Y(new_n2047));
  nor_4  g01671(.A(new_n2047), .B(new_n1716), .Y(new_n2048));
  xnor_3 g01672(.A(new_n2048), .B(new_n2046), .Y(new_n2049));
  nand_4 g01673(.A(new_n2049), .B(new_n2045), .Y(new_n2050));
  xnor_3 g01674(.A(new_n2050), .B(new_n2044), .Y(new_n2051));
  xnor_3 g01675(.A(new_n2051), .B(new_n2016), .Y(new_n2052));
  not_3  g01676(.A(new_n1699), .Y(new_n2053));
  nand_4 g01677(.A(new_n1729), .B(new_n2053), .Y(new_n2054));
  nand_4 g01678(.A(new_n1730), .B(new_n1697), .Y(new_n2055));
  nand_4 g01679(.A(new_n2055), .B(new_n2054), .Y(new_n2056));
  xnor_3 g01680(.A(new_n2056), .B(new_n2052), .Y(new_n2057));
  not_3  g01681(.A(new_n2057), .Y(new_n2058));
  not_3  g01682(.A(new_n1811), .Y(new_n2059));
  nand_4 g01683(.A(new_n1814), .B(new_n2059), .Y(new_n2060));
  not_3  g01684(.A(new_n1805), .Y(new_n2061));
  nand_4 g01685(.A(new_n2061), .B(new_n1801), .Y(new_n2062));
  not_3  g01686(.A(new_n1809), .Y(new_n2063));
  nand_4 g01687(.A(new_n2063), .B(new_n1806), .Y(new_n2064));
  nand_4 g01688(.A(new_n2064), .B(new_n2062), .Y(new_n2065));
  nand_4 g01689(.A(n5814), .B(n3992), .Y(new_n2066));
  not_3  g01690(.A(new_n2066), .Y(new_n2067));
  nand_4 g01691(.A(n12704), .B(n8384), .Y(new_n2068));
  nand_4 g01692(.A(n7236), .B(n4903), .Y(new_n2069));
  xnor_3 g01693(.A(new_n2069), .B(new_n2068), .Y(new_n2070));
  xor_3  g01694(.A(new_n2070), .B(new_n2067), .Y(new_n2071));
  not_3  g01695(.A(new_n2071), .Y(new_n2072));
  xnor_3 g01696(.A(new_n2072), .B(new_n2065), .Y(new_n2073));
  nor_4  g01697(.A(new_n1808), .B(new_n1807), .Y(new_n2074));
  nand_4 g01698(.A(n7294), .B(n6358), .Y(new_n2075));
  not_3  g01699(.A(new_n2075), .Y(new_n2076));
  xor_3  g01700(.A(new_n2076), .B(new_n2074), .Y(new_n2077));
  nand_4 g01701(.A(n10848), .B(n1471), .Y(new_n2078));
  nand_4 g01702(.A(n5198), .B(n1980), .Y(new_n2079));
  nand_4 g01703(.A(n8028), .B(n7646), .Y(new_n2080));
  not_3  g01704(.A(new_n2080), .Y(new_n2081));
  xor_3  g01705(.A(new_n2081), .B(new_n2079), .Y(new_n2082));
  xnor_3 g01706(.A(new_n2082), .B(new_n2078), .Y(new_n2083));
  not_3  g01707(.A(new_n2083), .Y(new_n2084));
  xnor_3 g01708(.A(new_n2084), .B(new_n2077), .Y(new_n2085));
  xnor_3 g01709(.A(new_n2085), .B(new_n2073), .Y(new_n2086));
  nand_4 g01710(.A(new_n1799), .B(new_n1796), .Y(new_n2087_1));
  nor_4  g01711(.A(new_n1798_1), .B(new_n1797), .Y(new_n2088));
  nor_4  g01712(.A(new_n1810), .B(new_n1800), .Y(new_n2089));
  xnor_3 g01713(.A(new_n2089), .B(new_n2088), .Y(new_n2090));
  nand_4 g01714(.A(new_n2090), .B(new_n2087_1), .Y(new_n2091));
  xnor_3 g01715(.A(new_n2091), .B(new_n2086), .Y(new_n2092));
  xnor_3 g01716(.A(new_n2092), .B(new_n2060), .Y(new_n2093));
  nand_4 g01717(.A(new_n1815), .B(new_n1791), .Y(new_n2094));
  not_3  g01718(.A(new_n2094), .Y(new_n2095));
  nor_4  g01719(.A(new_n1817), .B(new_n2095), .Y(new_n2096_1));
  xnor_3 g01720(.A(new_n2096_1), .B(new_n2093), .Y(new_n2097));
  not_3  g01721(.A(new_n1905), .Y(new_n2098));
  nand_4 g01722(.A(new_n1909), .B(new_n1877), .Y(new_n2099));
  nand_4 g01723(.A(new_n2099), .B(new_n2098), .Y(new_n2100));
  nor_4  g01724(.A(new_n1903), .B(new_n1902), .Y(new_n2101));
  not_3  g01725(.A(new_n2101), .Y(new_n2102));
  not_3  g01726(.A(new_n1883), .Y(new_n2103));
  nand_4 g01727(.A(new_n1891), .B(new_n1887), .Y(new_n2104));
  nand_4 g01728(.A(new_n2104), .B(new_n2103), .Y(new_n2105));
  nand_4 g01729(.A(n11478), .B(n5069), .Y(new_n2106));
  not_3  g01730(.A(new_n2106), .Y(new_n2107));
  nand_4 g01731(.A(n6806), .B(n5283), .Y(new_n2108));
  nand_4 g01732(.A(n12044), .B(n4805), .Y(new_n2109));
  nand_4 g01733(.A(new_n2109), .B(new_n2108), .Y(new_n2110));
  not_3  g01734(.A(new_n2108), .Y(new_n2111));
  not_3  g01735(.A(new_n2109), .Y(new_n2112));
  nand_4 g01736(.A(new_n2112), .B(new_n2111), .Y(new_n2113));
  nand_4 g01737(.A(new_n2113), .B(new_n2110), .Y(new_n2114));
  xor_3  g01738(.A(new_n2114), .B(new_n2107), .Y(new_n2115));
  xnor_3 g01739(.A(new_n2115), .B(new_n2105), .Y(new_n2116));
  nor_4  g01740(.A(new_n1881), .B(new_n1880), .Y(new_n2117));
  nand_4 g01741(.A(n2802), .B(n137), .Y(new_n2118));
  not_3  g01742(.A(new_n2118), .Y(new_n2119));
  xor_3  g01743(.A(new_n2119), .B(new_n2117), .Y(new_n2120));
  nand_4 g01744(.A(n6797), .B(n1512), .Y(new_n2121));
  not_3  g01745(.A(new_n2121), .Y(new_n2122));
  nand_4 g01746(.A(n6294), .B(n533), .Y(new_n2123));
  nand_4 g01747(.A(n3146), .B(n1564), .Y(new_n2124));
  xnor_3 g01748(.A(new_n2124), .B(new_n2123), .Y(new_n2125));
  xor_3  g01749(.A(new_n2125), .B(new_n2122), .Y(new_n2126));
  not_3  g01750(.A(new_n2126), .Y(new_n2127));
  nor_4  g01751(.A(new_n2127), .B(new_n2120), .Y(new_n2128));
  not_3  g01752(.A(new_n2120), .Y(new_n2129));
  nor_4  g01753(.A(new_n2126), .B(new_n2129), .Y(new_n2130));
  nor_4  g01754(.A(new_n2130), .B(new_n2128), .Y(new_n2131_1));
  xnor_3 g01755(.A(new_n2131_1), .B(new_n2116), .Y(new_n2132));
  nand_4 g01756(.A(new_n1896), .B(new_n1893), .Y(new_n2133));
  nor_4  g01757(.A(new_n1895), .B(new_n1894), .Y(new_n2134));
  xnor_3 g01758(.A(new_n1896), .B(new_n1892), .Y(new_n2135));
  not_3  g01759(.A(new_n1901), .Y(new_n2136));
  nand_4 g01760(.A(new_n2136), .B(new_n2135), .Y(new_n2137));
  not_3  g01761(.A(new_n2137), .Y(new_n2138));
  xnor_3 g01762(.A(new_n2138), .B(new_n2134), .Y(new_n2139));
  nand_4 g01763(.A(new_n2139), .B(new_n2133), .Y(new_n2140));
  xnor_3 g01764(.A(new_n2140), .B(new_n2132), .Y(new_n2141));
  xnor_3 g01765(.A(new_n2141), .B(new_n2102), .Y(new_n2142));
  xnor_3 g01766(.A(new_n2142), .B(new_n2100), .Y(new_n2143));
  xnor_3 g01767(.A(new_n2143), .B(new_n2097), .Y(new_n2144));
  not_3  g01768(.A(new_n1821), .Y(new_n2145));
  nand_4 g01769(.A(new_n1910), .B(new_n2145), .Y(new_n2146));
  not_3  g01770(.A(new_n1968), .Y(new_n2147));
  nand_4 g01771(.A(new_n2147), .B(new_n1911), .Y(new_n2148));
  nand_4 g01772(.A(new_n2148), .B(new_n2146), .Y(new_n2149));
  xnor_3 g01773(.A(new_n2149), .B(new_n2144), .Y(new_n2150));
  xnor_3 g01774(.A(new_n2150), .B(new_n2058), .Y(new_n2151));
  xnor_3 g01775(.A(new_n2151), .B(new_n2015), .Y(new_n2152));
  nand_4 g01776(.A(new_n2152), .B(new_n1641), .Y(new_n2153));
  xnor_3 g01777(.A(new_n2152), .B(new_n1640), .Y(new_n2154));
  xor_3  g01778(.A(new_n1637), .B(new_n1634), .Y(new_n2155));
  xnor_3 g01779(.A(new_n2013), .B(new_n1971), .Y(new_n2156));
  nand_4 g01780(.A(new_n2156), .B(new_n2155), .Y(new_n2157));
  not_3  g01781(.A(new_n1630), .Y(new_n2158));
  xor_3  g01782(.A(new_n1633), .B(new_n2158), .Y(new_n2159));
  not_3  g01783(.A(new_n2159), .Y(new_n2160));
  not_3  g01784(.A(new_n1980_1), .Y(new_n2161));
  xnor_3 g01785(.A(new_n2011), .B(new_n2161), .Y(new_n2162));
  nor_4  g01786(.A(new_n2162), .B(new_n2160), .Y(new_n2163));
  xnor_3 g01787(.A(new_n2162), .B(new_n2160), .Y(new_n2164));
  xor_3  g01788(.A(new_n1629), .B(new_n1626), .Y(new_n2165));
  not_3  g01789(.A(new_n1986), .Y(new_n2166));
  xnor_3 g01790(.A(new_n2009), .B(new_n2166), .Y(new_n2167));
  nor_4  g01791(.A(new_n2167), .B(new_n2165), .Y(new_n2168));
  xnor_3 g01792(.A(new_n2007), .B(new_n1996), .Y(new_n2169));
  not_3  g01793(.A(new_n1291), .Y(new_n2170));
  nor_4  g01794(.A(new_n1530), .B(new_n2170), .Y(new_n2171));
  nor_4  g01795(.A(new_n2171), .B(new_n1621), .Y(new_n2172));
  nor_4  g01796(.A(new_n1535), .B(new_n2170), .Y(new_n2173));
  nor_4  g01797(.A(new_n2173), .B(new_n2172), .Y(new_n2174));
  nor_4  g01798(.A(new_n2174), .B(new_n2169), .Y(new_n2175));
  xnor_3 g01799(.A(new_n2174), .B(new_n2169), .Y(new_n2176));
  nor_4  g01800(.A(new_n1298), .B(new_n1291), .Y(new_n2177));
  xor_3  g01801(.A(new_n1623), .B(new_n1622), .Y(new_n2178));
  nor_4  g01802(.A(new_n2178), .B(new_n2177), .Y(new_n2179));
  xnor_3 g01803(.A(new_n2005), .B(new_n2003), .Y(new_n2180));
  not_3  g01804(.A(new_n2178), .Y(new_n2181));
  xor_3  g01805(.A(new_n2181), .B(new_n2177), .Y(new_n2182));
  nor_4  g01806(.A(new_n2182), .B(new_n2180), .Y(new_n2183));
  nor_4  g01807(.A(new_n2183), .B(new_n2179), .Y(new_n2184));
  nor_4  g01808(.A(new_n2184), .B(new_n2176), .Y(new_n2185));
  nor_4  g01809(.A(new_n2185), .B(new_n2175), .Y(new_n2186));
  xnor_3 g01810(.A(new_n2167), .B(new_n2165), .Y(new_n2187));
  nor_4  g01811(.A(new_n2187), .B(new_n2186), .Y(new_n2188));
  nor_4  g01812(.A(new_n2188), .B(new_n2168), .Y(new_n2189));
  nor_4  g01813(.A(new_n2189), .B(new_n2164), .Y(new_n2190));
  nor_4  g01814(.A(new_n2190), .B(new_n2163), .Y(new_n2191));
  not_3  g01815(.A(new_n2155), .Y(new_n2192));
  xnor_3 g01816(.A(new_n2156), .B(new_n2192), .Y(new_n2193));
  nand_4 g01817(.A(new_n2193), .B(new_n2191), .Y(new_n2194));
  nand_4 g01818(.A(new_n2194), .B(new_n2157), .Y(new_n2195));
  nand_4 g01819(.A(new_n2195), .B(new_n2154), .Y(new_n2196));
  nand_4 g01820(.A(new_n2196), .B(new_n2153), .Y(new_n2197));
  nand_4 g01821(.A(new_n2076), .B(new_n2074), .Y(new_n2198));
  nand_4 g01822(.A(new_n2084), .B(new_n2077), .Y(new_n2199));
  nand_4 g01823(.A(new_n2199), .B(new_n2198), .Y(new_n2200));
  nand_4 g01824(.A(new_n2025), .B(new_n2022), .Y(new_n2201));
  nand_4 g01825(.A(new_n2201), .B(new_n2028), .Y(new_n2202));
  nand_4 g01826(.A(n6294), .B(n2802), .Y(new_n2203));
  nand_4 g01827(.A(n6797), .B(n533), .Y(new_n2204));
  xor_3  g01828(.A(new_n2204), .B(new_n2203), .Y(new_n2205));
  xor_3  g01829(.A(new_n2205), .B(new_n2202), .Y(new_n2206));
  xor_3  g01830(.A(new_n2206), .B(new_n2200), .Y(new_n2207));
  nand_4 g01831(.A(new_n2143), .B(new_n2097), .Y(new_n2208));
  not_3  g01832(.A(new_n2097), .Y(new_n2209));
  xnor_3 g01833(.A(new_n2143), .B(new_n2209), .Y(new_n2210));
  nand_4 g01834(.A(new_n2149), .B(new_n2210), .Y(new_n2211));
  nand_4 g01835(.A(new_n2211), .B(new_n2208), .Y(new_n2212));
  not_3  g01836(.A(new_n1581), .Y(new_n2213));
  nand_4 g01837(.A(new_n1614), .B(new_n2213), .Y(new_n2214));
  nand_4 g01838(.A(new_n1639), .B(new_n1615), .Y(new_n2215));
  nand_4 g01839(.A(new_n2215), .B(new_n2214), .Y(new_n2216));
  nand_4 g01840(.A(new_n2051), .B(new_n1726), .Y(new_n2217));
  nand_4 g01841(.A(new_n2056), .B(new_n2052), .Y(new_n2218));
  nand_4 g01842(.A(new_n2218), .B(new_n2217), .Y(new_n2219));
  xnor_3 g01843(.A(new_n2219), .B(new_n2216), .Y(new_n2220));
  xnor_3 g01844(.A(new_n2220), .B(new_n2212), .Y(new_n2221));
  not_3  g01845(.A(new_n2105), .Y(new_n2222));
  nand_4 g01846(.A(new_n2115), .B(new_n2222), .Y(new_n2223));
  not_3  g01847(.A(new_n2131_1), .Y(new_n2224));
  nand_4 g01848(.A(new_n2224), .B(new_n2116), .Y(new_n2225));
  nand_4 g01849(.A(new_n2225), .B(new_n2223), .Y(new_n2226_1));
  nand_4 g01850(.A(new_n2119), .B(new_n2117), .Y(new_n2227));
  nand_4 g01851(.A(new_n2127), .B(new_n2120), .Y(new_n2228));
  nand_4 g01852(.A(new_n2228), .B(new_n2227), .Y(new_n2229));
  nand_4 g01853(.A(n6826), .B(n6038), .Y(new_n2230));
  not_3  g01854(.A(new_n2230), .Y(new_n2231));
  nand_4 g01855(.A(new_n2110), .B(new_n2107), .Y(new_n2232));
  nand_4 g01856(.A(new_n2232), .B(new_n2113), .Y(new_n2233));
  xor_3  g01857(.A(new_n2233), .B(new_n2231), .Y(new_n2234));
  xor_3  g01858(.A(new_n2234), .B(new_n2229), .Y(new_n2235));
  xnor_3 g01859(.A(new_n2235), .B(new_n2226_1), .Y(new_n2236));
  nand_4 g01860(.A(new_n2030), .B(new_n2019), .Y(new_n2237));
  nand_4 g01861(.A(new_n2042), .B(new_n2031), .Y(new_n2238));
  nand_4 g01862(.A(new_n2238), .B(new_n2237), .Y(new_n2239));
  nand_4 g01863(.A(n5283), .B(n5069), .Y(new_n2240));
  nand_4 g01864(.A(n4928), .B(n2464), .Y(new_n2241));
  not_3  g01865(.A(new_n2241), .Y(new_n2242));
  xor_3  g01866(.A(new_n2242), .B(new_n2240), .Y(new_n2243));
  xnor_3 g01867(.A(new_n2243), .B(new_n2239), .Y(new_n2244));
  xnor_3 g01868(.A(new_n2244), .B(new_n2236), .Y(new_n2245));
  nand_4 g01869(.A(new_n2138), .B(new_n2134), .Y(new_n2246));
  not_3  g01870(.A(new_n2132), .Y(new_n2247));
  nand_4 g01871(.A(new_n2140), .B(new_n2247), .Y(new_n2248));
  nand_4 g01872(.A(new_n2248), .B(new_n2246), .Y(new_n2249));
  not_3  g01873(.A(new_n2079), .Y(new_n2250));
  nor_4  g01874(.A(new_n2081), .B(new_n2250), .Y(new_n2251));
  not_3  g01875(.A(new_n2078), .Y(new_n2252));
  nor_4  g01876(.A(new_n2082), .B(new_n2252), .Y(new_n2253_1));
  nor_4  g01877(.A(new_n2253_1), .B(new_n2251), .Y(new_n2254));
  nand_4 g01878(.A(n10848), .B(n7646), .Y(new_n2255));
  not_3  g01879(.A(new_n2255), .Y(new_n2256));
  nand_4 g01880(.A(n6806), .B(n137), .Y(new_n2257));
  nand_4 g01881(.A(n8384), .B(n5814), .Y(new_n2258));
  xor_3  g01882(.A(new_n2258), .B(new_n2257), .Y(new_n2259));
  xor_3  g01883(.A(new_n2259), .B(new_n2256), .Y(new_n2260));
  xnor_3 g01884(.A(new_n2260), .B(new_n2254), .Y(new_n2261));
  xnor_3 g01885(.A(new_n2261), .B(new_n2249), .Y(new_n2262));
  xnor_3 g01886(.A(new_n2262), .B(new_n2245), .Y(new_n2263));
  nand_4 g01887(.A(new_n2141), .B(new_n2101), .Y(new_n2264));
  nand_4 g01888(.A(new_n2142), .B(new_n2100), .Y(new_n2265));
  nand_4 g01889(.A(new_n2265), .B(new_n2264), .Y(new_n2266));
  nand_4 g01890(.A(new_n1584), .B(new_n1583), .Y(new_n2267));
  nand_4 g01891(.A(new_n1612), .B(new_n1586), .Y(new_n2268));
  nand_4 g01892(.A(new_n2268), .B(new_n2267), .Y(new_n2269));
  nand_4 g01893(.A(new_n2089), .B(new_n2088), .Y(new_n2270));
  nand_4 g01894(.A(new_n2091), .B(new_n2086), .Y(new_n2271));
  nand_4 g01895(.A(new_n2271), .B(new_n2270), .Y(new_n2272));
  xnor_3 g01896(.A(new_n2272), .B(new_n2269), .Y(new_n2273));
  nand_4 g01897(.A(new_n2048), .B(new_n2046), .Y(new_n2274));
  nand_4 g01898(.A(new_n2050), .B(new_n2043), .Y(new_n2275));
  nand_4 g01899(.A(new_n2275), .B(new_n2274), .Y(new_n2276));
  nor_4  g01900(.A(new_n1610), .B(new_n1601), .Y(new_n2277));
  nor_4  g01901(.A(new_n1611), .B(new_n1598), .Y(new_n2278_1));
  nor_4  g01902(.A(new_n2278_1), .B(new_n2277), .Y(new_n2279));
  and_4  g01903(.A(new_n1594), .B(new_n1593), .Y(new_n2280));
  nor_4  g01904(.A(new_n1595), .B(new_n1592), .Y(new_n2281));
  nor_4  g01905(.A(new_n2281), .B(new_n2280), .Y(new_n2282));
  nand_4 g01906(.A(n12706), .B(n1333), .Y(new_n2283));
  nand_4 g01907(.A(n5240), .B(n2508), .Y(new_n2284));
  nand_4 g01908(.A(n4005), .B(n3172), .Y(new_n2285));
  xnor_3 g01909(.A(new_n2285), .B(new_n2284), .Y(new_n2286));
  xnor_3 g01910(.A(new_n2286), .B(new_n2283), .Y(new_n2287));
  xnor_3 g01911(.A(new_n2287), .B(new_n2282), .Y(new_n2288));
  and_4  g01912(.A(new_n2038), .B(new_n2037), .Y(new_n2289));
  nor_4  g01913(.A(new_n2039), .B(new_n2036), .Y(new_n2290));
  nor_4  g01914(.A(new_n2290), .B(new_n2289), .Y(new_n2291));
  nand_4 g01915(.A(n4203), .B(n1209), .Y(new_n2292));
  nand_4 g01916(.A(n9400), .B(n8236), .Y(new_n2293));
  nand_4 g01917(.A(n5105), .B(n4187), .Y(new_n2294));
  xnor_3 g01918(.A(new_n2294), .B(new_n2293), .Y(new_n2295));
  xnor_3 g01919(.A(new_n2295), .B(new_n2292), .Y(new_n2296));
  xnor_3 g01920(.A(new_n2296), .B(new_n2291), .Y(new_n2297));
  xnor_3 g01921(.A(new_n2297), .B(new_n2288), .Y(new_n2298));
  nand_4 g01922(.A(n12720), .B(n11821), .Y(new_n2299));
  nand_4 g01923(.A(n6877), .B(n783), .Y(new_n2300));
  xnor_3 g01924(.A(new_n2300), .B(new_n2299), .Y(new_n2301_1));
  nand_4 g01925(.A(n9080), .B(n2509), .Y(new_n2302));
  nand_4 g01926(.A(n11757), .B(n2585), .Y(new_n2303));
  xnor_3 g01927(.A(new_n2303), .B(new_n2302), .Y(new_n2304));
  xnor_3 g01928(.A(new_n2304), .B(new_n2301_1), .Y(new_n2305));
  not_3  g01929(.A(new_n1602), .Y(new_n2306));
  nand_4 g01930(.A(new_n1605), .B(new_n2306), .Y(new_n2307));
  nand_4 g01931(.A(new_n2307), .B(new_n1608), .Y(new_n2308));
  nand_4 g01932(.A(n12753), .B(n7500), .Y(new_n2309));
  nand_4 g01933(.A(n10174), .B(n7354), .Y(new_n2310));
  xnor_3 g01934(.A(new_n2310), .B(new_n2309), .Y(new_n2311));
  xnor_3 g01935(.A(new_n2311), .B(new_n2308), .Y(new_n2312));
  xnor_3 g01936(.A(new_n2312), .B(new_n2305), .Y(new_n2313));
  xnor_3 g01937(.A(new_n2313), .B(new_n2298), .Y(new_n2314));
  and_4  g01938(.A(new_n2124), .B(new_n2123), .Y(new_n2315));
  nor_4  g01939(.A(new_n2125), .B(new_n2122), .Y(new_n2316_1));
  nor_4  g01940(.A(new_n2316_1), .B(new_n2315), .Y(new_n2317));
  nand_4 g01941(.A(n11311), .B(n4141), .Y(new_n2318));
  nand_4 g01942(.A(n12044), .B(n11478), .Y(new_n2319));
  nand_4 g01943(.A(n7862), .B(n615), .Y(new_n2320));
  xnor_3 g01944(.A(new_n2320), .B(new_n2319), .Y(new_n2321));
  xnor_3 g01945(.A(new_n2321), .B(new_n2318), .Y(new_n2322));
  xnor_3 g01946(.A(new_n2322), .B(new_n2317), .Y(new_n2323));
  nand_4 g01947(.A(n1980), .B(n1471), .Y(new_n2324));
  not_3  g01948(.A(new_n2033), .Y(new_n2325));
  nand_4 g01949(.A(new_n2325), .B(new_n2032), .Y(new_n2326));
  nand_4 g01950(.A(new_n2040), .B(new_n2034), .Y(new_n2327));
  nand_4 g01951(.A(new_n2327), .B(new_n2326), .Y(new_n2328));
  xnor_3 g01952(.A(new_n2328), .B(new_n2324), .Y(new_n2329));
  xnor_3 g01953(.A(new_n2329), .B(new_n2323), .Y(new_n2330));
  xnor_3 g01954(.A(new_n2330), .B(new_n2314), .Y(new_n2331));
  xnor_3 g01955(.A(new_n2331), .B(new_n2279), .Y(new_n2332));
  xnor_3 g01956(.A(new_n2332), .B(new_n2276), .Y(new_n2333));
  nand_4 g01957(.A(n8028), .B(n4722), .Y(new_n2334));
  not_3  g01958(.A(new_n2334), .Y(new_n2335));
  nand_4 g01959(.A(new_n2071), .B(new_n2065), .Y(new_n2336));
  nand_4 g01960(.A(new_n2085), .B(new_n2073), .Y(new_n2337));
  nand_4 g01961(.A(new_n2337), .B(new_n2336), .Y(new_n2338));
  nand_4 g01962(.A(n3146), .B(n1512), .Y(new_n2339));
  not_3  g01963(.A(new_n2339), .Y(new_n2340));
  nand_4 g01964(.A(n5694), .B(n4805), .Y(new_n2341));
  nand_4 g01965(.A(n4903), .B(n3992), .Y(new_n2342));
  xnor_3 g01966(.A(new_n2342), .B(new_n2341), .Y(new_n2343));
  nand_4 g01967(.A(n4938), .B(n1564), .Y(new_n2344));
  nand_4 g01968(.A(n12704), .B(n6358), .Y(new_n2345));
  xnor_3 g01969(.A(new_n2345), .B(new_n2344), .Y(new_n2346));
  xnor_3 g01970(.A(new_n2346), .B(new_n2343), .Y(new_n2347_1));
  xnor_3 g01971(.A(new_n2347_1), .B(new_n2340), .Y(new_n2348));
  nand_4 g01972(.A(n7294), .B(n5198), .Y(new_n2349));
  not_3  g01973(.A(new_n2349), .Y(new_n2350));
  and_4  g01974(.A(new_n2069), .B(new_n2068), .Y(new_n2351));
  nor_4  g01975(.A(new_n2070), .B(new_n2067), .Y(new_n2352));
  nor_4  g01976(.A(new_n2352), .B(new_n2351), .Y(new_n2353));
  xnor_3 g01977(.A(new_n2353), .B(new_n2350), .Y(new_n2354));
  xnor_3 g01978(.A(new_n2354), .B(new_n2348), .Y(new_n2355));
  nand_4 g01979(.A(n7236), .B(n1906), .Y(new_n2356));
  nand_4 g01980(.A(new_n1589), .B(new_n1587), .Y(new_n2357));
  nand_4 g01981(.A(new_n1596), .B(new_n1590), .Y(new_n2358));
  nand_4 g01982(.A(new_n2358), .B(new_n2357), .Y(new_n2359));
  xnor_3 g01983(.A(new_n2359), .B(new_n2356), .Y(new_n2360));
  xnor_3 g01984(.A(new_n2360), .B(new_n2355), .Y(new_n2361));
  xnor_3 g01985(.A(new_n2361), .B(new_n2338), .Y(new_n2362));
  xnor_3 g01986(.A(new_n2362), .B(new_n2335), .Y(new_n2363));
  xnor_3 g01987(.A(new_n2363), .B(new_n2333), .Y(new_n2364));
  xnor_3 g01988(.A(new_n2364), .B(new_n2273), .Y(new_n2365));
  xnor_3 g01989(.A(new_n2365), .B(new_n2266), .Y(new_n2366));
  xnor_3 g01990(.A(new_n2366), .B(new_n2263), .Y(new_n2367));
  xnor_3 g01991(.A(new_n2367), .B(new_n2221), .Y(new_n2368));
  xnor_3 g01992(.A(new_n2368), .B(new_n2207), .Y(new_n2369));
  nor_4  g01993(.A(new_n2092), .B(new_n2060), .Y(new_n2370));
  nor_4  g01994(.A(new_n2096_1), .B(new_n2093), .Y(new_n2371));
  nor_4  g01995(.A(new_n2371), .B(new_n2370), .Y(new_n2372));
  nand_4 g01996(.A(new_n2150), .B(new_n2057), .Y(new_n2373));
  nand_4 g01997(.A(new_n2151), .B(new_n2015), .Y(new_n2374));
  nand_4 g01998(.A(new_n2374), .B(new_n2373), .Y(new_n2375));
  xnor_3 g01999(.A(new_n2375), .B(new_n2372), .Y(new_n2376));
  xnor_3 g02000(.A(new_n2376), .B(new_n2369), .Y(new_n2377));
  xnor_3 g02001(.A(new_n2377), .B(new_n2197), .Y(n671));
  nand_4 g02002(.A(n5964), .B(n2577), .Y(new_n2379));
  nand_4 g02003(.A(n3842), .B(n1097), .Y(new_n2380));
  nor_4  g02004(.A(new_n2380), .B(new_n2379), .Y(new_n2381));
  nand_4 g02005(.A(n11917), .B(n4312), .Y(new_n2382));
  nand_4 g02006(.A(n12705), .B(n4921), .Y(new_n2383_1));
  nand_4 g02007(.A(n12025), .B(n9956), .Y(new_n2384));
  xnor_3 g02008(.A(new_n2384), .B(new_n2383_1), .Y(new_n2385));
  xnor_3 g02009(.A(new_n2385), .B(new_n2382), .Y(new_n2386));
  nand_4 g02010(.A(n12705), .B(n9956), .Y(new_n2387));
  not_3  g02011(.A(new_n2387), .Y(new_n2388));
  nand_4 g02012(.A(n11917), .B(n1097), .Y(new_n2389));
  not_3  g02013(.A(new_n2389), .Y(new_n2390));
  nor_4  g02014(.A(new_n2390), .B(new_n2388), .Y(new_n2391));
  nor_4  g02015(.A(new_n2389), .B(new_n2387), .Y(new_n2392));
  nand_4 g02016(.A(n4921), .B(n4312), .Y(new_n2393_1));
  not_3  g02017(.A(new_n2393_1), .Y(new_n2394));
  nor_4  g02018(.A(new_n2394), .B(new_n2392), .Y(new_n2395));
  nor_4  g02019(.A(new_n2395), .B(new_n2391), .Y(new_n2396));
  xnor_3 g02020(.A(new_n2396), .B(new_n2386), .Y(new_n2397));
  xor_3  g02021(.A(new_n2380), .B(new_n2379), .Y(new_n2398));
  xnor_3 g02022(.A(new_n2398), .B(new_n2397), .Y(new_n2399));
  nand_4 g02023(.A(n5964), .B(n3842), .Y(new_n2400));
  not_3  g02024(.A(new_n2400), .Y(new_n2401));
  nand_4 g02025(.A(n9956), .B(n4312), .Y(new_n2402));
  not_3  g02026(.A(new_n2402), .Y(new_n2403));
  nand_4 g02027(.A(n11917), .B(n5964), .Y(new_n2404));
  not_3  g02028(.A(new_n2404), .Y(new_n2405));
  nor_4  g02029(.A(new_n2405), .B(new_n2403), .Y(new_n2406));
  nor_4  g02030(.A(new_n2404), .B(new_n2402), .Y(new_n2407));
  nand_4 g02031(.A(n4921), .B(n1097), .Y(new_n2408));
  not_3  g02032(.A(new_n2408), .Y(new_n2409));
  nor_4  g02033(.A(new_n2409), .B(new_n2407), .Y(new_n2410));
  nor_4  g02034(.A(new_n2410), .B(new_n2406), .Y(new_n2411));
  nand_4 g02035(.A(new_n2411), .B(new_n2401), .Y(new_n2412));
  not_3  g02036(.A(new_n2412), .Y(new_n2413));
  nor_4  g02037(.A(new_n2411), .B(new_n2401), .Y(new_n2414));
  nor_4  g02038(.A(new_n2414), .B(new_n2413), .Y(new_n2415));
  not_3  g02039(.A(new_n2391), .Y(new_n2416));
  not_3  g02040(.A(new_n2392), .Y(new_n2417));
  nand_4 g02041(.A(new_n2417), .B(new_n2416), .Y(new_n2418));
  xnor_3 g02042(.A(new_n2418), .B(new_n2393_1), .Y(new_n2419));
  not_3  g02043(.A(new_n2419), .Y(new_n2420));
  nand_4 g02044(.A(new_n2420), .B(new_n2415), .Y(new_n2421));
  nand_4 g02045(.A(new_n2421), .B(new_n2412), .Y(new_n2422));
  not_3  g02046(.A(new_n2422), .Y(new_n2423));
  nor_4  g02047(.A(new_n2423), .B(new_n2399), .Y(new_n2424));
  and_4  g02048(.A(new_n2424), .B(new_n2381), .Y(new_n2425_1));
  nand_4 g02049(.A(new_n2385), .B(new_n2382), .Y(new_n2426));
  not_3  g02050(.A(new_n2386), .Y(new_n2427));
  not_3  g02051(.A(new_n2396), .Y(new_n2428));
  nand_4 g02052(.A(new_n2428), .B(new_n2427), .Y(new_n2429));
  and_4  g02053(.A(new_n2429), .B(new_n2426), .Y(new_n2430));
  nand_4 g02054(.A(n9637), .B(n5964), .Y(new_n2431_1));
  not_3  g02055(.A(new_n2431_1), .Y(new_n2432));
  nand_4 g02056(.A(n2577), .B(n1097), .Y(new_n2433_1));
  nand_4 g02057(.A(n5305), .B(n1835), .Y(new_n2434_1));
  xnor_3 g02058(.A(new_n2434_1), .B(new_n2433_1), .Y(new_n2435));
  xor_3  g02059(.A(new_n2435), .B(new_n2432), .Y(new_n2436));
  xnor_3 g02060(.A(new_n2436), .B(new_n2430), .Y(new_n2437));
  not_3  g02061(.A(new_n2437), .Y(new_n2438));
  nor_4  g02062(.A(new_n2384), .B(new_n2383_1), .Y(new_n2439));
  not_3  g02063(.A(new_n2439), .Y(new_n2440));
  nand_4 g02064(.A(n4312), .B(n3842), .Y(new_n2441));
  xor_3  g02065(.A(new_n2441), .B(new_n2440), .Y(new_n2442));
  not_3  g02066(.A(new_n2442), .Y(new_n2443));
  nand_4 g02067(.A(n12025), .B(n4921), .Y(new_n2444));
  not_3  g02068(.A(new_n2444), .Y(new_n2445));
  nand_4 g02069(.A(n12705), .B(n11917), .Y(new_n2446));
  nand_4 g02070(.A(n11257), .B(n9956), .Y(new_n2447));
  xnor_3 g02071(.A(new_n2447), .B(new_n2446), .Y(new_n2448));
  and_4  g02072(.A(new_n2448), .B(new_n2445), .Y(new_n2449));
  nor_4  g02073(.A(new_n2448), .B(new_n2445), .Y(new_n2450));
  nor_4  g02074(.A(new_n2450), .B(new_n2449), .Y(new_n2451));
  xnor_3 g02075(.A(new_n2451), .B(new_n2443), .Y(new_n2452));
  xnor_3 g02076(.A(new_n2452), .B(new_n2438), .Y(new_n2453));
  not_3  g02077(.A(new_n2453), .Y(new_n2454));
  nand_4 g02078(.A(new_n2398), .B(new_n2397), .Y(new_n2455));
  xnor_3 g02079(.A(new_n2424), .B(new_n2381), .Y(new_n2456));
  nand_4 g02080(.A(new_n2456), .B(new_n2455), .Y(new_n2457));
  and_4  g02081(.A(new_n2457), .B(new_n2454), .Y(new_n2458));
  nor_4  g02082(.A(new_n2458), .B(new_n2425_1), .Y(new_n2459));
  nand_4 g02083(.A(n8759), .B(n8065), .Y(new_n2460));
  not_3  g02084(.A(new_n2460), .Y(new_n2461));
  nand_4 g02085(.A(n7436), .B(n6126), .Y(new_n2462));
  nand_4 g02086(.A(n8276), .B(n3602), .Y(new_n2463));
  nand_4 g02087(.A(n9241), .B(n3719), .Y(new_n2464_1));
  xnor_3 g02088(.A(new_n2464_1), .B(new_n2463), .Y(new_n2465));
  nor_4  g02089(.A(new_n2465), .B(new_n2462), .Y(new_n2466));
  not_3  g02090(.A(new_n2462), .Y(new_n2467));
  not_3  g02091(.A(new_n2465), .Y(new_n2468));
  nor_4  g02092(.A(new_n2468), .B(new_n2467), .Y(new_n2469));
  nor_4  g02093(.A(new_n2469), .B(new_n2466), .Y(new_n2470));
  nand_4 g02094(.A(n8276), .B(n3719), .Y(new_n2471));
  not_3  g02095(.A(new_n2471), .Y(new_n2472));
  nand_4 g02096(.A(n12299), .B(n6126), .Y(new_n2473));
  not_3  g02097(.A(new_n2473), .Y(new_n2474));
  nor_4  g02098(.A(new_n2474), .B(new_n2472), .Y(new_n2475));
  nor_4  g02099(.A(new_n2473), .B(new_n2471), .Y(new_n2476));
  nand_4 g02100(.A(n7436), .B(n3602), .Y(new_n2477));
  not_3  g02101(.A(new_n2477), .Y(new_n2478));
  nor_4  g02102(.A(new_n2478), .B(new_n2476), .Y(new_n2479));
  nor_4  g02103(.A(new_n2479), .B(new_n2475), .Y(new_n2480));
  xnor_3 g02104(.A(new_n2480), .B(new_n2470), .Y(new_n2481));
  nand_4 g02105(.A(n10439), .B(n6776), .Y(new_n2482));
  nand_4 g02106(.A(n12299), .B(n8595), .Y(new_n2483));
  xor_3  g02107(.A(new_n2483), .B(new_n2482), .Y(new_n2484));
  xnor_3 g02108(.A(new_n2484), .B(new_n2481), .Y(new_n2485));
  nand_4 g02109(.A(n8595), .B(n6776), .Y(new_n2486));
  not_3  g02110(.A(new_n2486), .Y(new_n2487));
  nand_4 g02111(.A(n7436), .B(n3719), .Y(new_n2488));
  not_3  g02112(.A(new_n2488), .Y(new_n2489));
  nand_4 g02113(.A(n6776), .B(n6126), .Y(new_n2490));
  not_3  g02114(.A(new_n2490), .Y(new_n2491));
  nor_4  g02115(.A(new_n2491), .B(new_n2489), .Y(new_n2492));
  nor_4  g02116(.A(new_n2490), .B(new_n2488), .Y(new_n2493));
  nand_4 g02117(.A(n12299), .B(n3602), .Y(new_n2494));
  not_3  g02118(.A(new_n2494), .Y(new_n2495));
  nor_4  g02119(.A(new_n2495), .B(new_n2493), .Y(new_n2496));
  nor_4  g02120(.A(new_n2496), .B(new_n2492), .Y(new_n2497));
  nand_4 g02121(.A(new_n2497), .B(new_n2487), .Y(new_n2498_1));
  not_3  g02122(.A(new_n2498_1), .Y(new_n2499));
  xnor_3 g02123(.A(new_n2497), .B(new_n2487), .Y(new_n2500));
  nor_4  g02124(.A(new_n2476), .B(new_n2475), .Y(new_n2501));
  xnor_3 g02125(.A(new_n2501), .B(new_n2478), .Y(new_n2502));
  nor_4  g02126(.A(new_n2502), .B(new_n2500), .Y(new_n2503));
  nor_4  g02127(.A(new_n2503), .B(new_n2499), .Y(new_n2504));
  not_3  g02128(.A(new_n2504), .Y(new_n2505));
  nand_4 g02129(.A(new_n2505), .B(new_n2485), .Y(new_n2506));
  not_3  g02130(.A(new_n2506), .Y(new_n2507_1));
  nor_4  g02131(.A(new_n2505), .B(new_n2485), .Y(new_n2508_1));
  nor_4  g02132(.A(new_n2508_1), .B(new_n2507_1), .Y(new_n2509_1));
  not_3  g02133(.A(new_n2509_1), .Y(new_n2510));
  nand_4 g02134(.A(n10439), .B(n8759), .Y(new_n2511));
  not_3  g02135(.A(new_n2511), .Y(new_n2512_1));
  xnor_3 g02136(.A(new_n2502), .B(new_n2500), .Y(new_n2513));
  not_3  g02137(.A(new_n2513), .Y(new_n2514));
  nor_4  g02138(.A(new_n2514), .B(new_n2512_1), .Y(new_n2515_1));
  not_3  g02139(.A(new_n2515_1), .Y(new_n2516));
  nor_4  g02140(.A(new_n2513), .B(new_n2511), .Y(new_n2517));
  nor_4  g02141(.A(new_n2517), .B(new_n2515_1), .Y(new_n2518));
  nand_4 g02142(.A(n8759), .B(n8595), .Y(new_n2519));
  nand_4 g02143(.A(n12299), .B(n3719), .Y(new_n2520));
  not_3  g02144(.A(new_n2520), .Y(new_n2521));
  nand_4 g02145(.A(n8759), .B(n6126), .Y(new_n2522_1));
  not_3  g02146(.A(new_n2522_1), .Y(new_n2523));
  nand_4 g02147(.A(new_n2523), .B(new_n2521), .Y(new_n2524));
  nand_4 g02148(.A(new_n2522_1), .B(new_n2520), .Y(new_n2525));
  nand_4 g02149(.A(n6776), .B(n3602), .Y(new_n2526));
  not_3  g02150(.A(new_n2526), .Y(new_n2527));
  nand_4 g02151(.A(new_n2527), .B(new_n2525), .Y(new_n2528));
  nand_4 g02152(.A(new_n2528), .B(new_n2524), .Y(new_n2529));
  not_3  g02153(.A(new_n2529), .Y(new_n2530_1));
  nor_4  g02154(.A(new_n2530_1), .B(new_n2519), .Y(new_n2531));
  xor_3  g02155(.A(new_n2529), .B(new_n2519), .Y(new_n2532));
  nor_4  g02156(.A(new_n2493), .B(new_n2492), .Y(new_n2533));
  xor_3  g02157(.A(new_n2533), .B(new_n2494), .Y(new_n2534));
  nor_4  g02158(.A(new_n2534), .B(new_n2532), .Y(new_n2535));
  nor_4  g02159(.A(new_n2535), .B(new_n2531), .Y(new_n2536));
  nand_4 g02160(.A(new_n2536), .B(new_n2518), .Y(new_n2537));
  nand_4 g02161(.A(new_n2537), .B(new_n2516), .Y(new_n2538));
  nor_4  g02162(.A(new_n2538), .B(new_n2510), .Y(new_n2539));
  not_3  g02163(.A(new_n2538), .Y(new_n2540));
  nor_4  g02164(.A(new_n2540), .B(new_n2509_1), .Y(new_n2541));
  nor_4  g02165(.A(new_n2541), .B(new_n2539), .Y(new_n2542));
  nand_4 g02166(.A(new_n2542), .B(new_n2461), .Y(new_n2543));
  and_4  g02167(.A(new_n2525), .B(new_n2524), .Y(new_n2544));
  nand_4 g02168(.A(n6776), .B(n3719), .Y(new_n2545));
  nand_4 g02169(.A(n8759), .B(n3602), .Y(new_n2546));
  nor_4  g02170(.A(new_n2546), .B(new_n2545), .Y(new_n2547));
  not_3  g02171(.A(new_n2547), .Y(new_n2548));
  nor_4  g02172(.A(new_n2548), .B(new_n2544), .Y(new_n2549));
  not_3  g02173(.A(new_n2549), .Y(new_n2550));
  xnor_3 g02174(.A(new_n2534), .B(new_n2532), .Y(new_n2551_1));
  nor_4  g02175(.A(new_n2551_1), .B(new_n2550), .Y(new_n2552));
  not_3  g02176(.A(new_n2552), .Y(new_n2553));
  xnor_3 g02177(.A(new_n2536), .B(new_n2518), .Y(new_n2554));
  not_3  g02178(.A(new_n2554), .Y(new_n2555));
  nor_4  g02179(.A(new_n2555), .B(new_n2553), .Y(new_n2556));
  xnor_3 g02180(.A(new_n2542), .B(new_n2460), .Y(new_n2557));
  nand_4 g02181(.A(new_n2557), .B(new_n2556), .Y(new_n2558_1));
  nand_4 g02182(.A(new_n2558_1), .B(new_n2543), .Y(new_n2559));
  not_3  g02183(.A(new_n2466), .Y(new_n2560));
  nand_4 g02184(.A(new_n2480), .B(new_n2470), .Y(new_n2561));
  nand_4 g02185(.A(new_n2561), .B(new_n2560), .Y(new_n2562));
  nand_4 g02186(.A(n8065), .B(n6776), .Y(new_n2563));
  nand_4 g02187(.A(n12299), .B(n10439), .Y(new_n2564_1));
  nand_4 g02188(.A(n10391), .B(n8759), .Y(new_n2565));
  not_3  g02189(.A(new_n2565), .Y(new_n2566));
  xor_3  g02190(.A(new_n2566), .B(new_n2564_1), .Y(new_n2567));
  xnor_3 g02191(.A(new_n2567), .B(new_n2563), .Y(new_n2568));
  not_3  g02192(.A(new_n2568), .Y(new_n2569));
  xor_3  g02193(.A(new_n2569), .B(new_n2562), .Y(new_n2570));
  nor_4  g02194(.A(new_n2464_1), .B(new_n2463), .Y(new_n2571));
  not_3  g02195(.A(new_n2571), .Y(new_n2572));
  nand_4 g02196(.A(n8595), .B(n7436), .Y(new_n2573));
  xor_3  g02197(.A(new_n2573), .B(new_n2572), .Y(new_n2574));
  nand_4 g02198(.A(n9241), .B(n3602), .Y(new_n2575));
  not_3  g02199(.A(new_n2575), .Y(new_n2576));
  nand_4 g02200(.A(n8276), .B(n6126), .Y(new_n2577_1));
  nand_4 g02201(.A(n10510), .B(n3719), .Y(new_n2578));
  xor_3  g02202(.A(new_n2578), .B(new_n2577_1), .Y(new_n2579));
  xnor_3 g02203(.A(new_n2579), .B(new_n2576), .Y(new_n2580));
  xnor_3 g02204(.A(new_n2580), .B(new_n2574), .Y(new_n2581_1));
  xnor_3 g02205(.A(new_n2581_1), .B(new_n2570), .Y(new_n2582));
  not_3  g02206(.A(new_n2481), .Y(new_n2583));
  nand_4 g02207(.A(new_n2484), .B(new_n2583), .Y(new_n2584));
  nor_4  g02208(.A(new_n2483), .B(new_n2482), .Y(new_n2585_1));
  xnor_3 g02209(.A(new_n2507_1), .B(new_n2585_1), .Y(new_n2586));
  nand_4 g02210(.A(new_n2586), .B(new_n2584), .Y(new_n2587));
  xnor_3 g02211(.A(new_n2587), .B(new_n2582), .Y(new_n2588));
  xnor_3 g02212(.A(new_n2588), .B(new_n2539), .Y(new_n2589));
  xnor_3 g02213(.A(new_n2589), .B(new_n2559), .Y(new_n2590));
  nand_4 g02214(.A(n12648), .B(n4826), .Y(new_n2591));
  nand_4 g02215(.A(n10545), .B(n7733), .Y(new_n2592));
  nand_4 g02216(.A(n12925), .B(n7690), .Y(new_n2593));
  xnor_3 g02217(.A(new_n2593), .B(new_n2592), .Y(new_n2594));
  nor_4  g02218(.A(new_n2594), .B(new_n2591), .Y(new_n2595));
  not_3  g02219(.A(new_n2591), .Y(new_n2596));
  not_3  g02220(.A(new_n2594), .Y(new_n2597));
  nor_4  g02221(.A(new_n2597), .B(new_n2596), .Y(new_n2598));
  nor_4  g02222(.A(new_n2598), .B(new_n2595), .Y(new_n2599));
  nand_4 g02223(.A(n12925), .B(n10545), .Y(new_n2600));
  not_3  g02224(.A(new_n2600), .Y(new_n2601));
  nand_4 g02225(.A(n4826), .B(n2530), .Y(new_n2602));
  not_3  g02226(.A(new_n2602), .Y(new_n2603));
  nor_4  g02227(.A(new_n2603), .B(new_n2601), .Y(new_n2604));
  nand_4 g02228(.A(n12648), .B(n7733), .Y(new_n2605));
  not_3  g02229(.A(new_n2605), .Y(new_n2606));
  xnor_3 g02230(.A(new_n2602), .B(new_n2600), .Y(new_n2607));
  nor_4  g02231(.A(new_n2607), .B(new_n2606), .Y(new_n2608));
  nor_4  g02232(.A(new_n2608), .B(new_n2604), .Y(new_n2609));
  xnor_3 g02233(.A(new_n2609), .B(new_n2599), .Y(new_n2610));
  nand_4 g02234(.A(n8476), .B(n4970), .Y(new_n2611));
  nand_4 g02235(.A(n7610), .B(n2530), .Y(new_n2612));
  xor_3  g02236(.A(new_n2612), .B(new_n2611), .Y(new_n2613));
  xnor_3 g02237(.A(new_n2613), .B(new_n2610), .Y(new_n2614));
  nand_4 g02238(.A(n8476), .B(n7610), .Y(new_n2615));
  not_3  g02239(.A(new_n2615), .Y(new_n2616));
  nand_4 g02240(.A(n12925), .B(n12648), .Y(new_n2617));
  not_3  g02241(.A(new_n2617), .Y(new_n2618));
  nand_4 g02242(.A(n8476), .B(n4826), .Y(new_n2619));
  not_3  g02243(.A(new_n2619), .Y(new_n2620));
  nor_4  g02244(.A(new_n2620), .B(new_n2618), .Y(new_n2621));
  nand_4 g02245(.A(n7733), .B(n2530), .Y(new_n2622));
  not_3  g02246(.A(new_n2622), .Y(new_n2623));
  xnor_3 g02247(.A(new_n2619), .B(new_n2617), .Y(new_n2624_1));
  nor_4  g02248(.A(new_n2624_1), .B(new_n2623), .Y(new_n2625));
  nor_4  g02249(.A(new_n2625), .B(new_n2621), .Y(new_n2626));
  nand_4 g02250(.A(new_n2626), .B(new_n2616), .Y(new_n2627));
  not_3  g02251(.A(new_n2627), .Y(new_n2628));
  nor_4  g02252(.A(new_n2626), .B(new_n2616), .Y(new_n2629));
  nor_4  g02253(.A(new_n2629), .B(new_n2628), .Y(new_n2630));
  xnor_3 g02254(.A(new_n2607), .B(new_n2605), .Y(new_n2631));
  not_3  g02255(.A(new_n2631), .Y(new_n2632));
  nand_4 g02256(.A(new_n2632), .B(new_n2630), .Y(new_n2633));
  nand_4 g02257(.A(new_n2633), .B(new_n2627), .Y(new_n2634));
  xnor_3 g02258(.A(new_n2634), .B(new_n2614), .Y(new_n2635));
  nand_4 g02259(.A(n5331), .B(n4970), .Y(new_n2636));
  not_3  g02260(.A(new_n2636), .Y(new_n2637));
  nand_4 g02261(.A(n7610), .B(n5331), .Y(new_n2638));
  not_3  g02262(.A(new_n2638), .Y(new_n2639));
  nand_4 g02263(.A(n12925), .B(n2530), .Y(new_n2640));
  not_3  g02264(.A(new_n2640), .Y(new_n2641));
  nand_4 g02265(.A(n5331), .B(n4826), .Y(new_n2642));
  not_3  g02266(.A(new_n2642), .Y(new_n2643));
  nor_4  g02267(.A(new_n2643), .B(new_n2641), .Y(new_n2644));
  nor_4  g02268(.A(new_n2642), .B(new_n2640), .Y(new_n2645));
  nand_4 g02269(.A(n8476), .B(n7733), .Y(new_n2646));
  not_3  g02270(.A(new_n2646), .Y(new_n2647));
  nor_4  g02271(.A(new_n2647), .B(new_n2645), .Y(new_n2648));
  nor_4  g02272(.A(new_n2648), .B(new_n2644), .Y(new_n2649));
  nand_4 g02273(.A(new_n2649), .B(new_n2639), .Y(new_n2650));
  not_3  g02274(.A(new_n2650), .Y(new_n2651));
  nor_4  g02275(.A(new_n2649), .B(new_n2639), .Y(new_n2652));
  nor_4  g02276(.A(new_n2652), .B(new_n2651), .Y(new_n2653));
  xnor_3 g02277(.A(new_n2624_1), .B(new_n2622), .Y(new_n2654));
  not_3  g02278(.A(new_n2654), .Y(new_n2655));
  nand_4 g02279(.A(new_n2655), .B(new_n2653), .Y(new_n2656));
  nand_4 g02280(.A(new_n2656), .B(new_n2650), .Y(new_n2657));
  nor_4  g02281(.A(new_n2657), .B(new_n2637), .Y(new_n2658));
  not_3  g02282(.A(new_n2658), .Y(new_n2659));
  xnor_3 g02283(.A(new_n2632), .B(new_n2630), .Y(new_n2660));
  not_3  g02284(.A(new_n2657), .Y(new_n2661));
  nor_4  g02285(.A(new_n2661), .B(new_n2636), .Y(new_n2662));
  nor_4  g02286(.A(new_n2662), .B(new_n2658), .Y(new_n2663));
  nand_4 g02287(.A(new_n2663), .B(new_n2660), .Y(new_n2664));
  nand_4 g02288(.A(new_n2664), .B(new_n2659), .Y(new_n2665));
  nor_4  g02289(.A(new_n2665), .B(new_n2635), .Y(new_n2666));
  not_3  g02290(.A(new_n2610), .Y(new_n2667));
  nand_4 g02291(.A(new_n2613), .B(new_n2667), .Y(new_n2668));
  nor_4  g02292(.A(new_n2612), .B(new_n2611), .Y(new_n2669));
  nand_4 g02293(.A(new_n2634), .B(new_n2614), .Y(new_n2670));
  not_3  g02294(.A(new_n2670), .Y(new_n2671));
  xnor_3 g02295(.A(new_n2671), .B(new_n2669), .Y(new_n2672));
  nand_4 g02296(.A(new_n2672), .B(new_n2668), .Y(new_n2673));
  not_3  g02297(.A(new_n2595), .Y(new_n2674));
  nand_4 g02298(.A(new_n2609), .B(new_n2599), .Y(new_n2675));
  nand_4 g02299(.A(new_n2675), .B(new_n2674), .Y(new_n2676));
  nand_4 g02300(.A(n8476), .B(n503), .Y(new_n2677));
  nand_4 g02301(.A(n4970), .B(n2530), .Y(new_n2678));
  nand_4 g02302(.A(n10965), .B(n5331), .Y(new_n2679_1));
  xnor_3 g02303(.A(new_n2679_1), .B(new_n2678), .Y(new_n2680));
  xor_3  g02304(.A(new_n2680), .B(new_n2677), .Y(new_n2681));
  xnor_3 g02305(.A(new_n2681), .B(new_n2676), .Y(new_n2682));
  nor_4  g02306(.A(new_n2593), .B(new_n2592), .Y(new_n2683));
  nand_4 g02307(.A(n12648), .B(n7610), .Y(new_n2684));
  not_3  g02308(.A(new_n2684), .Y(new_n2685));
  xor_3  g02309(.A(new_n2685), .B(new_n2683), .Y(new_n2686));
  not_3  g02310(.A(new_n2686), .Y(new_n2687));
  nand_4 g02311(.A(n7733), .B(n7690), .Y(new_n2688));
  not_3  g02312(.A(new_n2688), .Y(new_n2689));
  nand_4 g02313(.A(n10545), .B(n4826), .Y(new_n2690));
  nand_4 g02314(.A(n12925), .B(n3616), .Y(new_n2691));
  xnor_3 g02315(.A(new_n2691), .B(new_n2690), .Y(new_n2692));
  xnor_3 g02316(.A(new_n2692), .B(new_n2689), .Y(new_n2693));
  not_3  g02317(.A(new_n2693), .Y(new_n2694));
  xor_3  g02318(.A(new_n2694), .B(new_n2687), .Y(new_n2695));
  xnor_3 g02319(.A(new_n2695), .B(new_n2682), .Y(new_n2696));
  xnor_3 g02320(.A(new_n2696), .B(new_n2673), .Y(new_n2697));
  xnor_3 g02321(.A(new_n2697), .B(new_n2666), .Y(new_n2698));
  nand_4 g02322(.A(n5331), .B(n503), .Y(new_n2699));
  not_3  g02323(.A(new_n2699), .Y(new_n2700));
  not_3  g02324(.A(new_n2665), .Y(new_n2701));
  xnor_3 g02325(.A(new_n2701), .B(new_n2635), .Y(new_n2702));
  nand_4 g02326(.A(new_n2702), .B(new_n2700), .Y(new_n2703));
  xnor_3 g02327(.A(new_n2649), .B(new_n2639), .Y(new_n2704));
  xnor_3 g02328(.A(new_n2654), .B(new_n2704), .Y(new_n2705));
  not_3  g02329(.A(new_n2644), .Y(new_n2706));
  nand_4 g02330(.A(n12925), .B(n5331), .Y(new_n2707));
  not_3  g02331(.A(new_n2707), .Y(new_n2708_1));
  nor_4  g02332(.A(new_n2708_1), .B(new_n2646), .Y(new_n2709));
  nor_4  g02333(.A(new_n2709), .B(new_n2706), .Y(new_n2710));
  nor_4  g02334(.A(new_n2710), .B(new_n2645), .Y(new_n2711));
  nor_4  g02335(.A(new_n2711), .B(new_n2646), .Y(new_n2712));
  not_3  g02336(.A(new_n2712), .Y(new_n2713));
  nor_4  g02337(.A(new_n2713), .B(new_n2705), .Y(new_n2714));
  xnor_3 g02338(.A(new_n2663), .B(new_n2660), .Y(new_n2715));
  nand_4 g02339(.A(new_n2715), .B(new_n2714), .Y(new_n2716));
  not_3  g02340(.A(new_n2716), .Y(new_n2717));
  xnor_3 g02341(.A(new_n2702), .B(new_n2699), .Y(new_n2718));
  nand_4 g02342(.A(new_n2718), .B(new_n2717), .Y(new_n2719));
  nand_4 g02343(.A(new_n2719), .B(new_n2703), .Y(new_n2720));
  xnor_3 g02344(.A(new_n2720), .B(new_n2698), .Y(new_n2721));
  nand_4 g02345(.A(n4086), .B(n2393), .Y(new_n2722));
  nand_4 g02346(.A(n5860), .B(n405), .Y(new_n2723));
  nand_4 g02347(.A(n8433), .B(n3986), .Y(new_n2724));
  xnor_3 g02348(.A(new_n2724), .B(new_n2723), .Y(new_n2725));
  nor_4  g02349(.A(new_n2725), .B(new_n2722), .Y(new_n2726));
  not_3  g02350(.A(new_n2722), .Y(new_n2727));
  not_3  g02351(.A(new_n2725), .Y(new_n2728));
  nor_4  g02352(.A(new_n2728), .B(new_n2727), .Y(new_n2729));
  nor_4  g02353(.A(new_n2729), .B(new_n2726), .Y(new_n2730));
  nand_4 g02354(.A(n8433), .B(n5860), .Y(new_n2731));
  not_3  g02355(.A(new_n2731), .Y(new_n2732));
  nand_4 g02356(.A(n11892), .B(n4086), .Y(new_n2733));
  not_3  g02357(.A(new_n2733), .Y(new_n2734));
  nor_4  g02358(.A(new_n2734), .B(new_n2732), .Y(new_n2735));
  nand_4 g02359(.A(n2393), .B(n405), .Y(new_n2736));
  not_3  g02360(.A(new_n2736), .Y(new_n2737));
  xnor_3 g02361(.A(new_n2733), .B(new_n2731), .Y(new_n2738));
  nor_4  g02362(.A(new_n2738), .B(new_n2737), .Y(new_n2739));
  nor_4  g02363(.A(new_n2739), .B(new_n2735), .Y(new_n2740));
  xnor_3 g02364(.A(new_n2740), .B(new_n2730), .Y(new_n2741));
  not_3  g02365(.A(new_n2741), .Y(new_n2742));
  nand_4 g02366(.A(n7388), .B(n6611), .Y(new_n2743));
  nand_4 g02367(.A(n11892), .B(n217), .Y(new_n2744));
  xor_3  g02368(.A(new_n2744), .B(new_n2743), .Y(new_n2745));
  xnor_3 g02369(.A(new_n2745), .B(new_n2742), .Y(new_n2746));
  nand_4 g02370(.A(n7388), .B(n217), .Y(new_n2747));
  not_3  g02371(.A(new_n2747), .Y(new_n2748));
  nand_4 g02372(.A(n8433), .B(n2393), .Y(new_n2749_1));
  not_3  g02373(.A(new_n2749_1), .Y(new_n2750));
  nand_4 g02374(.A(n7388), .B(n4086), .Y(new_n2751));
  not_3  g02375(.A(new_n2751), .Y(new_n2752));
  nor_4  g02376(.A(new_n2752), .B(new_n2750), .Y(new_n2753));
  nor_4  g02377(.A(new_n2751), .B(new_n2749_1), .Y(new_n2754));
  nand_4 g02378(.A(n11892), .B(n405), .Y(new_n2755));
  not_3  g02379(.A(new_n2755), .Y(new_n2756));
  nor_4  g02380(.A(new_n2756), .B(new_n2754), .Y(new_n2757));
  nor_4  g02381(.A(new_n2757), .B(new_n2753), .Y(new_n2758));
  nand_4 g02382(.A(new_n2758), .B(new_n2748), .Y(new_n2759));
  not_3  g02383(.A(new_n2759), .Y(new_n2760));
  xnor_3 g02384(.A(new_n2758), .B(new_n2748), .Y(new_n2761));
  xnor_3 g02385(.A(new_n2738), .B(new_n2736), .Y(new_n2762));
  nor_4  g02386(.A(new_n2762), .B(new_n2761), .Y(new_n2763));
  nor_4  g02387(.A(new_n2763), .B(new_n2760), .Y(new_n2764));
  xnor_3 g02388(.A(new_n2764), .B(new_n2746), .Y(new_n2765));
  nand_4 g02389(.A(n7965), .B(n6611), .Y(new_n2766));
  xnor_3 g02390(.A(new_n2762), .B(new_n2761), .Y(new_n2767));
  nor_4  g02391(.A(new_n2767), .B(new_n2766), .Y(new_n2768));
  xnor_3 g02392(.A(new_n2767), .B(new_n2766), .Y(new_n2769));
  nand_4 g02393(.A(n7965), .B(n217), .Y(new_n2770));
  nand_4 g02394(.A(n11892), .B(n8433), .Y(new_n2771));
  not_3  g02395(.A(new_n2771), .Y(new_n2772));
  nand_4 g02396(.A(n7965), .B(n4086), .Y(new_n2773));
  not_3  g02397(.A(new_n2773), .Y(new_n2774));
  nand_4 g02398(.A(new_n2774), .B(new_n2772), .Y(new_n2775));
  nand_4 g02399(.A(new_n2773), .B(new_n2771), .Y(new_n2776));
  nand_4 g02400(.A(n7388), .B(n405), .Y(new_n2777));
  not_3  g02401(.A(new_n2777), .Y(new_n2778));
  nand_4 g02402(.A(new_n2778), .B(new_n2776), .Y(new_n2779));
  nand_4 g02403(.A(new_n2779), .B(new_n2775), .Y(new_n2780));
  not_3  g02404(.A(new_n2780), .Y(new_n2781));
  nor_4  g02405(.A(new_n2781), .B(new_n2770), .Y(new_n2782));
  xnor_3 g02406(.A(new_n2781), .B(new_n2770), .Y(new_n2783));
  nor_4  g02407(.A(new_n2754), .B(new_n2753), .Y(new_n2784));
  xnor_3 g02408(.A(new_n2784), .B(new_n2756), .Y(new_n2785));
  nor_4  g02409(.A(new_n2785), .B(new_n2783), .Y(new_n2786));
  nor_4  g02410(.A(new_n2786), .B(new_n2782), .Y(new_n2787));
  nor_4  g02411(.A(new_n2787), .B(new_n2769), .Y(new_n2788));
  nor_4  g02412(.A(new_n2788), .B(new_n2768), .Y(new_n2789));
  nor_4  g02413(.A(new_n2789), .B(new_n2765), .Y(new_n2790));
  not_3  g02414(.A(new_n2790), .Y(new_n2791));
  nand_4 g02415(.A(new_n2745), .B(new_n2742), .Y(new_n2792));
  nor_4  g02416(.A(new_n2744), .B(new_n2743), .Y(new_n2793));
  xnor_3 g02417(.A(new_n2745), .B(new_n2741), .Y(new_n2794));
  not_3  g02418(.A(new_n2764), .Y(new_n2795));
  nand_4 g02419(.A(new_n2795), .B(new_n2794), .Y(new_n2796));
  not_3  g02420(.A(new_n2796), .Y(new_n2797));
  xnor_3 g02421(.A(new_n2797), .B(new_n2793), .Y(new_n2798));
  nand_4 g02422(.A(new_n2798), .B(new_n2792), .Y(new_n2799));
  nor_4  g02423(.A(new_n2724), .B(new_n2723), .Y(new_n2800));
  nand_4 g02424(.A(n2393), .B(n217), .Y(new_n2801));
  xor_3  g02425(.A(new_n2801), .B(new_n2800), .Y(new_n2802_1));
  nand_4 g02426(.A(n3986), .B(n405), .Y(new_n2803));
  not_3  g02427(.A(new_n2803), .Y(new_n2804));
  nand_4 g02428(.A(n5860), .B(n4086), .Y(new_n2805));
  nand_4 g02429(.A(n8433), .B(n5857), .Y(new_n2806));
  xnor_3 g02430(.A(new_n2806), .B(new_n2805), .Y(new_n2807));
  and_4  g02431(.A(new_n2807), .B(new_n2804), .Y(new_n2808));
  nor_4  g02432(.A(new_n2807), .B(new_n2804), .Y(new_n2809));
  nor_4  g02433(.A(new_n2809), .B(new_n2808), .Y(new_n2810));
  xnor_3 g02434(.A(new_n2810), .B(new_n2802_1), .Y(new_n2811));
  not_3  g02435(.A(new_n2811), .Y(new_n2812));
  nand_4 g02436(.A(new_n2740), .B(new_n2730), .Y(new_n2813));
  not_3  g02437(.A(new_n2813), .Y(new_n2814));
  nor_4  g02438(.A(new_n2814), .B(new_n2726), .Y(new_n2815));
  not_3  g02439(.A(new_n2815), .Y(new_n2816));
  nand_4 g02440(.A(n11296), .B(n7965), .Y(new_n2817));
  not_3  g02441(.A(new_n2817), .Y(new_n2818_1));
  nand_4 g02442(.A(n11892), .B(n6611), .Y(new_n2819));
  nand_4 g02443(.A(n7388), .B(n6359), .Y(new_n2820));
  xnor_3 g02444(.A(new_n2820), .B(new_n2819), .Y(new_n2821));
  xor_3  g02445(.A(new_n2821), .B(new_n2818_1), .Y(new_n2822));
  xnor_3 g02446(.A(new_n2822), .B(new_n2816), .Y(new_n2823));
  xnor_3 g02447(.A(new_n2823), .B(new_n2812), .Y(new_n2824));
  xnor_3 g02448(.A(new_n2824), .B(new_n2799), .Y(new_n2825));
  xnor_3 g02449(.A(new_n2825), .B(new_n2791), .Y(new_n2826));
  nand_4 g02450(.A(n7965), .B(n6359), .Y(new_n2827));
  not_3  g02451(.A(new_n2827), .Y(new_n2828));
  not_3  g02452(.A(new_n2765), .Y(new_n2829));
  xnor_3 g02453(.A(new_n2789), .B(new_n2829), .Y(new_n2830));
  nand_4 g02454(.A(new_n2830), .B(new_n2828), .Y(new_n2831));
  nand_4 g02455(.A(new_n2776), .B(new_n2775), .Y(new_n2832));
  not_3  g02456(.A(new_n2832), .Y(new_n2833));
  nand_4 g02457(.A(n8433), .B(n7388), .Y(new_n2834));
  nand_4 g02458(.A(n7965), .B(n405), .Y(new_n2835));
  nor_4  g02459(.A(new_n2835), .B(new_n2834), .Y(new_n2836));
  not_3  g02460(.A(new_n2836), .Y(new_n2837));
  nor_4  g02461(.A(new_n2837), .B(new_n2833), .Y(new_n2838));
  not_3  g02462(.A(new_n2838), .Y(new_n2839));
  xnor_3 g02463(.A(new_n2785), .B(new_n2783), .Y(new_n2840));
  nor_4  g02464(.A(new_n2840), .B(new_n2839), .Y(new_n2841));
  not_3  g02465(.A(new_n2841), .Y(new_n2842));
  xnor_3 g02466(.A(new_n2787), .B(new_n2769), .Y(new_n2843));
  nor_4  g02467(.A(new_n2843), .B(new_n2842), .Y(new_n2844));
  xnor_3 g02468(.A(new_n2830), .B(new_n2827), .Y(new_n2845));
  nand_4 g02469(.A(new_n2845), .B(new_n2844), .Y(new_n2846));
  nand_4 g02470(.A(new_n2846), .B(new_n2831), .Y(new_n2847));
  xnor_3 g02471(.A(new_n2847), .B(new_n2826), .Y(new_n2848));
  xnor_3 g02472(.A(new_n2848), .B(new_n2721), .Y(new_n2849));
  xnor_3 g02473(.A(new_n2702), .B(new_n2700), .Y(new_n2850));
  nor_4  g02474(.A(new_n2850), .B(new_n2716), .Y(new_n2851));
  nor_4  g02475(.A(new_n2718), .B(new_n2717), .Y(new_n2852));
  nor_4  g02476(.A(new_n2852), .B(new_n2851), .Y(new_n2853));
  not_3  g02477(.A(new_n2853), .Y(new_n2854));
  xnor_3 g02478(.A(new_n2845), .B(new_n2844), .Y(new_n2855));
  nand_4 g02479(.A(new_n2855), .B(new_n2854), .Y(new_n2856));
  xnor_3 g02480(.A(new_n2843), .B(new_n2842), .Y(new_n2857));
  not_3  g02481(.A(new_n2857), .Y(new_n2858));
  not_3  g02482(.A(new_n2705), .Y(new_n2859));
  nor_4  g02483(.A(new_n2712), .B(new_n2859), .Y(new_n2860));
  nor_4  g02484(.A(new_n2860), .B(new_n2714), .Y(new_n2861));
  xnor_3 g02485(.A(new_n2840), .B(new_n2839), .Y(new_n2862));
  not_3  g02486(.A(new_n2862), .Y(new_n2863));
  nor_4  g02487(.A(new_n2863), .B(new_n2861), .Y(new_n2864));
  not_3  g02488(.A(new_n2864), .Y(new_n2865));
  nand_4 g02489(.A(n8433), .B(n7965), .Y(new_n2866));
  nor_4  g02490(.A(new_n2866), .B(new_n2707), .Y(new_n2867));
  xnor_3 g02491(.A(new_n2835), .B(new_n2834), .Y(new_n2868));
  not_3  g02492(.A(new_n2868), .Y(new_n2869));
  nor_4  g02493(.A(new_n2869), .B(new_n2867), .Y(new_n2870));
  not_3  g02494(.A(new_n2870), .Y(new_n2871));
  not_3  g02495(.A(new_n2867), .Y(new_n2872));
  nor_4  g02496(.A(new_n2868), .B(new_n2872), .Y(new_n2873));
  nor_4  g02497(.A(new_n2873), .B(new_n2870), .Y(new_n2874));
  nand_4 g02498(.A(n12925), .B(n8476), .Y(new_n2875));
  nand_4 g02499(.A(n7733), .B(n5331), .Y(new_n2876));
  xnor_3 g02500(.A(new_n2876), .B(new_n2875), .Y(new_n2877));
  nand_4 g02501(.A(new_n2877), .B(new_n2874), .Y(new_n2878));
  nand_4 g02502(.A(new_n2878), .B(new_n2871), .Y(new_n2879_1));
  not_3  g02503(.A(new_n2879_1), .Y(new_n2880));
  not_3  g02504(.A(new_n2711), .Y(new_n2881));
  not_3  g02505(.A(new_n2709), .Y(new_n2882));
  nor_4  g02506(.A(new_n2882), .B(new_n2644), .Y(new_n2883));
  nor_4  g02507(.A(new_n2883), .B(new_n2881), .Y(new_n2884));
  nor_4  g02508(.A(new_n2884), .B(new_n2880), .Y(new_n2885));
  not_3  g02509(.A(new_n2885), .Y(new_n2886));
  not_3  g02510(.A(new_n2884), .Y(new_n2887));
  nor_4  g02511(.A(new_n2887), .B(new_n2879_1), .Y(new_n2888));
  nor_4  g02512(.A(new_n2888), .B(new_n2885), .Y(new_n2889));
  not_3  g02513(.A(new_n2866), .Y(new_n2890));
  nor_4  g02514(.A(new_n2890), .B(new_n2777), .Y(new_n2891));
  nor_4  g02515(.A(new_n2891), .B(new_n2833), .Y(new_n2892));
  nor_4  g02516(.A(new_n2890), .B(new_n2779), .Y(new_n2893));
  nor_4  g02517(.A(new_n2893), .B(new_n2892), .Y(new_n2894));
  not_3  g02518(.A(new_n2894), .Y(new_n2895));
  nand_4 g02519(.A(new_n2895), .B(new_n2889), .Y(new_n2896));
  nand_4 g02520(.A(new_n2896), .B(new_n2886), .Y(new_n2897));
  not_3  g02521(.A(new_n2861), .Y(new_n2898));
  nor_4  g02522(.A(new_n2862), .B(new_n2898), .Y(new_n2899));
  nor_4  g02523(.A(new_n2899), .B(new_n2864), .Y(new_n2900));
  nand_4 g02524(.A(new_n2900), .B(new_n2897), .Y(new_n2901));
  nand_4 g02525(.A(new_n2901), .B(new_n2865), .Y(new_n2902_1));
  not_3  g02526(.A(new_n2902_1), .Y(new_n2903));
  nor_4  g02527(.A(new_n2903), .B(new_n2858), .Y(new_n2904));
  nor_4  g02528(.A(new_n2715), .B(new_n2714), .Y(new_n2905));
  nor_4  g02529(.A(new_n2905), .B(new_n2717), .Y(new_n2906));
  xnor_3 g02530(.A(new_n2902_1), .B(new_n2857), .Y(new_n2907));
  nor_4  g02531(.A(new_n2907), .B(new_n2906), .Y(new_n2908));
  nor_4  g02532(.A(new_n2908), .B(new_n2904), .Y(new_n2909));
  not_3  g02533(.A(new_n2909), .Y(new_n2910));
  xnor_3 g02534(.A(new_n2855), .B(new_n2853), .Y(new_n2911));
  nand_4 g02535(.A(new_n2911), .B(new_n2910), .Y(new_n2912));
  nand_4 g02536(.A(new_n2912), .B(new_n2856), .Y(new_n2913));
  xnor_3 g02537(.A(new_n2913), .B(new_n2849), .Y(new_n2914));
  not_3  g02538(.A(new_n2914), .Y(new_n2915));
  nand_4 g02539(.A(new_n2915), .B(new_n2590), .Y(new_n2916));
  xnor_3 g02540(.A(new_n2914), .B(new_n2590), .Y(new_n2917));
  not_3  g02541(.A(new_n2556), .Y(new_n2918));
  xnor_3 g02542(.A(new_n2557), .B(new_n2918), .Y(new_n2919));
  xnor_3 g02543(.A(new_n2911), .B(new_n2910), .Y(new_n2920));
  nor_4  g02544(.A(new_n2920), .B(new_n2919), .Y(new_n2921));
  not_3  g02545(.A(new_n2921), .Y(new_n2922));
  not_3  g02546(.A(new_n2919), .Y(new_n2923));
  xnor_3 g02547(.A(new_n2911), .B(new_n2909), .Y(new_n2924));
  nor_4  g02548(.A(new_n2924), .B(new_n2923), .Y(new_n2925));
  nor_4  g02549(.A(new_n2925), .B(new_n2921), .Y(new_n2926));
  xnor_3 g02550(.A(new_n2554), .B(new_n2552), .Y(new_n2927));
  xnor_3 g02551(.A(new_n2907), .B(new_n2906), .Y(new_n2928));
  not_3  g02552(.A(new_n2928), .Y(new_n2929));
  nor_4  g02553(.A(new_n2929), .B(new_n2927), .Y(new_n2930));
  not_3  g02554(.A(new_n2930), .Y(new_n2931));
  xnor_3 g02555(.A(new_n2928), .B(new_n2927), .Y(new_n2932));
  not_3  g02556(.A(new_n2551_1), .Y(new_n2933));
  xor_3  g02557(.A(new_n2933), .B(new_n2550), .Y(new_n2934));
  not_3  g02558(.A(new_n2901), .Y(new_n2935));
  nor_4  g02559(.A(new_n2900), .B(new_n2897), .Y(new_n2936));
  nor_4  g02560(.A(new_n2936), .B(new_n2935), .Y(new_n2937));
  nor_4  g02561(.A(new_n2937), .B(new_n2934), .Y(new_n2938));
  not_3  g02562(.A(new_n2938), .Y(new_n2939));
  xnor_3 g02563(.A(new_n2937), .B(new_n2934), .Y(new_n2940));
  xnor_3 g02564(.A(new_n2895), .B(new_n2889), .Y(new_n2941));
  not_3  g02565(.A(new_n2941), .Y(new_n2942));
  not_3  g02566(.A(new_n2544), .Y(new_n2943));
  nand_4 g02567(.A(n8759), .B(n3719), .Y(new_n2944));
  not_3  g02568(.A(new_n2944), .Y(new_n2945));
  nor_4  g02569(.A(new_n2945), .B(new_n2526), .Y(new_n2946));
  not_3  g02570(.A(new_n2946), .Y(new_n2947));
  nand_4 g02571(.A(new_n2947), .B(new_n2943), .Y(new_n2948));
  nand_4 g02572(.A(new_n2946), .B(new_n2525), .Y(new_n2949));
  nand_4 g02573(.A(new_n2949), .B(new_n2948), .Y(new_n2950));
  nor_4  g02574(.A(new_n2950), .B(new_n2942), .Y(new_n2951));
  not_3  g02575(.A(new_n2950), .Y(new_n2952));
  nor_4  g02576(.A(new_n2952), .B(new_n2941), .Y(new_n2953));
  nor_4  g02577(.A(new_n2953), .B(new_n2951), .Y(new_n2954));
  not_3  g02578(.A(new_n2954), .Y(new_n2955));
  xor_3  g02579(.A(new_n2877), .B(new_n2874), .Y(new_n2956));
  xor_3  g02580(.A(new_n2546), .B(new_n2545), .Y(new_n2957));
  not_3  g02581(.A(new_n2957), .Y(new_n2958));
  nor_4  g02582(.A(new_n2958), .B(new_n2956), .Y(new_n2959));
  xor_3  g02583(.A(new_n2890), .B(new_n2707), .Y(new_n2960));
  nor_4  g02584(.A(new_n2960), .B(new_n2944), .Y(new_n2961));
  not_3  g02585(.A(new_n2961), .Y(new_n2962));
  not_3  g02586(.A(new_n2956), .Y(new_n2963));
  xor_3  g02587(.A(new_n2958), .B(new_n2963), .Y(new_n2964));
  nor_4  g02588(.A(new_n2964), .B(new_n2962), .Y(new_n2965));
  nor_4  g02589(.A(new_n2965), .B(new_n2959), .Y(new_n2966));
  nor_4  g02590(.A(new_n2966), .B(new_n2955), .Y(new_n2967));
  nor_4  g02591(.A(new_n2967), .B(new_n2951), .Y(new_n2968));
  nor_4  g02592(.A(new_n2968), .B(new_n2940), .Y(new_n2969));
  not_3  g02593(.A(new_n2969), .Y(new_n2970));
  nand_4 g02594(.A(new_n2970), .B(new_n2939), .Y(new_n2971));
  nand_4 g02595(.A(new_n2971), .B(new_n2932), .Y(new_n2972));
  nand_4 g02596(.A(new_n2972), .B(new_n2931), .Y(new_n2973));
  not_3  g02597(.A(new_n2973), .Y(new_n2974));
  nand_4 g02598(.A(new_n2974), .B(new_n2926), .Y(new_n2975));
  nand_4 g02599(.A(new_n2975), .B(new_n2922), .Y(new_n2976));
  not_3  g02600(.A(new_n2976), .Y(new_n2977));
  nand_4 g02601(.A(new_n2977), .B(new_n2917), .Y(new_n2978));
  nand_4 g02602(.A(new_n2978), .B(new_n2916), .Y(new_n2979));
  xnor_3 g02603(.A(new_n2979), .B(new_n2459), .Y(new_n2980));
  not_3  g02604(.A(new_n2980), .Y(new_n2981));
  xnor_3 g02605(.A(new_n2422), .B(new_n2399), .Y(new_n2982));
  not_3  g02606(.A(new_n2982), .Y(new_n2983));
  nand_4 g02607(.A(n5305), .B(n2577), .Y(new_n2984));
  not_3  g02608(.A(new_n2984), .Y(new_n2985));
  xnor_3 g02609(.A(new_n2420), .B(new_n2415), .Y(new_n2986));
  not_3  g02610(.A(new_n2986), .Y(new_n2987));
  nor_4  g02611(.A(new_n2987), .B(new_n2985), .Y(new_n2988));
  not_3  g02612(.A(new_n2988), .Y(new_n2989));
  nor_4  g02613(.A(new_n2986), .B(new_n2984), .Y(new_n2990));
  nor_4  g02614(.A(new_n2990), .B(new_n2988), .Y(new_n2991));
  nand_4 g02615(.A(n5305), .B(n3842), .Y(new_n2992));
  nand_4 g02616(.A(n9956), .B(n1097), .Y(new_n2993));
  not_3  g02617(.A(new_n2993), .Y(new_n2994));
  nand_4 g02618(.A(n11917), .B(n5305), .Y(new_n2995));
  not_3  g02619(.A(new_n2995), .Y(new_n2996));
  nand_4 g02620(.A(new_n2996), .B(new_n2994), .Y(new_n2997));
  nand_4 g02621(.A(new_n2995), .B(new_n2993), .Y(new_n2998));
  nand_4 g02622(.A(n5964), .B(n4921), .Y(new_n2999));
  not_3  g02623(.A(new_n2999), .Y(new_n3000));
  nand_4 g02624(.A(new_n3000), .B(new_n2998), .Y(new_n3001));
  nand_4 g02625(.A(new_n3001), .B(new_n2997), .Y(new_n3002));
  not_3  g02626(.A(new_n3002), .Y(new_n3003));
  nor_4  g02627(.A(new_n3003), .B(new_n2992), .Y(new_n3004));
  not_3  g02628(.A(new_n2992), .Y(new_n3005));
  xnor_3 g02629(.A(new_n3002), .B(new_n3005), .Y(new_n3006));
  nor_4  g02630(.A(new_n2407), .B(new_n2406), .Y(new_n3007));
  xnor_3 g02631(.A(new_n3007), .B(new_n2409), .Y(new_n3008));
  nor_4  g02632(.A(new_n3008), .B(new_n3006), .Y(new_n3009));
  nor_4  g02633(.A(new_n3009), .B(new_n3004), .Y(new_n3010));
  nand_4 g02634(.A(new_n3010), .B(new_n2991), .Y(new_n3011));
  nand_4 g02635(.A(new_n3011), .B(new_n2989), .Y(new_n3012));
  nor_4  g02636(.A(new_n3012), .B(new_n2983), .Y(new_n3013));
  not_3  g02637(.A(new_n3013), .Y(new_n3014));
  xnor_3 g02638(.A(new_n2457), .B(new_n2453), .Y(new_n3015));
  xnor_3 g02639(.A(new_n3015), .B(new_n3014), .Y(new_n3016));
  nand_4 g02640(.A(n9637), .B(n5305), .Y(new_n3017));
  not_3  g02641(.A(new_n3017), .Y(new_n3018));
  not_3  g02642(.A(new_n3012), .Y(new_n3019));
  nor_4  g02643(.A(new_n3019), .B(new_n2982), .Y(new_n3020));
  nor_4  g02644(.A(new_n3020), .B(new_n3013), .Y(new_n3021));
  nand_4 g02645(.A(new_n3021), .B(new_n3018), .Y(new_n3022_1));
  and_4  g02646(.A(new_n2998), .B(new_n2997), .Y(new_n3023));
  nand_4 g02647(.A(n9956), .B(n5964), .Y(new_n3024));
  nand_4 g02648(.A(n5305), .B(n4921), .Y(new_n3025));
  nor_4  g02649(.A(new_n3025), .B(new_n3024), .Y(new_n3026));
  not_3  g02650(.A(new_n3026), .Y(new_n3027));
  nor_4  g02651(.A(new_n3027), .B(new_n3023), .Y(new_n3028));
  xor_3  g02652(.A(new_n3008), .B(new_n3006), .Y(new_n3029));
  nand_4 g02653(.A(new_n3029), .B(new_n3028), .Y(new_n3030));
  not_3  g02654(.A(new_n3011), .Y(new_n3031));
  nor_4  g02655(.A(new_n3010), .B(new_n2991), .Y(new_n3032));
  nor_4  g02656(.A(new_n3032), .B(new_n3031), .Y(new_n3033));
  nor_4  g02657(.A(new_n3033), .B(new_n3030), .Y(new_n3034));
  xnor_3 g02658(.A(new_n3021), .B(new_n3017), .Y(new_n3035));
  nand_4 g02659(.A(new_n3035), .B(new_n3034), .Y(new_n3036));
  nand_4 g02660(.A(new_n3036), .B(new_n3022_1), .Y(new_n3037));
  xnor_3 g02661(.A(new_n3037), .B(new_n3016), .Y(new_n3038));
  not_3  g02662(.A(new_n3038), .Y(new_n3039));
  xnor_3 g02663(.A(new_n2976), .B(new_n2917), .Y(new_n3040));
  nor_4  g02664(.A(new_n3040), .B(new_n3039), .Y(new_n3041));
  not_3  g02665(.A(new_n3041), .Y(new_n3042));
  nand_4 g02666(.A(new_n3040), .B(new_n3039), .Y(new_n3043));
  xor_3  g02667(.A(new_n3035), .B(new_n3034), .Y(new_n3044));
  not_3  g02668(.A(new_n3044), .Y(new_n3045));
  xnor_3 g02669(.A(new_n2974), .B(new_n2926), .Y(new_n3046));
  not_3  g02670(.A(new_n3046), .Y(new_n3047));
  nand_4 g02671(.A(new_n3047), .B(new_n3045), .Y(new_n3048));
  nand_4 g02672(.A(new_n3046), .B(new_n3044), .Y(new_n3049));
  xor_3  g02673(.A(new_n3033), .B(new_n3030), .Y(new_n3050));
  not_3  g02674(.A(new_n3050), .Y(new_n3051));
  xnor_3 g02675(.A(new_n2971), .B(new_n2932), .Y(new_n3052));
  nand_4 g02676(.A(new_n3052), .B(new_n3051), .Y(new_n3053));
  not_3  g02677(.A(new_n3053), .Y(new_n3054));
  nor_4  g02678(.A(new_n3052), .B(new_n3051), .Y(new_n3055));
  nor_4  g02679(.A(new_n3055), .B(new_n3054), .Y(new_n3056));
  not_3  g02680(.A(new_n3029), .Y(new_n3057));
  xor_3  g02681(.A(new_n3057), .B(new_n3028), .Y(new_n3058));
  xnor_3 g02682(.A(new_n2968), .B(new_n2940), .Y(new_n3059));
  nand_4 g02683(.A(new_n3059), .B(new_n3058), .Y(new_n3060));
  xnor_3 g02684(.A(new_n2966), .B(new_n2955), .Y(new_n3061));
  not_3  g02685(.A(new_n3023), .Y(new_n3062));
  nand_4 g02686(.A(n9956), .B(n5305), .Y(new_n3063));
  not_3  g02687(.A(new_n3063), .Y(new_n3064));
  nor_4  g02688(.A(new_n3064), .B(new_n2999), .Y(new_n3065));
  not_3  g02689(.A(new_n3065), .Y(new_n3066));
  nand_4 g02690(.A(new_n3066), .B(new_n3062), .Y(new_n3067));
  nand_4 g02691(.A(new_n3065), .B(new_n2998), .Y(new_n3068));
  nand_4 g02692(.A(new_n3068), .B(new_n3067), .Y(new_n3069));
  nand_4 g02693(.A(new_n3069), .B(new_n3061), .Y(new_n3070));
  not_3  g02694(.A(new_n3070), .Y(new_n3071_1));
  nor_4  g02695(.A(new_n3069), .B(new_n3061), .Y(new_n3072));
  nor_4  g02696(.A(new_n3072), .B(new_n3071_1), .Y(new_n3073));
  xor_3  g02697(.A(new_n2960), .B(new_n2944), .Y(new_n3074));
  nand_4 g02698(.A(new_n3074), .B(new_n3064), .Y(new_n3075));
  not_3  g02699(.A(new_n3075), .Y(new_n3076));
  xor_3  g02700(.A(new_n3025), .B(new_n3024), .Y(new_n3077));
  or_4   g02701(.A(new_n3077), .B(new_n3076), .Y(new_n3078));
  xnor_3 g02702(.A(new_n2964), .B(new_n2962), .Y(new_n3079));
  xor_3  g02703(.A(new_n3077), .B(new_n3076), .Y(new_n3080));
  nand_4 g02704(.A(new_n3080), .B(new_n3079), .Y(new_n3081));
  nand_4 g02705(.A(new_n3081), .B(new_n3078), .Y(new_n3082));
  nand_4 g02706(.A(new_n3082), .B(new_n3073), .Y(new_n3083));
  nand_4 g02707(.A(new_n3083), .B(new_n3070), .Y(new_n3084));
  not_3  g02708(.A(new_n3060), .Y(new_n3085));
  nor_4  g02709(.A(new_n3059), .B(new_n3058), .Y(new_n3086));
  nor_4  g02710(.A(new_n3086), .B(new_n3085), .Y(new_n3087));
  nand_4 g02711(.A(new_n3087), .B(new_n3084), .Y(new_n3088));
  nand_4 g02712(.A(new_n3088), .B(new_n3060), .Y(new_n3089));
  nand_4 g02713(.A(new_n3089), .B(new_n3056), .Y(new_n3090));
  nand_4 g02714(.A(new_n3090), .B(new_n3053), .Y(new_n3091));
  nand_4 g02715(.A(new_n3091), .B(new_n3049), .Y(new_n3092));
  nand_4 g02716(.A(new_n3092), .B(new_n3048), .Y(new_n3093));
  nand_4 g02717(.A(new_n3093), .B(new_n3043), .Y(new_n3094));
  nand_4 g02718(.A(new_n3094), .B(new_n3042), .Y(new_n3095));
  xnor_3 g02719(.A(new_n3095), .B(new_n2981), .Y(new_n3096));
  nand_4 g02720(.A(n11536), .B(n5305), .Y(new_n3097));
  not_3  g02721(.A(new_n3097), .Y(new_n3098));
  nand_4 g02722(.A(n10545), .B(n7610), .Y(new_n3099));
  nand_4 g02723(.A(n7690), .B(n4826), .Y(new_n3100));
  not_3  g02724(.A(new_n3100), .Y(new_n3101));
  xor_3  g02725(.A(new_n3101), .B(new_n3099), .Y(new_n3102));
  nand_4 g02726(.A(new_n2848), .B(new_n2721), .Y(new_n3103));
  not_3  g02727(.A(new_n2849), .Y(new_n3104));
  nand_4 g02728(.A(new_n2913), .B(new_n3104), .Y(new_n3105));
  nand_4 g02729(.A(new_n3105), .B(new_n3103), .Y(new_n3106));
  nand_4 g02730(.A(n10510), .B(n3602), .Y(new_n3107));
  nand_4 g02731(.A(new_n2507_1), .B(new_n2585_1), .Y(new_n3108));
  not_3  g02732(.A(new_n2582), .Y(new_n3109));
  nand_4 g02733(.A(new_n2587), .B(new_n3109), .Y(new_n3110));
  nand_4 g02734(.A(new_n3110), .B(new_n3108), .Y(new_n3111));
  xnor_3 g02735(.A(new_n3111), .B(new_n3107), .Y(new_n3112));
  nor_4  g02736(.A(new_n2569), .B(new_n2562), .Y(new_n3113));
  not_3  g02737(.A(new_n2570), .Y(new_n3114));
  nor_4  g02738(.A(new_n2581_1), .B(new_n3114), .Y(new_n3115));
  nor_4  g02739(.A(new_n3115), .B(new_n3113), .Y(new_n3116));
  nor_4  g02740(.A(new_n2573), .B(new_n2572), .Y(new_n3117));
  not_3  g02741(.A(new_n2574), .Y(new_n3118));
  nor_4  g02742(.A(new_n2580), .B(new_n3118), .Y(new_n3119));
  nor_4  g02743(.A(new_n3119), .B(new_n3117), .Y(new_n3120));
  not_3  g02744(.A(new_n2564_1), .Y(new_n3121));
  nor_4  g02745(.A(new_n2566), .B(new_n3121), .Y(new_n3122));
  not_3  g02746(.A(new_n2563), .Y(new_n3123));
  nor_4  g02747(.A(new_n2567), .B(new_n3123), .Y(new_n3124_1));
  nor_4  g02748(.A(new_n3124_1), .B(new_n3122), .Y(new_n3125));
  nand_4 g02749(.A(n10439), .B(n7436), .Y(new_n3126));
  not_3  g02750(.A(new_n3126), .Y(new_n3127));
  nand_4 g02751(.A(n10391), .B(n6776), .Y(new_n3128));
  nand_4 g02752(.A(n8595), .B(n8276), .Y(new_n3129));
  xor_3  g02753(.A(new_n3129), .B(new_n3128), .Y(new_n3130));
  xnor_3 g02754(.A(new_n3130), .B(new_n3127), .Y(new_n3131));
  xnor_3 g02755(.A(new_n3131), .B(new_n3125), .Y(new_n3132));
  xnor_3 g02756(.A(new_n3132), .B(new_n3120), .Y(new_n3133));
  nor_4  g02757(.A(new_n2578), .B(new_n2577_1), .Y(new_n3134));
  nand_4 g02758(.A(new_n2578), .B(new_n2577_1), .Y(new_n3135));
  nand_4 g02759(.A(new_n3135), .B(new_n2576), .Y(new_n3136));
  not_3  g02760(.A(new_n3136), .Y(new_n3137));
  or_4   g02761(.A(new_n3137), .B(new_n3134), .Y(new_n3138));
  nand_4 g02762(.A(n9241), .B(n6126), .Y(new_n3139));
  nand_4 g02763(.A(n12299), .B(n8065), .Y(new_n3140));
  xor_3  g02764(.A(new_n3140), .B(new_n3139), .Y(new_n3141));
  nand_4 g02765(.A(n10644), .B(n3719), .Y(new_n3142));
  nand_4 g02766(.A(n8759), .B(n4190), .Y(new_n3143));
  xor_3  g02767(.A(new_n3143), .B(new_n3142), .Y(new_n3144));
  xnor_3 g02768(.A(new_n3144), .B(new_n3141), .Y(new_n3145));
  xnor_3 g02769(.A(new_n3145), .B(new_n3138), .Y(new_n3146_1));
  xnor_3 g02770(.A(new_n3146_1), .B(new_n3133), .Y(new_n3147));
  xnor_3 g02771(.A(new_n3147), .B(new_n3116), .Y(new_n3148));
  nand_4 g02772(.A(new_n2797), .B(new_n2793), .Y(new_n3149));
  not_3  g02773(.A(new_n2824), .Y(new_n3150));
  nand_4 g02774(.A(new_n3150), .B(new_n2799), .Y(new_n3151));
  nand_4 g02775(.A(new_n3151), .B(new_n3149), .Y(new_n3152));
  not_3  g02776(.A(new_n2430), .Y(new_n3153));
  nand_4 g02777(.A(new_n2436), .B(new_n3153), .Y(new_n3154));
  nand_4 g02778(.A(new_n2452), .B(new_n2437), .Y(new_n3155));
  nand_4 g02779(.A(new_n3155), .B(new_n3154), .Y(new_n3156));
  nand_4 g02780(.A(n11257), .B(n4921), .Y(new_n3157));
  nand_4 g02781(.A(n5964), .B(n1835), .Y(new_n3158));
  xor_3  g02782(.A(new_n3158), .B(new_n3157), .Y(new_n3159));
  nand_4 g02783(.A(n4312), .B(n2577), .Y(new_n3160));
  nand_4 g02784(.A(n12025), .B(n11917), .Y(new_n3161));
  xor_3  g02785(.A(new_n3161), .B(new_n3160), .Y(new_n3162));
  xnor_3 g02786(.A(new_n3162), .B(new_n3159), .Y(new_n3163));
  and_4  g02787(.A(new_n2447), .B(new_n2446), .Y(new_n3164));
  nor_4  g02788(.A(new_n2450), .B(new_n3164), .Y(new_n3165));
  and_4  g02789(.A(new_n2434_1), .B(new_n2433_1), .Y(new_n3166));
  nor_4  g02790(.A(new_n2435), .B(new_n2432), .Y(new_n3167));
  nor_4  g02791(.A(new_n3167), .B(new_n3166), .Y(new_n3168));
  xnor_3 g02792(.A(new_n3168), .B(new_n3165), .Y(new_n3169));
  xnor_3 g02793(.A(new_n3169), .B(new_n3163), .Y(new_n3170));
  nand_4 g02794(.A(new_n2441), .B(new_n2440), .Y(new_n3171));
  nand_4 g02795(.A(new_n2451), .B(new_n2442), .Y(new_n3172_1));
  nand_4 g02796(.A(new_n3172_1), .B(new_n3171), .Y(new_n3173));
  nand_4 g02797(.A(n9637), .B(n1097), .Y(new_n3174));
  xnor_3 g02798(.A(new_n3174), .B(new_n3173), .Y(new_n3175));
  xnor_3 g02799(.A(new_n3175), .B(new_n3170), .Y(new_n3176));
  xnor_3 g02800(.A(new_n3176), .B(new_n3156), .Y(new_n3177));
  nand_4 g02801(.A(n4086), .B(n3986), .Y(new_n3178));
  nand_4 g02802(.A(n12705), .B(n3842), .Y(new_n3179));
  not_3  g02803(.A(new_n3179), .Y(new_n3180));
  xor_3  g02804(.A(new_n3180), .B(new_n3178), .Y(new_n3181));
  xnor_3 g02805(.A(new_n3181), .B(new_n3177), .Y(new_n3182));
  xnor_3 g02806(.A(new_n3182), .B(new_n3152), .Y(new_n3183));
  xnor_3 g02807(.A(new_n3183), .B(new_n3148), .Y(new_n3184));
  xnor_3 g02808(.A(new_n3184), .B(new_n3112), .Y(new_n3185));
  xnor_3 g02809(.A(new_n3185), .B(new_n3106), .Y(new_n3186));
  nand_4 g02810(.A(new_n2588), .B(new_n2539), .Y(new_n3187));
  not_3  g02811(.A(new_n2589), .Y(new_n3188));
  nand_4 g02812(.A(new_n3188), .B(new_n2559), .Y(new_n3189));
  nand_4 g02813(.A(new_n3189), .B(new_n3187), .Y(new_n3190));
  not_3  g02814(.A(new_n2697), .Y(new_n3191));
  nand_4 g02815(.A(new_n3191), .B(new_n2666), .Y(new_n3192));
  nand_4 g02816(.A(new_n2720), .B(new_n2698), .Y(new_n3193));
  nand_4 g02817(.A(new_n3193), .B(new_n3192), .Y(new_n3194));
  xnor_3 g02818(.A(new_n3194), .B(new_n3190), .Y(new_n3195));
  nand_4 g02819(.A(n8433), .B(n45), .Y(new_n3196));
  not_3  g02820(.A(new_n3196), .Y(new_n3197));
  nand_4 g02821(.A(n5857), .B(n405), .Y(new_n3198));
  nand_4 g02822(.A(n7965), .B(n1357), .Y(new_n3199));
  xor_3  g02823(.A(new_n3199), .B(new_n3198), .Y(new_n3200));
  xor_3  g02824(.A(new_n3200), .B(new_n3197), .Y(new_n3201));
  and_4  g02825(.A(new_n2820), .B(new_n2819), .Y(new_n3202));
  nor_4  g02826(.A(new_n2821), .B(new_n2818_1), .Y(new_n3203));
  nor_4  g02827(.A(new_n3203), .B(new_n3202), .Y(new_n3204));
  and_4  g02828(.A(new_n2806), .B(new_n2805), .Y(new_n3205));
  nor_4  g02829(.A(new_n2809), .B(new_n3205), .Y(new_n3206));
  xnor_3 g02830(.A(new_n3206), .B(new_n3204), .Y(new_n3207));
  nand_4 g02831(.A(n10965), .B(n8476), .Y(new_n3208));
  and_4  g02832(.A(new_n2691), .B(new_n2690), .Y(new_n3209));
  nor_4  g02833(.A(new_n2692), .B(new_n2689), .Y(new_n3210));
  nor_4  g02834(.A(new_n3210), .B(new_n3209), .Y(new_n3211));
  xnor_3 g02835(.A(new_n3211), .B(new_n3208), .Y(new_n3212));
  xnor_3 g02836(.A(new_n3212), .B(new_n3207), .Y(new_n3213));
  nand_4 g02837(.A(new_n2685), .B(new_n2683), .Y(new_n3214_1));
  nand_4 g02838(.A(new_n2693), .B(new_n2686), .Y(new_n3215));
  nand_4 g02839(.A(new_n3215), .B(new_n3214_1), .Y(new_n3216));
  nand_4 g02840(.A(n5860), .B(n217), .Y(new_n3217));
  nand_4 g02841(.A(n6611), .B(n2393), .Y(new_n3218));
  not_3  g02842(.A(new_n3218), .Y(new_n3219));
  xor_3  g02843(.A(new_n3219), .B(new_n3217), .Y(new_n3220));
  nand_4 g02844(.A(n7546), .B(n5331), .Y(new_n3221));
  nand_4 g02845(.A(n12925), .B(n4499), .Y(new_n3222));
  xnor_3 g02846(.A(new_n3222), .B(new_n3221), .Y(new_n3223));
  nand_4 g02847(.A(n11892), .B(n6359), .Y(new_n3224));
  nand_4 g02848(.A(n11296), .B(n7388), .Y(new_n3225));
  xnor_3 g02849(.A(new_n3225), .B(new_n3224), .Y(new_n3226));
  xnor_3 g02850(.A(new_n3226), .B(new_n3223), .Y(new_n3227));
  xnor_3 g02851(.A(new_n3227), .B(new_n3220), .Y(new_n3228));
  xnor_3 g02852(.A(new_n3228), .B(new_n3216), .Y(new_n3229));
  xnor_3 g02853(.A(new_n3229), .B(new_n3213), .Y(new_n3230_1));
  nand_4 g02854(.A(n2530), .B(n503), .Y(new_n3231));
  not_3  g02855(.A(new_n2800), .Y(new_n3232));
  nor_4  g02856(.A(new_n2801), .B(new_n3232), .Y(new_n3233));
  nor_4  g02857(.A(new_n2810), .B(new_n2802_1), .Y(new_n3234));
  nor_4  g02858(.A(new_n3234), .B(new_n3233), .Y(new_n3235));
  and_4  g02859(.A(new_n2679_1), .B(new_n2678), .Y(new_n3236));
  not_3  g02860(.A(new_n2677), .Y(new_n3237));
  nor_4  g02861(.A(new_n2680), .B(new_n3237), .Y(new_n3238));
  nor_4  g02862(.A(new_n3238), .B(new_n3236), .Y(new_n3239));
  nand_4 g02863(.A(n7733), .B(n3616), .Y(new_n3240));
  nand_4 g02864(.A(n12648), .B(n4970), .Y(new_n3241));
  not_3  g02865(.A(new_n3241), .Y(new_n3242));
  xor_3  g02866(.A(new_n3242), .B(new_n3240), .Y(new_n3243));
  xnor_3 g02867(.A(new_n3243), .B(new_n3239), .Y(new_n3244));
  xnor_3 g02868(.A(new_n3244), .B(new_n3235), .Y(new_n3245));
  xnor_3 g02869(.A(new_n3245), .B(new_n3231), .Y(new_n3246));
  xnor_3 g02870(.A(new_n3246), .B(new_n3230_1), .Y(new_n3247));
  nand_4 g02871(.A(new_n2822), .B(new_n2815), .Y(new_n3248));
  nand_4 g02872(.A(new_n2823), .B(new_n2811), .Y(new_n3249));
  nand_4 g02873(.A(new_n3249), .B(new_n3248), .Y(new_n3250));
  nand_4 g02874(.A(new_n2681), .B(new_n2676), .Y(new_n3251));
  not_3  g02875(.A(new_n2682), .Y(new_n3252));
  nand_4 g02876(.A(new_n2695), .B(new_n3252), .Y(new_n3253));
  nand_4 g02877(.A(new_n3253), .B(new_n3251), .Y(new_n3254));
  xnor_3 g02878(.A(new_n3254), .B(new_n3250), .Y(new_n3255));
  xnor_3 g02879(.A(new_n3255), .B(new_n3247), .Y(new_n3256));
  nand_4 g02880(.A(new_n2671), .B(new_n2669), .Y(new_n3257));
  nand_4 g02881(.A(new_n2696), .B(new_n2673), .Y(new_n3258));
  nand_4 g02882(.A(new_n3258), .B(new_n3257), .Y(new_n3259));
  nand_4 g02883(.A(n10547), .B(n9956), .Y(new_n3260));
  not_3  g02884(.A(new_n3260), .Y(new_n3261));
  xnor_3 g02885(.A(new_n3261), .B(new_n3259), .Y(new_n3262));
  xnor_3 g02886(.A(new_n3262), .B(new_n3256), .Y(new_n3263));
  xnor_3 g02887(.A(new_n3263), .B(new_n3201), .Y(new_n3264));
  nand_4 g02888(.A(new_n3015), .B(new_n3013), .Y(new_n3265));
  nand_4 g02889(.A(new_n3037), .B(new_n3016), .Y(new_n3266));
  nand_4 g02890(.A(new_n3266), .B(new_n3265), .Y(new_n3267));
  nand_4 g02891(.A(new_n2825), .B(new_n2790), .Y(new_n3268));
  nand_4 g02892(.A(new_n2847), .B(new_n2826), .Y(new_n3269));
  nand_4 g02893(.A(new_n3269), .B(new_n3268), .Y(new_n3270));
  xnor_3 g02894(.A(new_n3270), .B(new_n3267), .Y(new_n3271));
  xnor_3 g02895(.A(new_n3271), .B(new_n3264), .Y(new_n3272_1));
  xnor_3 g02896(.A(new_n3272_1), .B(new_n3195), .Y(new_n3273));
  xnor_3 g02897(.A(new_n3273), .B(new_n3186), .Y(new_n3274));
  xnor_3 g02898(.A(new_n3274), .B(new_n3102), .Y(new_n3275));
  xnor_3 g02899(.A(new_n3275), .B(new_n3098), .Y(new_n3276));
  nand_4 g02900(.A(new_n3276), .B(new_n3096), .Y(new_n3277));
  xnor_3 g02901(.A(new_n3095), .B(new_n2980), .Y(new_n3278));
  xnor_3 g02902(.A(new_n3275), .B(new_n3097), .Y(new_n3279));
  nand_4 g02903(.A(new_n3279), .B(new_n3278), .Y(new_n3280));
  nand_4 g02904(.A(new_n3280), .B(new_n3277), .Y(n837));
  nand_4 g02905(.A(n11917), .B(n11757), .Y(new_n3282));
  not_3  g02906(.A(new_n3282), .Y(new_n3283));
  nand_4 g02907(.A(n9956), .B(n5240), .Y(new_n3284));
  nand_4 g02908(.A(n11757), .B(n4921), .Y(new_n3285));
  not_3  g02909(.A(new_n3285), .Y(new_n3286));
  nand_4 g02910(.A(n11917), .B(n3172), .Y(new_n3287_1));
  xnor_3 g02911(.A(new_n3287_1), .B(new_n3284), .Y(new_n3288));
  nor_4  g02912(.A(new_n3288), .B(new_n3286), .Y(new_n3289));
  nor_4  g02913(.A(new_n3289), .B(new_n3284), .Y(new_n3290));
  nor_4  g02914(.A(new_n3290), .B(new_n3283), .Y(new_n3291));
  nand_4 g02915(.A(n4921), .B(n3172), .Y(new_n3292));
  not_3  g02916(.A(new_n3292), .Y(new_n3293));
  nor_4  g02917(.A(new_n3293), .B(new_n3290), .Y(new_n3294));
  nor_4  g02918(.A(new_n3294), .B(new_n3282), .Y(new_n3295));
  nor_4  g02919(.A(new_n3295), .B(new_n3291), .Y(new_n3296));
  nand_4 g02920(.A(n5240), .B(n4921), .Y(new_n3297));
  nand_4 g02921(.A(n11821), .B(n9956), .Y(new_n3298));
  xor_3  g02922(.A(new_n3298), .B(new_n3297), .Y(new_n3299));
  xnor_3 g02923(.A(new_n3299), .B(new_n3296), .Y(new_n3300));
  not_3  g02924(.A(new_n3300), .Y(new_n3301));
  nand_4 g02925(.A(n2577), .B(n1333), .Y(new_n3302));
  nand_4 g02926(.A(n3842), .B(n3172), .Y(new_n3303));
  xor_3  g02927(.A(new_n3303), .B(new_n3302), .Y(new_n3304));
  xnor_3 g02928(.A(new_n3304), .B(new_n3301), .Y(new_n3305));
  nand_4 g02929(.A(n3842), .B(n1333), .Y(new_n3306));
  not_3  g02930(.A(new_n3306), .Y(new_n3307));
  nand_4 g02931(.A(n11757), .B(n9956), .Y(new_n3308));
  not_3  g02932(.A(new_n3308), .Y(new_n3309));
  nand_4 g02933(.A(n11917), .B(n1333), .Y(new_n3310));
  not_3  g02934(.A(new_n3310), .Y(new_n3311));
  nor_4  g02935(.A(new_n3311), .B(new_n3309), .Y(new_n3312));
  nor_4  g02936(.A(new_n3310), .B(new_n3308), .Y(new_n3313));
  nor_4  g02937(.A(new_n3313), .B(new_n3293), .Y(new_n3314));
  nor_4  g02938(.A(new_n3314), .B(new_n3312), .Y(new_n3315));
  and_4  g02939(.A(new_n3315), .B(new_n3307), .Y(new_n3316));
  not_3  g02940(.A(new_n3288), .Y(new_n3317));
  nor_4  g02941(.A(new_n3317), .B(new_n3285), .Y(new_n3318));
  nor_4  g02942(.A(new_n3318), .B(new_n3289), .Y(new_n3319));
  xnor_3 g02943(.A(new_n3315), .B(new_n3307), .Y(new_n3320));
  nor_4  g02944(.A(new_n3320), .B(new_n3319), .Y(new_n3321));
  nor_4  g02945(.A(new_n3321), .B(new_n3316), .Y(new_n3322));
  xnor_3 g02946(.A(new_n3322), .B(new_n3305), .Y(new_n3323));
  not_3  g02947(.A(new_n3323), .Y(new_n3324));
  nand_4 g02948(.A(n7862), .B(n2577), .Y(new_n3325));
  xnor_3 g02949(.A(new_n3320), .B(new_n3319), .Y(new_n3326));
  nor_4  g02950(.A(new_n3326), .B(new_n3325), .Y(new_n3327));
  not_3  g02951(.A(new_n3327), .Y(new_n3328));
  nand_4 g02952(.A(n7862), .B(n3842), .Y(new_n3329));
  nand_4 g02953(.A(n9956), .B(n3172), .Y(new_n3330));
  not_3  g02954(.A(new_n3330), .Y(new_n3331));
  nand_4 g02955(.A(n11917), .B(n7862), .Y(new_n3332));
  not_3  g02956(.A(new_n3332), .Y(new_n3333));
  nand_4 g02957(.A(new_n3333), .B(new_n3331), .Y(new_n3334));
  nand_4 g02958(.A(new_n3332), .B(new_n3330), .Y(new_n3335));
  nand_4 g02959(.A(n4921), .B(n1333), .Y(new_n3336));
  not_3  g02960(.A(new_n3336), .Y(new_n3337));
  nand_4 g02961(.A(new_n3337), .B(new_n3335), .Y(new_n3338));
  nand_4 g02962(.A(new_n3338), .B(new_n3334), .Y(new_n3339_1));
  not_3  g02963(.A(new_n3339_1), .Y(new_n3340));
  nor_4  g02964(.A(new_n3340), .B(new_n3329), .Y(new_n3341));
  not_3  g02965(.A(new_n3341), .Y(new_n3342_1));
  xor_3  g02966(.A(new_n3340), .B(new_n3329), .Y(new_n3343));
  nor_4  g02967(.A(new_n3313), .B(new_n3312), .Y(new_n3344));
  xor_3  g02968(.A(new_n3344), .B(new_n3293), .Y(new_n3345));
  nand_4 g02969(.A(new_n3345), .B(new_n3343), .Y(new_n3346));
  nand_4 g02970(.A(new_n3346), .B(new_n3342_1), .Y(new_n3347));
  xnor_3 g02971(.A(new_n3326), .B(new_n3325), .Y(new_n3348));
  not_3  g02972(.A(new_n3348), .Y(new_n3349));
  nand_4 g02973(.A(new_n3349), .B(new_n3347), .Y(new_n3350));
  nand_4 g02974(.A(new_n3350), .B(new_n3328), .Y(new_n3351));
  nand_4 g02975(.A(new_n3351), .B(new_n3324), .Y(new_n3352));
  not_3  g02976(.A(new_n3295), .Y(new_n3353));
  nand_4 g02977(.A(new_n3299), .B(new_n3296), .Y(new_n3354));
  nand_4 g02978(.A(new_n3354), .B(new_n3353), .Y(new_n3355));
  nand_4 g02979(.A(n9637), .B(n1333), .Y(new_n3356));
  not_3  g02980(.A(new_n3356), .Y(new_n3357));
  nand_4 g02981(.A(n3172), .B(n2577), .Y(new_n3358));
  nand_4 g02982(.A(n7862), .B(n1835), .Y(new_n3359));
  xor_3  g02983(.A(new_n3359), .B(new_n3358), .Y(new_n3360));
  xnor_3 g02984(.A(new_n3360), .B(new_n3357), .Y(new_n3361));
  xnor_3 g02985(.A(new_n3361), .B(new_n3355), .Y(new_n3362));
  nor_4  g02986(.A(new_n3298), .B(new_n3297), .Y(new_n3363));
  not_3  g02987(.A(new_n3363), .Y(new_n3364));
  nand_4 g02988(.A(n11757), .B(n3842), .Y(new_n3365));
  xor_3  g02989(.A(new_n3365), .B(new_n3364), .Y(new_n3366));
  nand_4 g02990(.A(n11821), .B(n4921), .Y(new_n3367));
  nand_4 g02991(.A(n9956), .B(n9080), .Y(new_n3368));
  nand_4 g02992(.A(n11917), .B(n5240), .Y(new_n3369));
  not_3  g02993(.A(new_n3369), .Y(new_n3370));
  xor_3  g02994(.A(new_n3370), .B(new_n3368), .Y(new_n3371));
  xnor_3 g02995(.A(new_n3371), .B(new_n3367), .Y(new_n3372));
  not_3  g02996(.A(new_n3372), .Y(new_n3373));
  nor_4  g02997(.A(new_n3373), .B(new_n3366), .Y(new_n3374));
  not_3  g02998(.A(new_n3366), .Y(new_n3375));
  nor_4  g02999(.A(new_n3372), .B(new_n3375), .Y(new_n3376));
  nor_4  g03000(.A(new_n3376), .B(new_n3374), .Y(new_n3377));
  xnor_3 g03001(.A(new_n3377), .B(new_n3362), .Y(new_n3378));
  nand_4 g03002(.A(new_n3304), .B(new_n3301), .Y(new_n3379));
  nor_4  g03003(.A(new_n3303), .B(new_n3302), .Y(new_n3380));
  nor_4  g03004(.A(new_n3322), .B(new_n3305), .Y(new_n3381));
  xnor_3 g03005(.A(new_n3381), .B(new_n3380), .Y(new_n3382));
  nand_4 g03006(.A(new_n3382), .B(new_n3379), .Y(new_n3383));
  xnor_3 g03007(.A(new_n3383), .B(new_n3378), .Y(new_n3384));
  xnor_3 g03008(.A(new_n3384), .B(new_n3352), .Y(new_n3385));
  nand_4 g03009(.A(n9637), .B(n7862), .Y(new_n3386));
  not_3  g03010(.A(new_n3386), .Y(new_n3387));
  xnor_3 g03011(.A(new_n3351), .B(new_n3324), .Y(new_n3388));
  not_3  g03012(.A(new_n3388), .Y(new_n3389));
  nand_4 g03013(.A(new_n3389), .B(new_n3387), .Y(new_n3390));
  and_4  g03014(.A(new_n3335), .B(new_n3334), .Y(new_n3391));
  nand_4 g03015(.A(n9956), .B(n1333), .Y(new_n3392));
  nand_4 g03016(.A(n7862), .B(n4921), .Y(new_n3393));
  nor_4  g03017(.A(new_n3393), .B(new_n3392), .Y(new_n3394));
  not_3  g03018(.A(new_n3394), .Y(new_n3395));
  nor_4  g03019(.A(new_n3395), .B(new_n3391), .Y(new_n3396));
  xor_3  g03020(.A(new_n3339_1), .B(new_n3329), .Y(new_n3397));
  xor_3  g03021(.A(new_n3344), .B(new_n3292), .Y(new_n3398));
  nor_4  g03022(.A(new_n3398), .B(new_n3397), .Y(new_n3399));
  nor_4  g03023(.A(new_n3345), .B(new_n3343), .Y(new_n3400));
  nor_4  g03024(.A(new_n3400), .B(new_n3399), .Y(new_n3401));
  nand_4 g03025(.A(new_n3401), .B(new_n3396), .Y(new_n3402));
  xnor_3 g03026(.A(new_n3349), .B(new_n3347), .Y(new_n3403));
  nor_4  g03027(.A(new_n3403), .B(new_n3402), .Y(new_n3404));
  xnor_3 g03028(.A(new_n3388), .B(new_n3387), .Y(new_n3405));
  nand_4 g03029(.A(new_n3405), .B(new_n3404), .Y(new_n3406));
  nand_4 g03030(.A(new_n3406), .B(new_n3390), .Y(new_n3407));
  xor_3  g03031(.A(new_n3407), .B(new_n3385), .Y(new_n3408));
  not_3  g03032(.A(new_n3405), .Y(new_n3409));
  xor_3  g03033(.A(new_n3409), .B(new_n3404), .Y(new_n3410));
  not_3  g03034(.A(new_n3410), .Y(new_n3411));
  nand_4 g03035(.A(n8595), .B(n6877), .Y(new_n3412));
  nand_4 g03036(.A(n6877), .B(n6126), .Y(new_n3413));
  not_3  g03037(.A(new_n3413), .Y(new_n3414));
  nand_4 g03038(.A(n3719), .B(n2464), .Y(new_n3415));
  not_3  g03039(.A(new_n3415), .Y(new_n3416));
  nor_4  g03040(.A(new_n3416), .B(new_n3414), .Y(new_n3417));
  nor_4  g03041(.A(new_n3415), .B(new_n3413), .Y(new_n3418));
  nand_4 g03042(.A(n9400), .B(n3602), .Y(new_n3419));
  not_3  g03043(.A(new_n3419), .Y(new_n3420));
  nor_4  g03044(.A(new_n3420), .B(new_n3418), .Y(new_n3421));
  nor_4  g03045(.A(new_n3421), .B(new_n3417), .Y(new_n3422));
  xor_3  g03046(.A(new_n3422), .B(new_n3412), .Y(new_n3423));
  nand_4 g03047(.A(n3602), .B(n2464), .Y(new_n3424));
  nand_4 g03048(.A(n9400), .B(n6126), .Y(new_n3425));
  not_3  g03049(.A(new_n3425), .Y(new_n3426));
  nand_4 g03050(.A(n11311), .B(n3719), .Y(new_n3427));
  not_3  g03051(.A(new_n3427), .Y(new_n3428));
  nor_4  g03052(.A(new_n3428), .B(new_n3426), .Y(new_n3429));
  nor_4  g03053(.A(new_n3427), .B(new_n3425), .Y(new_n3430));
  nor_4  g03054(.A(new_n3430), .B(new_n3429), .Y(new_n3431));
  xor_3  g03055(.A(new_n3431), .B(new_n3424), .Y(new_n3432));
  xnor_3 g03056(.A(new_n3432), .B(new_n3423), .Y(new_n3433));
  nand_4 g03057(.A(n6877), .B(n3719), .Y(new_n3434));
  not_3  g03058(.A(new_n3434), .Y(new_n3435));
  nor_4  g03059(.A(new_n3435), .B(new_n3419), .Y(new_n3436));
  nor_4  g03060(.A(new_n3418), .B(new_n3417), .Y(new_n3437));
  nor_4  g03061(.A(new_n3437), .B(new_n3436), .Y(new_n3438));
  not_3  g03062(.A(new_n3438), .Y(new_n3439));
  nor_4  g03063(.A(new_n3439), .B(new_n3419), .Y(new_n3440));
  not_3  g03064(.A(new_n3440), .Y(new_n3441));
  nor_4  g03065(.A(new_n3441), .B(new_n3433), .Y(new_n3442));
  not_3  g03066(.A(new_n3442), .Y(new_n3443));
  nand_4 g03067(.A(n10439), .B(n6877), .Y(new_n3444));
  nand_4 g03068(.A(n9400), .B(n8595), .Y(new_n3445));
  not_3  g03069(.A(new_n3445), .Y(new_n3446));
  not_3  g03070(.A(new_n3424), .Y(new_n3447));
  nor_4  g03071(.A(new_n3430), .B(new_n3447), .Y(new_n3448));
  nor_4  g03072(.A(new_n3448), .B(new_n3429), .Y(new_n3449));
  xnor_3 g03073(.A(new_n3449), .B(new_n3446), .Y(new_n3450));
  nand_4 g03074(.A(n11311), .B(n3602), .Y(new_n3451));
  not_3  g03075(.A(new_n3451), .Y(new_n3452));
  nand_4 g03076(.A(n6126), .B(n2464), .Y(new_n3453));
  nand_4 g03077(.A(n4187), .B(n3719), .Y(new_n3454));
  xnor_3 g03078(.A(new_n3454), .B(new_n3453), .Y(new_n3455));
  xor_3  g03079(.A(new_n3455), .B(new_n3452), .Y(new_n3456_1));
  xnor_3 g03080(.A(new_n3456_1), .B(new_n3450), .Y(new_n3457));
  xnor_3 g03081(.A(new_n3457), .B(new_n3444), .Y(new_n3458));
  not_3  g03082(.A(new_n3412), .Y(new_n3459));
  and_4  g03083(.A(new_n3422), .B(new_n3459), .Y(new_n3460));
  nor_4  g03084(.A(new_n3432), .B(new_n3423), .Y(new_n3461));
  nor_4  g03085(.A(new_n3461), .B(new_n3460), .Y(new_n3462));
  xnor_3 g03086(.A(new_n3462), .B(new_n3458), .Y(new_n3463));
  nor_4  g03087(.A(new_n3463), .B(new_n3443), .Y(new_n3464));
  not_3  g03088(.A(new_n3464), .Y(new_n3465));
  nand_4 g03089(.A(n8065), .B(n6877), .Y(new_n3466));
  nand_4 g03090(.A(n11311), .B(n6126), .Y(new_n3467));
  nand_4 g03091(.A(n4203), .B(n3719), .Y(new_n3468));
  nand_4 g03092(.A(n4187), .B(n3602), .Y(new_n3469));
  xnor_3 g03093(.A(new_n3469), .B(new_n3468), .Y(new_n3470));
  nor_4  g03094(.A(new_n3470), .B(new_n3467), .Y(new_n3471));
  not_3  g03095(.A(new_n3467), .Y(new_n3472));
  not_3  g03096(.A(new_n3470), .Y(new_n3473));
  nor_4  g03097(.A(new_n3473), .B(new_n3472), .Y(new_n3474));
  nor_4  g03098(.A(new_n3474), .B(new_n3471), .Y(new_n3475));
  and_4  g03099(.A(new_n3454), .B(new_n3453), .Y(new_n3476));
  nor_4  g03100(.A(new_n3455), .B(new_n3452), .Y(new_n3477));
  nor_4  g03101(.A(new_n3477), .B(new_n3476), .Y(new_n3478));
  not_3  g03102(.A(new_n3478), .Y(new_n3479));
  xor_3  g03103(.A(new_n3479), .B(new_n3475), .Y(new_n3480));
  nand_4 g03104(.A(n10439), .B(n9400), .Y(new_n3481));
  nand_4 g03105(.A(n8595), .B(n2464), .Y(new_n3482));
  xor_3  g03106(.A(new_n3482), .B(new_n3481), .Y(new_n3483));
  not_3  g03107(.A(new_n3483), .Y(new_n3484));
  xnor_3 g03108(.A(new_n3484), .B(new_n3480), .Y(new_n3485));
  and_4  g03109(.A(new_n3449), .B(new_n3446), .Y(new_n3486));
  not_3  g03110(.A(new_n3486), .Y(new_n3487));
  not_3  g03111(.A(new_n3450), .Y(new_n3488));
  not_3  g03112(.A(new_n3456_1), .Y(new_n3489));
  nand_4 g03113(.A(new_n3489), .B(new_n3488), .Y(new_n3490));
  and_4  g03114(.A(new_n3490), .B(new_n3487), .Y(new_n3491));
  xnor_3 g03115(.A(new_n3491), .B(new_n3485), .Y(new_n3492));
  not_3  g03116(.A(new_n3444), .Y(new_n3493));
  not_3  g03117(.A(new_n3457), .Y(new_n3494));
  nand_4 g03118(.A(new_n3494), .B(new_n3493), .Y(new_n3495));
  xor_3  g03119(.A(new_n3494), .B(new_n3493), .Y(new_n3496));
  not_3  g03120(.A(new_n3462), .Y(new_n3497));
  nand_4 g03121(.A(new_n3497), .B(new_n3496), .Y(new_n3498));
  nand_4 g03122(.A(new_n3498), .B(new_n3495), .Y(new_n3499));
  not_3  g03123(.A(new_n3499), .Y(new_n3500));
  xnor_3 g03124(.A(new_n3500), .B(new_n3492), .Y(new_n3501));
  xnor_3 g03125(.A(new_n3501), .B(new_n3466), .Y(new_n3502));
  xnor_3 g03126(.A(new_n3502), .B(new_n3465), .Y(new_n3503));
  not_3  g03127(.A(new_n3463), .Y(new_n3504));
  xor_3  g03128(.A(new_n3504), .B(new_n3443), .Y(new_n3505));
  not_3  g03129(.A(new_n3505), .Y(new_n3506));
  not_3  g03130(.A(new_n3433), .Y(new_n3507));
  xor_3  g03131(.A(new_n3440), .B(new_n3507), .Y(new_n3508));
  not_3  g03132(.A(new_n3508), .Y(new_n3509));
  nand_4 g03133(.A(n8433), .B(n7236), .Y(new_n3510));
  nand_4 g03134(.A(n12925), .B(n4805), .Y(new_n3511));
  nor_4  g03135(.A(new_n3511), .B(new_n3510), .Y(new_n3512));
  nand_4 g03136(.A(n7733), .B(n4805), .Y(new_n3513));
  nand_4 g03137(.A(n12925), .B(n11478), .Y(new_n3514));
  xnor_3 g03138(.A(new_n3514), .B(new_n3513), .Y(new_n3515));
  not_3  g03139(.A(new_n3515), .Y(new_n3516));
  nor_4  g03140(.A(new_n3516), .B(new_n3512), .Y(new_n3517));
  not_3  g03141(.A(new_n3517), .Y(new_n3518));
  not_3  g03142(.A(new_n3512), .Y(new_n3519));
  nor_4  g03143(.A(new_n3515), .B(new_n3519), .Y(new_n3520));
  nor_4  g03144(.A(new_n3520), .B(new_n3517), .Y(new_n3521));
  nand_4 g03145(.A(n7236), .B(n405), .Y(new_n3522));
  nand_4 g03146(.A(n8433), .B(n3992), .Y(new_n3523));
  xnor_3 g03147(.A(new_n3523), .B(new_n3522), .Y(new_n3524));
  nand_4 g03148(.A(new_n3524), .B(new_n3521), .Y(new_n3525));
  nand_4 g03149(.A(new_n3525), .B(new_n3518), .Y(new_n3526));
  not_3  g03150(.A(new_n3510), .Y(new_n3527));
  nand_4 g03151(.A(n3992), .B(n405), .Y(new_n3528));
  nor_4  g03152(.A(new_n3528), .B(new_n3527), .Y(new_n3529));
  nand_4 g03153(.A(n8433), .B(n8384), .Y(new_n3530));
  not_3  g03154(.A(new_n3530), .Y(new_n3531));
  nand_4 g03155(.A(n7236), .B(n4086), .Y(new_n3532));
  not_3  g03156(.A(new_n3532), .Y(new_n3533));
  nor_4  g03157(.A(new_n3533), .B(new_n3531), .Y(new_n3534));
  not_3  g03158(.A(new_n3534), .Y(new_n3535));
  nor_4  g03159(.A(new_n3535), .B(new_n3529), .Y(new_n3536));
  nor_4  g03160(.A(new_n3532), .B(new_n3530), .Y(new_n3537));
  nor_4  g03161(.A(new_n3537), .B(new_n3536), .Y(new_n3538));
  not_3  g03162(.A(new_n3529), .Y(new_n3539));
  nor_4  g03163(.A(new_n3534), .B(new_n3539), .Y(new_n3540));
  not_3  g03164(.A(new_n3540), .Y(new_n3541));
  nand_4 g03165(.A(new_n3541), .B(new_n3538), .Y(new_n3542));
  xnor_3 g03166(.A(new_n3542), .B(new_n3526), .Y(new_n3543));
  not_3  g03167(.A(new_n3511), .Y(new_n3544));
  nand_4 g03168(.A(n11478), .B(n7733), .Y(new_n3545));
  nor_4  g03169(.A(new_n3545), .B(new_n3544), .Y(new_n3546));
  not_3  g03170(.A(new_n3546), .Y(new_n3547));
  nand_4 g03171(.A(n12925), .B(n5283), .Y(new_n3548));
  nand_4 g03172(.A(n4826), .B(n4805), .Y(new_n3549));
  nand_4 g03173(.A(new_n3549), .B(new_n3548), .Y(new_n3550));
  nor_4  g03174(.A(new_n3550), .B(new_n3547), .Y(new_n3551));
  not_3  g03175(.A(new_n3550), .Y(new_n3552));
  not_3  g03176(.A(new_n3548), .Y(new_n3553));
  not_3  g03177(.A(new_n3549), .Y(new_n3554));
  nand_4 g03178(.A(new_n3554), .B(new_n3553), .Y(new_n3555));
  not_3  g03179(.A(new_n3555), .Y(new_n3556));
  nor_4  g03180(.A(new_n3556), .B(new_n3552), .Y(new_n3557));
  not_3  g03181(.A(new_n3557), .Y(new_n3558));
  nor_4  g03182(.A(new_n3558), .B(new_n3546), .Y(new_n3559));
  nor_4  g03183(.A(new_n3559), .B(new_n3551), .Y(new_n3560));
  not_3  g03184(.A(new_n3560), .Y(new_n3561));
  xnor_3 g03185(.A(new_n3561), .B(new_n3543), .Y(new_n3562));
  not_3  g03186(.A(new_n3562), .Y(new_n3563));
  not_3  g03187(.A(new_n3417), .Y(new_n3564));
  nand_4 g03188(.A(new_n3436), .B(new_n3564), .Y(new_n3565));
  nand_4 g03189(.A(new_n3565), .B(new_n3439), .Y(new_n3566));
  nor_4  g03190(.A(new_n3566), .B(new_n3563), .Y(new_n3567));
  not_3  g03191(.A(new_n3566), .Y(new_n3568));
  nor_4  g03192(.A(new_n3568), .B(new_n3562), .Y(new_n3569));
  nor_4  g03193(.A(new_n3569), .B(new_n3567), .Y(new_n3570));
  not_3  g03194(.A(new_n3570), .Y(new_n3571));
  xnor_3 g03195(.A(new_n3524), .B(new_n3521), .Y(new_n3572));
  not_3  g03196(.A(new_n3572), .Y(new_n3573));
  nand_4 g03197(.A(n9400), .B(n3719), .Y(new_n3574));
  nand_4 g03198(.A(n6877), .B(n3602), .Y(new_n3575));
  not_3  g03199(.A(new_n3575), .Y(new_n3576));
  xor_3  g03200(.A(new_n3576), .B(new_n3574), .Y(new_n3577));
  nor_4  g03201(.A(new_n3577), .B(new_n3573), .Y(new_n3578));
  xor_3  g03202(.A(new_n3511), .B(new_n3510), .Y(new_n3579));
  nand_4 g03203(.A(new_n3579), .B(new_n3435), .Y(new_n3580));
  xnor_3 g03204(.A(new_n3577), .B(new_n3572), .Y(new_n3581));
  not_3  g03205(.A(new_n3581), .Y(new_n3582));
  nor_4  g03206(.A(new_n3582), .B(new_n3580), .Y(new_n3583));
  nor_4  g03207(.A(new_n3583), .B(new_n3578), .Y(new_n3584));
  nor_4  g03208(.A(new_n3584), .B(new_n3571), .Y(new_n3585));
  nor_4  g03209(.A(new_n3585), .B(new_n3567), .Y(new_n3586));
  nor_4  g03210(.A(new_n3586), .B(new_n3509), .Y(new_n3587));
  not_3  g03211(.A(new_n3587), .Y(new_n3588));
  nand_4 g03212(.A(new_n3586), .B(new_n3509), .Y(new_n3589));
  nand_4 g03213(.A(n7610), .B(n4805), .Y(new_n3590));
  not_3  g03214(.A(new_n3545), .Y(new_n3591));
  nand_4 g03215(.A(new_n3550), .B(new_n3591), .Y(new_n3592));
  nand_4 g03216(.A(new_n3592), .B(new_n3555), .Y(new_n3593));
  not_3  g03217(.A(new_n3593), .Y(new_n3594));
  xnor_3 g03218(.A(new_n3594), .B(new_n3590), .Y(new_n3595));
  nand_4 g03219(.A(n7733), .B(n5283), .Y(new_n3596));
  nand_4 g03220(.A(n12925), .B(n137), .Y(new_n3597));
  nand_4 g03221(.A(n11478), .B(n4826), .Y(new_n3598));
  xnor_3 g03222(.A(new_n3598), .B(new_n3597), .Y(new_n3599));
  xnor_3 g03223(.A(new_n3599), .B(new_n3596), .Y(new_n3600));
  xnor_3 g03224(.A(new_n3600), .B(new_n3595), .Y(new_n3601));
  not_3  g03225(.A(new_n3601), .Y(new_n3602_1));
  nor_4  g03226(.A(new_n3514), .B(new_n3513), .Y(new_n3603));
  not_3  g03227(.A(new_n3603), .Y(new_n3604));
  nor_4  g03228(.A(new_n3557), .B(new_n3604), .Y(new_n3605));
  nor_4  g03229(.A(new_n3605), .B(new_n3602_1), .Y(new_n3606));
  not_3  g03230(.A(new_n3605), .Y(new_n3607));
  nor_4  g03231(.A(new_n3607), .B(new_n3601), .Y(new_n3608));
  nor_4  g03232(.A(new_n3608), .B(new_n3606), .Y(new_n3609));
  nand_4 g03233(.A(n7236), .B(n217), .Y(new_n3610));
  not_3  g03234(.A(new_n3610), .Y(new_n3611));
  not_3  g03235(.A(new_n3528), .Y(new_n3612));
  nor_4  g03236(.A(new_n3537), .B(new_n3612), .Y(new_n3613));
  nor_4  g03237(.A(new_n3613), .B(new_n3534), .Y(new_n3614));
  xnor_3 g03238(.A(new_n3614), .B(new_n3611), .Y(new_n3615));
  nand_4 g03239(.A(n8384), .B(n405), .Y(new_n3616_1));
  nand_4 g03240(.A(n8433), .B(n6358), .Y(new_n3617));
  nand_4 g03241(.A(n4086), .B(n3992), .Y(new_n3618));
  xnor_3 g03242(.A(new_n3618), .B(new_n3617), .Y(new_n3619));
  xnor_3 g03243(.A(new_n3619), .B(new_n3616_1), .Y(new_n3620));
  xnor_3 g03244(.A(new_n3620), .B(new_n3615), .Y(new_n3621));
  not_3  g03245(.A(new_n3621), .Y(new_n3622));
  nor_4  g03246(.A(new_n3538), .B(new_n3528), .Y(new_n3623));
  nor_4  g03247(.A(new_n3623), .B(new_n3622), .Y(new_n3624));
  not_3  g03248(.A(new_n3623), .Y(new_n3625));
  nor_4  g03249(.A(new_n3625), .B(new_n3621), .Y(new_n3626));
  nor_4  g03250(.A(new_n3626), .B(new_n3624), .Y(new_n3627_1));
  xnor_3 g03251(.A(new_n3627_1), .B(new_n3609), .Y(new_n3628));
  not_3  g03252(.A(new_n3628), .Y(new_n3629));
  and_4  g03253(.A(new_n3542), .B(new_n3526), .Y(new_n3630));
  nor_4  g03254(.A(new_n3561), .B(new_n3543), .Y(new_n3631));
  nor_4  g03255(.A(new_n3631), .B(new_n3630), .Y(new_n3632));
  not_3  g03256(.A(new_n3632), .Y(new_n3633));
  nor_4  g03257(.A(new_n3633), .B(new_n3629), .Y(new_n3634));
  nor_4  g03258(.A(new_n3632), .B(new_n3628), .Y(new_n3635));
  nor_4  g03259(.A(new_n3635), .B(new_n3634), .Y(new_n3636));
  not_3  g03260(.A(new_n3636), .Y(new_n3637));
  nand_4 g03261(.A(new_n3637), .B(new_n3589), .Y(new_n3638));
  nand_4 g03262(.A(new_n3638), .B(new_n3588), .Y(new_n3639));
  nand_4 g03263(.A(new_n3639), .B(new_n3506), .Y(new_n3640));
  not_3  g03264(.A(new_n3586), .Y(new_n3641));
  nor_4  g03265(.A(new_n3641), .B(new_n3508), .Y(new_n3642));
  nor_4  g03266(.A(new_n3636), .B(new_n3642), .Y(new_n3643));
  nor_4  g03267(.A(new_n3643), .B(new_n3587), .Y(new_n3644));
  nand_4 g03268(.A(new_n3644), .B(new_n3505), .Y(new_n3645));
  nand_4 g03269(.A(n7236), .B(n6611), .Y(new_n3646));
  nand_4 g03270(.A(n3992), .B(n217), .Y(new_n3647));
  not_3  g03271(.A(new_n3647), .Y(new_n3648));
  not_3  g03272(.A(new_n3617), .Y(new_n3649));
  not_3  g03273(.A(new_n3618), .Y(new_n3650));
  nor_4  g03274(.A(new_n3650), .B(new_n3649), .Y(new_n3651));
  not_3  g03275(.A(new_n3616_1), .Y(new_n3652));
  nor_4  g03276(.A(new_n3619), .B(new_n3652), .Y(new_n3653));
  nor_4  g03277(.A(new_n3653), .B(new_n3651), .Y(new_n3654_1));
  xnor_3 g03278(.A(new_n3654_1), .B(new_n3648), .Y(new_n3655));
  nand_4 g03279(.A(n6358), .B(n405), .Y(new_n3656));
  nand_4 g03280(.A(n8384), .B(n4086), .Y(new_n3657));
  nand_4 g03281(.A(n8433), .B(n5198), .Y(new_n3658));
  xnor_3 g03282(.A(new_n3658), .B(new_n3657), .Y(new_n3659));
  xnor_3 g03283(.A(new_n3659), .B(new_n3656), .Y(new_n3660));
  xnor_3 g03284(.A(new_n3660), .B(new_n3655), .Y(new_n3661_1));
  nor_4  g03285(.A(new_n3661_1), .B(new_n3646), .Y(new_n3662));
  not_3  g03286(.A(new_n3646), .Y(new_n3663));
  not_3  g03287(.A(new_n3661_1), .Y(new_n3664));
  nor_4  g03288(.A(new_n3664), .B(new_n3663), .Y(new_n3665));
  nor_4  g03289(.A(new_n3665), .B(new_n3662), .Y(new_n3666));
  nand_4 g03290(.A(new_n3614), .B(new_n3611), .Y(new_n3667));
  not_3  g03291(.A(new_n3667), .Y(new_n3668));
  nor_4  g03292(.A(new_n3620), .B(new_n3615), .Y(new_n3669));
  nor_4  g03293(.A(new_n3669), .B(new_n3668), .Y(new_n3670));
  not_3  g03294(.A(new_n3670), .Y(new_n3671));
  nand_4 g03295(.A(new_n3671), .B(new_n3666), .Y(new_n3672));
  not_3  g03296(.A(new_n3672), .Y(new_n3673));
  nor_4  g03297(.A(new_n3671), .B(new_n3666), .Y(new_n3674));
  nor_4  g03298(.A(new_n3674), .B(new_n3673), .Y(new_n3675));
  nor_4  g03299(.A(new_n3675), .B(new_n3626), .Y(new_n3676));
  nand_4 g03300(.A(new_n3675), .B(new_n3626), .Y(new_n3677_1));
  not_3  g03301(.A(new_n3677_1), .Y(new_n3678));
  nor_4  g03302(.A(new_n3678), .B(new_n3676), .Y(new_n3679));
  nand_4 g03303(.A(n4970), .B(n4805), .Y(new_n3680));
  nand_4 g03304(.A(n11478), .B(n7610), .Y(new_n3681));
  not_3  g03305(.A(new_n3681), .Y(new_n3682));
  not_3  g03306(.A(new_n3597), .Y(new_n3683));
  not_3  g03307(.A(new_n3598), .Y(new_n3684));
  nor_4  g03308(.A(new_n3684), .B(new_n3683), .Y(new_n3685));
  not_3  g03309(.A(new_n3596), .Y(new_n3686));
  nor_4  g03310(.A(new_n3599), .B(new_n3686), .Y(new_n3687));
  nor_4  g03311(.A(new_n3687), .B(new_n3685), .Y(new_n3688));
  xnor_3 g03312(.A(new_n3688), .B(new_n3682), .Y(new_n3689));
  nand_4 g03313(.A(n7733), .B(n137), .Y(new_n3690));
  nand_4 g03314(.A(n5283), .B(n4826), .Y(new_n3691));
  nand_4 g03315(.A(n12925), .B(n6294), .Y(new_n3692));
  xnor_3 g03316(.A(new_n3692), .B(new_n3691), .Y(new_n3693));
  xnor_3 g03317(.A(new_n3693), .B(new_n3690), .Y(new_n3694));
  xnor_3 g03318(.A(new_n3694), .B(new_n3689), .Y(new_n3695));
  nor_4  g03319(.A(new_n3695), .B(new_n3680), .Y(new_n3696));
  not_3  g03320(.A(new_n3680), .Y(new_n3697));
  not_3  g03321(.A(new_n3695), .Y(new_n3698));
  nor_4  g03322(.A(new_n3698), .B(new_n3697), .Y(new_n3699));
  nor_4  g03323(.A(new_n3699), .B(new_n3696), .Y(new_n3700));
  nor_4  g03324(.A(new_n3594), .B(new_n3590), .Y(new_n3701));
  nor_4  g03325(.A(new_n3600), .B(new_n3595), .Y(new_n3702));
  nor_4  g03326(.A(new_n3702), .B(new_n3701), .Y(new_n3703));
  not_3  g03327(.A(new_n3703), .Y(new_n3704));
  xnor_3 g03328(.A(new_n3704), .B(new_n3700), .Y(new_n3705));
  not_3  g03329(.A(new_n3705), .Y(new_n3706));
  nor_4  g03330(.A(new_n3706), .B(new_n3608), .Y(new_n3707));
  not_3  g03331(.A(new_n3608), .Y(new_n3708));
  nor_4  g03332(.A(new_n3705), .B(new_n3708), .Y(new_n3709));
  nor_4  g03333(.A(new_n3709), .B(new_n3707), .Y(new_n3710));
  nor_4  g03334(.A(new_n3627_1), .B(new_n3609), .Y(new_n3711));
  nor_4  g03335(.A(new_n3635), .B(new_n3711), .Y(new_n3712));
  xnor_3 g03336(.A(new_n3712), .B(new_n3710), .Y(new_n3713));
  xnor_3 g03337(.A(new_n3713), .B(new_n3679), .Y(new_n3714));
  nand_4 g03338(.A(new_n3714), .B(new_n3645), .Y(new_n3715));
  nand_4 g03339(.A(new_n3715), .B(new_n3640), .Y(new_n3716));
  xnor_3 g03340(.A(new_n3716), .B(new_n3503), .Y(new_n3717));
  nand_4 g03341(.A(n7236), .B(n6359), .Y(new_n3718));
  not_3  g03342(.A(new_n3718), .Y(new_n3719_1));
  nand_4 g03343(.A(n6358), .B(n4086), .Y(new_n3720));
  not_3  g03344(.A(new_n3720), .Y(new_n3721));
  not_3  g03345(.A(new_n3657), .Y(new_n3722));
  not_3  g03346(.A(new_n3658), .Y(new_n3723));
  nor_4  g03347(.A(new_n3723), .B(new_n3722), .Y(new_n3724));
  not_3  g03348(.A(new_n3656), .Y(new_n3725));
  nor_4  g03349(.A(new_n3659), .B(new_n3725), .Y(new_n3726));
  nor_4  g03350(.A(new_n3726), .B(new_n3724), .Y(new_n3727));
  xnor_3 g03351(.A(new_n3727), .B(new_n3721), .Y(new_n3728));
  nand_4 g03352(.A(n5198), .B(n405), .Y(new_n3729));
  nand_4 g03353(.A(n8433), .B(n1471), .Y(new_n3730));
  xnor_3 g03354(.A(new_n3730), .B(new_n3729), .Y(new_n3731));
  xnor_3 g03355(.A(new_n3731), .B(new_n3728), .Y(new_n3732));
  not_3  g03356(.A(new_n3732), .Y(new_n3733));
  nand_4 g03357(.A(n8384), .B(n217), .Y(new_n3734));
  nand_4 g03358(.A(n6611), .B(n3992), .Y(new_n3735));
  xor_3  g03359(.A(new_n3735), .B(new_n3734), .Y(new_n3736));
  xnor_3 g03360(.A(new_n3736), .B(new_n3733), .Y(new_n3737));
  not_3  g03361(.A(new_n3737), .Y(new_n3738));
  and_4  g03362(.A(new_n3654_1), .B(new_n3648), .Y(new_n3739));
  nor_4  g03363(.A(new_n3660), .B(new_n3655), .Y(new_n3740));
  nor_4  g03364(.A(new_n3740), .B(new_n3739), .Y(new_n3741));
  xnor_3 g03365(.A(new_n3741), .B(new_n3738), .Y(new_n3742));
  not_3  g03366(.A(new_n3662), .Y(new_n3743));
  nand_4 g03367(.A(new_n3672), .B(new_n3743), .Y(new_n3744));
  xnor_3 g03368(.A(new_n3744), .B(new_n3742), .Y(new_n3745));
  xnor_3 g03369(.A(new_n3745), .B(new_n3719_1), .Y(new_n3746));
  nor_4  g03370(.A(new_n3746), .B(new_n3677_1), .Y(new_n3747));
  nand_4 g03371(.A(new_n3746), .B(new_n3677_1), .Y(new_n3748));
  not_3  g03372(.A(new_n3748), .Y(new_n3749));
  nor_4  g03373(.A(new_n3749), .B(new_n3747), .Y(new_n3750));
  nand_4 g03374(.A(n4805), .B(n503), .Y(new_n3751));
  not_3  g03375(.A(new_n3751), .Y(new_n3752));
  nand_4 g03376(.A(n4826), .B(n137), .Y(new_n3753));
  nand_4 g03377(.A(n7733), .B(n6294), .Y(new_n3754_1));
  nand_4 g03378(.A(n12925), .B(n6797), .Y(new_n3755));
  xnor_3 g03379(.A(new_n3755), .B(new_n3754_1), .Y(new_n3756));
  nor_4  g03380(.A(new_n3756), .B(new_n3753), .Y(new_n3757));
  not_3  g03381(.A(new_n3753), .Y(new_n3758));
  not_3  g03382(.A(new_n3756), .Y(new_n3759));
  nor_4  g03383(.A(new_n3759), .B(new_n3758), .Y(new_n3760));
  nor_4  g03384(.A(new_n3760), .B(new_n3757), .Y(new_n3761));
  and_4  g03385(.A(new_n3692), .B(new_n3691), .Y(new_n3762));
  not_3  g03386(.A(new_n3690), .Y(new_n3763));
  nor_4  g03387(.A(new_n3693), .B(new_n3763), .Y(new_n3764));
  nor_4  g03388(.A(new_n3764), .B(new_n3762), .Y(new_n3765));
  xnor_3 g03389(.A(new_n3765), .B(new_n3761), .Y(new_n3766));
  nand_4 g03390(.A(n11478), .B(n4970), .Y(new_n3767));
  nand_4 g03391(.A(n7610), .B(n5283), .Y(new_n3768));
  xor_3  g03392(.A(new_n3768), .B(new_n3767), .Y(new_n3769));
  xnor_3 g03393(.A(new_n3769), .B(new_n3766), .Y(new_n3770));
  nand_4 g03394(.A(new_n3688), .B(new_n3682), .Y(new_n3771));
  not_3  g03395(.A(new_n3771), .Y(new_n3772));
  nor_4  g03396(.A(new_n3694), .B(new_n3689), .Y(new_n3773));
  nor_4  g03397(.A(new_n3773), .B(new_n3772), .Y(new_n3774));
  not_3  g03398(.A(new_n3774), .Y(new_n3775));
  xnor_3 g03399(.A(new_n3775), .B(new_n3770), .Y(new_n3776));
  not_3  g03400(.A(new_n3696), .Y(new_n3777));
  nand_4 g03401(.A(new_n3704), .B(new_n3700), .Y(new_n3778));
  nand_4 g03402(.A(new_n3778), .B(new_n3777), .Y(new_n3779));
  xnor_3 g03403(.A(new_n3779), .B(new_n3776), .Y(new_n3780));
  xnor_3 g03404(.A(new_n3780), .B(new_n3752), .Y(new_n3781));
  xnor_3 g03405(.A(new_n3781), .B(new_n3709), .Y(new_n3782));
  xnor_3 g03406(.A(new_n3782), .B(new_n3750), .Y(new_n3783));
  nor_4  g03407(.A(new_n3712), .B(new_n3710), .Y(new_n3784));
  not_3  g03408(.A(new_n3784), .Y(new_n3785));
  not_3  g03409(.A(new_n3679), .Y(new_n3786));
  not_3  g03410(.A(new_n3713), .Y(new_n3787));
  nand_4 g03411(.A(new_n3787), .B(new_n3786), .Y(new_n3788));
  nand_4 g03412(.A(new_n3788), .B(new_n3785), .Y(new_n3789));
  xnor_3 g03413(.A(new_n3789), .B(new_n3783), .Y(new_n3790));
  xnor_3 g03414(.A(new_n3790), .B(new_n3717), .Y(new_n3791));
  not_3  g03415(.A(new_n3791), .Y(new_n3792));
  nor_4  g03416(.A(new_n3792), .B(new_n3411), .Y(new_n3793));
  nor_4  g03417(.A(new_n3791), .B(new_n3410), .Y(new_n3794));
  xor_3  g03418(.A(new_n3403), .B(new_n3402), .Y(new_n3795));
  nand_4 g03419(.A(new_n3645), .B(new_n3640), .Y(new_n3796));
  xnor_3 g03420(.A(new_n3796), .B(new_n3714), .Y(new_n3797));
  nand_4 g03421(.A(new_n3797), .B(new_n3795), .Y(new_n3798));
  not_3  g03422(.A(new_n3798), .Y(new_n3799));
  nor_4  g03423(.A(new_n3797), .B(new_n3795), .Y(new_n3800));
  nor_4  g03424(.A(new_n3800), .B(new_n3799), .Y(new_n3801));
  not_3  g03425(.A(new_n3401), .Y(new_n3802));
  xor_3  g03426(.A(new_n3802), .B(new_n3396), .Y(new_n3803));
  nand_4 g03427(.A(new_n3589), .B(new_n3588), .Y(new_n3804));
  xnor_3 g03428(.A(new_n3804), .B(new_n3636), .Y(new_n3805));
  nor_4  g03429(.A(new_n3805), .B(new_n3803), .Y(new_n3806));
  not_3  g03430(.A(new_n3806), .Y(new_n3807));
  not_3  g03431(.A(new_n3584), .Y(new_n3808));
  nor_4  g03432(.A(new_n3808), .B(new_n3570), .Y(new_n3809));
  nor_4  g03433(.A(new_n3809), .B(new_n3585), .Y(new_n3810));
  not_3  g03434(.A(new_n3391), .Y(new_n3811));
  nand_4 g03435(.A(n9956), .B(n7862), .Y(new_n3812));
  not_3  g03436(.A(new_n3812), .Y(new_n3813));
  nor_4  g03437(.A(new_n3813), .B(new_n3336), .Y(new_n3814));
  not_3  g03438(.A(new_n3814), .Y(new_n3815));
  nand_4 g03439(.A(new_n3815), .B(new_n3811), .Y(new_n3816));
  nand_4 g03440(.A(new_n3814), .B(new_n3335), .Y(new_n3817));
  nand_4 g03441(.A(new_n3817), .B(new_n3816), .Y(new_n3818));
  not_3  g03442(.A(new_n3818), .Y(new_n3819));
  nor_4  g03443(.A(new_n3819), .B(new_n3810), .Y(new_n3820));
  not_3  g03444(.A(new_n3810), .Y(new_n3821));
  nor_4  g03445(.A(new_n3818), .B(new_n3821), .Y(new_n3822));
  nor_4  g03446(.A(new_n3822), .B(new_n3820), .Y(new_n3823));
  not_3  g03447(.A(new_n3823), .Y(new_n3824));
  xor_3  g03448(.A(new_n3579), .B(new_n3434), .Y(new_n3825));
  nor_4  g03449(.A(new_n3825), .B(new_n3812), .Y(new_n3826));
  xor_3  g03450(.A(new_n3393), .B(new_n3392), .Y(new_n3827));
  nor_4  g03451(.A(new_n3827), .B(new_n3826), .Y(new_n3828));
  xor_3  g03452(.A(new_n3582), .B(new_n3580), .Y(new_n3829));
  xnor_3 g03453(.A(new_n3827), .B(new_n3826), .Y(new_n3830));
  nor_4  g03454(.A(new_n3830), .B(new_n3829), .Y(new_n3831));
  nor_4  g03455(.A(new_n3831), .B(new_n3828), .Y(new_n3832));
  nor_4  g03456(.A(new_n3832), .B(new_n3824), .Y(new_n3833));
  nor_4  g03457(.A(new_n3833), .B(new_n3820), .Y(new_n3834));
  not_3  g03458(.A(new_n3803), .Y(new_n3835));
  not_3  g03459(.A(new_n3805), .Y(new_n3836));
  nor_4  g03460(.A(new_n3836), .B(new_n3835), .Y(new_n3837));
  nor_4  g03461(.A(new_n3837), .B(new_n3806), .Y(new_n3838));
  nand_4 g03462(.A(new_n3838), .B(new_n3834), .Y(new_n3839));
  nand_4 g03463(.A(new_n3839), .B(new_n3807), .Y(new_n3840));
  nand_4 g03464(.A(new_n3840), .B(new_n3801), .Y(new_n3841));
  nand_4 g03465(.A(new_n3841), .B(new_n3798), .Y(new_n3842_1));
  nor_4  g03466(.A(new_n3842_1), .B(new_n3794), .Y(new_n3843));
  nor_4  g03467(.A(new_n3843), .B(new_n3793), .Y(new_n3844));
  nor_4  g03468(.A(new_n3844), .B(new_n3408), .Y(new_n3845));
  not_3  g03469(.A(new_n3408), .Y(new_n3846));
  not_3  g03470(.A(new_n3844), .Y(new_n3847));
  nor_4  g03471(.A(new_n3847), .B(new_n3846), .Y(new_n3848));
  nor_4  g03472(.A(new_n3848), .B(new_n3845), .Y(new_n3849_1));
  nor_4  g03473(.A(new_n3500), .B(new_n3492), .Y(new_n3850));
  not_3  g03474(.A(new_n3850), .Y(new_n3851));
  not_3  g03475(.A(new_n3471), .Y(new_n3852));
  nand_4 g03476(.A(new_n3478), .B(new_n3475), .Y(new_n3853));
  nand_4 g03477(.A(new_n3853), .B(new_n3852), .Y(new_n3854));
  nand_4 g03478(.A(n9400), .B(n8065), .Y(new_n3855));
  not_3  g03479(.A(new_n3855), .Y(new_n3856));
  nand_4 g03480(.A(n10439), .B(n2464), .Y(new_n3857));
  nand_4 g03481(.A(n10391), .B(n6877), .Y(new_n3858));
  xor_3  g03482(.A(new_n3858), .B(new_n3857), .Y(new_n3859));
  xnor_3 g03483(.A(new_n3859), .B(new_n3856), .Y(new_n3860));
  xnor_3 g03484(.A(new_n3860), .B(new_n3854), .Y(new_n3861));
  not_3  g03485(.A(new_n3861), .Y(new_n3862));
  nor_4  g03486(.A(new_n3469), .B(new_n3468), .Y(new_n3863));
  nand_4 g03487(.A(n11311), .B(n8595), .Y(new_n3864));
  not_3  g03488(.A(new_n3864), .Y(new_n3865_1));
  xor_3  g03489(.A(new_n3865_1), .B(new_n3863), .Y(new_n3866));
  nand_4 g03490(.A(n4203), .B(n3602), .Y(new_n3867));
  not_3  g03491(.A(new_n3867), .Y(new_n3868));
  nand_4 g03492(.A(n6126), .B(n4187), .Y(new_n3869));
  nand_4 g03493(.A(n12753), .B(n3719), .Y(new_n3870));
  xnor_3 g03494(.A(new_n3870), .B(new_n3869), .Y(new_n3871));
  xnor_3 g03495(.A(new_n3871), .B(new_n3868), .Y(new_n3872));
  xnor_3 g03496(.A(new_n3872), .B(new_n3866), .Y(new_n3873));
  not_3  g03497(.A(new_n3873), .Y(new_n3874));
  xor_3  g03498(.A(new_n3874), .B(new_n3862), .Y(new_n3875));
  nor_4  g03499(.A(new_n3484), .B(new_n3480), .Y(new_n3876));
  nor_4  g03500(.A(new_n3482), .B(new_n3481), .Y(new_n3877));
  not_3  g03501(.A(new_n3877), .Y(new_n3878));
  not_3  g03502(.A(new_n3485), .Y(new_n3879));
  not_3  g03503(.A(new_n3491), .Y(new_n3880));
  nand_4 g03504(.A(new_n3880), .B(new_n3879), .Y(new_n3881));
  nor_4  g03505(.A(new_n3881), .B(new_n3878), .Y(new_n3882));
  nor_4  g03506(.A(new_n3491), .B(new_n3485), .Y(new_n3883));
  nor_4  g03507(.A(new_n3883), .B(new_n3877), .Y(new_n3884));
  nor_4  g03508(.A(new_n3884), .B(new_n3882), .Y(new_n3885));
  nor_4  g03509(.A(new_n3885), .B(new_n3876), .Y(new_n3886));
  xnor_3 g03510(.A(new_n3886), .B(new_n3875), .Y(new_n3887));
  xnor_3 g03511(.A(new_n3887), .B(new_n3851), .Y(new_n3888));
  nand_4 g03512(.A(new_n3501), .B(new_n3466), .Y(new_n3889));
  not_3  g03513(.A(new_n3889), .Y(new_n3890));
  nor_4  g03514(.A(new_n3502), .B(new_n3464), .Y(new_n3891));
  nor_4  g03515(.A(new_n3891), .B(new_n3890), .Y(new_n3892));
  xnor_3 g03516(.A(new_n3892), .B(new_n3888), .Y(new_n3893));
  not_3  g03517(.A(new_n3779), .Y(new_n3894));
  nor_4  g03518(.A(new_n3894), .B(new_n3776), .Y(new_n3895));
  not_3  g03519(.A(new_n3895), .Y(new_n3896));
  nand_4 g03520(.A(n10965), .B(n4805), .Y(new_n3897));
  not_3  g03521(.A(new_n3897), .Y(new_n3898));
  nand_4 g03522(.A(n5283), .B(n4970), .Y(new_n3899));
  nand_4 g03523(.A(n11478), .B(n503), .Y(new_n3900));
  not_3  g03524(.A(new_n3900), .Y(new_n3901));
  xor_3  g03525(.A(new_n3901), .B(new_n3899), .Y(new_n3902));
  xnor_3 g03526(.A(new_n3902), .B(new_n3898), .Y(new_n3903));
  not_3  g03527(.A(new_n3757), .Y(new_n3904));
  nand_4 g03528(.A(new_n3765), .B(new_n3761), .Y(new_n3905));
  nand_4 g03529(.A(new_n3905), .B(new_n3904), .Y(new_n3906));
  xnor_3 g03530(.A(new_n3906), .B(new_n3903), .Y(new_n3907));
  nor_4  g03531(.A(new_n3755), .B(new_n3754_1), .Y(new_n3908));
  nand_4 g03532(.A(n7610), .B(n137), .Y(new_n3909));
  not_3  g03533(.A(new_n3909), .Y(new_n3910));
  xor_3  g03534(.A(new_n3910), .B(new_n3908), .Y(new_n3911));
  nand_4 g03535(.A(n7733), .B(n6797), .Y(new_n3912));
  nand_4 g03536(.A(n6294), .B(n4826), .Y(new_n3913));
  not_3  g03537(.A(new_n3913), .Y(new_n3914));
  nand_4 g03538(.A(n12925), .B(n3146), .Y(new_n3915));
  not_3  g03539(.A(new_n3915), .Y(new_n3916));
  nor_4  g03540(.A(new_n3916), .B(new_n3914), .Y(new_n3917));
  nor_4  g03541(.A(new_n3915), .B(new_n3913), .Y(new_n3918));
  nor_4  g03542(.A(new_n3918), .B(new_n3917), .Y(new_n3919));
  xor_3  g03543(.A(new_n3919), .B(new_n3912), .Y(new_n3920));
  xnor_3 g03544(.A(new_n3920), .B(new_n3911), .Y(new_n3921));
  xnor_3 g03545(.A(new_n3921), .B(new_n3907), .Y(new_n3922));
  not_3  g03546(.A(new_n3766), .Y(new_n3923));
  nand_4 g03547(.A(new_n3769), .B(new_n3923), .Y(new_n3924));
  nor_4  g03548(.A(new_n3768), .B(new_n3767), .Y(new_n3925));
  nand_4 g03549(.A(new_n3775), .B(new_n3770), .Y(new_n3926));
  not_3  g03550(.A(new_n3926), .Y(new_n3927));
  xnor_3 g03551(.A(new_n3927), .B(new_n3925), .Y(new_n3928));
  nand_4 g03552(.A(new_n3928), .B(new_n3924), .Y(new_n3929));
  xnor_3 g03553(.A(new_n3929), .B(new_n3922), .Y(new_n3930));
  xnor_3 g03554(.A(new_n3930), .B(new_n3896), .Y(new_n3931));
  nor_4  g03555(.A(new_n3780), .B(new_n3752), .Y(new_n3932_1));
  not_3  g03556(.A(new_n3932_1), .Y(new_n3933));
  not_3  g03557(.A(new_n3709), .Y(new_n3934));
  not_3  g03558(.A(new_n3780), .Y(new_n3935));
  nor_4  g03559(.A(new_n3935), .B(new_n3751), .Y(new_n3936));
  nor_4  g03560(.A(new_n3932_1), .B(new_n3936), .Y(new_n3937));
  nand_4 g03561(.A(new_n3937), .B(new_n3934), .Y(new_n3938));
  nand_4 g03562(.A(new_n3938), .B(new_n3933), .Y(new_n3939));
  xnor_3 g03563(.A(new_n3939), .B(new_n3931), .Y(new_n3940));
  not_3  g03564(.A(new_n3742), .Y(new_n3941));
  not_3  g03565(.A(new_n3744), .Y(new_n3942));
  nor_4  g03566(.A(new_n3942), .B(new_n3941), .Y(new_n3943));
  nand_4 g03567(.A(n11296), .B(n7236), .Y(new_n3944));
  nand_4 g03568(.A(n8384), .B(n6611), .Y(new_n3945));
  nand_4 g03569(.A(n6359), .B(n3992), .Y(new_n3946));
  not_3  g03570(.A(new_n3946), .Y(new_n3947));
  xor_3  g03571(.A(new_n3947), .B(new_n3945), .Y(new_n3948));
  xnor_3 g03572(.A(new_n3948), .B(new_n3944), .Y(new_n3949));
  nand_4 g03573(.A(new_n3727), .B(new_n3721), .Y(new_n3950));
  not_3  g03574(.A(new_n3728), .Y(new_n3951));
  not_3  g03575(.A(new_n3731), .Y(new_n3952));
  nand_4 g03576(.A(new_n3952), .B(new_n3951), .Y(new_n3953));
  nand_4 g03577(.A(new_n3953), .B(new_n3950), .Y(new_n3954));
  xnor_3 g03578(.A(new_n3954), .B(new_n3949), .Y(new_n3955));
  nor_4  g03579(.A(new_n3730), .B(new_n3729), .Y(new_n3956));
  not_3  g03580(.A(new_n3956), .Y(new_n3957));
  nand_4 g03581(.A(n6358), .B(n217), .Y(new_n3958));
  xor_3  g03582(.A(new_n3958), .B(new_n3957), .Y(new_n3959));
  nand_4 g03583(.A(n1471), .B(n405), .Y(new_n3960));
  not_3  g03584(.A(new_n3960), .Y(new_n3961));
  nand_4 g03585(.A(n5198), .B(n4086), .Y(new_n3962));
  nand_4 g03586(.A(n8433), .B(n7646), .Y(new_n3963));
  xor_3  g03587(.A(new_n3963), .B(new_n3962), .Y(new_n3964));
  xnor_3 g03588(.A(new_n3964), .B(new_n3961), .Y(new_n3965));
  xnor_3 g03589(.A(new_n3965), .B(new_n3959), .Y(new_n3966));
  xnor_3 g03590(.A(new_n3966), .B(new_n3955), .Y(new_n3967));
  nand_4 g03591(.A(new_n3736), .B(new_n3733), .Y(new_n3968));
  nor_4  g03592(.A(new_n3735), .B(new_n3734), .Y(new_n3969));
  nor_4  g03593(.A(new_n3741), .B(new_n3737), .Y(new_n3970));
  xnor_3 g03594(.A(new_n3970), .B(new_n3969), .Y(new_n3971));
  nand_4 g03595(.A(new_n3971), .B(new_n3968), .Y(new_n3972));
  xnor_3 g03596(.A(new_n3972), .B(new_n3967), .Y(new_n3973));
  xnor_3 g03597(.A(new_n3973), .B(new_n3943), .Y(new_n3974));
  nand_4 g03598(.A(new_n3745), .B(new_n3718), .Y(new_n3975));
  nand_4 g03599(.A(new_n3748), .B(new_n3975), .Y(new_n3976));
  xnor_3 g03600(.A(new_n3976), .B(new_n3974), .Y(new_n3977));
  xnor_3 g03601(.A(new_n3977), .B(new_n3940), .Y(new_n3978));
  not_3  g03602(.A(new_n3782), .Y(new_n3979));
  nand_4 g03603(.A(new_n3979), .B(new_n3750), .Y(new_n3980));
  nand_4 g03604(.A(new_n3789), .B(new_n3783), .Y(new_n3981));
  nand_4 g03605(.A(new_n3981), .B(new_n3980), .Y(new_n3982));
  xnor_3 g03606(.A(new_n3982), .B(new_n3978), .Y(new_n3983));
  xnor_3 g03607(.A(new_n3983), .B(new_n3893), .Y(new_n3984));
  not_3  g03608(.A(new_n3984), .Y(new_n3985));
  not_3  g03609(.A(new_n3716), .Y(new_n3986_1));
  nand_4 g03610(.A(new_n3986_1), .B(new_n3503), .Y(new_n3987));
  not_3  g03611(.A(new_n3790), .Y(new_n3988));
  nand_4 g03612(.A(new_n3988), .B(new_n3717), .Y(new_n3989));
  nand_4 g03613(.A(new_n3989), .B(new_n3987), .Y(new_n3990));
  xnor_3 g03614(.A(new_n3990), .B(new_n3985), .Y(new_n3991));
  xnor_3 g03615(.A(new_n3991), .B(new_n3849_1), .Y(n844));
  nand_4 g03616(.A(n7456), .B(n6687), .Y(new_n3993));
  not_3  g03617(.A(new_n3993), .Y(new_n3994));
  nand_4 g03618(.A(n12591), .B(n6687), .Y(new_n3995));
  not_3  g03619(.A(new_n3995), .Y(new_n3996));
  nand_4 g03620(.A(n4189), .B(n1798), .Y(new_n3997));
  not_3  g03621(.A(new_n3997), .Y(new_n3998));
  nor_4  g03622(.A(new_n3998), .B(new_n3996), .Y(new_n3999));
  nor_4  g03623(.A(new_n3997), .B(new_n3995), .Y(new_n4000));
  nand_4 g03624(.A(n3932), .B(n2564), .Y(new_n4001));
  not_3  g03625(.A(new_n4001), .Y(new_n4002));
  nor_4  g03626(.A(new_n4002), .B(new_n4000), .Y(new_n4003));
  nor_4  g03627(.A(new_n4003), .B(new_n3999), .Y(new_n4004));
  nand_4 g03628(.A(new_n4004), .B(new_n3994), .Y(new_n4005_1));
  not_3  g03629(.A(new_n4005_1), .Y(new_n4006));
  nor_4  g03630(.A(new_n4004), .B(new_n3994), .Y(new_n4007));
  nor_4  g03631(.A(new_n4007), .B(new_n4006), .Y(new_n4008));
  nand_4 g03632(.A(n4189), .B(n3932), .Y(new_n4009));
  nand_4 g03633(.A(n12591), .B(n2564), .Y(new_n4010));
  not_3  g03634(.A(new_n4010), .Y(new_n4011));
  nand_4 g03635(.A(n6770), .B(n1798), .Y(new_n4012));
  not_3  g03636(.A(new_n4012), .Y(new_n4013));
  nor_4  g03637(.A(new_n4013), .B(new_n4011), .Y(new_n4014));
  nor_4  g03638(.A(new_n4012), .B(new_n4010), .Y(new_n4015));
  nor_4  g03639(.A(new_n4015), .B(new_n4014), .Y(new_n4016));
  xnor_3 g03640(.A(new_n4016), .B(new_n4009), .Y(new_n4017));
  xor_3  g03641(.A(new_n4017), .B(new_n4008), .Y(new_n4018));
  not_3  g03642(.A(new_n4018), .Y(new_n4019));
  nand_4 g03643(.A(n6687), .B(n1798), .Y(new_n4020));
  not_3  g03644(.A(new_n4020), .Y(new_n4021));
  nor_4  g03645(.A(new_n4021), .B(new_n4001), .Y(new_n4022));
  nor_4  g03646(.A(new_n4000), .B(new_n3999), .Y(new_n4023));
  nor_4  g03647(.A(new_n4023), .B(new_n4022), .Y(new_n4024));
  not_3  g03648(.A(new_n4024), .Y(new_n4025));
  nor_4  g03649(.A(new_n4025), .B(new_n4001), .Y(new_n4026));
  not_3  g03650(.A(new_n4026), .Y(new_n4027));
  xor_3  g03651(.A(new_n4027), .B(new_n4019), .Y(new_n4028));
  not_3  g03652(.A(new_n4028), .Y(new_n4029));
  nand_4 g03653(.A(n8336), .B(n6703), .Y(new_n4030));
  nand_4 g03654(.A(n11876), .B(n11222), .Y(new_n4031));
  not_3  g03655(.A(new_n4031), .Y(new_n4032));
  nand_4 g03656(.A(n12069), .B(n5645), .Y(new_n4033));
  xor_3  g03657(.A(new_n4033), .B(new_n4032), .Y(new_n4034));
  nor_4  g03658(.A(new_n4034), .B(new_n4030), .Y(new_n4035));
  nand_4 g03659(.A(n9640), .B(n8336), .Y(new_n4036));
  nand_4 g03660(.A(n10928), .B(n6703), .Y(new_n4037));
  not_3  g03661(.A(new_n4037), .Y(new_n4038));
  xor_3  g03662(.A(new_n4038), .B(new_n4036), .Y(new_n4039));
  not_3  g03663(.A(new_n4039), .Y(new_n4040));
  nand_4 g03664(.A(new_n4040), .B(new_n4035), .Y(new_n4041));
  not_3  g03665(.A(new_n4041), .Y(new_n4042));
  nor_4  g03666(.A(new_n4033), .B(new_n4031), .Y(new_n4043));
  not_3  g03667(.A(new_n4043), .Y(new_n4044));
  nand_4 g03668(.A(n12391), .B(n5645), .Y(new_n4045));
  nand_4 g03669(.A(n12069), .B(n1067), .Y(new_n4046));
  xnor_3 g03670(.A(new_n4046), .B(new_n4045), .Y(new_n4047));
  nor_4  g03671(.A(new_n4047), .B(new_n4044), .Y(new_n4048));
  not_3  g03672(.A(new_n4047), .Y(new_n4049));
  nor_4  g03673(.A(new_n4049), .B(new_n4043), .Y(new_n4050));
  nor_4  g03674(.A(new_n4050), .B(new_n4048), .Y(new_n4051));
  not_3  g03675(.A(new_n4051), .Y(new_n4052));
  nand_4 g03676(.A(n11222), .B(n10898), .Y(new_n4053));
  nand_4 g03677(.A(n11876), .B(n11153), .Y(new_n4054));
  xor_3  g03678(.A(new_n4054), .B(new_n4053), .Y(new_n4055));
  xnor_3 g03679(.A(new_n4055), .B(new_n4052), .Y(new_n4056));
  not_3  g03680(.A(new_n4056), .Y(new_n4057));
  not_3  g03681(.A(new_n4035), .Y(new_n4058));
  xor_3  g03682(.A(new_n4040), .B(new_n4058), .Y(new_n4059));
  nor_4  g03683(.A(new_n4059), .B(new_n4057), .Y(new_n4060));
  nor_4  g03684(.A(new_n4060), .B(new_n4042), .Y(new_n4061));
  not_3  g03685(.A(new_n4030), .Y(new_n4062));
  nand_4 g03686(.A(n10928), .B(n9640), .Y(new_n4063));
  nor_4  g03687(.A(new_n4063), .B(new_n4062), .Y(new_n4064));
  nand_4 g03688(.A(n6986), .B(n6703), .Y(new_n4065));
  nand_4 g03689(.A(n8336), .B(n3022), .Y(new_n4066));
  nand_4 g03690(.A(new_n4066), .B(new_n4065), .Y(new_n4067));
  and_4  g03691(.A(new_n4067), .B(new_n4064), .Y(new_n4068));
  nor_4  g03692(.A(new_n4066), .B(new_n4065), .Y(new_n4069));
  nor_4  g03693(.A(new_n4067), .B(new_n4064), .Y(new_n4070));
  nor_4  g03694(.A(new_n4070), .B(new_n4069), .Y(new_n4071));
  not_3  g03695(.A(new_n4071), .Y(new_n4072));
  nor_4  g03696(.A(new_n4072), .B(new_n4068), .Y(new_n4073));
  not_3  g03697(.A(new_n4073), .Y(new_n4074));
  xnor_3 g03698(.A(new_n4074), .B(new_n4061), .Y(new_n4075));
  nor_4  g03699(.A(new_n4046), .B(new_n4045), .Y(new_n4076));
  nand_4 g03700(.A(n12069), .B(n8665), .Y(new_n4077));
  not_3  g03701(.A(new_n4077), .Y(new_n4078));
  nand_4 g03702(.A(n12391), .B(n1067), .Y(new_n4079));
  nand_4 g03703(.A(n7891), .B(n5645), .Y(new_n4080));
  xnor_3 g03704(.A(new_n4080), .B(new_n4079), .Y(new_n4081));
  xor_3  g03705(.A(new_n4081), .B(new_n4078), .Y(new_n4082));
  not_3  g03706(.A(new_n4082), .Y(new_n4083));
  xor_3  g03707(.A(new_n4083), .B(new_n4076), .Y(new_n4084));
  nor_4  g03708(.A(new_n4055), .B(new_n4052), .Y(new_n4085));
  nor_4  g03709(.A(new_n4085), .B(new_n4050), .Y(new_n4086_1));
  nand_4 g03710(.A(n11876), .B(n5314), .Y(new_n4087));
  nand_4 g03711(.A(n11222), .B(n3754), .Y(new_n4088_1));
  nor_4  g03712(.A(new_n4088_1), .B(new_n4087), .Y(new_n4089));
  nand_4 g03713(.A(new_n4088_1), .B(new_n4087), .Y(new_n4090));
  nand_4 g03714(.A(n11153), .B(n10898), .Y(new_n4091));
  nor_4  g03715(.A(new_n4091), .B(new_n4032), .Y(new_n4092));
  nor_4  g03716(.A(new_n4092), .B(new_n4090), .Y(new_n4093));
  nor_4  g03717(.A(new_n4093), .B(new_n4089), .Y(new_n4094_1));
  not_3  g03718(.A(new_n4094_1), .Y(new_n4095));
  not_3  g03719(.A(new_n4090), .Y(new_n4096));
  not_3  g03720(.A(new_n4092), .Y(new_n4097));
  nor_4  g03721(.A(new_n4097), .B(new_n4096), .Y(new_n4098));
  nor_4  g03722(.A(new_n4098), .B(new_n4095), .Y(new_n4099));
  xnor_3 g03723(.A(new_n4099), .B(new_n4086_1), .Y(new_n4100));
  xnor_3 g03724(.A(new_n4100), .B(new_n4084), .Y(new_n4101));
  xnor_3 g03725(.A(new_n4101), .B(new_n4075), .Y(new_n4102));
  not_3  g03726(.A(new_n3999), .Y(new_n4103));
  nand_4 g03727(.A(new_n4022), .B(new_n4103), .Y(new_n4104));
  nand_4 g03728(.A(new_n4104), .B(new_n4025), .Y(new_n4105));
  not_3  g03729(.A(new_n4105), .Y(new_n4106));
  nand_4 g03730(.A(new_n4106), .B(new_n4102), .Y(new_n4107));
  xor_3  g03731(.A(new_n4033), .B(new_n4031), .Y(new_n4108));
  xor_3  g03732(.A(new_n4108), .B(new_n4062), .Y(new_n4109));
  nand_4 g03733(.A(new_n4109), .B(new_n4021), .Y(new_n4110));
  not_3  g03734(.A(new_n4110), .Y(new_n4111));
  nand_4 g03735(.A(n2564), .B(n1798), .Y(new_n4112));
  nand_4 g03736(.A(n6687), .B(n3932), .Y(new_n4113));
  xor_3  g03737(.A(new_n4113), .B(new_n4112), .Y(new_n4114));
  nor_4  g03738(.A(new_n4114), .B(new_n4111), .Y(new_n4115));
  and_4  g03739(.A(new_n4059), .B(new_n4057), .Y(new_n4116));
  nor_4  g03740(.A(new_n4116), .B(new_n4060), .Y(new_n4117));
  not_3  g03741(.A(new_n4114), .Y(new_n4118));
  xor_3  g03742(.A(new_n4118), .B(new_n4111), .Y(new_n4119));
  nor_4  g03743(.A(new_n4119), .B(new_n4117), .Y(new_n4120));
  nor_4  g03744(.A(new_n4120), .B(new_n4115), .Y(new_n4121));
  xnor_3 g03745(.A(new_n4105), .B(new_n4102), .Y(new_n4122));
  nand_4 g03746(.A(new_n4122), .B(new_n4121), .Y(new_n4123));
  nand_4 g03747(.A(new_n4123), .B(new_n4107), .Y(new_n4124));
  xnor_3 g03748(.A(new_n4124), .B(new_n4029), .Y(new_n4125));
  not_3  g03749(.A(new_n4076), .Y(new_n4126));
  nor_4  g03750(.A(new_n4082), .B(new_n4126), .Y(new_n4127));
  nand_4 g03751(.A(n12069), .B(n11922), .Y(new_n4128));
  not_3  g03752(.A(new_n4128), .Y(new_n4129));
  not_3  g03753(.A(new_n4079), .Y(new_n4130));
  not_3  g03754(.A(new_n4080), .Y(new_n4131));
  nor_4  g03755(.A(new_n4131), .B(new_n4130), .Y(new_n4132));
  nor_4  g03756(.A(new_n4081), .B(new_n4078), .Y(new_n4133));
  nor_4  g03757(.A(new_n4133), .B(new_n4132), .Y(new_n4134));
  xnor_3 g03758(.A(new_n4134), .B(new_n4129), .Y(new_n4135));
  nand_4 g03759(.A(n7160), .B(n5645), .Y(new_n4136));
  nand_4 g03760(.A(n7891), .B(n1067), .Y(new_n4137));
  nand_4 g03761(.A(n12391), .B(n8665), .Y(new_n4138));
  nand_4 g03762(.A(new_n4138), .B(new_n4137), .Y(new_n4139));
  nor_4  g03763(.A(new_n4138), .B(new_n4137), .Y(new_n4140));
  not_3  g03764(.A(new_n4140), .Y(new_n4141_1));
  nand_4 g03765(.A(new_n4141_1), .B(new_n4139), .Y(new_n4142));
  xnor_3 g03766(.A(new_n4142), .B(new_n4136), .Y(new_n4143));
  xnor_3 g03767(.A(new_n4143), .B(new_n4135), .Y(new_n4144));
  xnor_3 g03768(.A(new_n4144), .B(new_n4127), .Y(new_n4145));
  nand_4 g03769(.A(n11222), .B(n2749), .Y(new_n4146));
  not_3  g03770(.A(new_n4146), .Y(new_n4147));
  not_3  g03771(.A(new_n4091), .Y(new_n4148));
  nor_4  g03772(.A(new_n4148), .B(new_n4089), .Y(new_n4149));
  nor_4  g03773(.A(new_n4149), .B(new_n4096), .Y(new_n4150));
  xnor_3 g03774(.A(new_n4150), .B(new_n4147), .Y(new_n4151));
  nand_4 g03775(.A(n10898), .B(n5314), .Y(new_n4152));
  nand_4 g03776(.A(n11153), .B(n3754), .Y(new_n4153));
  not_3  g03777(.A(new_n4153), .Y(new_n4154));
  nand_4 g03778(.A(n11876), .B(n996), .Y(new_n4155_1));
  not_3  g03779(.A(new_n4155_1), .Y(new_n4156));
  nor_4  g03780(.A(new_n4156), .B(new_n4154), .Y(new_n4157));
  nor_4  g03781(.A(new_n4155_1), .B(new_n4153), .Y(new_n4158));
  nor_4  g03782(.A(new_n4158), .B(new_n4157), .Y(new_n4159_1));
  xnor_3 g03783(.A(new_n4159_1), .B(new_n4152), .Y(new_n4160));
  not_3  g03784(.A(new_n4160), .Y(new_n4161));
  xnor_3 g03785(.A(new_n4161), .B(new_n4151), .Y(new_n4162));
  nor_4  g03786(.A(new_n4094_1), .B(new_n4091), .Y(new_n4163));
  not_3  g03787(.A(new_n4163), .Y(new_n4164));
  nor_4  g03788(.A(new_n4164), .B(new_n4162), .Y(new_n4165));
  not_3  g03789(.A(new_n4162), .Y(new_n4166));
  nor_4  g03790(.A(new_n4163), .B(new_n4166), .Y(new_n4167));
  nor_4  g03791(.A(new_n4167), .B(new_n4165), .Y(new_n4168));
  nor_4  g03792(.A(new_n4168), .B(new_n4145), .Y(new_n4169));
  not_3  g03793(.A(new_n4144), .Y(new_n4170));
  xnor_3 g03794(.A(new_n4170), .B(new_n4127), .Y(new_n4171));
  not_3  g03795(.A(new_n4168), .Y(new_n4172));
  nor_4  g03796(.A(new_n4172), .B(new_n4171), .Y(new_n4173));
  nor_4  g03797(.A(new_n4173), .B(new_n4169), .Y(new_n4174));
  nor_4  g03798(.A(new_n4099), .B(new_n4086_1), .Y(new_n4175));
  nor_4  g03799(.A(new_n4100), .B(new_n4084), .Y(new_n4176));
  nor_4  g03800(.A(new_n4176), .B(new_n4175), .Y(new_n4177));
  not_3  g03801(.A(new_n4177), .Y(new_n4178));
  nor_4  g03802(.A(new_n4178), .B(new_n4174), .Y(new_n4179));
  nand_4 g03803(.A(new_n4178), .B(new_n4174), .Y(new_n4180));
  not_3  g03804(.A(new_n4180), .Y(new_n4181));
  nor_4  g03805(.A(new_n4181), .B(new_n4179), .Y(new_n4182));
  not_3  g03806(.A(new_n4182), .Y(new_n4183));
  nand_4 g03807(.A(n11023), .B(n8336), .Y(new_n4184));
  not_3  g03808(.A(new_n4069), .Y(new_n4185));
  not_3  g03809(.A(new_n4063), .Y(new_n4186));
  nand_4 g03810(.A(new_n4067), .B(new_n4186), .Y(new_n4187_1));
  nand_4 g03811(.A(new_n4187_1), .B(new_n4185), .Y(new_n4188));
  not_3  g03812(.A(new_n4188), .Y(new_n4189_1));
  xor_3  g03813(.A(new_n4189_1), .B(new_n4184), .Y(new_n4190_1));
  nand_4 g03814(.A(n9640), .B(n6986), .Y(new_n4191));
  not_3  g03815(.A(new_n4191), .Y(new_n4192));
  nand_4 g03816(.A(n10928), .B(n3022), .Y(new_n4193));
  not_3  g03817(.A(new_n4193), .Y(new_n4194));
  nand_4 g03818(.A(n6703), .B(n2226), .Y(new_n4195));
  not_3  g03819(.A(new_n4195), .Y(new_n4196));
  nor_4  g03820(.A(new_n4196), .B(new_n4194), .Y(new_n4197));
  nor_4  g03821(.A(new_n4195), .B(new_n4193), .Y(new_n4198));
  nor_4  g03822(.A(new_n4198), .B(new_n4197), .Y(new_n4199));
  xor_3  g03823(.A(new_n4199), .B(new_n4192), .Y(new_n4200));
  xnor_3 g03824(.A(new_n4200), .B(new_n4190_1), .Y(new_n4201));
  not_3  g03825(.A(new_n4201), .Y(new_n4202));
  nor_4  g03826(.A(new_n4071), .B(new_n4063), .Y(new_n4203_1));
  xor_3  g03827(.A(new_n4203_1), .B(new_n4202), .Y(new_n4204));
  nand_4 g03828(.A(new_n4074), .B(new_n4061), .Y(new_n4205));
  not_3  g03829(.A(new_n4205), .Y(new_n4206));
  nor_4  g03830(.A(new_n4101), .B(new_n4075), .Y(new_n4207));
  nor_4  g03831(.A(new_n4207), .B(new_n4206), .Y(new_n4208));
  nand_4 g03832(.A(new_n4208), .B(new_n4204), .Y(new_n4209));
  not_3  g03833(.A(new_n4209), .Y(new_n4210));
  nor_4  g03834(.A(new_n4208), .B(new_n4204), .Y(new_n4211));
  nor_4  g03835(.A(new_n4211), .B(new_n4210), .Y(new_n4212));
  nor_4  g03836(.A(new_n4212), .B(new_n4183), .Y(new_n4213));
  nand_4 g03837(.A(new_n4212), .B(new_n4183), .Y(new_n4214));
  not_3  g03838(.A(new_n4214), .Y(new_n4215));
  nor_4  g03839(.A(new_n4215), .B(new_n4213), .Y(new_n4216));
  xor_3  g03840(.A(new_n4216), .B(new_n4125), .Y(n911));
  nand_4 g03841(.A(n9956), .B(n4189), .Y(new_n4218));
  nand_4 g03842(.A(n11917), .B(n6687), .Y(new_n4219));
  nand_4 g03843(.A(new_n4219), .B(new_n4218), .Y(new_n4220));
  nor_4  g03844(.A(new_n4219), .B(new_n4218), .Y(new_n4221));
  not_3  g03845(.A(new_n4221), .Y(new_n4222));
  and_4  g03846(.A(new_n4222), .B(new_n4220), .Y(new_n4223));
  nand_4 g03847(.A(n9956), .B(n2564), .Y(new_n4224));
  nand_4 g03848(.A(n6687), .B(n4921), .Y(new_n4225));
  nor_4  g03849(.A(new_n4225), .B(new_n4224), .Y(new_n4226_1));
  not_3  g03850(.A(new_n4226_1), .Y(new_n4227));
  nor_4  g03851(.A(new_n4227), .B(new_n4223), .Y(new_n4228));
  not_3  g03852(.A(new_n4228), .Y(new_n4229));
  nand_4 g03853(.A(n6687), .B(n3842), .Y(new_n4230_1));
  nand_4 g03854(.A(n4921), .B(n2564), .Y(new_n4231));
  not_3  g03855(.A(new_n4231), .Y(new_n4232));
  nand_4 g03856(.A(new_n4232), .B(new_n4220), .Y(new_n4233));
  nand_4 g03857(.A(new_n4233), .B(new_n4222), .Y(new_n4234));
  not_3  g03858(.A(new_n4234), .Y(new_n4235));
  xor_3  g03859(.A(new_n4235), .B(new_n4230_1), .Y(new_n4236));
  nand_4 g03860(.A(n4921), .B(n4189), .Y(new_n4237));
  not_3  g03861(.A(new_n4237), .Y(new_n4238));
  nand_4 g03862(.A(n11917), .B(n2564), .Y(new_n4239));
  not_3  g03863(.A(new_n4239), .Y(new_n4240));
  nand_4 g03864(.A(n9956), .B(n6770), .Y(new_n4241));
  not_3  g03865(.A(new_n4241), .Y(new_n4242));
  nor_4  g03866(.A(new_n4242), .B(new_n4240), .Y(new_n4243));
  nor_4  g03867(.A(new_n4241), .B(new_n4239), .Y(new_n4244));
  nor_4  g03868(.A(new_n4244), .B(new_n4243), .Y(new_n4245));
  xor_3  g03869(.A(new_n4245), .B(new_n4238), .Y(new_n4246));
  xnor_3 g03870(.A(new_n4246), .B(new_n4236), .Y(new_n4247));
  nor_4  g03871(.A(new_n4247), .B(new_n4229), .Y(new_n4248));
  not_3  g03872(.A(new_n4248), .Y(new_n4249));
  nand_4 g03873(.A(n6687), .B(n2577), .Y(new_n4250));
  nor_4  g03874(.A(new_n4235), .B(new_n4230_1), .Y(new_n4251));
  not_3  g03875(.A(new_n4251), .Y(new_n4252));
  nand_4 g03876(.A(new_n4246), .B(new_n4236), .Y(new_n4253));
  nand_4 g03877(.A(new_n4253), .B(new_n4252), .Y(new_n4254));
  not_3  g03878(.A(new_n4254), .Y(new_n4255));
  xor_3  g03879(.A(new_n4255), .B(new_n4250), .Y(new_n4256));
  nand_4 g03880(.A(n3842), .B(n2564), .Y(new_n4257));
  nor_4  g03881(.A(new_n4244), .B(new_n4238), .Y(new_n4258));
  nor_4  g03882(.A(new_n4258), .B(new_n4243), .Y(new_n4259));
  xor_3  g03883(.A(new_n4259), .B(new_n4257), .Y(new_n4260));
  not_3  g03884(.A(new_n4260), .Y(new_n4261));
  nand_4 g03885(.A(n6770), .B(n4921), .Y(new_n4262));
  nand_4 g03886(.A(n11917), .B(n4189), .Y(new_n4263));
  nand_4 g03887(.A(n9956), .B(n9920), .Y(new_n4264));
  not_3  g03888(.A(new_n4264), .Y(new_n4265));
  xor_3  g03889(.A(new_n4265), .B(new_n4263), .Y(new_n4266));
  xnor_3 g03890(.A(new_n4266), .B(new_n4262), .Y(new_n4267));
  not_3  g03891(.A(new_n4267), .Y(new_n4268));
  xor_3  g03892(.A(new_n4268), .B(new_n4261), .Y(new_n4269));
  xnor_3 g03893(.A(new_n4269), .B(new_n4256), .Y(new_n4270));
  xnor_3 g03894(.A(new_n4270), .B(new_n4249), .Y(new_n4271));
  not_3  g03895(.A(new_n4247), .Y(new_n4272));
  xor_3  g03896(.A(new_n4272), .B(new_n4229), .Y(new_n4273));
  not_3  g03897(.A(new_n4273), .Y(new_n4274));
  nand_4 g03898(.A(n8595), .B(n8336), .Y(new_n4275));
  not_3  g03899(.A(new_n4275), .Y(new_n4276));
  nand_4 g03900(.A(n8336), .B(n6126), .Y(new_n4277));
  not_3  g03901(.A(new_n4277), .Y(new_n4278));
  nand_4 g03902(.A(n6986), .B(n3719), .Y(new_n4279));
  not_3  g03903(.A(new_n4279), .Y(new_n4280));
  nor_4  g03904(.A(new_n4280), .B(new_n4278), .Y(new_n4281));
  nor_4  g03905(.A(new_n4279), .B(new_n4277), .Y(new_n4282));
  nand_4 g03906(.A(n10928), .B(n3602), .Y(new_n4283));
  not_3  g03907(.A(new_n4283), .Y(new_n4284));
  nor_4  g03908(.A(new_n4284), .B(new_n4282), .Y(new_n4285));
  nor_4  g03909(.A(new_n4285), .B(new_n4281), .Y(new_n4286));
  nand_4 g03910(.A(new_n4286), .B(new_n4276), .Y(new_n4287));
  not_3  g03911(.A(new_n4287), .Y(new_n4288));
  nor_4  g03912(.A(new_n4286), .B(new_n4276), .Y(new_n4289));
  nor_4  g03913(.A(new_n4289), .B(new_n4288), .Y(new_n4290));
  nand_4 g03914(.A(n6986), .B(n3602), .Y(new_n4291));
  not_3  g03915(.A(new_n4291), .Y(new_n4292));
  nand_4 g03916(.A(n10928), .B(n6126), .Y(new_n4293));
  nand_4 g03917(.A(n3719), .B(n2226), .Y(new_n4294));
  not_3  g03918(.A(new_n4294), .Y(new_n4295));
  xor_3  g03919(.A(new_n4295), .B(new_n4293), .Y(new_n4296));
  xnor_3 g03920(.A(new_n4296), .B(new_n4292), .Y(new_n4297));
  nand_4 g03921(.A(new_n4297), .B(new_n4290), .Y(new_n4298));
  not_3  g03922(.A(new_n4290), .Y(new_n4299));
  xnor_3 g03923(.A(new_n4296), .B(new_n4291), .Y(new_n4300_1));
  nand_4 g03924(.A(new_n4300_1), .B(new_n4299), .Y(new_n4301));
  nand_4 g03925(.A(new_n4301), .B(new_n4298), .Y(new_n4302));
  nand_4 g03926(.A(n8336), .B(n3719), .Y(new_n4303));
  not_3  g03927(.A(new_n4303), .Y(new_n4304));
  nor_4  g03928(.A(new_n4304), .B(new_n4283), .Y(new_n4305));
  nor_4  g03929(.A(new_n4282), .B(new_n4281), .Y(new_n4306));
  nor_4  g03930(.A(new_n4306), .B(new_n4305), .Y(new_n4307));
  not_3  g03931(.A(new_n4307), .Y(new_n4308));
  nor_4  g03932(.A(new_n4308), .B(new_n4283), .Y(new_n4309));
  xnor_3 g03933(.A(new_n4309), .B(new_n4302), .Y(new_n4310));
  nand_4 g03934(.A(n12925), .B(n7891), .Y(new_n4311));
  nand_4 g03935(.A(n12069), .B(n4826), .Y(new_n4312_1));
  nand_4 g03936(.A(new_n4312_1), .B(new_n4311), .Y(new_n4313));
  not_3  g03937(.A(new_n4313), .Y(new_n4314));
  not_3  g03938(.A(new_n4311), .Y(new_n4315));
  not_3  g03939(.A(new_n4312_1), .Y(new_n4316));
  nand_4 g03940(.A(new_n4316), .B(new_n4315), .Y(new_n4317));
  not_3  g03941(.A(new_n4317), .Y(new_n4318));
  nor_4  g03942(.A(new_n4318), .B(new_n4314), .Y(new_n4319));
  nand_4 g03943(.A(n12069), .B(n7733), .Y(new_n4320));
  nand_4 g03944(.A(n12925), .B(n12391), .Y(new_n4321));
  nor_4  g03945(.A(new_n4321), .B(new_n4320), .Y(new_n4322));
  not_3  g03946(.A(new_n4322), .Y(new_n4323));
  nor_4  g03947(.A(new_n4323), .B(new_n4319), .Y(new_n4324));
  not_3  g03948(.A(new_n4324), .Y(new_n4325));
  nand_4 g03949(.A(n12069), .B(n7610), .Y(new_n4326_1));
  nand_4 g03950(.A(n12391), .B(n7733), .Y(new_n4327));
  not_3  g03951(.A(new_n4327), .Y(new_n4328));
  nand_4 g03952(.A(new_n4328), .B(new_n4313), .Y(new_n4329));
  nand_4 g03953(.A(new_n4329), .B(new_n4317), .Y(new_n4330));
  not_3  g03954(.A(new_n4330), .Y(new_n4331));
  xnor_3 g03955(.A(new_n4331), .B(new_n4326_1), .Y(new_n4332));
  nand_4 g03956(.A(n12925), .B(n7160), .Y(new_n4333_1));
  not_3  g03957(.A(new_n4333_1), .Y(new_n4334));
  nand_4 g03958(.A(n12391), .B(n4826), .Y(new_n4335));
  not_3  g03959(.A(new_n4335), .Y(new_n4336));
  nand_4 g03960(.A(n7891), .B(n7733), .Y(new_n4337));
  not_3  g03961(.A(new_n4337), .Y(new_n4338));
  nor_4  g03962(.A(new_n4338), .B(new_n4336), .Y(new_n4339));
  nor_4  g03963(.A(new_n4337), .B(new_n4335), .Y(new_n4340));
  nor_4  g03964(.A(new_n4340), .B(new_n4339), .Y(new_n4341));
  xnor_3 g03965(.A(new_n4341), .B(new_n4334), .Y(new_n4342));
  xnor_3 g03966(.A(new_n4342), .B(new_n4332), .Y(new_n4343));
  nor_4  g03967(.A(new_n4343), .B(new_n4325), .Y(new_n4344));
  not_3  g03968(.A(new_n4343), .Y(new_n4345));
  nor_4  g03969(.A(new_n4345), .B(new_n4324), .Y(new_n4346));
  nor_4  g03970(.A(new_n4346), .B(new_n4344), .Y(new_n4347));
  nand_4 g03971(.A(n11222), .B(n217), .Y(new_n4348));
  not_3  g03972(.A(new_n4348), .Y(new_n4349));
  nand_4 g03973(.A(n8433), .B(n5314), .Y(new_n4350));
  not_3  g03974(.A(new_n4350), .Y(new_n4351));
  nand_4 g03975(.A(n11222), .B(n4086), .Y(new_n4352));
  not_3  g03976(.A(new_n4352), .Y(new_n4353));
  nor_4  g03977(.A(new_n4353), .B(new_n4351), .Y(new_n4354));
  nor_4  g03978(.A(new_n4352), .B(new_n4350), .Y(new_n4355));
  nand_4 g03979(.A(n11153), .B(n405), .Y(new_n4356));
  not_3  g03980(.A(new_n4356), .Y(new_n4357));
  nor_4  g03981(.A(new_n4357), .B(new_n4355), .Y(new_n4358));
  nor_4  g03982(.A(new_n4358), .B(new_n4354), .Y(new_n4359));
  xnor_3 g03983(.A(new_n4359), .B(new_n4349), .Y(new_n4360));
  nand_4 g03984(.A(n5314), .B(n405), .Y(new_n4361));
  nand_4 g03985(.A(n8433), .B(n996), .Y(new_n4362));
  nand_4 g03986(.A(n11153), .B(n4086), .Y(new_n4363));
  xnor_3 g03987(.A(new_n4363), .B(new_n4362), .Y(new_n4364));
  xnor_3 g03988(.A(new_n4364), .B(new_n4361), .Y(new_n4365));
  xnor_3 g03989(.A(new_n4365), .B(new_n4360), .Y(new_n4366));
  not_3  g03990(.A(new_n4355), .Y(new_n4367));
  nand_4 g03991(.A(n11222), .B(n8433), .Y(new_n4368));
  nand_4 g03992(.A(new_n4368), .B(new_n4357), .Y(new_n4369));
  nand_4 g03993(.A(new_n4369), .B(new_n4354), .Y(new_n4370_1));
  nand_4 g03994(.A(new_n4370_1), .B(new_n4367), .Y(new_n4371));
  not_3  g03995(.A(new_n4371), .Y(new_n4372));
  nor_4  g03996(.A(new_n4372), .B(new_n4356), .Y(new_n4373));
  not_3  g03997(.A(new_n4373), .Y(new_n4374));
  nor_4  g03998(.A(new_n4374), .B(new_n4366), .Y(new_n4375));
  not_3  g03999(.A(new_n4366), .Y(new_n4376));
  nor_4  g04000(.A(new_n4373), .B(new_n4376), .Y(new_n4377));
  nor_4  g04001(.A(new_n4377), .B(new_n4375), .Y(new_n4378_1));
  not_3  g04002(.A(new_n4378_1), .Y(new_n4379));
  xnor_3 g04003(.A(new_n4379), .B(new_n4347), .Y(new_n4380));
  nand_4 g04004(.A(n12925), .B(n12069), .Y(new_n4381));
  nor_4  g04005(.A(new_n4381), .B(new_n4368), .Y(new_n4382));
  not_3  g04006(.A(new_n4382), .Y(new_n4383));
  nand_4 g04007(.A(n11153), .B(n8433), .Y(new_n4384));
  nand_4 g04008(.A(n11222), .B(n405), .Y(new_n4385));
  xnor_3 g04009(.A(new_n4385), .B(new_n4384), .Y(new_n4386));
  nand_4 g04010(.A(new_n4386), .B(new_n4383), .Y(new_n4387));
  not_3  g04011(.A(new_n4387), .Y(new_n4388));
  nor_4  g04012(.A(new_n4386), .B(new_n4383), .Y(new_n4389));
  nor_4  g04013(.A(new_n4389), .B(new_n4388), .Y(new_n4390));
  xnor_3 g04014(.A(new_n4321), .B(new_n4320), .Y(new_n4391));
  nand_4 g04015(.A(new_n4391), .B(new_n4390), .Y(new_n4392));
  nand_4 g04016(.A(new_n4392), .B(new_n4387), .Y(new_n4393));
  not_3  g04017(.A(new_n4393), .Y(new_n4394));
  nor_4  g04018(.A(new_n4369), .B(new_n4354), .Y(new_n4395));
  nor_4  g04019(.A(new_n4395), .B(new_n4371), .Y(new_n4396));
  nor_4  g04020(.A(new_n4396), .B(new_n4394), .Y(new_n4397_1));
  not_3  g04021(.A(new_n4397_1), .Y(new_n4398));
  not_3  g04022(.A(new_n4396), .Y(new_n4399));
  nor_4  g04023(.A(new_n4399), .B(new_n4393), .Y(new_n4400));
  nor_4  g04024(.A(new_n4400), .B(new_n4397_1), .Y(new_n4401));
  not_3  g04025(.A(new_n4319), .Y(new_n4402));
  not_3  g04026(.A(new_n4381), .Y(new_n4403));
  nor_4  g04027(.A(new_n4403), .B(new_n4327), .Y(new_n4404));
  not_3  g04028(.A(new_n4404), .Y(new_n4405));
  nand_4 g04029(.A(new_n4405), .B(new_n4402), .Y(new_n4406));
  nand_4 g04030(.A(new_n4404), .B(new_n4313), .Y(new_n4407));
  nand_4 g04031(.A(new_n4407), .B(new_n4406), .Y(new_n4408));
  nand_4 g04032(.A(new_n4408), .B(new_n4401), .Y(new_n4409));
  nand_4 g04033(.A(new_n4409), .B(new_n4398), .Y(new_n4410));
  xnor_3 g04034(.A(new_n4410), .B(new_n4380), .Y(new_n4411));
  xnor_3 g04035(.A(new_n4411), .B(new_n4310), .Y(new_n4412));
  xnor_3 g04036(.A(new_n4408), .B(new_n4401), .Y(new_n4413));
  not_3  g04037(.A(new_n4413), .Y(new_n4414));
  not_3  g04038(.A(new_n4281), .Y(new_n4415));
  nand_4 g04039(.A(new_n4305), .B(new_n4415), .Y(new_n4416));
  nand_4 g04040(.A(new_n4416), .B(new_n4308), .Y(new_n4417));
  nor_4  g04041(.A(new_n4417), .B(new_n4414), .Y(new_n4418));
  xnor_3 g04042(.A(new_n4417), .B(new_n4414), .Y(new_n4419));
  xnor_3 g04043(.A(new_n4391), .B(new_n4390), .Y(new_n4420));
  not_3  g04044(.A(new_n4420), .Y(new_n4421));
  nand_4 g04045(.A(n10928), .B(n3719), .Y(new_n4422));
  nand_4 g04046(.A(n8336), .B(n3602), .Y(new_n4423));
  not_3  g04047(.A(new_n4423), .Y(new_n4424));
  xor_3  g04048(.A(new_n4424), .B(new_n4422), .Y(new_n4425));
  nor_4  g04049(.A(new_n4425), .B(new_n4421), .Y(new_n4426));
  xor_3  g04050(.A(new_n4381), .B(new_n4368), .Y(new_n4427));
  nand_4 g04051(.A(new_n4427), .B(new_n4304), .Y(new_n4428));
  xnor_3 g04052(.A(new_n4425), .B(new_n4421), .Y(new_n4429));
  nor_4  g04053(.A(new_n4429), .B(new_n4428), .Y(new_n4430));
  nor_4  g04054(.A(new_n4430), .B(new_n4426), .Y(new_n4431));
  nor_4  g04055(.A(new_n4431), .B(new_n4419), .Y(new_n4432));
  nor_4  g04056(.A(new_n4432), .B(new_n4418), .Y(new_n4433));
  xnor_3 g04057(.A(new_n4433), .B(new_n4412), .Y(new_n4434));
  not_3  g04058(.A(new_n4434), .Y(new_n4435));
  nand_4 g04059(.A(new_n4435), .B(new_n4274), .Y(new_n4436_1));
  nand_4 g04060(.A(new_n4434), .B(new_n4273), .Y(new_n4437));
  xnor_3 g04061(.A(new_n4431), .B(new_n4419), .Y(new_n4438));
  not_3  g04062(.A(new_n4438), .Y(new_n4439));
  not_3  g04063(.A(new_n4223), .Y(new_n4440));
  nand_4 g04064(.A(n9956), .B(n6687), .Y(new_n4441));
  not_3  g04065(.A(new_n4441), .Y(new_n4442));
  nor_4  g04066(.A(new_n4442), .B(new_n4231), .Y(new_n4443));
  not_3  g04067(.A(new_n4443), .Y(new_n4444));
  nand_4 g04068(.A(new_n4444), .B(new_n4440), .Y(new_n4445));
  nand_4 g04069(.A(new_n4443), .B(new_n4220), .Y(new_n4446));
  nand_4 g04070(.A(new_n4446), .B(new_n4445), .Y(new_n4447));
  not_3  g04071(.A(new_n4447), .Y(new_n4448));
  nor_4  g04072(.A(new_n4448), .B(new_n4439), .Y(new_n4449));
  xnor_3 g04073(.A(new_n4447), .B(new_n4438), .Y(new_n4450));
  not_3  g04074(.A(new_n4428), .Y(new_n4451));
  nor_4  g04075(.A(new_n4427), .B(new_n4304), .Y(new_n4452));
  nor_4  g04076(.A(new_n4452), .B(new_n4451), .Y(new_n4453));
  nand_4 g04077(.A(new_n4453), .B(new_n4442), .Y(new_n4454));
  not_3  g04078(.A(new_n4454), .Y(new_n4455));
  xor_3  g04079(.A(new_n4225), .B(new_n4224), .Y(new_n4456));
  nor_4  g04080(.A(new_n4456), .B(new_n4455), .Y(new_n4457));
  not_3  g04081(.A(new_n4429), .Y(new_n4458));
  nor_4  g04082(.A(new_n4458), .B(new_n4451), .Y(new_n4459));
  nor_4  g04083(.A(new_n4459), .B(new_n4430), .Y(new_n4460));
  xnor_3 g04084(.A(new_n4456), .B(new_n4455), .Y(new_n4461));
  nor_4  g04085(.A(new_n4461), .B(new_n4460), .Y(new_n4462));
  nor_4  g04086(.A(new_n4462), .B(new_n4457), .Y(new_n4463));
  nor_4  g04087(.A(new_n4463), .B(new_n4450), .Y(new_n4464));
  nor_4  g04088(.A(new_n4464), .B(new_n4449), .Y(new_n4465));
  nand_4 g04089(.A(new_n4465), .B(new_n4437), .Y(new_n4466));
  nand_4 g04090(.A(new_n4466), .B(new_n4436_1), .Y(new_n4467));
  xnor_3 g04091(.A(new_n4467), .B(new_n4271), .Y(new_n4468));
  not_3  g04092(.A(new_n4309), .Y(new_n4469));
  nor_4  g04093(.A(new_n4469), .B(new_n4302), .Y(new_n4470));
  nand_4 g04094(.A(n10439), .B(n8336), .Y(new_n4471));
  not_3  g04095(.A(new_n4471), .Y(new_n4472));
  nand_4 g04096(.A(new_n4298), .B(new_n4287), .Y(new_n4473));
  xnor_3 g04097(.A(new_n4473), .B(new_n4472), .Y(new_n4474));
  nand_4 g04098(.A(n10928), .B(n8595), .Y(new_n4475));
  not_3  g04099(.A(new_n4475), .Y(new_n4476));
  not_3  g04100(.A(new_n4293), .Y(new_n4477));
  nor_4  g04101(.A(new_n4295), .B(new_n4477), .Y(new_n4478));
  nor_4  g04102(.A(new_n4294), .B(new_n4293), .Y(new_n4479));
  nor_4  g04103(.A(new_n4479), .B(new_n4292), .Y(new_n4480));
  nor_4  g04104(.A(new_n4480), .B(new_n4478), .Y(new_n4481));
  xor_3  g04105(.A(new_n4481), .B(new_n4476), .Y(new_n4482));
  not_3  g04106(.A(new_n4482), .Y(new_n4483));
  nand_4 g04107(.A(n3602), .B(n2226), .Y(new_n4484));
  not_3  g04108(.A(new_n4484), .Y(new_n4485));
  nand_4 g04109(.A(n6986), .B(n6126), .Y(new_n4486));
  nand_4 g04110(.A(n3719), .B(n1094), .Y(new_n4487));
  xnor_3 g04111(.A(new_n4487), .B(new_n4486), .Y(new_n4488));
  xor_3  g04112(.A(new_n4488), .B(new_n4485), .Y(new_n4489));
  not_3  g04113(.A(new_n4489), .Y(new_n4490));
  xor_3  g04114(.A(new_n4490), .B(new_n4483), .Y(new_n4491));
  nor_4  g04115(.A(new_n4491), .B(new_n4474), .Y(new_n4492));
  xnor_3 g04116(.A(new_n4473), .B(new_n4471), .Y(new_n4493));
  not_3  g04117(.A(new_n4491), .Y(new_n4494));
  nor_4  g04118(.A(new_n4494), .B(new_n4493), .Y(new_n4495));
  nor_4  g04119(.A(new_n4495), .B(new_n4492), .Y(new_n4496));
  xnor_3 g04120(.A(new_n4496), .B(new_n4470), .Y(new_n4497));
  not_3  g04121(.A(new_n4375), .Y(new_n4498));
  nand_4 g04122(.A(n11222), .B(n6611), .Y(new_n4499_1));
  not_3  g04123(.A(new_n4499_1), .Y(new_n4500));
  nand_4 g04124(.A(n11153), .B(n217), .Y(new_n4501));
  nand_4 g04125(.A(n996), .B(n405), .Y(new_n4502));
  nand_4 g04126(.A(n5314), .B(n4086), .Y(new_n4503));
  not_3  g04127(.A(new_n4503), .Y(new_n4504));
  nand_4 g04128(.A(n8433), .B(n5767), .Y(new_n4505));
  not_3  g04129(.A(new_n4505), .Y(new_n4506));
  nor_4  g04130(.A(new_n4506), .B(new_n4504), .Y(new_n4507));
  nor_4  g04131(.A(new_n4505), .B(new_n4503), .Y(new_n4508));
  nor_4  g04132(.A(new_n4508), .B(new_n4507), .Y(new_n4509));
  xnor_3 g04133(.A(new_n4509), .B(new_n4502), .Y(new_n4510));
  xnor_3 g04134(.A(new_n4510), .B(new_n4501), .Y(new_n4511));
  not_3  g04135(.A(new_n4511), .Y(new_n4512));
  and_4  g04136(.A(new_n4363), .B(new_n4362), .Y(new_n4513));
  not_3  g04137(.A(new_n4361), .Y(new_n4514));
  nor_4  g04138(.A(new_n4363), .B(new_n4362), .Y(new_n4515));
  nor_4  g04139(.A(new_n4515), .B(new_n4514), .Y(new_n4516_1));
  nor_4  g04140(.A(new_n4516_1), .B(new_n4513), .Y(new_n4517));
  xnor_3 g04141(.A(new_n4517), .B(new_n4512), .Y(new_n4518));
  nand_4 g04142(.A(new_n4518), .B(new_n4500), .Y(new_n4519));
  xnor_3 g04143(.A(new_n4517), .B(new_n4511), .Y(new_n4520));
  nand_4 g04144(.A(new_n4520), .B(new_n4499_1), .Y(new_n4521));
  nand_4 g04145(.A(new_n4521), .B(new_n4519), .Y(new_n4522));
  nand_4 g04146(.A(new_n4359), .B(new_n4349), .Y(new_n4523));
  not_3  g04147(.A(new_n4523), .Y(new_n4524));
  nor_4  g04148(.A(new_n4365), .B(new_n4360), .Y(new_n4525));
  nor_4  g04149(.A(new_n4525), .B(new_n4524), .Y(new_n4526));
  xnor_3 g04150(.A(new_n4526), .B(new_n4522), .Y(new_n4527));
  nor_4  g04151(.A(new_n4527), .B(new_n4498), .Y(new_n4528));
  not_3  g04152(.A(new_n4527), .Y(new_n4529));
  nor_4  g04153(.A(new_n4529), .B(new_n4375), .Y(new_n4530));
  nor_4  g04154(.A(new_n4530), .B(new_n4528), .Y(new_n4531));
  not_3  g04155(.A(new_n4344), .Y(new_n4532));
  nand_4 g04156(.A(n12069), .B(n4970), .Y(new_n4533));
  nand_4 g04157(.A(n12391), .B(n7610), .Y(new_n4534));
  not_3  g04158(.A(new_n4534), .Y(new_n4535));
  nor_4  g04159(.A(new_n4340), .B(new_n4334), .Y(new_n4536));
  nor_4  g04160(.A(new_n4536), .B(new_n4339), .Y(new_n4537));
  xnor_3 g04161(.A(new_n4537), .B(new_n4535), .Y(new_n4538));
  nand_4 g04162(.A(n7733), .B(n7160), .Y(new_n4539));
  nand_4 g04163(.A(n7891), .B(n4826), .Y(new_n4540));
  nand_4 g04164(.A(n12925), .B(n4828), .Y(new_n4541));
  xnor_3 g04165(.A(new_n4541), .B(new_n4540), .Y(new_n4542));
  xnor_3 g04166(.A(new_n4542), .B(new_n4539), .Y(new_n4543));
  xnor_3 g04167(.A(new_n4543), .B(new_n4538), .Y(new_n4544));
  xnor_3 g04168(.A(new_n4544), .B(new_n4533), .Y(new_n4545));
  nor_4  g04169(.A(new_n4331), .B(new_n4326_1), .Y(new_n4546));
  nor_4  g04170(.A(new_n4342), .B(new_n4332), .Y(new_n4547));
  nor_4  g04171(.A(new_n4547), .B(new_n4546), .Y(new_n4548));
  xnor_3 g04172(.A(new_n4548), .B(new_n4545), .Y(new_n4549));
  xnor_3 g04173(.A(new_n4549), .B(new_n4532), .Y(new_n4550));
  nor_4  g04174(.A(new_n4378_1), .B(new_n4347), .Y(new_n4551));
  not_3  g04175(.A(new_n4551), .Y(new_n4552));
  nand_4 g04176(.A(new_n4410), .B(new_n4380), .Y(new_n4553_1));
  nand_4 g04177(.A(new_n4553_1), .B(new_n4552), .Y(new_n4554));
  xnor_3 g04178(.A(new_n4554), .B(new_n4550), .Y(new_n4555));
  xnor_3 g04179(.A(new_n4555), .B(new_n4531), .Y(new_n4556));
  not_3  g04180(.A(new_n4556), .Y(new_n4557));
  xnor_3 g04181(.A(new_n4557), .B(new_n4497), .Y(new_n4558));
  nand_4 g04182(.A(new_n4411), .B(new_n4310), .Y(new_n4559));
  not_3  g04183(.A(new_n4412), .Y(new_n4560));
  not_3  g04184(.A(new_n4433), .Y(new_n4561));
  nand_4 g04185(.A(new_n4561), .B(new_n4560), .Y(new_n4562));
  nand_4 g04186(.A(new_n4562), .B(new_n4559), .Y(new_n4563));
  xnor_3 g04187(.A(new_n4563), .B(new_n4558), .Y(new_n4564));
  xor_3  g04188(.A(new_n4564), .B(new_n4468), .Y(n992));
  nand_4 g04189(.A(n7265), .B(n6687), .Y(new_n4566));
  not_3  g04190(.A(new_n4566), .Y(new_n4567));
  nand_4 g04191(.A(n8336), .B(n7946), .Y(new_n4568));
  not_3  g04192(.A(new_n4568), .Y(new_n4569));
  nand_4 g04193(.A(n11222), .B(n9763), .Y(new_n4570));
  nand_4 g04194(.A(n12069), .B(n2558), .Y(new_n4571));
  xor_3  g04195(.A(new_n4571), .B(new_n4570), .Y(new_n4572));
  xor_3  g04196(.A(new_n4572), .B(new_n4569), .Y(new_n4573));
  xor_3  g04197(.A(new_n4573), .B(new_n4567), .Y(n1020));
  not_3  g04198(.A(new_n2193), .Y(new_n4575));
  xnor_3 g04199(.A(new_n4575), .B(new_n2191), .Y(n1136));
  and_4  g04200(.A(new_n4437), .B(new_n4436_1), .Y(new_n4577));
  xor_3  g04201(.A(new_n4577), .B(new_n4465), .Y(n1138));
  nand_4 g04202(.A(n12591), .B(n11757), .Y(new_n4579));
  nand_4 g04203(.A(n5240), .B(n3932), .Y(new_n4580));
  nand_4 g04204(.A(n11821), .B(n1798), .Y(new_n4581));
  xnor_3 g04205(.A(new_n4581), .B(new_n4580), .Y(new_n4582));
  nor_4  g04206(.A(new_n4582), .B(new_n4579), .Y(new_n4583));
  not_3  g04207(.A(new_n4579), .Y(new_n4584));
  not_3  g04208(.A(new_n4582), .Y(new_n4585));
  nor_4  g04209(.A(new_n4585), .B(new_n4584), .Y(new_n4586));
  nor_4  g04210(.A(new_n4586), .B(new_n4583), .Y(new_n4587));
  nand_4 g04211(.A(n5240), .B(n1798), .Y(new_n4588));
  not_3  g04212(.A(new_n4588), .Y(new_n4589));
  nand_4 g04213(.A(n12591), .B(n3172), .Y(new_n4590));
  not_3  g04214(.A(new_n4590), .Y(new_n4591));
  nor_4  g04215(.A(new_n4591), .B(new_n4589), .Y(new_n4592));
  nor_4  g04216(.A(new_n4590), .B(new_n4588), .Y(new_n4593));
  nand_4 g04217(.A(n11757), .B(n3932), .Y(new_n4594));
  not_3  g04218(.A(new_n4594), .Y(new_n4595));
  nor_4  g04219(.A(new_n4595), .B(new_n4593), .Y(new_n4596));
  nor_4  g04220(.A(new_n4596), .B(new_n4592), .Y(new_n4597));
  xnor_3 g04221(.A(new_n4597), .B(new_n4587), .Y(new_n4598));
  nand_4 g04222(.A(n7456), .B(n1333), .Y(new_n4599));
  not_3  g04223(.A(new_n4599), .Y(new_n4600));
  nand_4 g04224(.A(n11757), .B(n1798), .Y(new_n4601));
  not_3  g04225(.A(new_n4601), .Y(new_n4602));
  nand_4 g04226(.A(n12591), .B(n1333), .Y(new_n4603));
  not_3  g04227(.A(new_n4603), .Y(new_n4604));
  nor_4  g04228(.A(new_n4604), .B(new_n4602), .Y(new_n4605));
  nor_4  g04229(.A(new_n4603), .B(new_n4601), .Y(new_n4606));
  nand_4 g04230(.A(n3932), .B(n3172), .Y(new_n4607));
  not_3  g04231(.A(new_n4607), .Y(new_n4608));
  nor_4  g04232(.A(new_n4608), .B(new_n4606), .Y(new_n4609));
  nor_4  g04233(.A(new_n4609), .B(new_n4605), .Y(new_n4610));
  nand_4 g04234(.A(new_n4610), .B(new_n4600), .Y(new_n4611));
  xnor_3 g04235(.A(new_n4610), .B(new_n4599), .Y(new_n4612));
  nor_4  g04236(.A(new_n4593), .B(new_n4592), .Y(new_n4613));
  xnor_3 g04237(.A(new_n4613), .B(new_n4594), .Y(new_n4614));
  nand_4 g04238(.A(new_n4614), .B(new_n4612), .Y(new_n4615));
  nand_4 g04239(.A(new_n4615), .B(new_n4611), .Y(new_n4616));
  nand_4 g04240(.A(n11662), .B(n1333), .Y(new_n4617));
  nand_4 g04241(.A(n7456), .B(n3172), .Y(new_n4618));
  xor_3  g04242(.A(new_n4618), .B(new_n4617), .Y(new_n4619));
  xnor_3 g04243(.A(new_n4619), .B(new_n4616), .Y(new_n4620));
  xnor_3 g04244(.A(new_n4620), .B(new_n4598), .Y(new_n4621));
  nand_4 g04245(.A(n11662), .B(n7862), .Y(new_n4622));
  not_3  g04246(.A(new_n4622), .Y(new_n4623));
  xnor_3 g04247(.A(new_n4614), .B(new_n4612), .Y(new_n4624));
  not_3  g04248(.A(new_n4624), .Y(new_n4625));
  nor_4  g04249(.A(new_n4625), .B(new_n4623), .Y(new_n4626));
  not_3  g04250(.A(new_n4626), .Y(new_n4627));
  nor_4  g04251(.A(new_n4624), .B(new_n4622), .Y(new_n4628));
  nor_4  g04252(.A(new_n4628), .B(new_n4626), .Y(new_n4629));
  nand_4 g04253(.A(n7862), .B(n7456), .Y(new_n4630));
  nand_4 g04254(.A(n3172), .B(n1798), .Y(new_n4631));
  not_3  g04255(.A(new_n4631), .Y(new_n4632));
  nand_4 g04256(.A(n12591), .B(n7862), .Y(new_n4633));
  not_3  g04257(.A(new_n4633), .Y(new_n4634_1));
  nand_4 g04258(.A(new_n4634_1), .B(new_n4632), .Y(new_n4635));
  nand_4 g04259(.A(new_n4633), .B(new_n4631), .Y(new_n4636));
  nand_4 g04260(.A(n3932), .B(n1333), .Y(new_n4637));
  not_3  g04261(.A(new_n4637), .Y(new_n4638));
  nand_4 g04262(.A(new_n4638), .B(new_n4636), .Y(new_n4639));
  nand_4 g04263(.A(new_n4639), .B(new_n4635), .Y(new_n4640));
  not_3  g04264(.A(new_n4640), .Y(new_n4641));
  nor_4  g04265(.A(new_n4641), .B(new_n4630), .Y(new_n4642));
  xnor_3 g04266(.A(new_n4641), .B(new_n4630), .Y(new_n4643));
  nor_4  g04267(.A(new_n4606), .B(new_n4605), .Y(new_n4644));
  xnor_3 g04268(.A(new_n4644), .B(new_n4608), .Y(new_n4645));
  nor_4  g04269(.A(new_n4645), .B(new_n4643), .Y(new_n4646));
  nor_4  g04270(.A(new_n4646), .B(new_n4642), .Y(new_n4647));
  nand_4 g04271(.A(new_n4647), .B(new_n4629), .Y(new_n4648));
  nand_4 g04272(.A(new_n4648), .B(new_n4627), .Y(new_n4649));
  nor_4  g04273(.A(new_n4649), .B(new_n4621), .Y(new_n4650));
  not_3  g04274(.A(new_n4650), .Y(new_n4651));
  not_3  g04275(.A(new_n4587), .Y(new_n4652));
  not_3  g04276(.A(new_n4597), .Y(new_n4653));
  nor_4  g04277(.A(new_n4653), .B(new_n4652), .Y(new_n4654));
  nor_4  g04278(.A(new_n4654), .B(new_n4583), .Y(new_n4655));
  not_3  g04279(.A(new_n4655), .Y(new_n4656));
  nand_4 g04280(.A(n10327), .B(n1333), .Y(new_n4657));
  nand_4 g04281(.A(n11662), .B(n3172), .Y(new_n4658));
  nand_4 g04282(.A(n9583), .B(n7862), .Y(new_n4659));
  not_3  g04283(.A(new_n4659), .Y(new_n4660));
  xor_3  g04284(.A(new_n4660), .B(new_n4658), .Y(new_n4661));
  xnor_3 g04285(.A(new_n4661), .B(new_n4657), .Y(new_n4662));
  xnor_3 g04286(.A(new_n4662), .B(new_n4656), .Y(new_n4663));
  nor_4  g04287(.A(new_n4581), .B(new_n4580), .Y(new_n4664));
  nand_4 g04288(.A(n11757), .B(n7456), .Y(new_n4665));
  not_3  g04289(.A(new_n4665), .Y(new_n4666));
  xor_3  g04290(.A(new_n4666), .B(new_n4664), .Y(new_n4667));
  not_3  g04291(.A(new_n4667), .Y(new_n4668));
  nand_4 g04292(.A(n11821), .B(n3932), .Y(new_n4669));
  nand_4 g04293(.A(n12591), .B(n5240), .Y(new_n4670));
  nand_4 g04294(.A(n9080), .B(n1798), .Y(new_n4671));
  not_3  g04295(.A(new_n4671), .Y(new_n4672));
  xor_3  g04296(.A(new_n4672), .B(new_n4670), .Y(new_n4673));
  xnor_3 g04297(.A(new_n4673), .B(new_n4669), .Y(new_n4674));
  not_3  g04298(.A(new_n4674), .Y(new_n4675));
  xor_3  g04299(.A(new_n4675), .B(new_n4668), .Y(new_n4676));
  xnor_3 g04300(.A(new_n4676), .B(new_n4663), .Y(new_n4677));
  not_3  g04301(.A(new_n4677), .Y(new_n4678));
  nand_4 g04302(.A(new_n4619), .B(new_n4616), .Y(new_n4679));
  nor_4  g04303(.A(new_n4618), .B(new_n4617), .Y(new_n4680));
  nor_4  g04304(.A(new_n4620), .B(new_n4598), .Y(new_n4681));
  xnor_3 g04305(.A(new_n4681), .B(new_n4680), .Y(new_n4682));
  nand_4 g04306(.A(new_n4682), .B(new_n4679), .Y(new_n4683));
  xnor_3 g04307(.A(new_n4683), .B(new_n4678), .Y(new_n4684));
  xnor_3 g04308(.A(new_n4684), .B(new_n4651), .Y(new_n4685));
  nand_4 g04309(.A(n10327), .B(n7862), .Y(new_n4686_1));
  xnor_3 g04310(.A(new_n4649), .B(new_n4621), .Y(new_n4687));
  nor_4  g04311(.A(new_n4687), .B(new_n4686_1), .Y(new_n4688));
  not_3  g04312(.A(new_n4688), .Y(new_n4689_1));
  and_4  g04313(.A(new_n4636), .B(new_n4635), .Y(new_n4690));
  nand_4 g04314(.A(n1798), .B(n1333), .Y(new_n4691));
  nand_4 g04315(.A(n7862), .B(n3932), .Y(new_n4692));
  nor_4  g04316(.A(new_n4692), .B(new_n4691), .Y(new_n4693));
  not_3  g04317(.A(new_n4693), .Y(new_n4694));
  nor_4  g04318(.A(new_n4694), .B(new_n4690), .Y(new_n4695));
  xor_3  g04319(.A(new_n4645), .B(new_n4643), .Y(new_n4696));
  nand_4 g04320(.A(new_n4696), .B(new_n4695), .Y(new_n4697));
  not_3  g04321(.A(new_n4648), .Y(new_n4698));
  nor_4  g04322(.A(new_n4647), .B(new_n4629), .Y(new_n4699));
  nor_4  g04323(.A(new_n4699), .B(new_n4698), .Y(new_n4700));
  nor_4  g04324(.A(new_n4700), .B(new_n4697), .Y(new_n4701));
  not_3  g04325(.A(new_n4686_1), .Y(new_n4702));
  not_3  g04326(.A(new_n4687), .Y(new_n4703));
  nor_4  g04327(.A(new_n4703), .B(new_n4702), .Y(new_n4704));
  nor_4  g04328(.A(new_n4704), .B(new_n4688), .Y(new_n4705));
  nand_4 g04329(.A(new_n4705), .B(new_n4701), .Y(new_n4706));
  nand_4 g04330(.A(new_n4706), .B(new_n4689_1), .Y(new_n4707));
  xnor_3 g04331(.A(new_n4707), .B(new_n4685), .Y(new_n4708));
  nand_4 g04332(.A(n11311), .B(n3022), .Y(new_n4709));
  not_3  g04333(.A(new_n4709), .Y(new_n4710));
  nand_4 g04334(.A(n9640), .B(n4187), .Y(new_n4711));
  nand_4 g04335(.A(n6703), .B(n4203), .Y(new_n4712));
  not_3  g04336(.A(new_n4712), .Y(new_n4713));
  xor_3  g04337(.A(new_n4713), .B(new_n4711), .Y(new_n4714));
  xnor_3 g04338(.A(new_n4714), .B(new_n4710), .Y(new_n4715));
  not_3  g04339(.A(new_n4715), .Y(new_n4716));
  nand_4 g04340(.A(n6703), .B(n4187), .Y(new_n4717));
  not_3  g04341(.A(new_n4717), .Y(new_n4718));
  nand_4 g04342(.A(n3022), .B(n2464), .Y(new_n4719));
  not_3  g04343(.A(new_n4719), .Y(new_n4720));
  nor_4  g04344(.A(new_n4720), .B(new_n4718), .Y(new_n4721));
  nor_4  g04345(.A(new_n4719), .B(new_n4717), .Y(new_n4722_1));
  nand_4 g04346(.A(n11311), .B(n9640), .Y(new_n4723));
  not_3  g04347(.A(new_n4723), .Y(new_n4724));
  nor_4  g04348(.A(new_n4724), .B(new_n4722_1), .Y(new_n4725));
  nor_4  g04349(.A(new_n4725), .B(new_n4721), .Y(new_n4726));
  xor_3  g04350(.A(new_n4726), .B(new_n4716), .Y(new_n4727));
  nand_4 g04351(.A(n10451), .B(n9400), .Y(new_n4728));
  nand_4 g04352(.A(n11023), .B(n2464), .Y(new_n4729));
  xor_3  g04353(.A(new_n4729), .B(new_n4728), .Y(new_n4730));
  xnor_3 g04354(.A(new_n4730), .B(new_n4727), .Y(new_n4731));
  nand_4 g04355(.A(n11023), .B(n9400), .Y(new_n4732));
  not_3  g04356(.A(new_n4732), .Y(new_n4733_1));
  nand_4 g04357(.A(n11311), .B(n6703), .Y(new_n4734));
  not_3  g04358(.A(new_n4734), .Y(new_n4735));
  nand_4 g04359(.A(n9400), .B(n3022), .Y(new_n4736));
  not_3  g04360(.A(new_n4736), .Y(new_n4737));
  nor_4  g04361(.A(new_n4737), .B(new_n4735), .Y(new_n4738));
  nor_4  g04362(.A(new_n4736), .B(new_n4734), .Y(new_n4739));
  nand_4 g04363(.A(n9640), .B(n2464), .Y(new_n4740));
  not_3  g04364(.A(new_n4740), .Y(new_n4741));
  nor_4  g04365(.A(new_n4741), .B(new_n4739), .Y(new_n4742));
  nor_4  g04366(.A(new_n4742), .B(new_n4738), .Y(new_n4743));
  and_4  g04367(.A(new_n4743), .B(new_n4733_1), .Y(new_n4744));
  xnor_3 g04368(.A(new_n4743), .B(new_n4733_1), .Y(new_n4745));
  nor_4  g04369(.A(new_n4722_1), .B(new_n4721), .Y(new_n4746));
  xnor_3 g04370(.A(new_n4746), .B(new_n4724), .Y(new_n4747));
  nor_4  g04371(.A(new_n4747), .B(new_n4745), .Y(new_n4748));
  nor_4  g04372(.A(new_n4748), .B(new_n4744), .Y(new_n4749));
  xnor_3 g04373(.A(new_n4749), .B(new_n4731), .Y(new_n4750));
  nand_4 g04374(.A(n10451), .B(n6877), .Y(new_n4751));
  not_3  g04375(.A(new_n4751), .Y(new_n4752));
  xnor_3 g04376(.A(new_n4747), .B(new_n4745), .Y(new_n4753));
  not_3  g04377(.A(new_n4753), .Y(new_n4754));
  nand_4 g04378(.A(new_n4754), .B(new_n4752), .Y(new_n4755));
  nand_4 g04379(.A(n11023), .B(n6877), .Y(new_n4756));
  not_3  g04380(.A(new_n4756), .Y(new_n4757_1));
  nand_4 g04381(.A(n6703), .B(n2464), .Y(new_n4758));
  not_3  g04382(.A(new_n4758), .Y(new_n4759));
  nand_4 g04383(.A(n6877), .B(n3022), .Y(new_n4760));
  not_3  g04384(.A(new_n4760), .Y(new_n4761));
  nor_4  g04385(.A(new_n4761), .B(new_n4759), .Y(new_n4762));
  nor_4  g04386(.A(new_n4760), .B(new_n4758), .Y(new_n4763));
  nand_4 g04387(.A(n9640), .B(n9400), .Y(new_n4764));
  not_3  g04388(.A(new_n4764), .Y(new_n4765));
  nor_4  g04389(.A(new_n4765), .B(new_n4763), .Y(new_n4766));
  nor_4  g04390(.A(new_n4766), .B(new_n4762), .Y(new_n4767));
  and_4  g04391(.A(new_n4767), .B(new_n4757_1), .Y(new_n4768));
  not_3  g04392(.A(new_n4768), .Y(new_n4769));
  xor_3  g04393(.A(new_n4767), .B(new_n4756), .Y(new_n4770));
  not_3  g04394(.A(new_n4770), .Y(new_n4771));
  nor_4  g04395(.A(new_n4739), .B(new_n4738), .Y(new_n4772));
  xor_3  g04396(.A(new_n4772), .B(new_n4740), .Y(new_n4773));
  not_3  g04397(.A(new_n4773), .Y(new_n4774));
  nand_4 g04398(.A(new_n4774), .B(new_n4771), .Y(new_n4775));
  nand_4 g04399(.A(new_n4775), .B(new_n4769), .Y(new_n4776));
  xor_3  g04400(.A(new_n4754), .B(new_n4752), .Y(new_n4777));
  nand_4 g04401(.A(new_n4777), .B(new_n4776), .Y(new_n4778));
  nand_4 g04402(.A(new_n4778), .B(new_n4755), .Y(new_n4779));
  nand_4 g04403(.A(new_n4779), .B(new_n4750), .Y(new_n4780));
  not_3  g04404(.A(new_n4714), .Y(new_n4781));
  nand_4 g04405(.A(new_n4781), .B(new_n4710), .Y(new_n4782));
  nand_4 g04406(.A(new_n4726), .B(new_n4715), .Y(new_n4783));
  nand_4 g04407(.A(new_n4783), .B(new_n4782), .Y(new_n4784));
  nand_4 g04408(.A(n10278), .B(n9400), .Y(new_n4785));
  not_3  g04409(.A(new_n4785), .Y(new_n4786));
  nand_4 g04410(.A(n10451), .B(n2464), .Y(new_n4787));
  not_3  g04411(.A(new_n4787), .Y(new_n4788));
  nand_4 g04412(.A(n11423), .B(n6877), .Y(new_n4789));
  not_3  g04413(.A(new_n4789), .Y(new_n4790));
  nand_4 g04414(.A(new_n4790), .B(new_n4788), .Y(new_n4791));
  nand_4 g04415(.A(new_n4789), .B(new_n4787), .Y(new_n4792));
  nand_4 g04416(.A(new_n4792), .B(new_n4791), .Y(new_n4793));
  xor_3  g04417(.A(new_n4793), .B(new_n4786), .Y(new_n4794));
  xnor_3 g04418(.A(new_n4794), .B(new_n4784), .Y(new_n4795));
  nor_4  g04419(.A(new_n4712), .B(new_n4711), .Y(new_n4796));
  nand_4 g04420(.A(n11311), .B(n11023), .Y(new_n4797));
  not_3  g04421(.A(new_n4797), .Y(new_n4798));
  xor_3  g04422(.A(new_n4798), .B(new_n4796), .Y(new_n4799));
  nand_4 g04423(.A(n9640), .B(n4203), .Y(new_n4800));
  not_3  g04424(.A(new_n4800), .Y(new_n4801));
  nand_4 g04425(.A(n4187), .B(n3022), .Y(new_n4802));
  not_3  g04426(.A(new_n4802), .Y(new_n4803));
  nand_4 g04427(.A(n12753), .B(n6703), .Y(new_n4804));
  not_3  g04428(.A(new_n4804), .Y(new_n4805_1));
  nor_4  g04429(.A(new_n4805_1), .B(new_n4803), .Y(new_n4806));
  nor_4  g04430(.A(new_n4804), .B(new_n4802), .Y(new_n4807));
  nor_4  g04431(.A(new_n4807), .B(new_n4806), .Y(new_n4808));
  xor_3  g04432(.A(new_n4808), .B(new_n4801), .Y(new_n4809));
  not_3  g04433(.A(new_n4809), .Y(new_n4810));
  xnor_3 g04434(.A(new_n4810), .B(new_n4799), .Y(new_n4811));
  xnor_3 g04435(.A(new_n4811), .B(new_n4795), .Y(new_n4812));
  not_3  g04436(.A(new_n4730), .Y(new_n4813));
  nor_4  g04437(.A(new_n4813), .B(new_n4727), .Y(new_n4814));
  not_3  g04438(.A(new_n4814), .Y(new_n4815));
  nor_4  g04439(.A(new_n4729), .B(new_n4728), .Y(new_n4816));
  not_3  g04440(.A(new_n4816), .Y(new_n4817_1));
  not_3  g04441(.A(new_n4749), .Y(new_n4818));
  nand_4 g04442(.A(new_n4818), .B(new_n4731), .Y(new_n4819));
  xnor_3 g04443(.A(new_n4819), .B(new_n4817_1), .Y(new_n4820));
  nand_4 g04444(.A(new_n4820), .B(new_n4815), .Y(new_n4821));
  not_3  g04445(.A(new_n4821), .Y(new_n4822));
  xnor_3 g04446(.A(new_n4822), .B(new_n4812), .Y(new_n4823));
  xnor_3 g04447(.A(new_n4823), .B(new_n4780), .Y(new_n4824));
  nand_4 g04448(.A(n10278), .B(n6877), .Y(new_n4825));
  xnor_3 g04449(.A(new_n4779), .B(new_n4750), .Y(new_n4826_1));
  nor_4  g04450(.A(new_n4826_1), .B(new_n4825), .Y(new_n4827));
  xnor_3 g04451(.A(new_n4773), .B(new_n4770), .Y(new_n4828_1));
  not_3  g04452(.A(new_n4762), .Y(new_n4829));
  nand_4 g04453(.A(n6877), .B(n6703), .Y(new_n4830));
  not_3  g04454(.A(new_n4830), .Y(new_n4831));
  nor_4  g04455(.A(new_n4831), .B(new_n4764), .Y(new_n4832));
  nor_4  g04456(.A(new_n4832), .B(new_n4829), .Y(new_n4833));
  nor_4  g04457(.A(new_n4833), .B(new_n4763), .Y(new_n4834));
  nor_4  g04458(.A(new_n4834), .B(new_n4764), .Y(new_n4835));
  not_3  g04459(.A(new_n4835), .Y(new_n4836));
  nor_4  g04460(.A(new_n4836), .B(new_n4828_1), .Y(new_n4837));
  not_3  g04461(.A(new_n4837), .Y(new_n4838));
  xnor_3 g04462(.A(new_n4777), .B(new_n4776), .Y(new_n4839));
  nor_4  g04463(.A(new_n4839), .B(new_n4838), .Y(new_n4840));
  not_3  g04464(.A(new_n4840), .Y(new_n4841));
  xnor_3 g04465(.A(new_n4826_1), .B(new_n4825), .Y(new_n4842));
  nor_4  g04466(.A(new_n4842), .B(new_n4841), .Y(new_n4843));
  nor_4  g04467(.A(new_n4843), .B(new_n4827), .Y(new_n4844));
  xnor_3 g04468(.A(new_n4844), .B(new_n4824), .Y(new_n4845));
  nand_4 g04469(.A(n12826), .B(n4805), .Y(new_n4846));
  nand_4 g04470(.A(n8665), .B(n137), .Y(new_n4847));
  nand_4 g04471(.A(n6294), .B(n1067), .Y(new_n4848));
  nand_4 g04472(.A(n6797), .B(n5645), .Y(new_n4849));
  xnor_3 g04473(.A(new_n4849), .B(new_n4848), .Y(new_n4850));
  nor_4  g04474(.A(new_n4850), .B(new_n4847), .Y(new_n4851));
  not_3  g04475(.A(new_n4847), .Y(new_n4852));
  not_3  g04476(.A(new_n4850), .Y(new_n4853));
  nor_4  g04477(.A(new_n4853), .B(new_n4852), .Y(new_n4854));
  nor_4  g04478(.A(new_n4854), .B(new_n4851), .Y(new_n4855));
  nand_4 g04479(.A(n6294), .B(n5645), .Y(new_n4856));
  nand_4 g04480(.A(n8665), .B(n5283), .Y(new_n4857));
  and_4  g04481(.A(new_n4857), .B(new_n4856), .Y(new_n4858));
  nand_4 g04482(.A(n1067), .B(n137), .Y(new_n4859));
  not_3  g04483(.A(new_n4859), .Y(new_n4860));
  xnor_3 g04484(.A(new_n4857), .B(new_n4856), .Y(new_n4861));
  nor_4  g04485(.A(new_n4861), .B(new_n4860), .Y(new_n4862));
  nor_4  g04486(.A(new_n4862), .B(new_n4858), .Y(new_n4863));
  xnor_3 g04487(.A(new_n4863), .B(new_n4855), .Y(new_n4864));
  nand_4 g04488(.A(n11922), .B(n11478), .Y(new_n4865));
  not_3  g04489(.A(new_n4865), .Y(new_n4866));
  nand_4 g04490(.A(n11478), .B(n8665), .Y(new_n4867));
  not_3  g04491(.A(new_n4867), .Y(new_n4868));
  nand_4 g04492(.A(n5283), .B(n1067), .Y(new_n4869));
  not_3  g04493(.A(new_n4869), .Y(new_n4870));
  nor_4  g04494(.A(new_n4870), .B(new_n4868), .Y(new_n4871));
  nor_4  g04495(.A(new_n4869), .B(new_n4867), .Y(new_n4872));
  nand_4 g04496(.A(n5645), .B(n137), .Y(new_n4873));
  not_3  g04497(.A(new_n4873), .Y(new_n4874));
  nor_4  g04498(.A(new_n4874), .B(new_n4872), .Y(new_n4875));
  nor_4  g04499(.A(new_n4875), .B(new_n4871), .Y(new_n4876));
  nand_4 g04500(.A(new_n4876), .B(new_n4866), .Y(new_n4877));
  xnor_3 g04501(.A(new_n4861), .B(new_n4859), .Y(new_n4878));
  not_3  g04502(.A(new_n4878), .Y(new_n4879));
  xnor_3 g04503(.A(new_n4876), .B(new_n4865), .Y(new_n4880));
  nand_4 g04504(.A(new_n4880), .B(new_n4879), .Y(new_n4881));
  nand_4 g04505(.A(new_n4881), .B(new_n4877), .Y(new_n4882));
  nand_4 g04506(.A(n11478), .B(n2551), .Y(new_n4883));
  nand_4 g04507(.A(n11922), .B(n5283), .Y(new_n4884));
  xor_3  g04508(.A(new_n4884), .B(new_n4883), .Y(new_n4885));
  xnor_3 g04509(.A(new_n4885), .B(new_n4882), .Y(new_n4886));
  xnor_3 g04510(.A(new_n4886), .B(new_n4864), .Y(new_n4887));
  nand_4 g04511(.A(n4805), .B(n2551), .Y(new_n4888));
  not_3  g04512(.A(new_n4888), .Y(new_n4889));
  nand_4 g04513(.A(n11922), .B(n4805), .Y(new_n4890));
  not_3  g04514(.A(new_n4890), .Y(new_n4891));
  nand_4 g04515(.A(n5645), .B(n5283), .Y(new_n4892));
  not_3  g04516(.A(new_n4892), .Y(new_n4893));
  nand_4 g04517(.A(n8665), .B(n4805), .Y(new_n4894));
  not_3  g04518(.A(new_n4894), .Y(new_n4895));
  nand_4 g04519(.A(new_n4895), .B(new_n4893), .Y(new_n4896));
  nand_4 g04520(.A(n11478), .B(n1067), .Y(new_n4897));
  not_3  g04521(.A(new_n4897), .Y(new_n4898));
  nand_4 g04522(.A(new_n4894), .B(new_n4892), .Y(new_n4899));
  nand_4 g04523(.A(new_n4899), .B(new_n4898), .Y(new_n4900));
  nand_4 g04524(.A(new_n4900), .B(new_n4896), .Y(new_n4901));
  nand_4 g04525(.A(new_n4901), .B(new_n4891), .Y(new_n4902));
  not_3  g04526(.A(new_n4902), .Y(new_n4903_1));
  nor_4  g04527(.A(new_n4901), .B(new_n4891), .Y(new_n4904));
  nor_4  g04528(.A(new_n4904), .B(new_n4903_1), .Y(new_n4905));
  xnor_3 g04529(.A(new_n4869), .B(new_n4867), .Y(new_n4906));
  xnor_3 g04530(.A(new_n4906), .B(new_n4873), .Y(new_n4907));
  not_3  g04531(.A(new_n4907), .Y(new_n4908));
  nand_4 g04532(.A(new_n4908), .B(new_n4905), .Y(new_n4909));
  nand_4 g04533(.A(new_n4909), .B(new_n4902), .Y(new_n4910));
  nor_4  g04534(.A(new_n4910), .B(new_n4889), .Y(new_n4911));
  xnor_3 g04535(.A(new_n4880), .B(new_n4878), .Y(new_n4912));
  xnor_3 g04536(.A(new_n4910), .B(new_n4889), .Y(new_n4913));
  nor_4  g04537(.A(new_n4913), .B(new_n4912), .Y(new_n4914));
  nor_4  g04538(.A(new_n4914), .B(new_n4911), .Y(new_n4915));
  not_3  g04539(.A(new_n4915), .Y(new_n4916));
  xnor_3 g04540(.A(new_n4916), .B(new_n4887), .Y(new_n4917));
  nor_4  g04541(.A(new_n4917), .B(new_n4846), .Y(new_n4918));
  nand_4 g04542(.A(new_n4899), .B(new_n4896), .Y(new_n4919));
  nand_4 g04543(.A(n4805), .B(n1067), .Y(new_n4920));
  nand_4 g04544(.A(n11478), .B(n5645), .Y(new_n4921_1));
  nor_4  g04545(.A(new_n4921_1), .B(new_n4920), .Y(new_n4922));
  nand_4 g04546(.A(new_n4922), .B(new_n4919), .Y(new_n4923));
  xnor_3 g04547(.A(new_n4908), .B(new_n4905), .Y(new_n4924));
  nor_4  g04548(.A(new_n4924), .B(new_n4923), .Y(new_n4925));
  not_3  g04549(.A(new_n4925), .Y(new_n4926));
  not_3  g04550(.A(new_n4912), .Y(new_n4927));
  xnor_3 g04551(.A(new_n4913), .B(new_n4927), .Y(new_n4928_1));
  nor_4  g04552(.A(new_n4928_1), .B(new_n4926), .Y(new_n4929));
  not_3  g04553(.A(new_n4929), .Y(new_n4930));
  xnor_3 g04554(.A(new_n4917), .B(new_n4846), .Y(new_n4931));
  nor_4  g04555(.A(new_n4931), .B(new_n4930), .Y(new_n4932));
  nor_4  g04556(.A(new_n4932), .B(new_n4918), .Y(new_n4933));
  nor_4  g04557(.A(new_n4916), .B(new_n4887), .Y(new_n4934));
  not_3  g04558(.A(new_n4851), .Y(new_n4935));
  nand_4 g04559(.A(new_n4863), .B(new_n4855), .Y(new_n4936));
  nand_4 g04560(.A(new_n4936), .B(new_n4935), .Y(new_n4937));
  nand_4 g04561(.A(n12826), .B(n11478), .Y(new_n4938_1));
  not_3  g04562(.A(new_n4938_1), .Y(new_n4939));
  nand_4 g04563(.A(n5283), .B(n2551), .Y(new_n4940));
  nand_4 g04564(.A(n4805), .B(n4094), .Y(new_n4941));
  nand_4 g04565(.A(new_n4941), .B(new_n4940), .Y(new_n4942));
  not_3  g04566(.A(new_n4940), .Y(new_n4943));
  not_3  g04567(.A(new_n4941), .Y(new_n4944));
  nand_4 g04568(.A(new_n4944), .B(new_n4943), .Y(new_n4945));
  nand_4 g04569(.A(new_n4945), .B(new_n4942), .Y(new_n4946));
  xor_3  g04570(.A(new_n4946), .B(new_n4939), .Y(new_n4947));
  xnor_3 g04571(.A(new_n4947), .B(new_n4937), .Y(new_n4948));
  nor_4  g04572(.A(new_n4849), .B(new_n4848), .Y(new_n4949));
  nand_4 g04573(.A(n11922), .B(n137), .Y(new_n4950));
  not_3  g04574(.A(new_n4950), .Y(new_n4951));
  xor_3  g04575(.A(new_n4951), .B(new_n4949), .Y(new_n4952));
  not_3  g04576(.A(new_n4952), .Y(new_n4953));
  nand_4 g04577(.A(n6797), .B(n1067), .Y(new_n4954));
  not_3  g04578(.A(new_n4954), .Y(new_n4955));
  nand_4 g04579(.A(n8665), .B(n6294), .Y(new_n4956));
  nand_4 g04580(.A(n5645), .B(n3146), .Y(new_n4957));
  not_3  g04581(.A(new_n4957), .Y(new_n4958));
  xor_3  g04582(.A(new_n4958), .B(new_n4956), .Y(new_n4959));
  xnor_3 g04583(.A(new_n4959), .B(new_n4955), .Y(new_n4960));
  xnor_3 g04584(.A(new_n4960), .B(new_n4953), .Y(new_n4961));
  xnor_3 g04585(.A(new_n4961), .B(new_n4948), .Y(new_n4962));
  nand_4 g04586(.A(new_n4885), .B(new_n4882), .Y(new_n4963));
  nor_4  g04587(.A(new_n4884), .B(new_n4883), .Y(new_n4964));
  nor_4  g04588(.A(new_n4886), .B(new_n4864), .Y(new_n4965));
  xnor_3 g04589(.A(new_n4965), .B(new_n4964), .Y(new_n4966));
  nand_4 g04590(.A(new_n4966), .B(new_n4963), .Y(new_n4967));
  xnor_3 g04591(.A(new_n4967), .B(new_n4962), .Y(new_n4968));
  xnor_3 g04592(.A(new_n4968), .B(new_n4934), .Y(new_n4969));
  xnor_3 g04593(.A(new_n4969), .B(new_n4933), .Y(new_n4970_1));
  nand_4 g04594(.A(n3992), .B(n2749), .Y(new_n4971_1));
  not_3  g04595(.A(new_n4971_1), .Y(new_n4972));
  nand_4 g04596(.A(n11876), .B(n6358), .Y(new_n4973));
  not_3  g04597(.A(new_n4973), .Y(new_n4974));
  nand_4 g04598(.A(n3992), .B(n3754), .Y(new_n4975));
  not_3  g04599(.A(new_n4975), .Y(new_n4976));
  nor_4  g04600(.A(new_n4976), .B(new_n4974), .Y(new_n4977));
  nor_4  g04601(.A(new_n4975), .B(new_n4973), .Y(new_n4978));
  nand_4 g04602(.A(n10898), .B(n8384), .Y(new_n4979));
  not_3  g04603(.A(new_n4979), .Y(new_n4980));
  nor_4  g04604(.A(new_n4980), .B(new_n4978), .Y(new_n4981));
  nor_4  g04605(.A(new_n4981), .B(new_n4977), .Y(new_n4982));
  nand_4 g04606(.A(new_n4982), .B(new_n4972), .Y(new_n4983));
  xnor_3 g04607(.A(new_n4982), .B(new_n4971_1), .Y(new_n4984));
  nand_4 g04608(.A(n10898), .B(n6358), .Y(new_n4985));
  not_3  g04609(.A(new_n4985), .Y(new_n4986));
  nand_4 g04610(.A(n8384), .B(n3754), .Y(new_n4987));
  nand_4 g04611(.A(n11876), .B(n5198), .Y(new_n4988));
  xnor_3 g04612(.A(new_n4988), .B(new_n4987), .Y(new_n4989));
  xnor_3 g04613(.A(new_n4989), .B(new_n4986), .Y(new_n4990));
  nand_4 g04614(.A(new_n4990), .B(new_n4984), .Y(new_n4991));
  nand_4 g04615(.A(new_n4991), .B(new_n4983), .Y(new_n4992));
  nand_4 g04616(.A(n8384), .B(n2749), .Y(new_n4993));
  nand_4 g04617(.A(n3992), .B(n159), .Y(new_n4994));
  xor_3  g04618(.A(new_n4994), .B(new_n4993), .Y(new_n4995));
  xnor_3 g04619(.A(new_n4995), .B(new_n4992), .Y(new_n4996));
  nand_4 g04620(.A(n6358), .B(n3754), .Y(new_n4997));
  not_3  g04621(.A(new_n4997), .Y(new_n4998));
  nand_4 g04622(.A(n10898), .B(n5198), .Y(new_n4999));
  nand_4 g04623(.A(n11876), .B(n1471), .Y(new_n5000));
  xnor_3 g04624(.A(new_n5000), .B(new_n4999), .Y(new_n5001));
  not_3  g04625(.A(new_n5001), .Y(new_n5002));
  nor_4  g04626(.A(new_n5002), .B(new_n4998), .Y(new_n5003));
  nor_4  g04627(.A(new_n5001), .B(new_n4997), .Y(new_n5004));
  nor_4  g04628(.A(new_n5004), .B(new_n5003), .Y(new_n5005));
  not_3  g04629(.A(new_n5005), .Y(new_n5006));
  and_4  g04630(.A(new_n4988), .B(new_n4987), .Y(new_n5007));
  nor_4  g04631(.A(new_n4989), .B(new_n4986), .Y(new_n5008));
  nor_4  g04632(.A(new_n5008), .B(new_n5007), .Y(new_n5009));
  nor_4  g04633(.A(new_n5009), .B(new_n5006), .Y(new_n5010));
  not_3  g04634(.A(new_n5009), .Y(new_n5011));
  nor_4  g04635(.A(new_n5011), .B(new_n5005), .Y(new_n5012));
  nor_4  g04636(.A(new_n5012), .B(new_n5010), .Y(new_n5013));
  xnor_3 g04637(.A(new_n5013), .B(new_n4996), .Y(new_n5014));
  nand_4 g04638(.A(n7236), .B(n159), .Y(new_n5015));
  not_3  g04639(.A(new_n5015), .Y(new_n5016));
  nand_4 g04640(.A(n7236), .B(n2749), .Y(new_n5017));
  not_3  g04641(.A(new_n5017), .Y(new_n5018));
  nand_4 g04642(.A(n11876), .B(n8384), .Y(new_n5019));
  not_3  g04643(.A(new_n5019), .Y(new_n5020));
  nand_4 g04644(.A(n7236), .B(n3754), .Y(new_n5021));
  not_3  g04645(.A(new_n5021), .Y(new_n5022));
  nor_4  g04646(.A(new_n5022), .B(new_n5020), .Y(new_n5023));
  nand_4 g04647(.A(n11876), .B(n7236), .Y(new_n5024));
  nor_4  g04648(.A(new_n5024), .B(new_n4987), .Y(new_n5025));
  nand_4 g04649(.A(n10898), .B(n3992), .Y(new_n5026));
  not_3  g04650(.A(new_n5026), .Y(new_n5027));
  nor_4  g04651(.A(new_n5027), .B(new_n5025), .Y(new_n5028));
  nor_4  g04652(.A(new_n5028), .B(new_n5023), .Y(new_n5029));
  nand_4 g04653(.A(new_n5029), .B(new_n5018), .Y(new_n5030_1));
  not_3  g04654(.A(new_n5030_1), .Y(new_n5031));
  nor_4  g04655(.A(new_n5029), .B(new_n5018), .Y(new_n5032));
  nor_4  g04656(.A(new_n5032), .B(new_n5031), .Y(new_n5033));
  xnor_3 g04657(.A(new_n4975), .B(new_n4973), .Y(new_n5034_1));
  xnor_3 g04658(.A(new_n5034_1), .B(new_n4979), .Y(new_n5035));
  not_3  g04659(.A(new_n5035), .Y(new_n5036));
  nand_4 g04660(.A(new_n5036), .B(new_n5033), .Y(new_n5037));
  nand_4 g04661(.A(new_n5037), .B(new_n5030_1), .Y(new_n5038));
  nor_4  g04662(.A(new_n5038), .B(new_n5016), .Y(new_n5039));
  not_3  g04663(.A(new_n5039), .Y(new_n5040));
  xnor_3 g04664(.A(new_n4990), .B(new_n4984), .Y(new_n5041));
  not_3  g04665(.A(new_n5038), .Y(new_n5042));
  nor_4  g04666(.A(new_n5042), .B(new_n5015), .Y(new_n5043));
  nor_4  g04667(.A(new_n5043), .B(new_n5039), .Y(new_n5044));
  nand_4 g04668(.A(new_n5044), .B(new_n5041), .Y(new_n5045));
  nand_4 g04669(.A(new_n5045), .B(new_n5040), .Y(new_n5046));
  nor_4  g04670(.A(new_n5046), .B(new_n5014), .Y(new_n5047));
  not_3  g04671(.A(new_n5047), .Y(new_n5048));
  nor_4  g04672(.A(new_n5000), .B(new_n4999), .Y(new_n5049));
  not_3  g04673(.A(new_n5049), .Y(new_n5050));
  nand_4 g04674(.A(n6358), .B(n2749), .Y(new_n5051));
  xor_3  g04675(.A(new_n5051), .B(new_n5050), .Y(new_n5052));
  nand_4 g04676(.A(n10898), .B(n1471), .Y(new_n5053));
  nand_4 g04677(.A(n5198), .B(n3754), .Y(new_n5054));
  nand_4 g04678(.A(n11876), .B(n7646), .Y(new_n5055));
  not_3  g04679(.A(new_n5055), .Y(new_n5056));
  xor_3  g04680(.A(new_n5056), .B(new_n5054), .Y(new_n5057));
  xnor_3 g04681(.A(new_n5057), .B(new_n5053), .Y(new_n5058));
  xnor_3 g04682(.A(new_n5058), .B(new_n5052), .Y(new_n5059));
  nor_4  g04683(.A(new_n5010), .B(new_n5003), .Y(new_n5060));
  nand_4 g04684(.A(n3992), .B(n1510), .Y(new_n5061));
  nand_4 g04685(.A(n8384), .B(n159), .Y(new_n5062));
  nand_4 g04686(.A(n12247), .B(n7236), .Y(new_n5063));
  not_3  g04687(.A(new_n5063), .Y(new_n5064));
  xor_3  g04688(.A(new_n5064), .B(new_n5062), .Y(new_n5065));
  xnor_3 g04689(.A(new_n5065), .B(new_n5061), .Y(new_n5066));
  xnor_3 g04690(.A(new_n5066), .B(new_n5060), .Y(new_n5067));
  xnor_3 g04691(.A(new_n5067), .B(new_n5059), .Y(new_n5068));
  nand_4 g04692(.A(new_n4995), .B(new_n4992), .Y(new_n5069_1));
  nor_4  g04693(.A(new_n4994), .B(new_n4993), .Y(new_n5070));
  nor_4  g04694(.A(new_n5013), .B(new_n4996), .Y(new_n5071));
  xnor_3 g04695(.A(new_n5071), .B(new_n5070), .Y(new_n5072));
  nand_4 g04696(.A(new_n5072), .B(new_n5069_1), .Y(new_n5073));
  xnor_3 g04697(.A(new_n5073), .B(new_n5068), .Y(new_n5074));
  xnor_3 g04698(.A(new_n5074), .B(new_n5048), .Y(new_n5075));
  nand_4 g04699(.A(n7236), .B(n1510), .Y(new_n5076));
  not_3  g04700(.A(new_n5076), .Y(new_n5077));
  not_3  g04701(.A(new_n5046), .Y(new_n5078));
  xnor_3 g04702(.A(new_n5078), .B(new_n5014), .Y(new_n5079));
  nand_4 g04703(.A(new_n5079), .B(new_n5077), .Y(new_n5080));
  nor_4  g04704(.A(new_n5025), .B(new_n5023), .Y(new_n5081));
  nand_4 g04705(.A(n11876), .B(n3992), .Y(new_n5082));
  nand_4 g04706(.A(n10898), .B(n7236), .Y(new_n5083));
  nor_4  g04707(.A(new_n5083), .B(new_n5082), .Y(new_n5084));
  not_3  g04708(.A(new_n5084), .Y(new_n5085));
  nor_4  g04709(.A(new_n5085), .B(new_n5081), .Y(new_n5086));
  not_3  g04710(.A(new_n5086), .Y(new_n5087));
  xnor_3 g04711(.A(new_n5036), .B(new_n5033), .Y(new_n5088));
  nor_4  g04712(.A(new_n5088), .B(new_n5087), .Y(new_n5089));
  xnor_3 g04713(.A(new_n5044), .B(new_n5041), .Y(new_n5090));
  nand_4 g04714(.A(new_n5090), .B(new_n5089), .Y(new_n5091));
  not_3  g04715(.A(new_n5091), .Y(new_n5092));
  xnor_3 g04716(.A(new_n5079), .B(new_n5076), .Y(new_n5093));
  nand_4 g04717(.A(new_n5093), .B(new_n5092), .Y(new_n5094_1));
  nand_4 g04718(.A(new_n5094_1), .B(new_n5080), .Y(new_n5095));
  xnor_3 g04719(.A(new_n5095), .B(new_n5075), .Y(new_n5096));
  xnor_3 g04720(.A(new_n5096), .B(new_n4970_1), .Y(new_n5097));
  not_3  g04721(.A(new_n4846), .Y(new_n5098));
  xnor_3 g04722(.A(new_n4917), .B(new_n5098), .Y(new_n5099));
  nor_4  g04723(.A(new_n5099), .B(new_n4929), .Y(new_n5100));
  nor_4  g04724(.A(new_n5100), .B(new_n4932), .Y(new_n5101));
  not_3  g04725(.A(new_n5101), .Y(new_n5102));
  xnor_3 g04726(.A(new_n5093), .B(new_n5092), .Y(new_n5103));
  nand_4 g04727(.A(new_n5103), .B(new_n5102), .Y(new_n5104));
  xnor_3 g04728(.A(new_n5103), .B(new_n5101), .Y(new_n5105_1));
  nor_4  g04729(.A(new_n5090), .B(new_n5089), .Y(new_n5106));
  nor_4  g04730(.A(new_n5106), .B(new_n5092), .Y(new_n5107));
  not_3  g04731(.A(new_n4923), .Y(new_n5108));
  not_3  g04732(.A(new_n4924), .Y(new_n5109));
  nor_4  g04733(.A(new_n5109), .B(new_n5108), .Y(new_n5110));
  nor_4  g04734(.A(new_n5110), .B(new_n4925), .Y(new_n5111));
  not_3  g04735(.A(new_n5088), .Y(new_n5112));
  nor_4  g04736(.A(new_n5112), .B(new_n5086), .Y(new_n5113));
  nor_4  g04737(.A(new_n5113), .B(new_n5089), .Y(new_n5114));
  nor_4  g04738(.A(new_n5114), .B(new_n5111), .Y(new_n5115));
  not_3  g04739(.A(new_n5115), .Y(new_n5116));
  xnor_3 g04740(.A(new_n5083), .B(new_n5082), .Y(new_n5117));
  xnor_3 g04741(.A(new_n4921_1), .B(new_n4920), .Y(new_n5118));
  nand_4 g04742(.A(new_n5118), .B(new_n5117), .Y(new_n5119));
  not_3  g04743(.A(new_n5119), .Y(new_n5120));
  nand_4 g04744(.A(n5645), .B(n4805), .Y(new_n5121));
  nor_4  g04745(.A(new_n5121), .B(new_n5024), .Y(new_n5122));
  xnor_3 g04746(.A(new_n5118), .B(new_n5117), .Y(new_n5123));
  nor_4  g04747(.A(new_n5123), .B(new_n5122), .Y(new_n5124));
  nor_4  g04748(.A(new_n5124), .B(new_n5120), .Y(new_n5125));
  not_3  g04749(.A(new_n5121), .Y(new_n5126));
  nor_4  g04750(.A(new_n5126), .B(new_n4897), .Y(new_n5127));
  not_3  g04751(.A(new_n5127), .Y(new_n5128));
  nand_4 g04752(.A(new_n5128), .B(new_n4919), .Y(new_n5129));
  nand_4 g04753(.A(new_n5127), .B(new_n4899), .Y(new_n5130));
  nand_4 g04754(.A(new_n5130), .B(new_n5129), .Y(new_n5131));
  not_3  g04755(.A(new_n5131), .Y(new_n5132_1));
  nor_4  g04756(.A(new_n5132_1), .B(new_n5125), .Y(new_n5133));
  xnor_3 g04757(.A(new_n5132_1), .B(new_n5125), .Y(new_n5134));
  not_3  g04758(.A(new_n5024), .Y(new_n5135));
  nor_4  g04759(.A(new_n5026), .B(new_n5135), .Y(new_n5136));
  nor_4  g04760(.A(new_n5136), .B(new_n5081), .Y(new_n5137));
  not_3  g04761(.A(new_n5136), .Y(new_n5138));
  nor_4  g04762(.A(new_n5138), .B(new_n5023), .Y(new_n5139));
  nor_4  g04763(.A(new_n5139), .B(new_n5137), .Y(new_n5140));
  nor_4  g04764(.A(new_n5140), .B(new_n5134), .Y(new_n5141));
  nor_4  g04765(.A(new_n5141), .B(new_n5133), .Y(new_n5142));
  xnor_3 g04766(.A(new_n5114), .B(new_n5111), .Y(new_n5143));
  nor_4  g04767(.A(new_n5143), .B(new_n5142), .Y(new_n5144));
  not_3  g04768(.A(new_n5144), .Y(new_n5145));
  nand_4 g04769(.A(new_n5145), .B(new_n5116), .Y(new_n5146));
  not_3  g04770(.A(new_n5146), .Y(new_n5147));
  nor_4  g04771(.A(new_n5147), .B(new_n5107), .Y(new_n5148));
  not_3  g04772(.A(new_n5148), .Y(new_n5149));
  not_3  g04773(.A(new_n4928_1), .Y(new_n5150));
  xor_3  g04774(.A(new_n5150), .B(new_n4926), .Y(new_n5151));
  xnor_3 g04775(.A(new_n5146), .B(new_n5107), .Y(new_n5152));
  nand_4 g04776(.A(new_n5152), .B(new_n5151), .Y(new_n5153_1));
  nand_4 g04777(.A(new_n5153_1), .B(new_n5149), .Y(new_n5154));
  nand_4 g04778(.A(new_n5154), .B(new_n5105_1), .Y(new_n5155));
  nand_4 g04779(.A(new_n5155), .B(new_n5104), .Y(new_n5156));
  xnor_3 g04780(.A(new_n5156), .B(new_n5097), .Y(new_n5157));
  nand_4 g04781(.A(new_n5157), .B(new_n4845), .Y(new_n5158));
  not_3  g04782(.A(new_n4824), .Y(new_n5159));
  xnor_3 g04783(.A(new_n4844), .B(new_n5159), .Y(new_n5160));
  not_3  g04784(.A(new_n4918), .Y(new_n5161));
  nand_4 g04785(.A(new_n5099), .B(new_n4929), .Y(new_n5162));
  nand_4 g04786(.A(new_n5162), .B(new_n5161), .Y(new_n5163));
  xnor_3 g04787(.A(new_n4969), .B(new_n5163), .Y(new_n5164));
  xnor_3 g04788(.A(new_n5096), .B(new_n5164), .Y(new_n5165));
  xnor_3 g04789(.A(new_n5156), .B(new_n5165), .Y(new_n5166));
  nand_4 g04790(.A(new_n5166), .B(new_n5160), .Y(new_n5167));
  nand_4 g04791(.A(new_n5167), .B(new_n5158), .Y(new_n5168));
  xnor_3 g04792(.A(new_n4842), .B(new_n4840), .Y(new_n5169));
  xnor_3 g04793(.A(new_n5154), .B(new_n5105_1), .Y(new_n5170));
  nand_4 g04794(.A(new_n5170), .B(new_n5169), .Y(new_n5171));
  xnor_3 g04795(.A(new_n4842), .B(new_n4841), .Y(new_n5172));
  xor_3  g04796(.A(new_n5150), .B(new_n4925), .Y(new_n5173));
  not_3  g04797(.A(new_n5152), .Y(new_n5174));
  nor_4  g04798(.A(new_n5174), .B(new_n5173), .Y(new_n5175));
  nor_4  g04799(.A(new_n5175), .B(new_n5148), .Y(new_n5176));
  xnor_3 g04800(.A(new_n5176), .B(new_n5105_1), .Y(new_n5177));
  nand_4 g04801(.A(new_n5177), .B(new_n5172), .Y(new_n5178));
  not_3  g04802(.A(new_n4839), .Y(new_n5179));
  nor_4  g04803(.A(new_n5179), .B(new_n4837), .Y(new_n5180));
  nor_4  g04804(.A(new_n5180), .B(new_n4840), .Y(new_n5181));
  not_3  g04805(.A(new_n4828_1), .Y(new_n5182));
  xor_3  g04806(.A(new_n4835), .B(new_n5182), .Y(new_n5183));
  xnor_3 g04807(.A(new_n5143), .B(new_n5142), .Y(new_n5184));
  nand_4 g04808(.A(new_n5184), .B(new_n5183), .Y(new_n5185));
  not_3  g04809(.A(new_n5184), .Y(new_n5186));
  xnor_3 g04810(.A(new_n5186), .B(new_n5183), .Y(new_n5187));
  xnor_3 g04811(.A(new_n5140), .B(new_n5134), .Y(new_n5188));
  not_3  g04812(.A(new_n4834), .Y(new_n5189));
  not_3  g04813(.A(new_n4832), .Y(new_n5190));
  nor_4  g04814(.A(new_n5190), .B(new_n4762), .Y(new_n5191_1));
  nor_4  g04815(.A(new_n5191_1), .B(new_n5189), .Y(new_n5192));
  nand_4 g04816(.A(new_n5192), .B(new_n5188), .Y(new_n5193));
  not_3  g04817(.A(new_n5193), .Y(new_n5194));
  nor_4  g04818(.A(new_n5192), .B(new_n5188), .Y(new_n5195));
  nor_4  g04819(.A(new_n5195), .B(new_n5194), .Y(new_n5196));
  not_3  g04820(.A(new_n5123), .Y(new_n5197));
  xor_3  g04821(.A(new_n5197), .B(new_n5122), .Y(new_n5198_1));
  nand_4 g04822(.A(n9400), .B(n6703), .Y(new_n5199));
  nand_4 g04823(.A(n9640), .B(n6877), .Y(new_n5200));
  xor_3  g04824(.A(new_n5200), .B(new_n5199), .Y(new_n5201));
  nand_4 g04825(.A(new_n5201), .B(new_n5198_1), .Y(new_n5202));
  xor_3  g04826(.A(new_n5126), .B(new_n5024), .Y(new_n5203));
  nor_4  g04827(.A(new_n5203), .B(new_n4830), .Y(new_n5204));
  not_3  g04828(.A(new_n5202), .Y(new_n5205));
  nor_4  g04829(.A(new_n5201), .B(new_n5198_1), .Y(new_n5206));
  nor_4  g04830(.A(new_n5206), .B(new_n5205), .Y(new_n5207));
  nand_4 g04831(.A(new_n5207), .B(new_n5204), .Y(new_n5208));
  nand_4 g04832(.A(new_n5208), .B(new_n5202), .Y(new_n5209));
  nand_4 g04833(.A(new_n5209), .B(new_n5196), .Y(new_n5210));
  nand_4 g04834(.A(new_n5210), .B(new_n5193), .Y(new_n5211));
  nand_4 g04835(.A(new_n5211), .B(new_n5187), .Y(new_n5212_1));
  nand_4 g04836(.A(new_n5212_1), .B(new_n5185), .Y(new_n5213));
  nor_4  g04837(.A(new_n5213), .B(new_n5181), .Y(new_n5214));
  xnor_3 g04838(.A(new_n5174), .B(new_n5173), .Y(new_n5215));
  xnor_3 g04839(.A(new_n5213), .B(new_n5181), .Y(new_n5216));
  nor_4  g04840(.A(new_n5216), .B(new_n5215), .Y(new_n5217));
  nor_4  g04841(.A(new_n5217), .B(new_n5214), .Y(new_n5218));
  nand_4 g04842(.A(new_n5218), .B(new_n5178), .Y(new_n5219));
  nand_4 g04843(.A(new_n5219), .B(new_n5171), .Y(new_n5220));
  xnor_3 g04844(.A(new_n5220), .B(new_n5168), .Y(new_n5221));
  not_3  g04845(.A(new_n5221), .Y(new_n5222));
  nand_4 g04846(.A(new_n5222), .B(new_n4708), .Y(new_n5223));
  not_3  g04847(.A(new_n4708), .Y(new_n5224));
  nand_4 g04848(.A(new_n5221), .B(new_n5224), .Y(new_n5225));
  xor_3  g04849(.A(new_n4705), .B(new_n4701), .Y(new_n5226));
  not_3  g04850(.A(new_n5226), .Y(new_n5227));
  nand_4 g04851(.A(new_n5178), .B(new_n5171), .Y(new_n5228));
  xnor_3 g04852(.A(new_n5228), .B(new_n5218), .Y(new_n5229));
  not_3  g04853(.A(new_n5229), .Y(new_n5230));
  nand_4 g04854(.A(new_n5230), .B(new_n5227), .Y(new_n5231));
  nand_4 g04855(.A(new_n5229), .B(new_n5226), .Y(new_n5232));
  not_3  g04856(.A(new_n4697), .Y(new_n5233));
  xor_3  g04857(.A(new_n4700), .B(new_n5233), .Y(new_n5234));
  not_3  g04858(.A(new_n5215), .Y(new_n5235));
  xnor_3 g04859(.A(new_n5216), .B(new_n5235), .Y(new_n5236));
  nand_4 g04860(.A(new_n5236), .B(new_n5234), .Y(new_n5237));
  not_3  g04861(.A(new_n5237), .Y(new_n5238));
  nor_4  g04862(.A(new_n5236), .B(new_n5234), .Y(new_n5239));
  nor_4  g04863(.A(new_n5239), .B(new_n5238), .Y(new_n5240_1));
  not_3  g04864(.A(new_n4696), .Y(new_n5241));
  xor_3  g04865(.A(new_n5241), .B(new_n4695), .Y(new_n5242));
  not_3  g04866(.A(new_n5242), .Y(new_n5243));
  xnor_3 g04867(.A(new_n5211), .B(new_n5187), .Y(new_n5244));
  not_3  g04868(.A(new_n5244), .Y(new_n5245));
  nor_4  g04869(.A(new_n5245), .B(new_n5243), .Y(new_n5246));
  not_3  g04870(.A(new_n5246), .Y(new_n5247));
  xnor_3 g04871(.A(new_n5209), .B(new_n5196), .Y(new_n5248));
  not_3  g04872(.A(new_n4690), .Y(new_n5249));
  nand_4 g04873(.A(n7862), .B(n1798), .Y(new_n5250));
  not_3  g04874(.A(new_n5250), .Y(new_n5251));
  nor_4  g04875(.A(new_n5251), .B(new_n4637), .Y(new_n5252));
  not_3  g04876(.A(new_n5252), .Y(new_n5253));
  nand_4 g04877(.A(new_n5253), .B(new_n5249), .Y(new_n5254));
  nand_4 g04878(.A(new_n5252), .B(new_n4636), .Y(new_n5255));
  nand_4 g04879(.A(new_n5255), .B(new_n5254), .Y(new_n5256));
  nand_4 g04880(.A(new_n5256), .B(new_n5248), .Y(new_n5257_1));
  not_3  g04881(.A(new_n5257_1), .Y(new_n5258));
  nor_4  g04882(.A(new_n5256), .B(new_n5248), .Y(new_n5259));
  nor_4  g04883(.A(new_n5259), .B(new_n5258), .Y(new_n5260));
  xor_3  g04884(.A(new_n5203), .B(new_n4830), .Y(new_n5261));
  nand_4 g04885(.A(new_n5261), .B(new_n5251), .Y(new_n5262));
  not_3  g04886(.A(new_n5262), .Y(new_n5263));
  xor_3  g04887(.A(new_n4692), .B(new_n4691), .Y(new_n5264));
  or_4   g04888(.A(new_n5264), .B(new_n5263), .Y(new_n5265));
  xnor_3 g04889(.A(new_n5207), .B(new_n5204), .Y(new_n5266));
  xor_3  g04890(.A(new_n5264), .B(new_n5263), .Y(new_n5267));
  nand_4 g04891(.A(new_n5267), .B(new_n5266), .Y(new_n5268));
  nand_4 g04892(.A(new_n5268), .B(new_n5265), .Y(new_n5269));
  nand_4 g04893(.A(new_n5269), .B(new_n5260), .Y(new_n5270));
  nand_4 g04894(.A(new_n5270), .B(new_n5257_1), .Y(new_n5271));
  nor_4  g04895(.A(new_n5244), .B(new_n5242), .Y(new_n5272));
  nor_4  g04896(.A(new_n5272), .B(new_n5246), .Y(new_n5273));
  nand_4 g04897(.A(new_n5273), .B(new_n5271), .Y(new_n5274));
  nand_4 g04898(.A(new_n5274), .B(new_n5247), .Y(new_n5275));
  nand_4 g04899(.A(new_n5275), .B(new_n5240_1), .Y(new_n5276));
  nand_4 g04900(.A(new_n5276), .B(new_n5237), .Y(new_n5277));
  nand_4 g04901(.A(new_n5277), .B(new_n5232), .Y(new_n5278));
  nand_4 g04902(.A(new_n5278), .B(new_n5231), .Y(new_n5279));
  nand_4 g04903(.A(new_n5279), .B(new_n5225), .Y(new_n5280));
  nand_4 g04904(.A(new_n5280), .B(new_n5223), .Y(new_n5281));
  nand_4 g04905(.A(new_n4662), .B(new_n4655), .Y(new_n5282));
  nand_4 g04906(.A(new_n4676), .B(new_n4663), .Y(new_n5283_1));
  nand_4 g04907(.A(new_n5283_1), .B(new_n5282), .Y(new_n5284));
  not_3  g04908(.A(new_n4658), .Y(new_n5285));
  nor_4  g04909(.A(new_n4660), .B(new_n5285), .Y(new_n5286));
  not_3  g04910(.A(new_n4657), .Y(new_n5287));
  nor_4  g04911(.A(new_n4661), .B(new_n5287), .Y(new_n5288));
  nor_4  g04912(.A(new_n5288), .B(new_n5286), .Y(new_n5289));
  xor_3  g04913(.A(new_n5289), .B(new_n5284), .Y(new_n5290));
  xnor_3 g04914(.A(new_n5290), .B(new_n5281), .Y(new_n5291));
  nor_4  g04915(.A(new_n4823), .B(new_n4780), .Y(new_n5292));
  nor_4  g04916(.A(new_n4844), .B(new_n4824), .Y(new_n5293));
  nor_4  g04917(.A(new_n5293), .B(new_n5292), .Y(new_n5294));
  nand_4 g04918(.A(new_n4968), .B(new_n4934), .Y(new_n5295));
  not_3  g04919(.A(new_n4969), .Y(new_n5296));
  nand_4 g04920(.A(new_n5296), .B(new_n5163), .Y(new_n5297));
  nand_4 g04921(.A(new_n5297), .B(new_n5295), .Y(new_n5298));
  xnor_3 g04922(.A(new_n5298), .B(new_n5294), .Y(new_n5299));
  nand_4 g04923(.A(n10327), .B(n3172), .Y(new_n5300));
  nand_4 g04924(.A(n4203), .B(n3022), .Y(new_n5301));
  xor_3  g04925(.A(new_n5301), .B(new_n5300), .Y(new_n5302));
  or_4   g04926(.A(new_n4806), .B(new_n4800), .Y(new_n5303));
  not_3  g04927(.A(new_n5303), .Y(new_n5304));
  nor_4  g04928(.A(new_n5304), .B(new_n4807), .Y(new_n5305_1));
  nand_4 g04929(.A(n10278), .B(n2464), .Y(new_n5306));
  not_3  g04930(.A(new_n5306), .Y(new_n5307));
  nand_4 g04931(.A(n11023), .B(n4187), .Y(new_n5308));
  nand_4 g04932(.A(n11311), .B(n10451), .Y(new_n5309));
  xor_3  g04933(.A(new_n5309), .B(new_n5308), .Y(new_n5310));
  xor_3  g04934(.A(new_n5310), .B(new_n5307), .Y(new_n5311));
  xnor_3 g04935(.A(new_n5311), .B(new_n5305_1), .Y(new_n5312));
  nand_4 g04936(.A(new_n4798), .B(new_n4796), .Y(new_n5313));
  nand_4 g04937(.A(new_n4809), .B(new_n4799), .Y(new_n5314_1));
  nand_4 g04938(.A(new_n5314_1), .B(new_n5313), .Y(new_n5315));
  nand_4 g04939(.A(n11423), .B(n9400), .Y(new_n5316));
  not_3  g04940(.A(new_n5316), .Y(new_n5317));
  xor_3  g04941(.A(new_n5317), .B(new_n5315), .Y(new_n5318));
  xnor_3 g04942(.A(new_n5318), .B(new_n5312), .Y(new_n5319_1));
  xnor_3 g04943(.A(new_n5319_1), .B(new_n5302), .Y(new_n5320_1));
  not_3  g04944(.A(new_n4794), .Y(new_n5321));
  nor_4  g04945(.A(new_n5321), .B(new_n4784), .Y(new_n5322));
  not_3  g04946(.A(new_n4795), .Y(new_n5323));
  nor_4  g04947(.A(new_n4811), .B(new_n5323), .Y(new_n5324));
  nor_4  g04948(.A(new_n5324), .B(new_n5322), .Y(new_n5325));
  nand_4 g04949(.A(new_n5074), .B(new_n5047), .Y(new_n5326));
  nand_4 g04950(.A(new_n5095), .B(new_n5075), .Y(new_n5327));
  nand_4 g04951(.A(new_n5327), .B(new_n5326), .Y(new_n5328));
  xnor_3 g04952(.A(new_n5328), .B(new_n5325), .Y(new_n5329));
  xnor_3 g04953(.A(new_n5329), .B(new_n5320_1), .Y(new_n5330));
  xnor_3 g04954(.A(new_n5330), .B(new_n5299), .Y(new_n5331_1));
  nand_4 g04955(.A(new_n5220), .B(new_n5158), .Y(new_n5332));
  nand_4 g04956(.A(new_n5332), .B(new_n5167), .Y(new_n5333));
  xnor_3 g04957(.A(new_n5333), .B(new_n5331_1), .Y(new_n5334));
  nand_4 g04958(.A(new_n4666), .B(new_n4664), .Y(new_n5335));
  nor_4  g04959(.A(new_n4674), .B(new_n4668), .Y(new_n5336));
  not_3  g04960(.A(new_n5336), .Y(new_n5337));
  nand_4 g04961(.A(new_n5337), .B(new_n5335), .Y(new_n5338));
  nand_4 g04962(.A(n12591), .B(n11821), .Y(new_n5339));
  nand_4 g04963(.A(n9080), .B(n3932), .Y(new_n5340));
  xor_3  g04964(.A(new_n5340), .B(new_n5339), .Y(new_n5341));
  nand_4 g04965(.A(n10174), .B(n6703), .Y(new_n5342));
  nand_4 g04966(.A(n12753), .B(n9640), .Y(new_n5343));
  not_3  g04967(.A(new_n5343), .Y(new_n5344));
  xor_3  g04968(.A(new_n5344), .B(new_n5342), .Y(new_n5345));
  nand_4 g04969(.A(n9583), .B(n1333), .Y(new_n5346));
  nand_4 g04970(.A(n6877), .B(n2278), .Y(new_n5347));
  xor_3  g04971(.A(new_n5347), .B(new_n5346), .Y(new_n5348));
  xor_3  g04972(.A(new_n5348), .B(new_n5345), .Y(new_n5349));
  xnor_3 g04973(.A(new_n5349), .B(new_n5341), .Y(new_n5350));
  xnor_3 g04974(.A(new_n5350), .B(new_n5338), .Y(new_n5351));
  nand_4 g04975(.A(new_n4684), .B(new_n4650), .Y(new_n5352));
  nand_4 g04976(.A(new_n4707), .B(new_n4685), .Y(new_n5353));
  nand_4 g04977(.A(new_n5353), .B(new_n5352), .Y(new_n5354));
  nand_4 g04978(.A(new_n4965), .B(new_n4964), .Y(new_n5355));
  not_3  g04979(.A(new_n4962), .Y(new_n5356));
  nand_4 g04980(.A(new_n4967), .B(new_n5356), .Y(new_n5357));
  nand_4 g04981(.A(new_n5357), .B(new_n5355), .Y(new_n5358));
  nand_4 g04982(.A(n11922), .B(n6294), .Y(new_n5359));
  nand_4 g04983(.A(new_n4951), .B(new_n4949), .Y(new_n5360));
  nand_4 g04984(.A(new_n4960), .B(new_n4952), .Y(new_n5361));
  nand_4 g04985(.A(new_n5361), .B(new_n5360), .Y(new_n5362));
  nand_4 g04986(.A(n11478), .B(n4094), .Y(new_n5363));
  not_3  g04987(.A(new_n5363), .Y(new_n5364));
  xnor_3 g04988(.A(new_n5364), .B(new_n5362), .Y(new_n5365));
  nor_4  g04989(.A(new_n5051), .B(new_n5050), .Y(new_n5366));
  not_3  g04990(.A(new_n5052), .Y(new_n5367));
  nor_4  g04991(.A(new_n5058), .B(new_n5367), .Y(new_n5368));
  nor_4  g04992(.A(new_n5368), .B(new_n5366), .Y(new_n5369));
  not_3  g04993(.A(new_n5062), .Y(new_n5370));
  nor_4  g04994(.A(new_n5064), .B(new_n5370), .Y(new_n5371));
  not_3  g04995(.A(new_n5061), .Y(new_n5372));
  nor_4  g04996(.A(new_n5065), .B(new_n5372), .Y(new_n5373));
  nor_4  g04997(.A(new_n5373), .B(new_n5371), .Y(new_n5374));
  nand_4 g04998(.A(n12247), .B(n3992), .Y(new_n5375));
  nand_4 g04999(.A(n8384), .B(n1510), .Y(new_n5376));
  not_3  g05000(.A(new_n5376), .Y(new_n5377));
  xor_3  g05001(.A(new_n5377), .B(new_n5375), .Y(new_n5378));
  xnor_3 g05002(.A(new_n5378), .B(new_n5374), .Y(new_n5379));
  xnor_3 g05003(.A(new_n5379), .B(new_n5369), .Y(new_n5380));
  xnor_3 g05004(.A(new_n5380), .B(new_n5365), .Y(new_n5381));
  xnor_3 g05005(.A(new_n5381), .B(new_n5359), .Y(new_n5382));
  xnor_3 g05006(.A(new_n5382), .B(new_n5358), .Y(new_n5383));
  xnor_3 g05007(.A(new_n5383), .B(new_n5354), .Y(new_n5384));
  nand_4 g05008(.A(new_n5071), .B(new_n5070), .Y(new_n5385));
  not_3  g05009(.A(new_n5068), .Y(new_n5386));
  nand_4 g05010(.A(new_n5073), .B(new_n5386), .Y(new_n5387));
  nand_4 g05011(.A(new_n5387), .B(new_n5385), .Y(new_n5388));
  not_3  g05012(.A(new_n5060), .Y(new_n5389));
  nand_4 g05013(.A(new_n5066), .B(new_n5389), .Y(new_n5390));
  not_3  g05014(.A(new_n5059), .Y(new_n5391));
  nand_4 g05015(.A(new_n5067), .B(new_n5391), .Y(new_n5392));
  nand_4 g05016(.A(new_n5392), .B(new_n5390), .Y(new_n5393));
  not_3  g05017(.A(new_n4947), .Y(new_n5394));
  nor_4  g05018(.A(new_n5394), .B(new_n4937), .Y(new_n5395));
  not_3  g05019(.A(new_n4948), .Y(new_n5396));
  nor_4  g05020(.A(new_n4961), .B(new_n5396), .Y(new_n5397));
  nor_4  g05021(.A(new_n5397), .B(new_n5395), .Y(new_n5398));
  xnor_3 g05022(.A(new_n5398), .B(new_n5393), .Y(new_n5399));
  xnor_3 g05023(.A(new_n5399), .B(new_n5388), .Y(new_n5400));
  not_3  g05024(.A(new_n4956), .Y(new_n5401));
  nor_4  g05025(.A(new_n4958), .B(new_n5401), .Y(new_n5402));
  nor_4  g05026(.A(new_n4959), .B(new_n4955), .Y(new_n5403));
  nor_4  g05027(.A(new_n5403), .B(new_n5402), .Y(new_n5404));
  nand_4 g05028(.A(n7862), .B(n753), .Y(new_n5405));
  nand_4 g05029(.A(n12511), .B(n7236), .Y(new_n5406));
  not_3  g05030(.A(new_n5406), .Y(new_n5407));
  xor_3  g05031(.A(new_n5407), .B(new_n5405), .Y(new_n5408));
  xnor_3 g05032(.A(new_n5408), .B(new_n5404), .Y(new_n5409));
  nand_4 g05033(.A(new_n4792), .B(new_n4786), .Y(new_n5410));
  nand_4 g05034(.A(new_n5410), .B(new_n4791), .Y(new_n5411_1));
  nand_4 g05035(.A(n10898), .B(n7646), .Y(new_n5412));
  nand_4 g05036(.A(n6826), .B(n1798), .Y(new_n5413));
  xor_3  g05037(.A(new_n5413), .B(new_n5412), .Y(new_n5414));
  nand_4 g05038(.A(n11876), .B(n4722), .Y(new_n5415));
  nand_4 g05039(.A(n3754), .B(n1471), .Y(new_n5416));
  xor_3  g05040(.A(new_n5416), .B(new_n5415), .Y(new_n5417));
  xnor_3 g05041(.A(new_n5417), .B(new_n5414), .Y(new_n5418));
  xnor_3 g05042(.A(new_n5418), .B(new_n5411_1), .Y(new_n5419));
  xnor_3 g05043(.A(new_n5419), .B(new_n5409), .Y(new_n5420));
  nand_4 g05044(.A(n3146), .B(n1067), .Y(new_n5421));
  nand_4 g05045(.A(n2551), .B(n137), .Y(new_n5422));
  xor_3  g05046(.A(new_n5422), .B(new_n5421), .Y(new_n5423));
  nand_4 g05047(.A(n8665), .B(n6797), .Y(new_n5424));
  nand_4 g05048(.A(n12826), .B(n5283), .Y(new_n5425));
  xor_3  g05049(.A(new_n5425), .B(new_n5424), .Y(new_n5426));
  xnor_3 g05050(.A(new_n5426), .B(new_n5423), .Y(new_n5427));
  nand_4 g05051(.A(new_n4942), .B(new_n4939), .Y(new_n5428));
  nand_4 g05052(.A(new_n5428), .B(new_n4945), .Y(new_n5429));
  nand_4 g05053(.A(n10685), .B(n4805), .Y(new_n5430));
  nand_4 g05054(.A(n5645), .B(n4938), .Y(new_n5431));
  xor_3  g05055(.A(new_n5431), .B(new_n5430), .Y(new_n5432));
  xnor_3 g05056(.A(new_n5432), .B(new_n5429), .Y(new_n5433));
  xnor_3 g05057(.A(new_n5433), .B(new_n5427), .Y(new_n5434));
  not_3  g05058(.A(new_n5054), .Y(new_n5435_1));
  nor_4  g05059(.A(new_n5056), .B(new_n5435_1), .Y(new_n5436));
  not_3  g05060(.A(new_n5053), .Y(new_n5437));
  nor_4  g05061(.A(new_n5057), .B(new_n5437), .Y(new_n5438));
  nor_4  g05062(.A(new_n5438), .B(new_n5436), .Y(new_n5439));
  nand_4 g05063(.A(n6358), .B(n159), .Y(new_n5440));
  nand_4 g05064(.A(n5198), .B(n2749), .Y(new_n5441));
  xor_3  g05065(.A(new_n5441), .B(new_n5440), .Y(new_n5442));
  xnor_3 g05066(.A(new_n5442), .B(new_n5439), .Y(new_n5443));
  xnor_3 g05067(.A(new_n5443), .B(new_n5434), .Y(new_n5444));
  xnor_3 g05068(.A(new_n5444), .B(new_n5420), .Y(new_n5445));
  nand_4 g05069(.A(new_n4681), .B(new_n4680), .Y(new_n5446));
  nand_4 g05070(.A(new_n4683), .B(new_n4677), .Y(new_n5447));
  nand_4 g05071(.A(new_n5447), .B(new_n5446), .Y(new_n5448));
  xnor_3 g05072(.A(new_n5448), .B(new_n5445), .Y(new_n5449));
  xnor_3 g05073(.A(new_n5449), .B(new_n5400), .Y(new_n5450));
  xnor_3 g05074(.A(new_n5450), .B(new_n5384), .Y(new_n5451));
  xnor_3 g05075(.A(new_n5451), .B(new_n5351), .Y(new_n5452));
  nor_4  g05076(.A(new_n4819), .B(new_n4817_1), .Y(new_n5453));
  nor_4  g05077(.A(new_n4822), .B(new_n4812), .Y(new_n5454));
  nor_4  g05078(.A(new_n5454), .B(new_n5453), .Y(new_n5455));
  nand_4 g05079(.A(new_n5096), .B(new_n4970_1), .Y(new_n5456));
  nand_4 g05080(.A(new_n5156), .B(new_n5165), .Y(new_n5457));
  nand_4 g05081(.A(new_n5457), .B(new_n5456), .Y(new_n5458));
  xnor_3 g05082(.A(new_n5458), .B(new_n5455), .Y(new_n5459));
  xnor_3 g05083(.A(new_n5459), .B(new_n5452), .Y(new_n5460));
  nor_4  g05084(.A(new_n4671), .B(new_n4670), .Y(new_n5461));
  not_3  g05085(.A(new_n4670), .Y(new_n5462));
  nor_4  g05086(.A(new_n4672), .B(new_n5462), .Y(new_n5463));
  or_4   g05087(.A(new_n5463), .B(new_n4669), .Y(new_n5464));
  not_3  g05088(.A(new_n5464), .Y(new_n5465));
  or_4   g05089(.A(new_n5465), .B(new_n5461), .Y(new_n5466));
  nand_4 g05090(.A(n11757), .B(n11662), .Y(new_n5467));
  nand_4 g05091(.A(n7456), .B(n5240), .Y(new_n5468));
  xor_3  g05092(.A(new_n5468), .B(new_n5467), .Y(new_n5469));
  xor_3  g05093(.A(new_n5469), .B(new_n5466), .Y(new_n5470));
  not_3  g05094(.A(new_n5470), .Y(new_n5471));
  xnor_3 g05095(.A(new_n5471), .B(new_n5460), .Y(new_n5472));
  xnor_3 g05096(.A(new_n5472), .B(new_n5334), .Y(new_n5473));
  nand_4 g05097(.A(new_n5473), .B(new_n5291), .Y(new_n5474));
  not_3  g05098(.A(new_n5290), .Y(new_n5475));
  xnor_3 g05099(.A(new_n5475), .B(new_n5281), .Y(new_n5476));
  xnor_3 g05100(.A(new_n5470), .B(new_n5460), .Y(new_n5477));
  xnor_3 g05101(.A(new_n5477), .B(new_n5334), .Y(new_n5478));
  nand_4 g05102(.A(new_n5478), .B(new_n5476), .Y(new_n5479));
  nand_4 g05103(.A(new_n5479), .B(new_n5474), .Y(n1269));
  nand_4 g05104(.A(n10223), .B(n4312), .Y(new_n5481));
  not_3  g05105(.A(new_n5481), .Y(new_n5482));
  nand_4 g05106(.A(n12705), .B(n7265), .Y(new_n5483));
  nand_4 g05107(.A(n4312), .B(n2879), .Y(new_n5484));
  not_3  g05108(.A(new_n5484), .Y(new_n5485));
  nand_4 g05109(.A(n10223), .B(n1097), .Y(new_n5486));
  xnor_3 g05110(.A(new_n5486), .B(new_n5483), .Y(new_n5487));
  nor_4  g05111(.A(new_n5487), .B(new_n5485), .Y(new_n5488));
  nor_4  g05112(.A(new_n5488), .B(new_n5483), .Y(new_n5489));
  nor_4  g05113(.A(new_n5489), .B(new_n5482), .Y(new_n5490));
  nor_4  g05114(.A(new_n5489), .B(new_n1087), .Y(new_n5491));
  nor_4  g05115(.A(new_n5491), .B(new_n5481), .Y(new_n5492));
  nor_4  g05116(.A(new_n5492), .B(new_n5490), .Y(new_n5493));
  nand_4 g05117(.A(n12025), .B(n7265), .Y(new_n5494));
  nand_4 g05118(.A(n12705), .B(n2879), .Y(new_n5495));
  xor_3  g05119(.A(new_n5495), .B(new_n5494), .Y(new_n5496));
  xnor_3 g05120(.A(new_n5496), .B(new_n5493), .Y(new_n5497));
  not_3  g05121(.A(new_n5497), .Y(new_n5498));
  nand_4 g05122(.A(n9195), .B(n5964), .Y(new_n5499));
  nand_4 g05123(.A(n4634), .B(n1097), .Y(new_n5500));
  xor_3  g05124(.A(new_n5500), .B(new_n5499), .Y(new_n5501));
  xnor_3 g05125(.A(new_n5501), .B(new_n5498), .Y(new_n5502));
  nand_4 g05126(.A(n5964), .B(n4634), .Y(new_n5503));
  not_3  g05127(.A(new_n5503), .Y(new_n5504));
  not_3  g05128(.A(new_n1088), .Y(new_n5505));
  not_3  g05129(.A(new_n1089), .Y(new_n5506));
  nor_4  g05130(.A(new_n5506), .B(new_n5505), .Y(new_n5507));
  nor_4  g05131(.A(new_n1089), .B(new_n1088), .Y(new_n5508));
  nor_4  g05132(.A(new_n5508), .B(new_n1087), .Y(new_n5509));
  nor_4  g05133(.A(new_n5509), .B(new_n5507), .Y(new_n5510));
  and_4  g05134(.A(new_n5510), .B(new_n5504), .Y(new_n5511));
  xor_3  g05135(.A(new_n5487), .B(new_n5485), .Y(new_n5512));
  xor_3  g05136(.A(new_n5510), .B(new_n5503), .Y(new_n5513));
  nor_4  g05137(.A(new_n5513), .B(new_n5512), .Y(new_n5514));
  nor_4  g05138(.A(new_n5514), .B(new_n5511), .Y(new_n5515));
  xnor_3 g05139(.A(new_n5515), .B(new_n5502), .Y(new_n5516));
  not_3  g05140(.A(new_n5516), .Y(new_n5517));
  nand_4 g05141(.A(n9195), .B(n5305), .Y(new_n5518));
  not_3  g05142(.A(new_n5518), .Y(new_n5519));
  nand_4 g05143(.A(new_n1091), .B(new_n1085), .Y(new_n5520));
  nand_4 g05144(.A(new_n5520), .B(new_n1082), .Y(new_n5521));
  nor_4  g05145(.A(new_n5521), .B(new_n5519), .Y(new_n5522));
  xor_3  g05146(.A(new_n5510), .B(new_n5504), .Y(new_n5523));
  xnor_3 g05147(.A(new_n5523), .B(new_n5512), .Y(new_n5524));
  xnor_3 g05148(.A(new_n5521), .B(new_n5519), .Y(new_n5525));
  nor_4  g05149(.A(new_n5525), .B(new_n5524), .Y(new_n5526));
  nor_4  g05150(.A(new_n5526), .B(new_n5522), .Y(new_n5527));
  nand_4 g05151(.A(new_n5527), .B(new_n5517), .Y(new_n5528));
  not_3  g05152(.A(new_n5492), .Y(new_n5529));
  nand_4 g05153(.A(new_n5496), .B(new_n5493), .Y(new_n5530));
  nand_4 g05154(.A(new_n5530), .B(new_n5529), .Y(new_n5531));
  nand_4 g05155(.A(n5964), .B(n2253), .Y(new_n5532));
  nand_4 g05156(.A(n9195), .B(n1097), .Y(new_n5533));
  nand_4 g05157(.A(n5305), .B(n3865), .Y(new_n5534));
  not_3  g05158(.A(new_n5534), .Y(new_n5535));
  xor_3  g05159(.A(new_n5535), .B(new_n5533), .Y(new_n5536));
  xnor_3 g05160(.A(new_n5536), .B(new_n5532), .Y(new_n5537));
  xnor_3 g05161(.A(new_n5537), .B(new_n5531), .Y(new_n5538));
  nor_4  g05162(.A(new_n5495), .B(new_n5494), .Y(new_n5539));
  not_3  g05163(.A(new_n5539), .Y(new_n5540));
  nand_4 g05164(.A(n4634), .B(n4312), .Y(new_n5541));
  xor_3  g05165(.A(new_n5541), .B(new_n5540), .Y(new_n5542));
  nand_4 g05166(.A(n12025), .B(n2879), .Y(new_n5543));
  nand_4 g05167(.A(n11257), .B(n7265), .Y(new_n5544));
  nand_4 g05168(.A(n12705), .B(n10223), .Y(new_n5545));
  not_3  g05169(.A(new_n5545), .Y(new_n5546));
  xor_3  g05170(.A(new_n5546), .B(new_n5544), .Y(new_n5547));
  xnor_3 g05171(.A(new_n5547), .B(new_n5543), .Y(new_n5548));
  xnor_3 g05172(.A(new_n5548), .B(new_n5542), .Y(new_n5549));
  xnor_3 g05173(.A(new_n5549), .B(new_n5538), .Y(new_n5550));
  nand_4 g05174(.A(new_n5501), .B(new_n5498), .Y(new_n5551));
  nor_4  g05175(.A(new_n5500), .B(new_n5499), .Y(new_n5552));
  nor_4  g05176(.A(new_n5515), .B(new_n5502), .Y(new_n5553));
  xnor_3 g05177(.A(new_n5553), .B(new_n5552), .Y(new_n5554));
  nand_4 g05178(.A(new_n5554), .B(new_n5551), .Y(new_n5555));
  xnor_3 g05179(.A(new_n5555), .B(new_n5550), .Y(new_n5556));
  xnor_3 g05180(.A(new_n5556), .B(new_n5528), .Y(new_n5557));
  not_3  g05181(.A(new_n5557), .Y(new_n5558));
  nand_4 g05182(.A(n5305), .B(n2253), .Y(new_n5559));
  not_3  g05183(.A(new_n5559), .Y(new_n5560));
  xnor_3 g05184(.A(new_n5527), .B(new_n5516), .Y(new_n5561));
  nand_4 g05185(.A(new_n5561), .B(new_n5560), .Y(new_n5562));
  nor_4  g05186(.A(new_n1101), .B(new_n1093), .Y(new_n5563));
  not_3  g05187(.A(new_n5563), .Y(new_n5564));
  not_3  g05188(.A(new_n5525), .Y(new_n5565));
  xnor_3 g05189(.A(new_n5565), .B(new_n5524), .Y(new_n5566));
  nor_4  g05190(.A(new_n5566), .B(new_n5564), .Y(new_n5567));
  xnor_3 g05191(.A(new_n5561), .B(new_n5559), .Y(new_n5568));
  nand_4 g05192(.A(new_n5568), .B(new_n5567), .Y(new_n5569));
  nand_4 g05193(.A(new_n5569), .B(new_n5562), .Y(new_n5570));
  xor_3  g05194(.A(new_n5570), .B(new_n5558), .Y(new_n5571));
  not_3  g05195(.A(new_n5569), .Y(new_n5572));
  nor_4  g05196(.A(new_n5568), .B(new_n5567), .Y(new_n5573));
  nor_4  g05197(.A(new_n5573), .B(new_n5572), .Y(new_n5574));
  not_3  g05198(.A(new_n5574), .Y(new_n5575));
  nor_4  g05199(.A(new_n1229), .B(new_n1226), .Y(new_n5576));
  not_3  g05200(.A(new_n5576), .Y(new_n5577));
  nand_4 g05201(.A(n12145), .B(n8759), .Y(new_n5578));
  not_3  g05202(.A(new_n1216), .Y(new_n5579_1));
  nand_4 g05203(.A(new_n1217), .B(new_n5579_1), .Y(new_n5580));
  nand_4 g05204(.A(new_n1225), .B(new_n1218), .Y(new_n5581));
  nand_4 g05205(.A(new_n5581), .B(new_n5580), .Y(new_n5582));
  not_3  g05206(.A(new_n5582), .Y(new_n5583));
  xnor_3 g05207(.A(new_n5583), .B(new_n5578), .Y(new_n5584));
  nand_4 g05208(.A(n6776), .B(n2522), .Y(new_n5585));
  not_3  g05209(.A(new_n1222), .Y(new_n5586));
  not_3  g05210(.A(new_n1223), .Y(new_n5587));
  nor_4  g05211(.A(new_n5587), .B(new_n5586), .Y(new_n5588));
  nor_4  g05212(.A(new_n1223), .B(new_n1222), .Y(new_n5589));
  nor_4  g05213(.A(new_n5589), .B(new_n1221), .Y(new_n5590));
  nor_4  g05214(.A(new_n5590), .B(new_n5588), .Y(new_n5591));
  xnor_3 g05215(.A(new_n5591), .B(new_n5585), .Y(new_n5592));
  nand_4 g05216(.A(n7436), .B(n2024), .Y(new_n5593));
  not_3  g05217(.A(new_n5593), .Y(new_n5594));
  nand_4 g05218(.A(n12299), .B(n9189), .Y(new_n5595));
  nand_4 g05219(.A(n8276), .B(n7946), .Y(new_n5596));
  xnor_3 g05220(.A(new_n5596), .B(new_n5595), .Y(new_n5597));
  xnor_3 g05221(.A(new_n5597), .B(new_n5594), .Y(new_n5598));
  xnor_3 g05222(.A(new_n5598), .B(new_n5592), .Y(new_n5599));
  not_3  g05223(.A(new_n5599), .Y(new_n5600));
  xor_3  g05224(.A(new_n5600), .B(new_n5584), .Y(new_n5601));
  nor_4  g05225(.A(new_n5601), .B(new_n5577), .Y(new_n5602));
  not_3  g05226(.A(new_n5602), .Y(new_n5603));
  nand_4 g05227(.A(n12221), .B(n8759), .Y(new_n5604));
  not_3  g05228(.A(new_n5585), .Y(new_n5605));
  nand_4 g05229(.A(new_n5591), .B(new_n5605), .Y(new_n5606));
  nand_4 g05230(.A(new_n5598), .B(new_n5592), .Y(new_n5607));
  nand_4 g05231(.A(new_n5607), .B(new_n5606), .Y(new_n5608));
  nand_4 g05232(.A(n12145), .B(n6776), .Y(new_n5609));
  nand_4 g05233(.A(n12299), .B(n2522), .Y(new_n5610));
  xor_3  g05234(.A(new_n5610), .B(new_n5609), .Y(new_n5611));
  xnor_3 g05235(.A(new_n5611), .B(new_n5608), .Y(new_n5612));
  nand_4 g05236(.A(n9189), .B(n7436), .Y(new_n5613));
  not_3  g05237(.A(new_n5613), .Y(new_n5614));
  nor_4  g05238(.A(new_n5597), .B(new_n5594), .Y(new_n5615));
  nor_4  g05239(.A(new_n5615), .B(new_n5596), .Y(new_n5616));
  nor_4  g05240(.A(new_n5616), .B(new_n5614), .Y(new_n5617));
  nor_4  g05241(.A(new_n5616), .B(new_n1221), .Y(new_n5618));
  nor_4  g05242(.A(new_n5618), .B(new_n5613), .Y(new_n5619));
  nor_4  g05243(.A(new_n5619), .B(new_n5617), .Y(new_n5620));
  nand_4 g05244(.A(n8276), .B(n2024), .Y(new_n5621));
  nand_4 g05245(.A(n9241), .B(n7946), .Y(new_n5622));
  xor_3  g05246(.A(new_n5622), .B(new_n5621), .Y(new_n5623));
  xnor_3 g05247(.A(new_n5623), .B(new_n5620), .Y(new_n5624));
  xnor_3 g05248(.A(new_n5624), .B(new_n5612), .Y(new_n5625));
  nor_4  g05249(.A(new_n5583), .B(new_n5578), .Y(new_n5626));
  nor_4  g05250(.A(new_n5599), .B(new_n5584), .Y(new_n5627));
  nor_4  g05251(.A(new_n5627), .B(new_n5626), .Y(new_n5628));
  xnor_3 g05252(.A(new_n5628), .B(new_n5625), .Y(new_n5629));
  nor_4  g05253(.A(new_n5629), .B(new_n5604), .Y(new_n5630));
  not_3  g05254(.A(new_n5604), .Y(new_n5631));
  not_3  g05255(.A(new_n5629), .Y(new_n5632));
  nor_4  g05256(.A(new_n5632), .B(new_n5631), .Y(new_n5633));
  nor_4  g05257(.A(new_n5633), .B(new_n5630), .Y(new_n5634));
  xnor_3 g05258(.A(new_n5634), .B(new_n5603), .Y(new_n5635));
  xnor_3 g05259(.A(new_n5601), .B(new_n5576), .Y(new_n5636));
  nand_4 g05260(.A(n6016), .B(n5331), .Y(new_n5637));
  nand_4 g05261(.A(n8476), .B(n521), .Y(new_n5638));
  not_3  g05262(.A(new_n5638), .Y(new_n5639));
  not_3  g05263(.A(new_n1241), .Y(new_n5640));
  nor_4  g05264(.A(new_n1247), .B(new_n5640), .Y(new_n5641_1));
  nor_4  g05265(.A(new_n5641_1), .B(new_n1246), .Y(new_n5642));
  xnor_3 g05266(.A(new_n5642), .B(new_n5639), .Y(new_n5643));
  nand_4 g05267(.A(n12648), .B(n2498), .Y(new_n5644));
  not_3  g05268(.A(new_n5644), .Y(new_n5645_1));
  nand_4 g05269(.A(n5579), .B(n2530), .Y(new_n5646));
  not_3  g05270(.A(new_n5646), .Y(new_n5647));
  nand_4 g05271(.A(n10545), .B(n2558), .Y(new_n5648));
  not_3  g05272(.A(new_n5648), .Y(new_n5649));
  nor_4  g05273(.A(new_n5649), .B(new_n5647), .Y(new_n5650));
  nor_4  g05274(.A(new_n5648), .B(new_n5646), .Y(new_n5651));
  nor_4  g05275(.A(new_n5651), .B(new_n5650), .Y(new_n5652));
  xnor_3 g05276(.A(new_n5652), .B(new_n5645_1), .Y(new_n5653));
  xnor_3 g05277(.A(new_n5653), .B(new_n5643), .Y(new_n5654));
  nor_4  g05278(.A(new_n5654), .B(new_n5637), .Y(new_n5655));
  not_3  g05279(.A(new_n5637), .Y(new_n5656));
  not_3  g05280(.A(new_n5654), .Y(new_n5657));
  nor_4  g05281(.A(new_n5657), .B(new_n5656), .Y(new_n5658));
  nor_4  g05282(.A(new_n5658), .B(new_n5655), .Y(new_n5659));
  nor_4  g05283(.A(new_n1239), .B(new_n1235), .Y(new_n5660));
  nor_4  g05284(.A(new_n1250), .B(new_n1240), .Y(new_n5661));
  nor_4  g05285(.A(new_n5661), .B(new_n5660), .Y(new_n5662));
  not_3  g05286(.A(new_n5662), .Y(new_n5663));
  xnor_3 g05287(.A(new_n5663), .B(new_n5659), .Y(new_n5664));
  xnor_3 g05288(.A(new_n5664), .B(new_n1255), .Y(new_n5665));
  not_3  g05289(.A(new_n1277), .Y(new_n5666));
  nand_4 g05290(.A(n7965), .B(n7270), .Y(new_n5667));
  nand_4 g05291(.A(n7388), .B(n806), .Y(new_n5668));
  not_3  g05292(.A(new_n5668), .Y(new_n5669));
  not_3  g05293(.A(new_n1263), .Y(new_n5670_1));
  nor_4  g05294(.A(new_n1269_1), .B(new_n5670_1), .Y(new_n5671));
  nor_4  g05295(.A(new_n5671), .B(new_n1268), .Y(new_n5672));
  xnor_3 g05296(.A(new_n5672), .B(new_n5669), .Y(new_n5673));
  nand_4 g05297(.A(n9111), .B(n2393), .Y(new_n5674));
  not_3  g05298(.A(new_n5674), .Y(new_n5675));
  nand_4 g05299(.A(n11892), .B(n3342), .Y(new_n5676));
  not_3  g05300(.A(new_n5676), .Y(new_n5677));
  nand_4 g05301(.A(n9763), .B(n5860), .Y(new_n5678));
  not_3  g05302(.A(new_n5678), .Y(new_n5679));
  nor_4  g05303(.A(new_n5679), .B(new_n5677), .Y(new_n5680));
  nor_4  g05304(.A(new_n5678), .B(new_n5676), .Y(new_n5681));
  nor_4  g05305(.A(new_n5681), .B(new_n5680), .Y(new_n5682));
  xnor_3 g05306(.A(new_n5682), .B(new_n5675), .Y(new_n5683));
  xnor_3 g05307(.A(new_n5683), .B(new_n5673), .Y(new_n5684));
  nor_4  g05308(.A(new_n5684), .B(new_n5667), .Y(new_n5685));
  not_3  g05309(.A(new_n5667), .Y(new_n5686));
  not_3  g05310(.A(new_n5684), .Y(new_n5687));
  nor_4  g05311(.A(new_n5687), .B(new_n5686), .Y(new_n5688));
  nor_4  g05312(.A(new_n5688), .B(new_n5685), .Y(new_n5689));
  nor_4  g05313(.A(new_n1261), .B(new_n1259), .Y(new_n5690));
  nor_4  g05314(.A(new_n1272), .B(new_n1262), .Y(new_n5691));
  nor_4  g05315(.A(new_n5691), .B(new_n5690), .Y(new_n5692));
  not_3  g05316(.A(new_n5692), .Y(new_n5693_1));
  xnor_3 g05317(.A(new_n5693_1), .B(new_n5689), .Y(new_n5694_1));
  nor_4  g05318(.A(new_n5694_1), .B(new_n5666), .Y(new_n5695));
  not_3  g05319(.A(new_n5694_1), .Y(new_n5696));
  nor_4  g05320(.A(new_n5696), .B(new_n1277), .Y(new_n5697));
  nor_4  g05321(.A(new_n5697), .B(new_n5695), .Y(new_n5698));
  xnor_3 g05322(.A(new_n5698), .B(new_n5665), .Y(new_n5699));
  nor_4  g05323(.A(new_n1280), .B(new_n1258), .Y(new_n5700));
  nor_4  g05324(.A(new_n1287), .B(new_n5700), .Y(new_n5701));
  xnor_3 g05325(.A(new_n5701), .B(new_n5699), .Y(new_n5702));
  nor_4  g05326(.A(new_n5702), .B(new_n5636), .Y(new_n5703));
  not_3  g05327(.A(new_n5703), .Y(new_n5704));
  nand_4 g05328(.A(new_n5702), .B(new_n5636), .Y(new_n5705));
  nor_4  g05329(.A(new_n1233), .B(new_n1230), .Y(new_n5706));
  nor_4  g05330(.A(new_n1288), .B(new_n1234), .Y(new_n5707));
  nor_4  g05331(.A(new_n5707), .B(new_n5706), .Y(new_n5708));
  nand_4 g05332(.A(new_n5708), .B(new_n5705), .Y(new_n5709));
  nand_4 g05333(.A(new_n5709), .B(new_n5704), .Y(new_n5710));
  xnor_3 g05334(.A(new_n5710), .B(new_n5635), .Y(new_n5711));
  not_3  g05335(.A(new_n1255), .Y(new_n5712));
  nor_4  g05336(.A(new_n5664), .B(new_n5712), .Y(new_n5713));
  nand_4 g05337(.A(n5798), .B(n5331), .Y(new_n5714));
  nand_4 g05338(.A(n12648), .B(n5579), .Y(new_n5715));
  nand_4 g05339(.A(n10545), .B(n2498), .Y(new_n5716));
  nand_4 g05340(.A(n7690), .B(n2558), .Y(new_n5717));
  xnor_3 g05341(.A(new_n5717), .B(new_n5716), .Y(new_n5718));
  nor_4  g05342(.A(new_n5718), .B(new_n5715), .Y(new_n5719));
  not_3  g05343(.A(new_n5715), .Y(new_n5720));
  not_3  g05344(.A(new_n5718), .Y(new_n5721));
  nor_4  g05345(.A(new_n5721), .B(new_n5720), .Y(new_n5722));
  nor_4  g05346(.A(new_n5722), .B(new_n5719), .Y(new_n5723));
  nor_4  g05347(.A(new_n5651), .B(new_n5645_1), .Y(new_n5724));
  nor_4  g05348(.A(new_n5724), .B(new_n5650), .Y(new_n5725));
  xnor_3 g05349(.A(new_n5725), .B(new_n5723), .Y(new_n5726));
  nand_4 g05350(.A(n8476), .B(n6016), .Y(new_n5727));
  nand_4 g05351(.A(n2530), .B(n521), .Y(new_n5728));
  xor_3  g05352(.A(new_n5728), .B(new_n5727), .Y(new_n5729));
  xnor_3 g05353(.A(new_n5729), .B(new_n5726), .Y(new_n5730));
  and_4  g05354(.A(new_n5642), .B(new_n5639), .Y(new_n5731));
  nor_4  g05355(.A(new_n5653), .B(new_n5643), .Y(new_n5732));
  nor_4  g05356(.A(new_n5732), .B(new_n5731), .Y(new_n5733));
  xnor_3 g05357(.A(new_n5733), .B(new_n5730), .Y(new_n5734));
  not_3  g05358(.A(new_n5655), .Y(new_n5735));
  nand_4 g05359(.A(new_n5663), .B(new_n5659), .Y(new_n5736));
  nand_4 g05360(.A(new_n5736), .B(new_n5735), .Y(new_n5737));
  xnor_3 g05361(.A(new_n5737), .B(new_n5734), .Y(new_n5738));
  nor_4  g05362(.A(new_n5738), .B(new_n5714), .Y(new_n5739));
  not_3  g05363(.A(new_n5714), .Y(new_n5740));
  not_3  g05364(.A(new_n5738), .Y(new_n5741));
  nor_4  g05365(.A(new_n5741), .B(new_n5740), .Y(new_n5742));
  nor_4  g05366(.A(new_n5742), .B(new_n5739), .Y(new_n5743));
  xnor_3 g05367(.A(new_n5743), .B(new_n5713), .Y(new_n5744));
  not_3  g05368(.A(new_n5695), .Y(new_n5745));
  nand_4 g05369(.A(n7965), .B(n5153), .Y(new_n5746));
  nand_4 g05370(.A(n3342), .B(n2393), .Y(new_n5747));
  nand_4 g05371(.A(n9763), .B(n3986), .Y(new_n5748));
  nand_4 g05372(.A(n9111), .B(n5860), .Y(new_n5749));
  xnor_3 g05373(.A(new_n5749), .B(new_n5748), .Y(new_n5750));
  nor_4  g05374(.A(new_n5750), .B(new_n5747), .Y(new_n5751));
  not_3  g05375(.A(new_n5747), .Y(new_n5752));
  not_3  g05376(.A(new_n5750), .Y(new_n5753));
  nor_4  g05377(.A(new_n5753), .B(new_n5752), .Y(new_n5754));
  nor_4  g05378(.A(new_n5754), .B(new_n5751), .Y(new_n5755));
  nor_4  g05379(.A(new_n5681), .B(new_n5675), .Y(new_n5756));
  nor_4  g05380(.A(new_n5756), .B(new_n5680), .Y(new_n5757));
  xnor_3 g05381(.A(new_n5757), .B(new_n5755), .Y(new_n5758));
  nand_4 g05382(.A(n7388), .B(n7270), .Y(new_n5759));
  nand_4 g05383(.A(n11892), .B(n806), .Y(new_n5760_1));
  xor_3  g05384(.A(new_n5760_1), .B(new_n5759), .Y(new_n5761));
  xnor_3 g05385(.A(new_n5761), .B(new_n5758), .Y(new_n5762));
  and_4  g05386(.A(new_n5672), .B(new_n5669), .Y(new_n5763));
  nor_4  g05387(.A(new_n5683), .B(new_n5673), .Y(new_n5764));
  nor_4  g05388(.A(new_n5764), .B(new_n5763), .Y(new_n5765));
  xnor_3 g05389(.A(new_n5765), .B(new_n5762), .Y(new_n5766));
  not_3  g05390(.A(new_n5685), .Y(new_n5767_1));
  nand_4 g05391(.A(new_n5693_1), .B(new_n5689), .Y(new_n5768));
  nand_4 g05392(.A(new_n5768), .B(new_n5767_1), .Y(new_n5769));
  xnor_3 g05393(.A(new_n5769), .B(new_n5766), .Y(new_n5770));
  nor_4  g05394(.A(new_n5770), .B(new_n5746), .Y(new_n5771));
  not_3  g05395(.A(new_n5746), .Y(new_n5772));
  not_3  g05396(.A(new_n5770), .Y(new_n5773));
  nor_4  g05397(.A(new_n5773), .B(new_n5772), .Y(new_n5774));
  nor_4  g05398(.A(new_n5774), .B(new_n5771), .Y(new_n5775));
  nor_4  g05399(.A(new_n5775), .B(new_n5745), .Y(new_n5776));
  xnor_3 g05400(.A(new_n5770), .B(new_n5746), .Y(new_n5777));
  nor_4  g05401(.A(new_n5777), .B(new_n5695), .Y(new_n5778));
  nor_4  g05402(.A(new_n5778), .B(new_n5776), .Y(new_n5779));
  not_3  g05403(.A(new_n5779), .Y(new_n5780));
  xnor_3 g05404(.A(new_n5780), .B(new_n5744), .Y(new_n5781));
  nor_4  g05405(.A(new_n5698), .B(new_n5665), .Y(new_n5782));
  nor_4  g05406(.A(new_n5701), .B(new_n5699), .Y(new_n5783));
  nor_4  g05407(.A(new_n5783), .B(new_n5782), .Y(new_n5784));
  not_3  g05408(.A(new_n5784), .Y(new_n5785));
  xnor_3 g05409(.A(new_n5785), .B(new_n5781), .Y(new_n5786));
  xnor_3 g05410(.A(new_n5786), .B(new_n5711), .Y(new_n5787));
  nor_4  g05411(.A(new_n5787), .B(new_n5575), .Y(new_n5788));
  not_3  g05412(.A(new_n5787), .Y(new_n5789));
  nor_4  g05413(.A(new_n5789), .B(new_n5574), .Y(new_n5790));
  xor_3  g05414(.A(new_n5566), .B(new_n5563), .Y(new_n5791));
  not_3  g05415(.A(new_n5708), .Y(new_n5792));
  nand_4 g05416(.A(new_n5705), .B(new_n5704), .Y(new_n5793));
  xnor_3 g05417(.A(new_n5793), .B(new_n5792), .Y(new_n5794));
  not_3  g05418(.A(new_n5794), .Y(new_n5795));
  nor_4  g05419(.A(new_n5795), .B(new_n5791), .Y(new_n5796));
  not_3  g05420(.A(new_n5791), .Y(new_n5797));
  nor_4  g05421(.A(new_n5794), .B(new_n5797), .Y(new_n5798_1));
  nand_4 g05422(.A(new_n1214), .B(new_n1102), .Y(new_n5799));
  not_3  g05423(.A(new_n5799), .Y(new_n5800));
  nor_4  g05424(.A(new_n1289), .B(new_n1215), .Y(new_n5801));
  nor_4  g05425(.A(new_n5801), .B(new_n5800), .Y(new_n5802));
  nor_4  g05426(.A(new_n5802), .B(new_n5798_1), .Y(new_n5803));
  nor_4  g05427(.A(new_n5803), .B(new_n5796), .Y(new_n5804));
  nor_4  g05428(.A(new_n5804), .B(new_n5790), .Y(new_n5805));
  nor_4  g05429(.A(new_n5805), .B(new_n5788), .Y(new_n5806));
  xnor_3 g05430(.A(new_n5806), .B(new_n5571), .Y(new_n5807));
  not_3  g05431(.A(new_n5630), .Y(new_n5808));
  nand_4 g05432(.A(new_n5634), .B(new_n5602), .Y(new_n5809));
  nand_4 g05433(.A(new_n5809), .B(new_n5808), .Y(new_n5810));
  nor_4  g05434(.A(new_n5628), .B(new_n5625), .Y(new_n5811));
  not_3  g05435(.A(new_n5619), .Y(new_n5812));
  nand_4 g05436(.A(new_n5623), .B(new_n5620), .Y(new_n5813));
  nand_4 g05437(.A(new_n5813), .B(new_n5812), .Y(new_n5814_1));
  nand_4 g05438(.A(n12221), .B(n6776), .Y(new_n5815));
  nand_4 g05439(.A(n12299), .B(n12145), .Y(new_n5816));
  nand_4 g05440(.A(n10217), .B(n8759), .Y(new_n5817));
  not_3  g05441(.A(new_n5817), .Y(new_n5818));
  xor_3  g05442(.A(new_n5818), .B(new_n5816), .Y(new_n5819));
  xnor_3 g05443(.A(new_n5819), .B(new_n5815), .Y(new_n5820));
  xnor_3 g05444(.A(new_n5820), .B(new_n5814_1), .Y(new_n5821));
  nor_4  g05445(.A(new_n5622), .B(new_n5621), .Y(new_n5822));
  nand_4 g05446(.A(n7436), .B(n2522), .Y(new_n5823));
  not_3  g05447(.A(new_n5823), .Y(new_n5824));
  xor_3  g05448(.A(new_n5824), .B(new_n5822), .Y(new_n5825));
  nand_4 g05449(.A(n9241), .B(n2024), .Y(new_n5826));
  nand_4 g05450(.A(n10510), .B(n7946), .Y(new_n5827));
  nand_4 g05451(.A(n9189), .B(n8276), .Y(new_n5828));
  nand_4 g05452(.A(new_n5828), .B(new_n5827), .Y(new_n5829));
  not_3  g05453(.A(new_n5827), .Y(new_n5830));
  not_3  g05454(.A(new_n5828), .Y(new_n5831));
  nand_4 g05455(.A(new_n5831), .B(new_n5830), .Y(new_n5832));
  nand_4 g05456(.A(new_n5832), .B(new_n5829), .Y(new_n5833));
  xor_3  g05457(.A(new_n5833), .B(new_n5826), .Y(new_n5834));
  xnor_3 g05458(.A(new_n5834), .B(new_n5825), .Y(new_n5835));
  xnor_3 g05459(.A(new_n5835), .B(new_n5821), .Y(new_n5836));
  nand_4 g05460(.A(new_n5611), .B(new_n5608), .Y(new_n5837));
  nor_4  g05461(.A(new_n5610), .B(new_n5609), .Y(new_n5838));
  nor_4  g05462(.A(new_n5624), .B(new_n5612), .Y(new_n5839));
  xnor_3 g05463(.A(new_n5839), .B(new_n5838), .Y(new_n5840));
  nand_4 g05464(.A(new_n5840), .B(new_n5837), .Y(new_n5841));
  xnor_3 g05465(.A(new_n5841), .B(new_n5836), .Y(new_n5842));
  not_3  g05466(.A(new_n5842), .Y(new_n5843));
  xor_3  g05467(.A(new_n5843), .B(new_n5811), .Y(new_n5844));
  xnor_3 g05468(.A(new_n5844), .B(new_n5810), .Y(new_n5845));
  not_3  g05469(.A(new_n5710), .Y(new_n5846));
  nand_4 g05470(.A(new_n5846), .B(new_n5635), .Y(new_n5847));
  nand_4 g05471(.A(new_n5786), .B(new_n5711), .Y(new_n5848));
  nand_4 g05472(.A(new_n5848), .B(new_n5847), .Y(new_n5849));
  xnor_3 g05473(.A(new_n5849), .B(new_n5845), .Y(new_n5850));
  not_3  g05474(.A(new_n5734), .Y(new_n5851));
  not_3  g05475(.A(new_n5737), .Y(new_n5852));
  nor_4  g05476(.A(new_n5852), .B(new_n5851), .Y(new_n5853));
  not_3  g05477(.A(new_n5719), .Y(new_n5854));
  nand_4 g05478(.A(new_n5725), .B(new_n5723), .Y(new_n5855));
  nand_4 g05479(.A(new_n5855), .B(new_n5854), .Y(new_n5856));
  nand_4 g05480(.A(n8476), .B(n5798), .Y(new_n5857_1));
  nand_4 g05481(.A(n6016), .B(n2530), .Y(new_n5858));
  nand_4 g05482(.A(n5331), .B(n2347), .Y(new_n5859));
  xnor_3 g05483(.A(new_n5859), .B(new_n5858), .Y(new_n5860_1));
  xnor_3 g05484(.A(new_n5860_1), .B(new_n5857_1), .Y(new_n5861));
  xnor_3 g05485(.A(new_n5861), .B(new_n5856), .Y(new_n5862));
  nor_4  g05486(.A(new_n5717), .B(new_n5716), .Y(new_n5863));
  nand_4 g05487(.A(n12648), .B(n521), .Y(new_n5864));
  xnor_3 g05488(.A(new_n5864), .B(new_n5863), .Y(new_n5865));
  nand_4 g05489(.A(n7690), .B(n2498), .Y(new_n5866));
  not_3  g05490(.A(new_n5866), .Y(new_n5867));
  nand_4 g05491(.A(n10545), .B(n5579), .Y(new_n5868));
  nand_4 g05492(.A(n3616), .B(n2558), .Y(new_n5869));
  xnor_3 g05493(.A(new_n5869), .B(new_n5868), .Y(new_n5870));
  xnor_3 g05494(.A(new_n5870), .B(new_n5867), .Y(new_n5871));
  not_3  g05495(.A(new_n5871), .Y(new_n5872));
  xor_3  g05496(.A(new_n5872), .B(new_n5865), .Y(new_n5873));
  xnor_3 g05497(.A(new_n5873), .B(new_n5862), .Y(new_n5874));
  not_3  g05498(.A(new_n5874), .Y(new_n5875));
  not_3  g05499(.A(new_n5726), .Y(new_n5876));
  nand_4 g05500(.A(new_n5729), .B(new_n5876), .Y(new_n5877));
  nor_4  g05501(.A(new_n5728), .B(new_n5727), .Y(new_n5878));
  not_3  g05502(.A(new_n5730), .Y(new_n5879));
  nor_4  g05503(.A(new_n5733), .B(new_n5879), .Y(new_n5880));
  xnor_3 g05504(.A(new_n5880), .B(new_n5878), .Y(new_n5881));
  nand_4 g05505(.A(new_n5881), .B(new_n5877), .Y(new_n5882));
  xnor_3 g05506(.A(new_n5882), .B(new_n5875), .Y(new_n5883));
  xnor_3 g05507(.A(new_n5883), .B(new_n5853), .Y(new_n5884));
  not_3  g05508(.A(new_n5739), .Y(new_n5885));
  nand_4 g05509(.A(new_n5743), .B(new_n5713), .Y(new_n5886));
  nand_4 g05510(.A(new_n5886), .B(new_n5885), .Y(new_n5887));
  xnor_3 g05511(.A(new_n5887), .B(new_n5884), .Y(new_n5888));
  not_3  g05512(.A(new_n5888), .Y(new_n5889));
  not_3  g05513(.A(new_n5766), .Y(new_n5890));
  not_3  g05514(.A(new_n5769), .Y(new_n5891));
  nor_4  g05515(.A(new_n5891), .B(new_n5890), .Y(new_n5892));
  not_3  g05516(.A(new_n5892), .Y(new_n5893));
  not_3  g05517(.A(new_n5751), .Y(new_n5894));
  nand_4 g05518(.A(new_n5757), .B(new_n5755), .Y(new_n5895));
  nand_4 g05519(.A(new_n5895), .B(new_n5894), .Y(new_n5896));
  nand_4 g05520(.A(n7388), .B(n5153), .Y(new_n5897));
  nand_4 g05521(.A(n11892), .B(n7270), .Y(new_n5898));
  nand_4 g05522(.A(n7965), .B(n2507), .Y(new_n5899));
  xnor_3 g05523(.A(new_n5899), .B(new_n5898), .Y(new_n5900));
  xnor_3 g05524(.A(new_n5900), .B(new_n5897), .Y(new_n5901));
  xnor_3 g05525(.A(new_n5901), .B(new_n5896), .Y(new_n5902));
  nor_4  g05526(.A(new_n5749), .B(new_n5748), .Y(new_n5903));
  nand_4 g05527(.A(n2393), .B(n806), .Y(new_n5904));
  xnor_3 g05528(.A(new_n5904), .B(new_n5903), .Y(new_n5905));
  nand_4 g05529(.A(n9111), .B(n3986), .Y(new_n5906));
  not_3  g05530(.A(new_n5906), .Y(new_n5907));
  nand_4 g05531(.A(n5860), .B(n3342), .Y(new_n5908));
  nand_4 g05532(.A(n9763), .B(n5857), .Y(new_n5909));
  xnor_3 g05533(.A(new_n5909), .B(new_n5908), .Y(new_n5910));
  xnor_3 g05534(.A(new_n5910), .B(new_n5907), .Y(new_n5911));
  not_3  g05535(.A(new_n5911), .Y(new_n5912));
  xor_3  g05536(.A(new_n5912), .B(new_n5905), .Y(new_n5913));
  not_3  g05537(.A(new_n5913), .Y(new_n5914));
  xor_3  g05538(.A(new_n5914), .B(new_n5902), .Y(new_n5915));
  not_3  g05539(.A(new_n5915), .Y(new_n5916));
  not_3  g05540(.A(new_n5758), .Y(new_n5917));
  nand_4 g05541(.A(new_n5761), .B(new_n5917), .Y(new_n5918));
  nor_4  g05542(.A(new_n5760_1), .B(new_n5759), .Y(new_n5919));
  not_3  g05543(.A(new_n5762), .Y(new_n5920));
  nor_4  g05544(.A(new_n5765), .B(new_n5920), .Y(new_n5921));
  xnor_3 g05545(.A(new_n5921), .B(new_n5919), .Y(new_n5922));
  nand_4 g05546(.A(new_n5922), .B(new_n5918), .Y(new_n5923));
  xnor_3 g05547(.A(new_n5923), .B(new_n5916), .Y(new_n5924));
  xnor_3 g05548(.A(new_n5924), .B(new_n5893), .Y(new_n5925));
  nor_4  g05549(.A(new_n5778), .B(new_n5774), .Y(new_n5926));
  not_3  g05550(.A(new_n5926), .Y(new_n5927));
  xnor_3 g05551(.A(new_n5927), .B(new_n5925), .Y(new_n5928));
  not_3  g05552(.A(new_n5928), .Y(new_n5929));
  nor_4  g05553(.A(new_n5929), .B(new_n5889), .Y(new_n5930));
  nor_4  g05554(.A(new_n5928), .B(new_n5888), .Y(new_n5931));
  nor_4  g05555(.A(new_n5931), .B(new_n5930), .Y(new_n5932));
  not_3  g05556(.A(new_n5932), .Y(new_n5933));
  nor_4  g05557(.A(new_n5779), .B(new_n5744), .Y(new_n5934_1));
  not_3  g05558(.A(new_n5934_1), .Y(new_n5935));
  nand_4 g05559(.A(new_n5784), .B(new_n5781), .Y(new_n5936));
  nand_4 g05560(.A(new_n5936), .B(new_n5935), .Y(new_n5937));
  nor_4  g05561(.A(new_n5937), .B(new_n5933), .Y(new_n5938));
  not_3  g05562(.A(new_n5937), .Y(new_n5939));
  nor_4  g05563(.A(new_n5939), .B(new_n5932), .Y(new_n5940));
  nor_4  g05564(.A(new_n5940), .B(new_n5938), .Y(new_n5941));
  xnor_3 g05565(.A(new_n5941), .B(new_n5850), .Y(new_n5942));
  xnor_3 g05566(.A(new_n5942), .B(new_n5807), .Y(n1523));
  nand_4 g05567(.A(n7265), .B(n4189), .Y(new_n5944));
  nand_4 g05568(.A(n10223), .B(n6687), .Y(new_n5945));
  nand_4 g05569(.A(new_n5945), .B(new_n5944), .Y(new_n5946));
  not_3  g05570(.A(new_n5944), .Y(new_n5947));
  not_3  g05571(.A(new_n5945), .Y(new_n5948));
  nand_4 g05572(.A(new_n5948), .B(new_n5947), .Y(new_n5949));
  and_4  g05573(.A(new_n5949), .B(new_n5946), .Y(new_n5950));
  nand_4 g05574(.A(n6687), .B(n2879), .Y(new_n5951));
  nand_4 g05575(.A(n7265), .B(n2564), .Y(new_n5952));
  nor_4  g05576(.A(new_n5952), .B(new_n5951), .Y(new_n5953));
  not_3  g05577(.A(new_n5953), .Y(new_n5954));
  nor_4  g05578(.A(new_n5954), .B(new_n5950), .Y(new_n5955));
  nand_4 g05579(.A(n6687), .B(n4634), .Y(new_n5956));
  not_3  g05580(.A(new_n5956), .Y(new_n5957));
  nand_4 g05581(.A(n2879), .B(n2564), .Y(new_n5958));
  not_3  g05582(.A(new_n5958), .Y(new_n5959));
  nand_4 g05583(.A(new_n5959), .B(new_n5946), .Y(new_n5960));
  nand_4 g05584(.A(new_n5960), .B(new_n5949), .Y(new_n5961));
  xor_3  g05585(.A(new_n5961), .B(new_n5957), .Y(new_n5962));
  nand_4 g05586(.A(n4189), .B(n2879), .Y(new_n5963));
  nand_4 g05587(.A(n10223), .B(n2564), .Y(new_n5964_1));
  nand_4 g05588(.A(n7265), .B(n6770), .Y(new_n5965));
  xnor_3 g05589(.A(new_n5965), .B(new_n5964_1), .Y(new_n5966));
  xor_3  g05590(.A(new_n5966), .B(new_n5963), .Y(new_n5967));
  nand_4 g05591(.A(new_n5967), .B(new_n5962), .Y(new_n5968));
  not_3  g05592(.A(new_n5968), .Y(new_n5969));
  nor_4  g05593(.A(new_n5967), .B(new_n5962), .Y(new_n5970));
  nor_4  g05594(.A(new_n5970), .B(new_n5969), .Y(new_n5971));
  nand_4 g05595(.A(new_n5971), .B(new_n5955), .Y(new_n5972));
  not_3  g05596(.A(new_n5972), .Y(new_n5973));
  nand_4 g05597(.A(n9195), .B(n6687), .Y(new_n5974));
  nand_4 g05598(.A(n4634), .B(n2564), .Y(new_n5975));
  nand_4 g05599(.A(n6770), .B(n2879), .Y(new_n5976));
  nand_4 g05600(.A(n10223), .B(n4189), .Y(new_n5977));
  nand_4 g05601(.A(n9920), .B(n7265), .Y(new_n5978));
  xnor_3 g05602(.A(new_n5978), .B(new_n5977), .Y(new_n5979));
  xnor_3 g05603(.A(new_n5979), .B(new_n5976), .Y(new_n5980));
  xnor_3 g05604(.A(new_n5980), .B(new_n5975), .Y(new_n5981));
  nand_4 g05605(.A(new_n5965), .B(new_n5964_1), .Y(new_n5982));
  not_3  g05606(.A(new_n5982), .Y(new_n5983));
  not_3  g05607(.A(new_n5963), .Y(new_n5984));
  nor_4  g05608(.A(new_n5966), .B(new_n5984), .Y(new_n5985));
  nor_4  g05609(.A(new_n5985), .B(new_n5983), .Y(new_n5986));
  xnor_3 g05610(.A(new_n5986), .B(new_n5981), .Y(new_n5987));
  not_3  g05611(.A(new_n5987), .Y(new_n5988));
  nor_4  g05612(.A(new_n5988), .B(new_n5974), .Y(new_n5989));
  not_3  g05613(.A(new_n5974), .Y(new_n5990));
  nor_4  g05614(.A(new_n5987), .B(new_n5990), .Y(new_n5991));
  nor_4  g05615(.A(new_n5991), .B(new_n5989), .Y(new_n5992));
  not_3  g05616(.A(new_n5961), .Y(new_n5993));
  nor_4  g05617(.A(new_n5993), .B(new_n5956), .Y(new_n5994));
  not_3  g05618(.A(new_n5994), .Y(new_n5995));
  nand_4 g05619(.A(new_n5968), .B(new_n5995), .Y(new_n5996));
  nand_4 g05620(.A(new_n5996), .B(new_n5992), .Y(new_n5997));
  not_3  g05621(.A(new_n5997), .Y(new_n5998));
  nor_4  g05622(.A(new_n5996), .B(new_n5992), .Y(new_n5999));
  nor_4  g05623(.A(new_n5999), .B(new_n5998), .Y(new_n6000));
  xor_3  g05624(.A(new_n6000), .B(new_n5973), .Y(new_n6001));
  nand_4 g05625(.A(n8336), .B(n2522), .Y(new_n6002));
  nand_4 g05626(.A(n9189), .B(n8336), .Y(new_n6003));
  not_3  g05627(.A(new_n6003), .Y(new_n6004));
  nand_4 g05628(.A(n7946), .B(n6986), .Y(new_n6005));
  not_3  g05629(.A(new_n6005), .Y(new_n6006));
  nor_4  g05630(.A(new_n6006), .B(new_n6004), .Y(new_n6007));
  nand_4 g05631(.A(n10928), .B(n2024), .Y(new_n6008));
  not_3  g05632(.A(new_n6008), .Y(new_n6009));
  nor_4  g05633(.A(new_n6005), .B(new_n6003), .Y(new_n6010));
  nor_4  g05634(.A(new_n6010), .B(new_n6009), .Y(new_n6011));
  nor_4  g05635(.A(new_n6011), .B(new_n6007), .Y(new_n6012));
  xor_3  g05636(.A(new_n6012), .B(new_n6002), .Y(new_n6013));
  nand_4 g05637(.A(n6986), .B(n2024), .Y(new_n6014));
  nand_4 g05638(.A(n10928), .B(n9189), .Y(new_n6015));
  not_3  g05639(.A(new_n6015), .Y(new_n6016_1));
  nand_4 g05640(.A(n7946), .B(n2226), .Y(new_n6017));
  not_3  g05641(.A(new_n6017), .Y(new_n6018));
  nor_4  g05642(.A(new_n6018), .B(new_n6016_1), .Y(new_n6019));
  nor_4  g05643(.A(new_n6017), .B(new_n6015), .Y(new_n6020));
  nor_4  g05644(.A(new_n6020), .B(new_n6019), .Y(new_n6021));
  xor_3  g05645(.A(new_n6021), .B(new_n6014), .Y(new_n6022));
  xnor_3 g05646(.A(new_n6022), .B(new_n6013), .Y(new_n6023));
  not_3  g05647(.A(new_n6007), .Y(new_n6024));
  nor_4  g05648(.A(new_n6008), .B(new_n4569), .Y(new_n6025));
  nor_4  g05649(.A(new_n6025), .B(new_n6024), .Y(new_n6026));
  nor_4  g05650(.A(new_n6026), .B(new_n6010), .Y(new_n6027));
  nor_4  g05651(.A(new_n6027), .B(new_n6008), .Y(new_n6028));
  not_3  g05652(.A(new_n6028), .Y(new_n6029));
  nor_4  g05653(.A(new_n6029), .B(new_n6023), .Y(new_n6030));
  not_3  g05654(.A(new_n6030), .Y(new_n6031));
  nand_4 g05655(.A(n12145), .B(n8336), .Y(new_n6032));
  not_3  g05656(.A(new_n6032), .Y(new_n6033));
  nand_4 g05657(.A(n10928), .B(n2522), .Y(new_n6034));
  not_3  g05658(.A(new_n6014), .Y(new_n6035));
  nor_4  g05659(.A(new_n6020), .B(new_n6035), .Y(new_n6036));
  nor_4  g05660(.A(new_n6036), .B(new_n6019), .Y(new_n6037));
  xor_3  g05661(.A(new_n6037), .B(new_n6034), .Y(new_n6038_1));
  nand_4 g05662(.A(n2226), .B(n2024), .Y(new_n6039));
  not_3  g05663(.A(new_n6039), .Y(new_n6040));
  nand_4 g05664(.A(n9189), .B(n6986), .Y(new_n6041));
  nand_4 g05665(.A(n7946), .B(n1094), .Y(new_n6042));
  xnor_3 g05666(.A(new_n6042), .B(new_n6041), .Y(new_n6043));
  xor_3  g05667(.A(new_n6043), .B(new_n6040), .Y(new_n6044));
  xnor_3 g05668(.A(new_n6044), .B(new_n6038_1), .Y(new_n6045));
  not_3  g05669(.A(new_n6045), .Y(new_n6046));
  xor_3  g05670(.A(new_n6046), .B(new_n6033), .Y(new_n6047));
  not_3  g05671(.A(new_n6002), .Y(new_n6048));
  and_4  g05672(.A(new_n6012), .B(new_n6048), .Y(new_n6049));
  not_3  g05673(.A(new_n6049), .Y(new_n6050));
  nor_4  g05674(.A(new_n6022), .B(new_n6013), .Y(new_n6051));
  not_3  g05675(.A(new_n6051), .Y(new_n6052));
  nand_4 g05676(.A(new_n6052), .B(new_n6050), .Y(new_n6053));
  xnor_3 g05677(.A(new_n6053), .B(new_n6047), .Y(new_n6054));
  xnor_3 g05678(.A(new_n6054), .B(new_n6031), .Y(new_n6055));
  not_3  g05679(.A(new_n6023), .Y(new_n6056));
  xor_3  g05680(.A(new_n6028), .B(new_n6056), .Y(new_n6057));
  nand_4 g05681(.A(n7891), .B(n2558), .Y(new_n6058));
  nand_4 g05682(.A(n12069), .B(n5579), .Y(new_n6059));
  nand_4 g05683(.A(new_n6059), .B(new_n6058), .Y(new_n6060));
  not_3  g05684(.A(new_n6060), .Y(new_n6061));
  not_3  g05685(.A(new_n6058), .Y(new_n6062));
  not_3  g05686(.A(new_n6059), .Y(new_n6063));
  nand_4 g05687(.A(new_n6063), .B(new_n6062), .Y(new_n6064));
  not_3  g05688(.A(new_n6064), .Y(new_n6065));
  nor_4  g05689(.A(new_n6065), .B(new_n6061), .Y(new_n6066));
  nand_4 g05690(.A(n12391), .B(n2558), .Y(new_n6067));
  nand_4 g05691(.A(n12069), .B(n2498), .Y(new_n6068));
  nor_4  g05692(.A(new_n6068), .B(new_n6067), .Y(new_n6069));
  not_3  g05693(.A(new_n6069), .Y(new_n6070));
  nor_4  g05694(.A(new_n6070), .B(new_n6066), .Y(new_n6071));
  not_3  g05695(.A(new_n6071), .Y(new_n6072));
  nand_4 g05696(.A(n12069), .B(n521), .Y(new_n6073));
  nand_4 g05697(.A(n12391), .B(n2498), .Y(new_n6074));
  not_3  g05698(.A(new_n6074), .Y(new_n6075));
  nand_4 g05699(.A(new_n6075), .B(new_n6060), .Y(new_n6076));
  nand_4 g05700(.A(new_n6076), .B(new_n6064), .Y(new_n6077));
  not_3  g05701(.A(new_n6077), .Y(new_n6078));
  xnor_3 g05702(.A(new_n6078), .B(new_n6073), .Y(new_n6079));
  nand_4 g05703(.A(n7891), .B(n2498), .Y(new_n6080));
  not_3  g05704(.A(new_n6080), .Y(new_n6081));
  nand_4 g05705(.A(n12391), .B(n5579), .Y(new_n6082));
  not_3  g05706(.A(new_n6082), .Y(new_n6083));
  nand_4 g05707(.A(n7160), .B(n2558), .Y(new_n6084));
  not_3  g05708(.A(new_n6084), .Y(new_n6085));
  nor_4  g05709(.A(new_n6085), .B(new_n6083), .Y(new_n6086));
  nor_4  g05710(.A(new_n6084), .B(new_n6082), .Y(new_n6087));
  nor_4  g05711(.A(new_n6087), .B(new_n6086), .Y(new_n6088));
  xnor_3 g05712(.A(new_n6088), .B(new_n6081), .Y(new_n6089_1));
  xnor_3 g05713(.A(new_n6089_1), .B(new_n6079), .Y(new_n6090));
  nor_4  g05714(.A(new_n6090), .B(new_n6072), .Y(new_n6091));
  not_3  g05715(.A(new_n6090), .Y(new_n6092));
  nor_4  g05716(.A(new_n6092), .B(new_n6071), .Y(new_n6093));
  nor_4  g05717(.A(new_n6093), .B(new_n6091), .Y(new_n6094));
  nand_4 g05718(.A(n11222), .B(n806), .Y(new_n6095));
  not_3  g05719(.A(new_n6095), .Y(new_n6096));
  nand_4 g05720(.A(n11222), .B(n3342), .Y(new_n6097));
  nand_4 g05721(.A(n9763), .B(n5314), .Y(new_n6098));
  nand_4 g05722(.A(new_n6098), .B(new_n6097), .Y(new_n6099));
  not_3  g05723(.A(new_n6099), .Y(new_n6100));
  nand_4 g05724(.A(n11153), .B(n9111), .Y(new_n6101));
  not_3  g05725(.A(new_n6101), .Y(new_n6102));
  nor_4  g05726(.A(new_n6098), .B(new_n6097), .Y(new_n6103));
  nor_4  g05727(.A(new_n6103), .B(new_n6102), .Y(new_n6104));
  nor_4  g05728(.A(new_n6104), .B(new_n6100), .Y(new_n6105));
  nand_4 g05729(.A(new_n6105), .B(new_n6096), .Y(new_n6106));
  not_3  g05730(.A(new_n6106), .Y(new_n6107));
  nor_4  g05731(.A(new_n6105), .B(new_n6096), .Y(new_n6108));
  nor_4  g05732(.A(new_n6108), .B(new_n6107), .Y(new_n6109));
  nand_4 g05733(.A(n9111), .B(n5314), .Y(new_n6110));
  nand_4 g05734(.A(n11153), .B(n3342), .Y(new_n6111));
  nand_4 g05735(.A(n9763), .B(n996), .Y(new_n6112));
  xnor_3 g05736(.A(new_n6112), .B(new_n6111), .Y(new_n6113));
  xnor_3 g05737(.A(new_n6113), .B(new_n6110), .Y(new_n6114));
  not_3  g05738(.A(new_n6114), .Y(new_n6115));
  xnor_3 g05739(.A(new_n6115), .B(new_n6109), .Y(new_n6116));
  not_3  g05740(.A(new_n4570), .Y(new_n6117));
  nor_4  g05741(.A(new_n6101), .B(new_n6117), .Y(new_n6118));
  nor_4  g05742(.A(new_n6118), .B(new_n6099), .Y(new_n6119));
  nor_4  g05743(.A(new_n6119), .B(new_n6103), .Y(new_n6120));
  nor_4  g05744(.A(new_n6120), .B(new_n6101), .Y(new_n6121));
  not_3  g05745(.A(new_n6121), .Y(new_n6122));
  nor_4  g05746(.A(new_n6122), .B(new_n6116), .Y(new_n6123));
  not_3  g05747(.A(new_n6116), .Y(new_n6124));
  nor_4  g05748(.A(new_n6121), .B(new_n6124), .Y(new_n6125));
  nor_4  g05749(.A(new_n6125), .B(new_n6123), .Y(new_n6126_1));
  xnor_3 g05750(.A(new_n6126_1), .B(new_n6094), .Y(new_n6127));
  not_3  g05751(.A(new_n6127), .Y(new_n6128));
  nor_4  g05752(.A(new_n4571), .B(new_n4570), .Y(new_n6129));
  xnor_3 g05753(.A(new_n6068), .B(new_n6067), .Y(new_n6130));
  not_3  g05754(.A(new_n6130), .Y(new_n6131));
  nor_4  g05755(.A(new_n6131), .B(new_n6129), .Y(new_n6132));
  not_3  g05756(.A(new_n6132), .Y(new_n6133));
  not_3  g05757(.A(new_n6129), .Y(new_n6134));
  nor_4  g05758(.A(new_n6130), .B(new_n6134), .Y(new_n6135));
  nor_4  g05759(.A(new_n6135), .B(new_n6132), .Y(new_n6136));
  nand_4 g05760(.A(n11153), .B(n9763), .Y(new_n6137));
  nand_4 g05761(.A(n11222), .B(n9111), .Y(new_n6138));
  xnor_3 g05762(.A(new_n6138), .B(new_n6137), .Y(new_n6139));
  nand_4 g05763(.A(new_n6139), .B(new_n6136), .Y(new_n6140));
  nand_4 g05764(.A(new_n6140), .B(new_n6133), .Y(new_n6141));
  not_3  g05765(.A(new_n6141), .Y(new_n6142));
  not_3  g05766(.A(new_n6118), .Y(new_n6143));
  nor_4  g05767(.A(new_n6143), .B(new_n6100), .Y(new_n6144));
  not_3  g05768(.A(new_n6144), .Y(new_n6145));
  nand_4 g05769(.A(new_n6145), .B(new_n6120), .Y(new_n6146));
  not_3  g05770(.A(new_n6146), .Y(new_n6147));
  nor_4  g05771(.A(new_n6147), .B(new_n6142), .Y(new_n6148));
  xnor_3 g05772(.A(new_n6146), .B(new_n6141), .Y(new_n6149));
  not_3  g05773(.A(new_n4571), .Y(new_n6150));
  nor_4  g05774(.A(new_n6074), .B(new_n6150), .Y(new_n6151));
  not_3  g05775(.A(new_n6151), .Y(new_n6152));
  nor_4  g05776(.A(new_n6152), .B(new_n6060), .Y(new_n6153));
  not_3  g05777(.A(new_n6066), .Y(new_n6154));
  nor_4  g05778(.A(new_n6151), .B(new_n6154), .Y(new_n6155));
  nor_4  g05779(.A(new_n6155), .B(new_n6153), .Y(new_n6156));
  not_3  g05780(.A(new_n6156), .Y(new_n6157));
  nor_4  g05781(.A(new_n6157), .B(new_n6149), .Y(new_n6158));
  nor_4  g05782(.A(new_n6158), .B(new_n6148), .Y(new_n6159));
  not_3  g05783(.A(new_n6159), .Y(new_n6160));
  nor_4  g05784(.A(new_n6160), .B(new_n6128), .Y(new_n6161));
  nor_4  g05785(.A(new_n6159), .B(new_n6127), .Y(new_n6162));
  nor_4  g05786(.A(new_n6162), .B(new_n6161), .Y(new_n6163));
  not_3  g05787(.A(new_n6163), .Y(new_n6164));
  nand_4 g05788(.A(new_n6164), .B(new_n6057), .Y(new_n6165));
  xnor_3 g05789(.A(new_n6163), .B(new_n6057), .Y(new_n6166));
  xnor_3 g05790(.A(new_n6157), .B(new_n6149), .Y(new_n6167));
  not_3  g05791(.A(new_n6027), .Y(new_n6168));
  not_3  g05792(.A(new_n6025), .Y(new_n6169));
  nor_4  g05793(.A(new_n6169), .B(new_n6007), .Y(new_n6170));
  nor_4  g05794(.A(new_n6170), .B(new_n6168), .Y(new_n6171));
  nand_4 g05795(.A(new_n6171), .B(new_n6167), .Y(new_n6172));
  xnor_3 g05796(.A(new_n6171), .B(new_n6167), .Y(new_n6173));
  not_3  g05797(.A(new_n6173), .Y(new_n6174));
  xnor_3 g05798(.A(new_n6139), .B(new_n6136), .Y(new_n6175));
  not_3  g05799(.A(new_n6175), .Y(new_n6176));
  nand_4 g05800(.A(n10928), .B(n7946), .Y(new_n6177));
  nand_4 g05801(.A(n8336), .B(n2024), .Y(new_n6178));
  xor_3  g05802(.A(new_n6178), .B(new_n6177), .Y(new_n6179));
  not_3  g05803(.A(new_n6179), .Y(new_n6180));
  nor_4  g05804(.A(new_n6180), .B(new_n6176), .Y(new_n6181));
  nand_4 g05805(.A(new_n4572), .B(new_n4569), .Y(new_n6182));
  xnor_3 g05806(.A(new_n6179), .B(new_n6175), .Y(new_n6183));
  nor_4  g05807(.A(new_n6183), .B(new_n6182), .Y(new_n6184));
  nor_4  g05808(.A(new_n6184), .B(new_n6181), .Y(new_n6185));
  not_3  g05809(.A(new_n6185), .Y(new_n6186));
  nand_4 g05810(.A(new_n6186), .B(new_n6174), .Y(new_n6187));
  nand_4 g05811(.A(new_n6187), .B(new_n6172), .Y(new_n6188));
  nand_4 g05812(.A(new_n6188), .B(new_n6166), .Y(new_n6189));
  nand_4 g05813(.A(new_n6189), .B(new_n6165), .Y(new_n6190));
  xnor_3 g05814(.A(new_n6190), .B(new_n6055), .Y(new_n6191));
  nand_4 g05815(.A(n12069), .B(n6016), .Y(new_n6192_1));
  nand_4 g05816(.A(n12391), .B(n521), .Y(new_n6193));
  not_3  g05817(.A(new_n6193), .Y(new_n6194));
  nor_4  g05818(.A(new_n6087), .B(new_n6081), .Y(new_n6195));
  nor_4  g05819(.A(new_n6195), .B(new_n6086), .Y(new_n6196));
  xnor_3 g05820(.A(new_n6196), .B(new_n6194), .Y(new_n6197));
  nand_4 g05821(.A(n7160), .B(n2498), .Y(new_n6198));
  nand_4 g05822(.A(n7891), .B(n5579), .Y(new_n6199));
  nand_4 g05823(.A(n4828), .B(n2558), .Y(new_n6200));
  xnor_3 g05824(.A(new_n6200), .B(new_n6199), .Y(new_n6201));
  not_3  g05825(.A(new_n6201), .Y(new_n6202));
  nor_4  g05826(.A(new_n6202), .B(new_n6198), .Y(new_n6203));
  not_3  g05827(.A(new_n6198), .Y(new_n6204));
  nor_4  g05828(.A(new_n6201), .B(new_n6204), .Y(new_n6205));
  nor_4  g05829(.A(new_n6205), .B(new_n6203), .Y(new_n6206));
  xnor_3 g05830(.A(new_n6206), .B(new_n6197), .Y(new_n6207));
  xnor_3 g05831(.A(new_n6207), .B(new_n6192_1), .Y(new_n6208));
  nor_4  g05832(.A(new_n6078), .B(new_n6073), .Y(new_n6209));
  nor_4  g05833(.A(new_n6089_1), .B(new_n6079), .Y(new_n6210));
  nor_4  g05834(.A(new_n6210), .B(new_n6209), .Y(new_n6211));
  xnor_3 g05835(.A(new_n6211), .B(new_n6208), .Y(new_n6212));
  not_3  g05836(.A(new_n6212), .Y(new_n6213));
  xor_3  g05837(.A(new_n6213), .B(new_n6091), .Y(new_n6214));
  nand_4 g05838(.A(n11222), .B(n7270), .Y(new_n6215));
  nand_4 g05839(.A(n11153), .B(n806), .Y(new_n6216));
  not_3  g05840(.A(new_n6216), .Y(new_n6217));
  not_3  g05841(.A(new_n6111), .Y(new_n6218));
  not_3  g05842(.A(new_n6112), .Y(new_n6219));
  nor_4  g05843(.A(new_n6219), .B(new_n6218), .Y(new_n6220));
  not_3  g05844(.A(new_n6110), .Y(new_n6221));
  nor_4  g05845(.A(new_n6112), .B(new_n6111), .Y(new_n6222));
  nor_4  g05846(.A(new_n6222), .B(new_n6221), .Y(new_n6223));
  nor_4  g05847(.A(new_n6223), .B(new_n6220), .Y(new_n6224));
  xnor_3 g05848(.A(new_n6224), .B(new_n6217), .Y(new_n6225));
  nand_4 g05849(.A(n9111), .B(n996), .Y(new_n6226));
  not_3  g05850(.A(new_n6226), .Y(new_n6227));
  nand_4 g05851(.A(n5314), .B(n3342), .Y(new_n6228));
  not_3  g05852(.A(new_n6228), .Y(new_n6229));
  nand_4 g05853(.A(n9763), .B(n5767), .Y(new_n6230));
  not_3  g05854(.A(new_n6230), .Y(new_n6231));
  nor_4  g05855(.A(new_n6231), .B(new_n6229), .Y(new_n6232));
  nor_4  g05856(.A(new_n6230), .B(new_n6228), .Y(new_n6233));
  nor_4  g05857(.A(new_n6233), .B(new_n6232), .Y(new_n6234));
  xnor_3 g05858(.A(new_n6234), .B(new_n6227), .Y(new_n6235));
  xnor_3 g05859(.A(new_n6235), .B(new_n6225), .Y(new_n6236));
  nor_4  g05860(.A(new_n6236), .B(new_n6215), .Y(new_n6237));
  not_3  g05861(.A(new_n6215), .Y(new_n6238));
  not_3  g05862(.A(new_n6236), .Y(new_n6239));
  nor_4  g05863(.A(new_n6239), .B(new_n6238), .Y(new_n6240));
  nor_4  g05864(.A(new_n6240), .B(new_n6237), .Y(new_n6241));
  nand_4 g05865(.A(new_n6115), .B(new_n6109), .Y(new_n6242));
  nand_4 g05866(.A(new_n6242), .B(new_n6106), .Y(new_n6243));
  xnor_3 g05867(.A(new_n6243), .B(new_n6241), .Y(new_n6244));
  not_3  g05868(.A(new_n6244), .Y(new_n6245));
  nor_4  g05869(.A(new_n6245), .B(new_n6123), .Y(new_n6246));
  not_3  g05870(.A(new_n6123), .Y(new_n6247));
  nor_4  g05871(.A(new_n6244), .B(new_n6247), .Y(new_n6248));
  nor_4  g05872(.A(new_n6248), .B(new_n6246), .Y(new_n6249));
  xnor_3 g05873(.A(new_n6249), .B(new_n6214), .Y(new_n6250));
  nor_4  g05874(.A(new_n6126_1), .B(new_n6094), .Y(new_n6251));
  nor_4  g05875(.A(new_n6162), .B(new_n6251), .Y(new_n6252));
  xnor_3 g05876(.A(new_n6252), .B(new_n6250), .Y(new_n6253));
  xnor_3 g05877(.A(new_n6253), .B(new_n6191), .Y(new_n6254_1));
  xnor_3 g05878(.A(new_n6254_1), .B(new_n6001), .Y(new_n6255));
  not_3  g05879(.A(new_n6255), .Y(new_n6256));
  xor_3  g05880(.A(new_n5971), .B(new_n5955), .Y(new_n6257));
  not_3  g05881(.A(new_n6257), .Y(new_n6258));
  xnor_3 g05882(.A(new_n6188), .B(new_n6166), .Y(new_n6259));
  nand_4 g05883(.A(new_n6259), .B(new_n6258), .Y(new_n6260));
  xnor_3 g05884(.A(new_n6185), .B(new_n6173), .Y(new_n6261));
  not_3  g05885(.A(new_n6261), .Y(new_n6262));
  not_3  g05886(.A(new_n5950), .Y(new_n6263));
  nor_4  g05887(.A(new_n5958), .B(new_n4567), .Y(new_n6264));
  not_3  g05888(.A(new_n6264), .Y(new_n6265));
  nand_4 g05889(.A(new_n6265), .B(new_n6263), .Y(new_n6266));
  nand_4 g05890(.A(new_n6264), .B(new_n5946), .Y(new_n6267));
  nand_4 g05891(.A(new_n6267), .B(new_n6266), .Y(new_n6268));
  not_3  g05892(.A(new_n6268), .Y(new_n6269));
  nor_4  g05893(.A(new_n6269), .B(new_n6262), .Y(new_n6270));
  not_3  g05894(.A(new_n6270), .Y(new_n6271));
  xor_3  g05895(.A(new_n6269), .B(new_n6262), .Y(new_n6272));
  nand_4 g05896(.A(new_n4573), .B(new_n4567), .Y(new_n6273_1));
  xor_3  g05897(.A(new_n5952), .B(new_n5951), .Y(new_n6274));
  not_3  g05898(.A(new_n6274), .Y(new_n6275));
  nand_4 g05899(.A(new_n6275), .B(new_n6273_1), .Y(new_n6276));
  not_3  g05900(.A(new_n6183), .Y(new_n6277));
  xor_3  g05901(.A(new_n6277), .B(new_n6182), .Y(new_n6278));
  not_3  g05902(.A(new_n6273_1), .Y(new_n6279));
  xor_3  g05903(.A(new_n6274), .B(new_n6279), .Y(new_n6280));
  nand_4 g05904(.A(new_n6280), .B(new_n6278), .Y(new_n6281));
  nand_4 g05905(.A(new_n6281), .B(new_n6276), .Y(new_n6282));
  nand_4 g05906(.A(new_n6282), .B(new_n6272), .Y(new_n6283));
  nand_4 g05907(.A(new_n6283), .B(new_n6271), .Y(new_n6284));
  xnor_3 g05908(.A(new_n6259), .B(new_n6257), .Y(new_n6285));
  nand_4 g05909(.A(new_n6285), .B(new_n6284), .Y(new_n6286));
  nand_4 g05910(.A(new_n6286), .B(new_n6260), .Y(new_n6287));
  xor_3  g05911(.A(new_n6287), .B(new_n6256), .Y(n1658));
  nand_4 g05912(.A(n7862), .B(n4634), .Y(new_n6289));
  nand_4 g05913(.A(n10223), .B(n7862), .Y(new_n6290));
  not_3  g05914(.A(new_n6290), .Y(new_n6291));
  nand_4 g05915(.A(n7265), .B(n3172), .Y(new_n6292));
  not_3  g05916(.A(new_n6292), .Y(new_n6293));
  nor_4  g05917(.A(new_n6293), .B(new_n6291), .Y(new_n6294_1));
  nor_4  g05918(.A(new_n6292), .B(new_n6290), .Y(new_n6295));
  nand_4 g05919(.A(n2879), .B(n1333), .Y(new_n6296));
  not_3  g05920(.A(new_n6296), .Y(new_n6297));
  nor_4  g05921(.A(new_n6297), .B(new_n6295), .Y(new_n6298));
  nor_4  g05922(.A(new_n6298), .B(new_n6294_1), .Y(new_n6299));
  xor_3  g05923(.A(new_n6299), .B(new_n6289), .Y(new_n6300));
  nand_4 g05924(.A(n3172), .B(n2879), .Y(new_n6301));
  nand_4 g05925(.A(n10223), .B(n1333), .Y(new_n6302));
  not_3  g05926(.A(new_n6302), .Y(new_n6303));
  nand_4 g05927(.A(n11757), .B(n7265), .Y(new_n6304));
  not_3  g05928(.A(new_n6304), .Y(new_n6305));
  nor_4  g05929(.A(new_n6305), .B(new_n6303), .Y(new_n6306));
  nor_4  g05930(.A(new_n6304), .B(new_n6302), .Y(new_n6307));
  nor_4  g05931(.A(new_n6307), .B(new_n6306), .Y(new_n6308));
  xor_3  g05932(.A(new_n6308), .B(new_n6301), .Y(new_n6309));
  xnor_3 g05933(.A(new_n6309), .B(new_n6300), .Y(new_n6310));
  not_3  g05934(.A(new_n6310), .Y(new_n6311));
  nand_4 g05935(.A(n7862), .B(n7265), .Y(new_n6312));
  not_3  g05936(.A(new_n6312), .Y(new_n6313));
  nor_4  g05937(.A(new_n6313), .B(new_n6296), .Y(new_n6314));
  nor_4  g05938(.A(new_n6295), .B(new_n6294_1), .Y(new_n6315));
  nor_4  g05939(.A(new_n6315), .B(new_n6314), .Y(new_n6316));
  not_3  g05940(.A(new_n6316), .Y(new_n6317));
  nor_4  g05941(.A(new_n6317), .B(new_n6296), .Y(new_n6318));
  xor_3  g05942(.A(new_n6318), .B(new_n6311), .Y(new_n6319));
  nand_4 g05943(.A(n6877), .B(n2522), .Y(new_n6320));
  nand_4 g05944(.A(n2464), .B(n2024), .Y(new_n6321));
  nand_4 g05945(.A(n9400), .B(n9189), .Y(new_n6322));
  nand_4 g05946(.A(n11311), .B(n7946), .Y(new_n6323));
  xnor_3 g05947(.A(new_n6323), .B(new_n6322), .Y(new_n6324));
  not_3  g05948(.A(new_n6324), .Y(new_n6325));
  nor_4  g05949(.A(new_n6325), .B(new_n6321), .Y(new_n6326));
  not_3  g05950(.A(new_n6321), .Y(new_n6327));
  nor_4  g05951(.A(new_n6324), .B(new_n6327), .Y(new_n6328));
  nor_4  g05952(.A(new_n6328), .B(new_n6326), .Y(new_n6329));
  xnor_3 g05953(.A(new_n6329), .B(new_n6320), .Y(new_n6330));
  nand_4 g05954(.A(n9189), .B(n6877), .Y(new_n6331));
  not_3  g05955(.A(new_n6331), .Y(new_n6332));
  nand_4 g05956(.A(n7946), .B(n2464), .Y(new_n6333));
  not_3  g05957(.A(new_n6333), .Y(new_n6334));
  nor_4  g05958(.A(new_n6334), .B(new_n6332), .Y(new_n6335));
  nor_4  g05959(.A(new_n6333), .B(new_n6331), .Y(new_n6336));
  nand_4 g05960(.A(n9400), .B(n2024), .Y(new_n6337));
  not_3  g05961(.A(new_n6337), .Y(new_n6338));
  nor_4  g05962(.A(new_n6338), .B(new_n6336), .Y(new_n6339));
  nor_4  g05963(.A(new_n6339), .B(new_n6335), .Y(new_n6340));
  not_3  g05964(.A(new_n6340), .Y(new_n6341));
  nor_4  g05965(.A(new_n6341), .B(new_n6330), .Y(new_n6342));
  not_3  g05966(.A(new_n6330), .Y(new_n6343));
  nor_4  g05967(.A(new_n6340), .B(new_n6343), .Y(new_n6344));
  nor_4  g05968(.A(new_n6344), .B(new_n6342), .Y(new_n6345));
  not_3  g05969(.A(new_n6345), .Y(new_n6346));
  nand_4 g05970(.A(n7946), .B(n6877), .Y(new_n6347));
  not_3  g05971(.A(new_n6347), .Y(new_n6348));
  nor_4  g05972(.A(new_n6348), .B(new_n6337), .Y(new_n6349));
  nor_4  g05973(.A(new_n6336), .B(new_n6335), .Y(new_n6350));
  nor_4  g05974(.A(new_n6350), .B(new_n6349), .Y(new_n6351));
  not_3  g05975(.A(new_n6351), .Y(new_n6352));
  nor_4  g05976(.A(new_n6352), .B(new_n6337), .Y(new_n6353));
  not_3  g05977(.A(new_n6353), .Y(new_n6354));
  nor_4  g05978(.A(new_n6354), .B(new_n6346), .Y(new_n6355));
  nor_4  g05979(.A(new_n6353), .B(new_n6345), .Y(new_n6356));
  nor_4  g05980(.A(new_n6356), .B(new_n6355), .Y(new_n6357));
  not_3  g05981(.A(new_n6357), .Y(new_n6358_1));
  nand_4 g05982(.A(n4805), .B(n2558), .Y(new_n6359_1));
  nand_4 g05983(.A(n9763), .B(n7236), .Y(new_n6360));
  xnor_3 g05984(.A(new_n6360), .B(new_n6359_1), .Y(new_n6361));
  nor_4  g05985(.A(new_n6361), .B(new_n6347), .Y(new_n6362));
  not_3  g05986(.A(new_n6362), .Y(new_n6363));
  nand_4 g05987(.A(n9400), .B(n7946), .Y(new_n6364));
  nand_4 g05988(.A(n6877), .B(n2024), .Y(new_n6365));
  not_3  g05989(.A(new_n6365), .Y(new_n6366));
  xnor_3 g05990(.A(new_n6366), .B(new_n6364), .Y(new_n6367));
  not_3  g05991(.A(new_n6367), .Y(new_n6368));
  nor_4  g05992(.A(new_n6368), .B(new_n6363), .Y(new_n6369));
  not_3  g05993(.A(new_n6369), .Y(new_n6370));
  nor_4  g05994(.A(new_n6360), .B(new_n6359_1), .Y(new_n6371));
  nand_4 g05995(.A(n9111), .B(n7236), .Y(new_n6372));
  nand_4 g05996(.A(n9763), .B(n3992), .Y(new_n6373));
  xnor_3 g05997(.A(new_n6373), .B(new_n6372), .Y(new_n6374));
  xnor_3 g05998(.A(new_n6374), .B(new_n6371), .Y(new_n6375));
  nand_4 g05999(.A(n4805), .B(n2498), .Y(new_n6376));
  nand_4 g06000(.A(n11478), .B(n2558), .Y(new_n6377));
  not_3  g06001(.A(new_n6377), .Y(new_n6378));
  xnor_3 g06002(.A(new_n6378), .B(new_n6376), .Y(new_n6379));
  not_3  g06003(.A(new_n6379), .Y(new_n6380));
  xnor_3 g06004(.A(new_n6380), .B(new_n6375), .Y(new_n6381));
  nor_4  g06005(.A(new_n6367), .B(new_n6362), .Y(new_n6382));
  nor_4  g06006(.A(new_n6382), .B(new_n6369), .Y(new_n6383));
  nand_4 g06007(.A(new_n6383), .B(new_n6381), .Y(new_n6384));
  nand_4 g06008(.A(new_n6384), .B(new_n6370), .Y(new_n6385));
  not_3  g06009(.A(new_n6335), .Y(new_n6386));
  nand_4 g06010(.A(new_n6349), .B(new_n6386), .Y(new_n6387));
  nand_4 g06011(.A(new_n6387), .B(new_n6352), .Y(new_n6388));
  not_3  g06012(.A(new_n6388), .Y(new_n6389));
  nor_4  g06013(.A(new_n6389), .B(new_n6385), .Y(new_n6390));
  not_3  g06014(.A(new_n6390), .Y(new_n6391));
  not_3  g06015(.A(new_n6374), .Y(new_n6392));
  nor_4  g06016(.A(new_n6392), .B(new_n6371), .Y(new_n6393));
  not_3  g06017(.A(new_n6393), .Y(new_n6394));
  nand_4 g06018(.A(new_n6380), .B(new_n6375), .Y(new_n6395));
  nand_4 g06019(.A(new_n6395), .B(new_n6394), .Y(new_n6396));
  not_3  g06020(.A(new_n6359_1), .Y(new_n6397));
  nand_4 g06021(.A(n11478), .B(n2498), .Y(new_n6398));
  nor_4  g06022(.A(new_n6398), .B(new_n6397), .Y(new_n6399));
  not_3  g06023(.A(new_n6399), .Y(new_n6400));
  nand_4 g06024(.A(n5283), .B(n2558), .Y(new_n6401));
  nand_4 g06025(.A(n5579), .B(n4805), .Y(new_n6402));
  nand_4 g06026(.A(new_n6402), .B(new_n6401), .Y(new_n6403));
  not_3  g06027(.A(new_n6403), .Y(new_n6404));
  nor_4  g06028(.A(new_n6404), .B(new_n6400), .Y(new_n6405));
  not_3  g06029(.A(new_n6405), .Y(new_n6406));
  not_3  g06030(.A(new_n6401), .Y(new_n6407));
  not_3  g06031(.A(new_n6402), .Y(new_n6408));
  nand_4 g06032(.A(new_n6408), .B(new_n6407), .Y(new_n6409));
  not_3  g06033(.A(new_n6409), .Y(new_n6410));
  nor_4  g06034(.A(new_n6403), .B(new_n6399), .Y(new_n6411));
  nor_4  g06035(.A(new_n6411), .B(new_n6410), .Y(new_n6412));
  nand_4 g06036(.A(new_n6412), .B(new_n6406), .Y(new_n6413));
  xnor_3 g06037(.A(new_n6413), .B(new_n6396), .Y(new_n6414));
  not_3  g06038(.A(new_n6360), .Y(new_n6415));
  nand_4 g06039(.A(n9111), .B(n3992), .Y(new_n6416));
  nor_4  g06040(.A(new_n6416), .B(new_n6415), .Y(new_n6417));
  not_3  g06041(.A(new_n6417), .Y(new_n6418));
  nand_4 g06042(.A(n9763), .B(n8384), .Y(new_n6419));
  nand_4 g06043(.A(n7236), .B(n3342), .Y(new_n6420));
  nand_4 g06044(.A(new_n6420), .B(new_n6419), .Y(new_n6421));
  nor_4  g06045(.A(new_n6421), .B(new_n6418), .Y(new_n6422));
  not_3  g06046(.A(new_n6421), .Y(new_n6423));
  not_3  g06047(.A(new_n6419), .Y(new_n6424));
  not_3  g06048(.A(new_n6420), .Y(new_n6425));
  nand_4 g06049(.A(new_n6425), .B(new_n6424), .Y(new_n6426));
  not_3  g06050(.A(new_n6426), .Y(new_n6427));
  nor_4  g06051(.A(new_n6427), .B(new_n6423), .Y(new_n6428));
  not_3  g06052(.A(new_n6428), .Y(new_n6429_1));
  nor_4  g06053(.A(new_n6429_1), .B(new_n6417), .Y(new_n6430));
  nor_4  g06054(.A(new_n6430), .B(new_n6422), .Y(new_n6431_1));
  not_3  g06055(.A(new_n6431_1), .Y(new_n6432));
  nor_4  g06056(.A(new_n6432), .B(new_n6414), .Y(new_n6433));
  not_3  g06057(.A(new_n6414), .Y(new_n6434));
  nor_4  g06058(.A(new_n6431_1), .B(new_n6434), .Y(new_n6435));
  nor_4  g06059(.A(new_n6435), .B(new_n6433), .Y(new_n6436));
  not_3  g06060(.A(new_n6385), .Y(new_n6437));
  nor_4  g06061(.A(new_n6388), .B(new_n6437), .Y(new_n6438));
  nor_4  g06062(.A(new_n6438), .B(new_n6390), .Y(new_n6439));
  nand_4 g06063(.A(new_n6439), .B(new_n6436), .Y(new_n6440));
  nand_4 g06064(.A(new_n6440), .B(new_n6391), .Y(new_n6441_1));
  nor_4  g06065(.A(new_n6441_1), .B(new_n6358_1), .Y(new_n6442));
  not_3  g06066(.A(new_n6441_1), .Y(new_n6443));
  nor_4  g06067(.A(new_n6443), .B(new_n6357), .Y(new_n6444));
  nor_4  g06068(.A(new_n6444), .B(new_n6442), .Y(new_n6445_1));
  nand_4 g06069(.A(n4805), .B(n521), .Y(new_n6446));
  not_3  g06070(.A(new_n6398), .Y(new_n6447));
  nand_4 g06071(.A(new_n6403), .B(new_n6447), .Y(new_n6448));
  nand_4 g06072(.A(new_n6448), .B(new_n6409), .Y(new_n6449));
  not_3  g06073(.A(new_n6449), .Y(new_n6450));
  nor_4  g06074(.A(new_n6450), .B(new_n6446), .Y(new_n6451));
  not_3  g06075(.A(new_n6446), .Y(new_n6452));
  nor_4  g06076(.A(new_n6449), .B(new_n6452), .Y(new_n6453));
  nor_4  g06077(.A(new_n6453), .B(new_n6451), .Y(new_n6454));
  nand_4 g06078(.A(n5283), .B(n2498), .Y(new_n6455));
  nand_4 g06079(.A(n2558), .B(n137), .Y(new_n6456));
  nand_4 g06080(.A(n11478), .B(n5579), .Y(new_n6457));
  xnor_3 g06081(.A(new_n6457), .B(new_n6456), .Y(new_n6458));
  xnor_3 g06082(.A(new_n6458), .B(new_n6455), .Y(new_n6459));
  not_3  g06083(.A(new_n6459), .Y(new_n6460));
  xnor_3 g06084(.A(new_n6460), .B(new_n6454), .Y(new_n6461));
  not_3  g06085(.A(new_n6461), .Y(new_n6462));
  nor_4  g06086(.A(new_n6412), .B(new_n6398), .Y(new_n6463));
  nor_4  g06087(.A(new_n6463), .B(new_n6462), .Y(new_n6464));
  not_3  g06088(.A(new_n6463), .Y(new_n6465));
  nor_4  g06089(.A(new_n6465), .B(new_n6461), .Y(new_n6466));
  nor_4  g06090(.A(new_n6466), .B(new_n6464), .Y(new_n6467));
  nand_4 g06091(.A(n7236), .B(n806), .Y(new_n6468));
  not_3  g06092(.A(new_n6416), .Y(new_n6469));
  nand_4 g06093(.A(new_n6421), .B(new_n6469), .Y(new_n6470));
  nand_4 g06094(.A(new_n6470), .B(new_n6426), .Y(new_n6471));
  not_3  g06095(.A(new_n6471), .Y(new_n6472));
  nor_4  g06096(.A(new_n6472), .B(new_n6468), .Y(new_n6473));
  not_3  g06097(.A(new_n6468), .Y(new_n6474));
  nor_4  g06098(.A(new_n6471), .B(new_n6474), .Y(new_n6475));
  nor_4  g06099(.A(new_n6475), .B(new_n6473), .Y(new_n6476));
  nand_4 g06100(.A(n9111), .B(n8384), .Y(new_n6477));
  nand_4 g06101(.A(n9763), .B(n6358), .Y(new_n6478));
  nand_4 g06102(.A(n3992), .B(n3342), .Y(new_n6479));
  xnor_3 g06103(.A(new_n6479), .B(new_n6478), .Y(new_n6480));
  xnor_3 g06104(.A(new_n6480), .B(new_n6477), .Y(new_n6481));
  not_3  g06105(.A(new_n6481), .Y(new_n6482));
  xnor_3 g06106(.A(new_n6482), .B(new_n6476), .Y(new_n6483));
  not_3  g06107(.A(new_n6483), .Y(new_n6484));
  nor_4  g06108(.A(new_n6373), .B(new_n6372), .Y(new_n6485));
  not_3  g06109(.A(new_n6485), .Y(new_n6486));
  nor_4  g06110(.A(new_n6428), .B(new_n6486), .Y(new_n6487));
  nor_4  g06111(.A(new_n6487), .B(new_n6484), .Y(new_n6488));
  not_3  g06112(.A(new_n6487), .Y(new_n6489));
  nor_4  g06113(.A(new_n6489), .B(new_n6483), .Y(new_n6490));
  nor_4  g06114(.A(new_n6490), .B(new_n6488), .Y(new_n6491));
  xnor_3 g06115(.A(new_n6491), .B(new_n6467), .Y(new_n6492));
  and_4  g06116(.A(new_n6413), .B(new_n6396), .Y(new_n6493));
  nor_4  g06117(.A(new_n6433), .B(new_n6493), .Y(new_n6494));
  xnor_3 g06118(.A(new_n6494), .B(new_n6492), .Y(new_n6495));
  nor_4  g06119(.A(new_n6495), .B(new_n6445_1), .Y(new_n6496));
  nand_4 g06120(.A(new_n6495), .B(new_n6445_1), .Y(new_n6497));
  not_3  g06121(.A(new_n6497), .Y(new_n6498));
  nor_4  g06122(.A(new_n6498), .B(new_n6496), .Y(new_n6499));
  nor_4  g06123(.A(new_n6499), .B(new_n6319), .Y(new_n6500));
  not_3  g06124(.A(new_n6500), .Y(new_n6501));
  nand_4 g06125(.A(new_n6499), .B(new_n6319), .Y(new_n6502));
  nand_4 g06126(.A(new_n6502), .B(new_n6501), .Y(new_n6503));
  not_3  g06127(.A(new_n6440), .Y(new_n6504));
  nor_4  g06128(.A(new_n6439), .B(new_n6436), .Y(new_n6505));
  nor_4  g06129(.A(new_n6505), .B(new_n6504), .Y(new_n6506));
  not_3  g06130(.A(new_n6314), .Y(new_n6507));
  nor_4  g06131(.A(new_n6507), .B(new_n6294_1), .Y(new_n6508));
  or_4   g06132(.A(new_n6508), .B(new_n6316), .Y(new_n6509));
  nor_4  g06133(.A(new_n6509), .B(new_n6506), .Y(new_n6510));
  xor_3  g06134(.A(new_n6361), .B(new_n6347), .Y(new_n6511));
  nand_4 g06135(.A(new_n6511), .B(new_n6313), .Y(new_n6512));
  not_3  g06136(.A(new_n6512), .Y(new_n6513));
  nand_4 g06137(.A(n7265), .B(n1333), .Y(new_n6514));
  nand_4 g06138(.A(n7862), .B(n2879), .Y(new_n6515));
  xor_3  g06139(.A(new_n6515), .B(new_n6514), .Y(new_n6516));
  nor_4  g06140(.A(new_n6516), .B(new_n6513), .Y(new_n6517));
  not_3  g06141(.A(new_n6517), .Y(new_n6518));
  not_3  g06142(.A(new_n6381), .Y(new_n6519));
  xor_3  g06143(.A(new_n6383), .B(new_n6519), .Y(new_n6520));
  xor_3  g06144(.A(new_n6516), .B(new_n6513), .Y(new_n6521));
  nand_4 g06145(.A(new_n6521), .B(new_n6520), .Y(new_n6522));
  nand_4 g06146(.A(new_n6522), .B(new_n6518), .Y(new_n6523));
  xnor_3 g06147(.A(new_n6509), .B(new_n6506), .Y(new_n6524));
  nor_4  g06148(.A(new_n6524), .B(new_n6523), .Y(new_n6525));
  nor_4  g06149(.A(new_n6525), .B(new_n6510), .Y(new_n6526));
  xor_3  g06150(.A(new_n6526), .B(new_n6503), .Y(n1847));
  nand_4 g06151(.A(n5305), .B(n1798), .Y(new_n6528));
  nand_4 g06152(.A(n8759), .B(n6703), .Y(new_n6529));
  not_3  g06153(.A(new_n6529), .Y(new_n6530));
  nand_4 g06154(.A(n5645), .B(n5331), .Y(new_n6531));
  nand_4 g06155(.A(n11876), .B(n7965), .Y(new_n6532));
  xor_3  g06156(.A(new_n6532), .B(new_n6531), .Y(new_n6533));
  not_3  g06157(.A(new_n6533), .Y(new_n6534));
  xor_3  g06158(.A(new_n6534), .B(new_n6530), .Y(new_n6535));
  nor_4  g06159(.A(new_n6535), .B(new_n6528), .Y(new_n6536));
  nand_4 g06160(.A(n5305), .B(n3932), .Y(new_n6537));
  nand_4 g06161(.A(n5964), .B(n1798), .Y(new_n6538));
  xor_3  g06162(.A(new_n6538), .B(new_n6537), .Y(new_n6539));
  xor_3  g06163(.A(new_n6539), .B(new_n6536), .Y(new_n6540));
  nor_4  g06164(.A(new_n6534), .B(new_n6529), .Y(new_n6541));
  nand_4 g06165(.A(n9640), .B(n8759), .Y(new_n6542));
  nand_4 g06166(.A(n6776), .B(n6703), .Y(new_n6543));
  xor_3  g06167(.A(new_n6543), .B(new_n6542), .Y(new_n6544));
  xnor_3 g06168(.A(new_n6544), .B(new_n6541), .Y(new_n6545));
  nor_4  g06169(.A(new_n6532), .B(new_n6531), .Y(new_n6546));
  not_3  g06170(.A(new_n6546), .Y(new_n6547));
  nand_4 g06171(.A(n10898), .B(n7965), .Y(new_n6548));
  nand_4 g06172(.A(n11876), .B(n7388), .Y(new_n6549));
  xnor_3 g06173(.A(new_n6549), .B(new_n6548), .Y(new_n6550));
  nor_4  g06174(.A(new_n6550), .B(new_n6547), .Y(new_n6551));
  not_3  g06175(.A(new_n6550), .Y(new_n6552));
  nor_4  g06176(.A(new_n6552), .B(new_n6546), .Y(new_n6553));
  nor_4  g06177(.A(new_n6553), .B(new_n6551), .Y(new_n6554));
  nand_4 g06178(.A(n5331), .B(n1067), .Y(new_n6555));
  nand_4 g06179(.A(n8476), .B(n5645), .Y(new_n6556));
  xor_3  g06180(.A(new_n6556), .B(new_n6555), .Y(new_n6557));
  xnor_3 g06181(.A(new_n6557), .B(new_n6554), .Y(new_n6558));
  nor_4  g06182(.A(new_n6558), .B(new_n6545), .Y(new_n6559));
  and_4  g06183(.A(new_n6558), .B(new_n6545), .Y(new_n6560));
  nor_4  g06184(.A(new_n6560), .B(new_n6559), .Y(new_n6561));
  xor_3  g06185(.A(new_n6561), .B(new_n6540), .Y(n2096));
  xor_3  g06186(.A(new_n3840), .B(new_n3801), .Y(n2131));
  nand_4 g06187(.A(n7456), .B(n2564), .Y(new_n6564));
  not_3  g06188(.A(new_n6564), .Y(new_n6565));
  not_3  g06189(.A(new_n4009), .Y(new_n6566));
  nor_4  g06190(.A(new_n4015), .B(new_n6566), .Y(new_n6567));
  nor_4  g06191(.A(new_n6567), .B(new_n4014), .Y(new_n6568));
  nand_4 g06192(.A(new_n6568), .B(new_n6565), .Y(new_n6569));
  xnor_3 g06193(.A(new_n6568), .B(new_n6564), .Y(new_n6570));
  nand_4 g06194(.A(n6770), .B(n3932), .Y(new_n6571));
  nand_4 g06195(.A(n12591), .B(n4189), .Y(new_n6572));
  not_3  g06196(.A(new_n6572), .Y(new_n6573));
  nand_4 g06197(.A(n9920), .B(n1798), .Y(new_n6574));
  not_3  g06198(.A(new_n6574), .Y(new_n6575));
  nor_4  g06199(.A(new_n6575), .B(new_n6573), .Y(new_n6576));
  nor_4  g06200(.A(new_n6574), .B(new_n6572), .Y(new_n6577));
  nor_4  g06201(.A(new_n6577), .B(new_n6576), .Y(new_n6578_1));
  xnor_3 g06202(.A(new_n6578_1), .B(new_n6571), .Y(new_n6579));
  nand_4 g06203(.A(new_n6579), .B(new_n6570), .Y(new_n6580));
  nand_4 g06204(.A(new_n6580), .B(new_n6569), .Y(new_n6581));
  nand_4 g06205(.A(n11662), .B(n2564), .Y(new_n6582));
  nand_4 g06206(.A(n7456), .B(n4189), .Y(new_n6583));
  xor_3  g06207(.A(new_n6583), .B(new_n6582), .Y(new_n6584));
  xnor_3 g06208(.A(new_n6584), .B(new_n6581), .Y(new_n6585));
  nand_4 g06209(.A(n12591), .B(n6770), .Y(new_n6586));
  not_3  g06210(.A(new_n6586), .Y(new_n6587));
  nand_4 g06211(.A(n3627), .B(n1798), .Y(new_n6588));
  nand_4 g06212(.A(n9920), .B(n3932), .Y(new_n6589));
  xor_3  g06213(.A(new_n6589), .B(new_n6588), .Y(new_n6590));
  xnor_3 g06214(.A(new_n6590), .B(new_n6587), .Y(new_n6591));
  not_3  g06215(.A(new_n6591), .Y(new_n6592));
  not_3  g06216(.A(new_n6571), .Y(new_n6593));
  nor_4  g06217(.A(new_n6577), .B(new_n6593), .Y(new_n6594));
  nor_4  g06218(.A(new_n6594), .B(new_n6576), .Y(new_n6595));
  not_3  g06219(.A(new_n6595), .Y(new_n6596));
  xor_3  g06220(.A(new_n6596), .B(new_n6592), .Y(new_n6597));
  xnor_3 g06221(.A(new_n6597), .B(new_n6585), .Y(new_n6598));
  not_3  g06222(.A(new_n6598), .Y(new_n6599));
  nand_4 g06223(.A(n11662), .B(n6687), .Y(new_n6600));
  not_3  g06224(.A(new_n6600), .Y(new_n6601));
  nand_4 g06225(.A(new_n4017), .B(new_n4008), .Y(new_n6602));
  nand_4 g06226(.A(new_n6602), .B(new_n4005_1), .Y(new_n6603));
  nor_4  g06227(.A(new_n6603), .B(new_n6601), .Y(new_n6604_1));
  not_3  g06228(.A(new_n6604_1), .Y(new_n6605));
  not_3  g06229(.A(new_n6570), .Y(new_n6606));
  xor_3  g06230(.A(new_n6579), .B(new_n6606), .Y(new_n6607));
  not_3  g06231(.A(new_n6603), .Y(new_n6608));
  nor_4  g06232(.A(new_n6608), .B(new_n6600), .Y(new_n6609));
  nor_4  g06233(.A(new_n6609), .B(new_n6604_1), .Y(new_n6610));
  nand_4 g06234(.A(new_n6610), .B(new_n6607), .Y(new_n6611_1));
  nand_4 g06235(.A(new_n6611_1), .B(new_n6605), .Y(new_n6612));
  not_3  g06236(.A(new_n6612), .Y(new_n6613));
  nand_4 g06237(.A(new_n6613), .B(new_n6599), .Y(new_n6614));
  nand_4 g06238(.A(new_n6590), .B(new_n6587), .Y(new_n6615));
  not_3  g06239(.A(new_n6615), .Y(new_n6616));
  nor_4  g06240(.A(new_n6596), .B(new_n6591), .Y(new_n6617));
  nor_4  g06241(.A(new_n6617), .B(new_n6616), .Y(new_n6618));
  not_3  g06242(.A(new_n6618), .Y(new_n6619));
  nand_4 g06243(.A(n10327), .B(n2564), .Y(new_n6620));
  nand_4 g06244(.A(n11662), .B(n4189), .Y(new_n6621));
  nand_4 g06245(.A(n9583), .B(n6687), .Y(new_n6622));
  not_3  g06246(.A(new_n6622), .Y(new_n6623));
  xor_3  g06247(.A(new_n6623), .B(new_n6621), .Y(new_n6624));
  xnor_3 g06248(.A(new_n6624), .B(new_n6620), .Y(new_n6625));
  xnor_3 g06249(.A(new_n6625), .B(new_n6619), .Y(new_n6626));
  nor_4  g06250(.A(new_n6589), .B(new_n6588), .Y(new_n6627));
  nand_4 g06251(.A(n7456), .B(n6770), .Y(new_n6628));
  not_3  g06252(.A(new_n6628), .Y(new_n6629));
  xor_3  g06253(.A(new_n6629), .B(new_n6627), .Y(new_n6630));
  nand_4 g06254(.A(n3932), .B(n3627), .Y(new_n6631));
  nand_4 g06255(.A(n12591), .B(n9920), .Y(new_n6632));
  nand_4 g06256(.A(n4516), .B(n1798), .Y(new_n6633));
  nand_4 g06257(.A(new_n6633), .B(new_n6632), .Y(new_n6634));
  not_3  g06258(.A(new_n6632), .Y(new_n6635));
  not_3  g06259(.A(new_n6633), .Y(new_n6636));
  nand_4 g06260(.A(new_n6636), .B(new_n6635), .Y(new_n6637));
  nand_4 g06261(.A(new_n6637), .B(new_n6634), .Y(new_n6638));
  xor_3  g06262(.A(new_n6638), .B(new_n6631), .Y(new_n6639));
  xnor_3 g06263(.A(new_n6639), .B(new_n6630), .Y(new_n6640));
  not_3  g06264(.A(new_n6640), .Y(new_n6641));
  xnor_3 g06265(.A(new_n6641), .B(new_n6626), .Y(new_n6642));
  nand_4 g06266(.A(new_n6584), .B(new_n6581), .Y(new_n6643));
  nor_4  g06267(.A(new_n6583), .B(new_n6582), .Y(new_n6644));
  nor_4  g06268(.A(new_n6597), .B(new_n6585), .Y(new_n6645_1));
  xnor_3 g06269(.A(new_n6645_1), .B(new_n6644), .Y(new_n6646));
  nand_4 g06270(.A(new_n6646), .B(new_n6643), .Y(new_n6647));
  xnor_3 g06271(.A(new_n6647), .B(new_n6642), .Y(new_n6648));
  xnor_3 g06272(.A(new_n6648), .B(new_n6614), .Y(new_n6649));
  nand_4 g06273(.A(n10327), .B(n6687), .Y(new_n6650));
  not_3  g06274(.A(new_n6650), .Y(new_n6651));
  xnor_3 g06275(.A(new_n6612), .B(new_n6598), .Y(new_n6652));
  not_3  g06276(.A(new_n6652), .Y(new_n6653));
  nand_4 g06277(.A(new_n6653), .B(new_n6651), .Y(new_n6654));
  nor_4  g06278(.A(new_n4027), .B(new_n4019), .Y(new_n6655));
  not_3  g06279(.A(new_n6655), .Y(new_n6656));
  not_3  g06280(.A(new_n6611_1), .Y(new_n6657));
  nor_4  g06281(.A(new_n6610), .B(new_n6607), .Y(new_n6658));
  nor_4  g06282(.A(new_n6658), .B(new_n6657), .Y(new_n6659));
  nor_4  g06283(.A(new_n6659), .B(new_n6656), .Y(new_n6660));
  nor_4  g06284(.A(new_n6652), .B(new_n6650), .Y(new_n6661));
  nor_4  g06285(.A(new_n6653), .B(new_n6651), .Y(new_n6662));
  nor_4  g06286(.A(new_n6662), .B(new_n6661), .Y(new_n6663));
  nand_4 g06287(.A(new_n6663), .B(new_n6660), .Y(new_n6664));
  nand_4 g06288(.A(new_n6664), .B(new_n6654), .Y(new_n6665));
  xnor_3 g06289(.A(new_n6665), .B(new_n6649), .Y(new_n6666));
  nand_4 g06290(.A(n3022), .B(n2226), .Y(new_n6667));
  nand_4 g06291(.A(n9640), .B(n1094), .Y(new_n6668));
  nand_4 g06292(.A(n10678), .B(n6703), .Y(new_n6669));
  xnor_3 g06293(.A(new_n6669), .B(new_n6668), .Y(new_n6670));
  nor_4  g06294(.A(new_n6670), .B(new_n6667), .Y(new_n6671));
  not_3  g06295(.A(new_n6667), .Y(new_n6672));
  not_3  g06296(.A(new_n6670), .Y(new_n6673));
  nor_4  g06297(.A(new_n6673), .B(new_n6672), .Y(new_n6674));
  nor_4  g06298(.A(new_n6674), .B(new_n6671), .Y(new_n6675));
  nand_4 g06299(.A(n6986), .B(n3022), .Y(new_n6676));
  not_3  g06300(.A(new_n6676), .Y(new_n6677));
  nand_4 g06301(.A(n6703), .B(n1094), .Y(new_n6678));
  not_3  g06302(.A(new_n6678), .Y(new_n6679));
  nor_4  g06303(.A(new_n6679), .B(new_n6677), .Y(new_n6680));
  nor_4  g06304(.A(new_n6678), .B(new_n6676), .Y(new_n6681));
  nand_4 g06305(.A(n9640), .B(n2226), .Y(new_n6682));
  not_3  g06306(.A(new_n6682), .Y(new_n6683));
  nor_4  g06307(.A(new_n6683), .B(new_n6681), .Y(new_n6684));
  nor_4  g06308(.A(new_n6684), .B(new_n6680), .Y(new_n6685));
  xnor_3 g06309(.A(new_n6685), .B(new_n6675), .Y(new_n6686));
  nand_4 g06310(.A(n10928), .B(n10451), .Y(new_n6687_1));
  nand_4 g06311(.A(n11023), .B(n6986), .Y(new_n6688));
  xor_3  g06312(.A(new_n6688), .B(new_n6687_1), .Y(new_n6689_1));
  xnor_3 g06313(.A(new_n6689_1), .B(new_n6686), .Y(new_n6690));
  nand_4 g06314(.A(n11023), .B(n10928), .Y(new_n6691));
  not_3  g06315(.A(new_n6691), .Y(new_n6692));
  nor_4  g06316(.A(new_n4198), .B(new_n4192), .Y(new_n6693));
  nor_4  g06317(.A(new_n6693), .B(new_n4197), .Y(new_n6694));
  nand_4 g06318(.A(new_n6694), .B(new_n6692), .Y(new_n6695));
  xor_3  g06319(.A(new_n6694), .B(new_n6692), .Y(new_n6696));
  nor_4  g06320(.A(new_n6681), .B(new_n6680), .Y(new_n6697));
  xor_3  g06321(.A(new_n6697), .B(new_n6683), .Y(new_n6698));
  nand_4 g06322(.A(new_n6698), .B(new_n6696), .Y(new_n6699));
  nand_4 g06323(.A(new_n6699), .B(new_n6695), .Y(new_n6700));
  xnor_3 g06324(.A(new_n6700), .B(new_n6690), .Y(new_n6701));
  not_3  g06325(.A(new_n6701), .Y(new_n6702));
  nand_4 g06326(.A(n10451), .B(n8336), .Y(new_n6703_1));
  not_3  g06327(.A(new_n6703_1), .Y(new_n6704));
  xor_3  g06328(.A(new_n6694), .B(new_n6691), .Y(new_n6705));
  xor_3  g06329(.A(new_n6697), .B(new_n6682), .Y(new_n6706));
  nor_4  g06330(.A(new_n6706), .B(new_n6705), .Y(new_n6707));
  nor_4  g06331(.A(new_n6698), .B(new_n6696), .Y(new_n6708));
  nor_4  g06332(.A(new_n6708), .B(new_n6707), .Y(new_n6709));
  nand_4 g06333(.A(new_n6709), .B(new_n6704), .Y(new_n6710));
  nor_4  g06334(.A(new_n4189_1), .B(new_n4184), .Y(new_n6711));
  not_3  g06335(.A(new_n6711), .Y(new_n6712));
  nand_4 g06336(.A(new_n4200), .B(new_n4190_1), .Y(new_n6713));
  nand_4 g06337(.A(new_n6713), .B(new_n6712), .Y(new_n6714));
  xnor_3 g06338(.A(new_n6706), .B(new_n6705), .Y(new_n6715));
  xnor_3 g06339(.A(new_n6715), .B(new_n6704), .Y(new_n6716));
  nand_4 g06340(.A(new_n6716), .B(new_n6714), .Y(new_n6717));
  nand_4 g06341(.A(new_n6717), .B(new_n6710), .Y(new_n6718));
  nand_4 g06342(.A(new_n6718), .B(new_n6702), .Y(new_n6719));
  nand_4 g06343(.A(new_n6685), .B(new_n6675), .Y(new_n6720));
  not_3  g06344(.A(new_n6720), .Y(new_n6721));
  nor_4  g06345(.A(new_n6721), .B(new_n6671), .Y(new_n6722));
  not_3  g06346(.A(new_n6722), .Y(new_n6723));
  nand_4 g06347(.A(n10928), .B(n10278), .Y(new_n6724));
  nand_4 g06348(.A(n10451), .B(n6986), .Y(new_n6725));
  nand_4 g06349(.A(n11423), .B(n8336), .Y(new_n6726));
  not_3  g06350(.A(new_n6726), .Y(new_n6727));
  xor_3  g06351(.A(new_n6727), .B(new_n6725), .Y(new_n6728));
  xnor_3 g06352(.A(new_n6728), .B(new_n6724), .Y(new_n6729));
  xnor_3 g06353(.A(new_n6729), .B(new_n6723), .Y(new_n6730));
  nor_4  g06354(.A(new_n6669), .B(new_n6668), .Y(new_n6731));
  not_3  g06355(.A(new_n6731), .Y(new_n6732));
  nand_4 g06356(.A(n11023), .B(n2226), .Y(new_n6733));
  xor_3  g06357(.A(new_n6733), .B(new_n6732), .Y(new_n6734));
  not_3  g06358(.A(new_n6734), .Y(new_n6735));
  nand_4 g06359(.A(n10678), .B(n9640), .Y(new_n6736));
  nand_4 g06360(.A(n3022), .B(n1094), .Y(new_n6737));
  nand_4 g06361(.A(n7320), .B(n6703), .Y(new_n6738));
  not_3  g06362(.A(new_n6738), .Y(new_n6739));
  xor_3  g06363(.A(new_n6739), .B(new_n6737), .Y(new_n6740));
  xnor_3 g06364(.A(new_n6740), .B(new_n6736), .Y(new_n6741));
  xnor_3 g06365(.A(new_n6741), .B(new_n6735), .Y(new_n6742_1));
  xnor_3 g06366(.A(new_n6742_1), .B(new_n6730), .Y(new_n6743));
  not_3  g06367(.A(new_n6743), .Y(new_n6744));
  not_3  g06368(.A(new_n6686), .Y(new_n6745));
  nand_4 g06369(.A(new_n6689_1), .B(new_n6745), .Y(new_n6746));
  nor_4  g06370(.A(new_n6688), .B(new_n6687_1), .Y(new_n6747));
  nand_4 g06371(.A(new_n6700), .B(new_n6690), .Y(new_n6748));
  not_3  g06372(.A(new_n6748), .Y(new_n6749));
  xnor_3 g06373(.A(new_n6749), .B(new_n6747), .Y(new_n6750));
  nand_4 g06374(.A(new_n6750), .B(new_n6746), .Y(new_n6751));
  xnor_3 g06375(.A(new_n6751), .B(new_n6744), .Y(new_n6752));
  xnor_3 g06376(.A(new_n6752), .B(new_n6719), .Y(new_n6753));
  nand_4 g06377(.A(n10278), .B(n8336), .Y(new_n6754));
  not_3  g06378(.A(new_n6754), .Y(new_n6755));
  xnor_3 g06379(.A(new_n6718), .B(new_n6701), .Y(new_n6756));
  nor_4  g06380(.A(new_n6756), .B(new_n6755), .Y(new_n6757));
  not_3  g06381(.A(new_n4203_1), .Y(new_n6758));
  nor_4  g06382(.A(new_n6758), .B(new_n4201), .Y(new_n6759));
  not_3  g06383(.A(new_n6759), .Y(new_n6760));
  xnor_3 g06384(.A(new_n6716), .B(new_n6714), .Y(new_n6761));
  nor_4  g06385(.A(new_n6761), .B(new_n6760), .Y(new_n6762));
  not_3  g06386(.A(new_n6756), .Y(new_n6763));
  xor_3  g06387(.A(new_n6763), .B(new_n6755), .Y(new_n6764));
  nor_4  g06388(.A(new_n6764), .B(new_n6762), .Y(new_n6765));
  nor_4  g06389(.A(new_n6765), .B(new_n6757), .Y(new_n6766));
  not_3  g06390(.A(new_n6766), .Y(new_n6767));
  xnor_3 g06391(.A(new_n6767), .B(new_n6753), .Y(new_n6768));
  nand_4 g06392(.A(n8665), .B(n7160), .Y(new_n6769));
  nand_4 g06393(.A(n4828), .B(n1067), .Y(new_n6770_1));
  nand_4 g06394(.A(n5645), .B(n2515), .Y(new_n6771));
  xnor_3 g06395(.A(new_n6771), .B(new_n6770_1), .Y(new_n6772));
  nor_4  g06396(.A(new_n6772), .B(new_n6769), .Y(new_n6773));
  not_3  g06397(.A(new_n6769), .Y(new_n6774));
  not_3  g06398(.A(new_n6772), .Y(new_n6775));
  nor_4  g06399(.A(new_n6775), .B(new_n6774), .Y(new_n6776_1));
  nor_4  g06400(.A(new_n6776_1), .B(new_n6773), .Y(new_n6777));
  nand_4 g06401(.A(n8665), .B(n7891), .Y(new_n6778));
  nand_4 g06402(.A(n5645), .B(n4828), .Y(new_n6779));
  and_4  g06403(.A(new_n6779), .B(new_n6778), .Y(new_n6780));
  nand_4 g06404(.A(n7160), .B(n1067), .Y(new_n6781));
  not_3  g06405(.A(new_n6781), .Y(new_n6782));
  xnor_3 g06406(.A(new_n6779), .B(new_n6778), .Y(new_n6783));
  nor_4  g06407(.A(new_n6783), .B(new_n6782), .Y(new_n6784));
  nor_4  g06408(.A(new_n6784), .B(new_n6780), .Y(new_n6785));
  xnor_3 g06409(.A(new_n6785), .B(new_n6777), .Y(new_n6786));
  nand_4 g06410(.A(n12391), .B(n2551), .Y(new_n6787));
  nand_4 g06411(.A(n11922), .B(n7891), .Y(new_n6788));
  not_3  g06412(.A(new_n6788), .Y(new_n6789));
  xor_3  g06413(.A(new_n6789), .B(new_n6787), .Y(new_n6790));
  xnor_3 g06414(.A(new_n6790), .B(new_n6786), .Y(new_n6791));
  nand_4 g06415(.A(n12391), .B(n11922), .Y(new_n6792));
  not_3  g06416(.A(new_n4136), .Y(new_n6793));
  nand_4 g06417(.A(new_n4139), .B(new_n6793), .Y(new_n6794));
  nand_4 g06418(.A(new_n6794), .B(new_n4141_1), .Y(new_n6795));
  not_3  g06419(.A(new_n6795), .Y(new_n6796));
  nor_4  g06420(.A(new_n6796), .B(new_n6792), .Y(new_n6797_1));
  xnor_3 g06421(.A(new_n6783), .B(new_n6781), .Y(new_n6798));
  xnor_3 g06422(.A(new_n6796), .B(new_n6792), .Y(new_n6799));
  nor_4  g06423(.A(new_n6799), .B(new_n6798), .Y(new_n6800));
  nor_4  g06424(.A(new_n6800), .B(new_n6797_1), .Y(new_n6801));
  xnor_3 g06425(.A(new_n6801), .B(new_n6791), .Y(new_n6802));
  nand_4 g06426(.A(n12069), .B(n2551), .Y(new_n6803));
  xnor_3 g06427(.A(new_n6799), .B(new_n6798), .Y(new_n6804));
  nor_4  g06428(.A(new_n6804), .B(new_n6803), .Y(new_n6805));
  not_3  g06429(.A(new_n6805), .Y(new_n6806_1));
  nand_4 g06430(.A(new_n6804), .B(new_n6803), .Y(new_n6807));
  nand_4 g06431(.A(new_n4134), .B(new_n4129), .Y(new_n6808));
  nor_4  g06432(.A(new_n4143), .B(new_n4135), .Y(new_n6809_1));
  not_3  g06433(.A(new_n6809_1), .Y(new_n6810));
  nand_4 g06434(.A(new_n6810), .B(new_n6808), .Y(new_n6811));
  nand_4 g06435(.A(new_n6811), .B(new_n6807), .Y(new_n6812));
  nand_4 g06436(.A(new_n6812), .B(new_n6806_1), .Y(new_n6813));
  not_3  g06437(.A(new_n6813), .Y(new_n6814));
  nor_4  g06438(.A(new_n6814), .B(new_n6802), .Y(new_n6815));
  not_3  g06439(.A(new_n6815), .Y(new_n6816));
  nand_4 g06440(.A(new_n6785), .B(new_n6777), .Y(new_n6817));
  not_3  g06441(.A(new_n6817), .Y(new_n6818));
  nor_4  g06442(.A(new_n6818), .B(new_n6773), .Y(new_n6819));
  not_3  g06443(.A(new_n6819), .Y(new_n6820));
  nand_4 g06444(.A(n12826), .B(n12391), .Y(new_n6821));
  nand_4 g06445(.A(n7891), .B(n2551), .Y(new_n6822_1));
  nand_4 g06446(.A(n12069), .B(n4094), .Y(new_n6823));
  not_3  g06447(.A(new_n6823), .Y(new_n6824));
  xor_3  g06448(.A(new_n6824), .B(new_n6822_1), .Y(new_n6825));
  xnor_3 g06449(.A(new_n6825), .B(new_n6821), .Y(new_n6826_1));
  xnor_3 g06450(.A(new_n6826_1), .B(new_n6820), .Y(new_n6827));
  nor_4  g06451(.A(new_n6771), .B(new_n6770_1), .Y(new_n6828));
  not_3  g06452(.A(new_n6828), .Y(new_n6829));
  nand_4 g06453(.A(n11922), .B(n7160), .Y(new_n6830));
  xor_3  g06454(.A(new_n6830), .B(new_n6829), .Y(new_n6831));
  nand_4 g06455(.A(n2515), .B(n1067), .Y(new_n6832));
  not_3  g06456(.A(new_n6832), .Y(new_n6833));
  nand_4 g06457(.A(n8665), .B(n4828), .Y(new_n6834));
  nand_4 g06458(.A(n5645), .B(n1199), .Y(new_n6835));
  xor_3  g06459(.A(new_n6835), .B(new_n6834), .Y(new_n6836));
  xnor_3 g06460(.A(new_n6836), .B(new_n6833), .Y(new_n6837));
  xnor_3 g06461(.A(new_n6837), .B(new_n6831), .Y(new_n6838));
  xnor_3 g06462(.A(new_n6838), .B(new_n6827), .Y(new_n6839));
  not_3  g06463(.A(new_n6786), .Y(new_n6840));
  not_3  g06464(.A(new_n6790), .Y(new_n6841));
  nand_4 g06465(.A(new_n6841), .B(new_n6840), .Y(new_n6842));
  nor_4  g06466(.A(new_n6788), .B(new_n6787), .Y(new_n6843));
  nor_4  g06467(.A(new_n6801), .B(new_n6791), .Y(new_n6844));
  xnor_3 g06468(.A(new_n6844), .B(new_n6843), .Y(new_n6845));
  nand_4 g06469(.A(new_n6845), .B(new_n6842), .Y(new_n6846));
  xnor_3 g06470(.A(new_n6846), .B(new_n6839), .Y(new_n6847));
  xnor_3 g06471(.A(new_n6847), .B(new_n6816), .Y(new_n6848));
  nand_4 g06472(.A(n12826), .B(n12069), .Y(new_n6849));
  not_3  g06473(.A(new_n6849), .Y(new_n6850));
  not_3  g06474(.A(new_n6802), .Y(new_n6851));
  nor_4  g06475(.A(new_n6813), .B(new_n6851), .Y(new_n6852));
  nor_4  g06476(.A(new_n6852), .B(new_n6815), .Y(new_n6853));
  nor_4  g06477(.A(new_n6853), .B(new_n6850), .Y(new_n6854));
  nand_4 g06478(.A(new_n4170), .B(new_n4127), .Y(new_n6855));
  not_3  g06479(.A(new_n6807), .Y(new_n6856));
  nor_4  g06480(.A(new_n6856), .B(new_n6805), .Y(new_n6857));
  xnor_3 g06481(.A(new_n6857), .B(new_n6811), .Y(new_n6858));
  nor_4  g06482(.A(new_n6858), .B(new_n6855), .Y(new_n6859));
  xnor_3 g06483(.A(new_n6853), .B(new_n6850), .Y(new_n6860_1));
  nor_4  g06484(.A(new_n6860_1), .B(new_n6859), .Y(new_n6861));
  nor_4  g06485(.A(new_n6861), .B(new_n6854), .Y(new_n6862));
  xnor_3 g06486(.A(new_n6862), .B(new_n6848), .Y(new_n6863));
  nand_4 g06487(.A(n3754), .B(n996), .Y(new_n6864));
  nand_4 g06488(.A(n10898), .B(n5767), .Y(new_n6865));
  nand_4 g06489(.A(n11876), .B(n5319), .Y(new_n6866));
  xnor_3 g06490(.A(new_n6866), .B(new_n6865), .Y(new_n6867));
  nor_4  g06491(.A(new_n6867), .B(new_n6864), .Y(new_n6868));
  not_3  g06492(.A(new_n6864), .Y(new_n6869));
  not_3  g06493(.A(new_n6867), .Y(new_n6870));
  nor_4  g06494(.A(new_n6870), .B(new_n6869), .Y(new_n6871));
  nor_4  g06495(.A(new_n6871), .B(new_n6868), .Y(new_n6872));
  nand_4 g06496(.A(n5314), .B(n3754), .Y(new_n6873));
  nand_4 g06497(.A(n10898), .B(n996), .Y(new_n6874));
  and_4  g06498(.A(new_n6874), .B(new_n6873), .Y(new_n6875));
  nand_4 g06499(.A(n11876), .B(n5767), .Y(new_n6876));
  not_3  g06500(.A(new_n6876), .Y(new_n6877_1));
  xnor_3 g06501(.A(new_n6874), .B(new_n6873), .Y(new_n6878));
  nor_4  g06502(.A(new_n6878), .B(new_n6877_1), .Y(new_n6879));
  nor_4  g06503(.A(new_n6879), .B(new_n6875), .Y(new_n6880));
  xnor_3 g06504(.A(new_n6880), .B(new_n6872), .Y(new_n6881));
  nand_4 g06505(.A(n11153), .B(n159), .Y(new_n6882));
  nand_4 g06506(.A(n5314), .B(n2749), .Y(new_n6883));
  not_3  g06507(.A(new_n6883), .Y(new_n6884));
  xor_3  g06508(.A(new_n6884), .B(new_n6882), .Y(new_n6885));
  xnor_3 g06509(.A(new_n6885), .B(new_n6881), .Y(new_n6886));
  nand_4 g06510(.A(n11153), .B(n2749), .Y(new_n6887));
  not_3  g06511(.A(new_n6887), .Y(new_n6888));
  not_3  g06512(.A(new_n4152), .Y(new_n6889));
  nor_4  g06513(.A(new_n4158), .B(new_n6889), .Y(new_n6890));
  nor_4  g06514(.A(new_n6890), .B(new_n4157), .Y(new_n6891));
  and_4  g06515(.A(new_n6891), .B(new_n6888), .Y(new_n6892));
  xnor_3 g06516(.A(new_n6891), .B(new_n6887), .Y(new_n6893));
  not_3  g06517(.A(new_n6893), .Y(new_n6894));
  xnor_3 g06518(.A(new_n6878), .B(new_n6876), .Y(new_n6895));
  nor_4  g06519(.A(new_n6895), .B(new_n6894), .Y(new_n6896));
  nor_4  g06520(.A(new_n6896), .B(new_n6892), .Y(new_n6897));
  xnor_3 g06521(.A(new_n6897), .B(new_n6886), .Y(new_n6898));
  nand_4 g06522(.A(n11222), .B(n159), .Y(new_n6899));
  xnor_3 g06523(.A(new_n6895), .B(new_n6894), .Y(new_n6900));
  nor_4  g06524(.A(new_n6900), .B(new_n6899), .Y(new_n6901));
  not_3  g06525(.A(new_n6901), .Y(new_n6902));
  nand_4 g06526(.A(new_n6900), .B(new_n6899), .Y(new_n6903));
  nand_4 g06527(.A(new_n4150), .B(new_n4147), .Y(new_n6904));
  not_3  g06528(.A(new_n6904), .Y(new_n6905));
  nor_4  g06529(.A(new_n4161), .B(new_n4151), .Y(new_n6906));
  nor_4  g06530(.A(new_n6906), .B(new_n6905), .Y(new_n6907));
  not_3  g06531(.A(new_n6907), .Y(new_n6908));
  nand_4 g06532(.A(new_n6908), .B(new_n6903), .Y(new_n6909));
  nand_4 g06533(.A(new_n6909), .B(new_n6902), .Y(new_n6910));
  not_3  g06534(.A(new_n6910), .Y(new_n6911));
  nor_4  g06535(.A(new_n6911), .B(new_n6898), .Y(new_n6912));
  not_3  g06536(.A(new_n6881), .Y(new_n6913));
  not_3  g06537(.A(new_n6885), .Y(new_n6914));
  nand_4 g06538(.A(new_n6914), .B(new_n6913), .Y(new_n6915));
  nor_4  g06539(.A(new_n6883), .B(new_n6882), .Y(new_n6916));
  nor_4  g06540(.A(new_n6897), .B(new_n6886), .Y(new_n6917));
  xnor_3 g06541(.A(new_n6917), .B(new_n6916), .Y(new_n6918));
  nand_4 g06542(.A(new_n6918), .B(new_n6915), .Y(new_n6919));
  not_3  g06543(.A(new_n6868), .Y(new_n6920));
  nand_4 g06544(.A(new_n6880), .B(new_n6872), .Y(new_n6921));
  nand_4 g06545(.A(new_n6921), .B(new_n6920), .Y(new_n6922));
  nand_4 g06546(.A(n11153), .B(n1510), .Y(new_n6923));
  not_3  g06547(.A(new_n6923), .Y(new_n6924));
  nand_4 g06548(.A(n5314), .B(n159), .Y(new_n6925));
  nand_4 g06549(.A(n12247), .B(n11222), .Y(new_n6926));
  not_3  g06550(.A(new_n6926), .Y(new_n6927));
  xor_3  g06551(.A(new_n6927), .B(new_n6925), .Y(new_n6928));
  xnor_3 g06552(.A(new_n6928), .B(new_n6924), .Y(new_n6929));
  not_3  g06553(.A(new_n6929), .Y(new_n6930));
  xnor_3 g06554(.A(new_n6930), .B(new_n6922), .Y(new_n6931));
  nor_4  g06555(.A(new_n6866), .B(new_n6865), .Y(new_n6932));
  nand_4 g06556(.A(n2749), .B(n996), .Y(new_n6933));
  not_3  g06557(.A(new_n6933), .Y(new_n6934));
  xor_3  g06558(.A(new_n6934), .B(new_n6932), .Y(new_n6935));
  not_3  g06559(.A(new_n6935), .Y(new_n6936));
  nand_4 g06560(.A(n10898), .B(n5319), .Y(new_n6937));
  not_3  g06561(.A(new_n6937), .Y(new_n6938));
  nand_4 g06562(.A(n11876), .B(n9457), .Y(new_n6939));
  nand_4 g06563(.A(n5767), .B(n3754), .Y(new_n6940));
  not_3  g06564(.A(new_n6940), .Y(new_n6941));
  xor_3  g06565(.A(new_n6941), .B(new_n6939), .Y(new_n6942));
  xnor_3 g06566(.A(new_n6942), .B(new_n6938), .Y(new_n6943));
  xnor_3 g06567(.A(new_n6943), .B(new_n6936), .Y(new_n6944));
  not_3  g06568(.A(new_n6944), .Y(new_n6945));
  xnor_3 g06569(.A(new_n6945), .B(new_n6931), .Y(new_n6946));
  xnor_3 g06570(.A(new_n6946), .B(new_n6919), .Y(new_n6947));
  xnor_3 g06571(.A(new_n6947), .B(new_n6912), .Y(new_n6948));
  nand_4 g06572(.A(n11222), .B(n1510), .Y(new_n6949));
  not_3  g06573(.A(new_n6949), .Y(new_n6950));
  not_3  g06574(.A(new_n6898), .Y(new_n6951));
  nor_4  g06575(.A(new_n6910), .B(new_n6951), .Y(new_n6952));
  nor_4  g06576(.A(new_n6952), .B(new_n6912), .Y(new_n6953));
  nor_4  g06577(.A(new_n6953), .B(new_n6950), .Y(new_n6954));
  not_3  g06578(.A(new_n4165), .Y(new_n6955));
  nand_4 g06579(.A(new_n6903), .B(new_n6902), .Y(new_n6956));
  xnor_3 g06580(.A(new_n6956), .B(new_n6908), .Y(new_n6957));
  not_3  g06581(.A(new_n6957), .Y(new_n6958));
  nor_4  g06582(.A(new_n6958), .B(new_n6955), .Y(new_n6959));
  xnor_3 g06583(.A(new_n6953), .B(new_n6950), .Y(new_n6960));
  nor_4  g06584(.A(new_n6960), .B(new_n6959), .Y(new_n6961));
  nor_4  g06585(.A(new_n6961), .B(new_n6954), .Y(new_n6962));
  xnor_3 g06586(.A(new_n6962), .B(new_n6948), .Y(new_n6963));
  xnor_3 g06587(.A(new_n6960), .B(new_n6959), .Y(new_n6964));
  xnor_3 g06588(.A(new_n6860_1), .B(new_n6859), .Y(new_n6965));
  nor_4  g06589(.A(new_n6965), .B(new_n6964), .Y(new_n6966));
  not_3  g06590(.A(new_n6966), .Y(new_n6967));
  not_3  g06591(.A(new_n6959), .Y(new_n6968));
  xnor_3 g06592(.A(new_n6960), .B(new_n6968), .Y(new_n6969));
  not_3  g06593(.A(new_n6859), .Y(new_n6970));
  xnor_3 g06594(.A(new_n6860_1), .B(new_n6970), .Y(new_n6971));
  nor_4  g06595(.A(new_n6971), .B(new_n6969), .Y(new_n6972));
  xnor_3 g06596(.A(new_n6858), .B(new_n6855), .Y(new_n6973));
  not_3  g06597(.A(new_n6973), .Y(new_n6974));
  not_3  g06598(.A(new_n4169), .Y(new_n6975));
  nand_4 g06599(.A(new_n4180), .B(new_n6975), .Y(new_n6976));
  not_3  g06600(.A(new_n6976), .Y(new_n6977));
  nand_4 g06601(.A(new_n6977), .B(new_n6974), .Y(new_n6978));
  nand_4 g06602(.A(new_n6976), .B(new_n6973), .Y(new_n6979));
  nor_4  g06603(.A(new_n6957), .B(new_n4165), .Y(new_n6980));
  nor_4  g06604(.A(new_n6980), .B(new_n6959), .Y(new_n6981));
  nand_4 g06605(.A(new_n6981), .B(new_n6979), .Y(new_n6982));
  nand_4 g06606(.A(new_n6982), .B(new_n6978), .Y(new_n6983));
  nor_4  g06607(.A(new_n6983), .B(new_n6972), .Y(new_n6984));
  not_3  g06608(.A(new_n6984), .Y(new_n6985));
  nand_4 g06609(.A(new_n6985), .B(new_n6967), .Y(new_n6986_1));
  xnor_3 g06610(.A(new_n6986_1), .B(new_n6963), .Y(new_n6987));
  xnor_3 g06611(.A(new_n6987), .B(new_n6863), .Y(new_n6988));
  xnor_3 g06612(.A(new_n6988), .B(new_n6768), .Y(new_n6989));
  not_3  g06613(.A(new_n6762), .Y(new_n6990));
  not_3  g06614(.A(new_n6764), .Y(new_n6991));
  nor_4  g06615(.A(new_n6991), .B(new_n6990), .Y(new_n6992));
  nor_4  g06616(.A(new_n6992), .B(new_n6765), .Y(new_n6993));
  not_3  g06617(.A(new_n6993), .Y(new_n6994));
  not_3  g06618(.A(new_n6761), .Y(new_n6995));
  xor_3  g06619(.A(new_n6995), .B(new_n6760), .Y(new_n6996));
  not_3  g06620(.A(new_n6996), .Y(new_n6997));
  not_3  g06621(.A(new_n6981), .Y(new_n6998));
  xnor_3 g06622(.A(new_n6976), .B(new_n6974), .Y(new_n6999));
  xnor_3 g06623(.A(new_n6999), .B(new_n6998), .Y(new_n7000));
  nand_4 g06624(.A(new_n7000), .B(new_n6997), .Y(new_n7001));
  xnor_3 g06625(.A(new_n6999), .B(new_n6981), .Y(new_n7002));
  nand_4 g06626(.A(new_n7002), .B(new_n6996), .Y(new_n7003));
  nand_4 g06627(.A(new_n4214), .B(new_n4209), .Y(new_n7004));
  nand_4 g06628(.A(new_n7004), .B(new_n7003), .Y(new_n7005));
  nand_4 g06629(.A(new_n7005), .B(new_n7001), .Y(new_n7006));
  nand_4 g06630(.A(new_n7006), .B(new_n6994), .Y(new_n7007));
  xnor_3 g06631(.A(new_n7006), .B(new_n6993), .Y(new_n7008));
  not_3  g06632(.A(new_n6972), .Y(new_n7009));
  nand_4 g06633(.A(new_n7009), .B(new_n6967), .Y(new_n7010));
  xnor_3 g06634(.A(new_n7010), .B(new_n6983), .Y(new_n7011));
  nand_4 g06635(.A(new_n7011), .B(new_n7008), .Y(new_n7012));
  nand_4 g06636(.A(new_n7012), .B(new_n7007), .Y(new_n7013));
  xnor_3 g06637(.A(new_n7013), .B(new_n6989), .Y(new_n7014));
  nand_4 g06638(.A(new_n7014), .B(new_n6666), .Y(new_n7015));
  not_3  g06639(.A(new_n6666), .Y(new_n7016));
  not_3  g06640(.A(new_n7014), .Y(new_n7017));
  nand_4 g06641(.A(new_n7017), .B(new_n7016), .Y(new_n7018));
  nand_4 g06642(.A(new_n7018), .B(new_n7015), .Y(new_n7019));
  not_3  g06643(.A(new_n6663), .Y(new_n7020));
  xor_3  g06644(.A(new_n7020), .B(new_n6660), .Y(new_n7021));
  not_3  g06645(.A(new_n7021), .Y(new_n7022));
  xnor_3 g06646(.A(new_n7011), .B(new_n7008), .Y(new_n7023));
  not_3  g06647(.A(new_n7023), .Y(new_n7024));
  nand_4 g06648(.A(new_n7024), .B(new_n7022), .Y(new_n7025));
  nand_4 g06649(.A(new_n7023), .B(new_n7021), .Y(new_n7026));
  xor_3  g06650(.A(new_n6659), .B(new_n6655), .Y(new_n7027));
  not_3  g06651(.A(new_n7027), .Y(new_n7028));
  nand_4 g06652(.A(new_n7003), .B(new_n7001), .Y(new_n7029));
  xnor_3 g06653(.A(new_n7029), .B(new_n7004), .Y(new_n7030));
  nor_4  g06654(.A(new_n7030), .B(new_n7028), .Y(new_n7031));
  nand_4 g06655(.A(new_n4124), .B(new_n4028), .Y(new_n7032));
  nand_4 g06656(.A(new_n4216), .B(new_n4125), .Y(new_n7033));
  nand_4 g06657(.A(new_n7033), .B(new_n7032), .Y(new_n7034));
  xnor_3 g06658(.A(new_n7030), .B(new_n7028), .Y(new_n7035));
  nor_4  g06659(.A(new_n7035), .B(new_n7034), .Y(new_n7036));
  nor_4  g06660(.A(new_n7036), .B(new_n7031), .Y(new_n7037));
  nand_4 g06661(.A(new_n7037), .B(new_n7026), .Y(new_n7038));
  nand_4 g06662(.A(new_n7038), .B(new_n7025), .Y(new_n7039));
  xnor_3 g06663(.A(new_n7039), .B(new_n7019), .Y(n2301));
  xor_3  g06664(.A(new_n4122), .B(new_n4121), .Y(n2316));
  nand_4 g06665(.A(n4634), .B(n1333), .Y(new_n7042));
  not_3  g06666(.A(new_n7042), .Y(new_n7043));
  not_3  g06667(.A(new_n6301), .Y(new_n7044));
  nor_4  g06668(.A(new_n6307), .B(new_n7044), .Y(new_n7045));
  nor_4  g06669(.A(new_n7045), .B(new_n6306), .Y(new_n7046));
  nand_4 g06670(.A(new_n7046), .B(new_n7043), .Y(new_n7047));
  xnor_3 g06671(.A(new_n7046), .B(new_n7042), .Y(new_n7048));
  nand_4 g06672(.A(n11757), .B(n2879), .Y(new_n7049));
  not_3  g06673(.A(new_n7049), .Y(new_n7050));
  nand_4 g06674(.A(n10223), .B(n3172), .Y(new_n7051));
  not_3  g06675(.A(new_n7051), .Y(new_n7052));
  nand_4 g06676(.A(n7265), .B(n5240), .Y(new_n7053));
  not_3  g06677(.A(new_n7053), .Y(new_n7054));
  nor_4  g06678(.A(new_n7054), .B(new_n7052), .Y(new_n7055));
  not_3  g06679(.A(new_n7055), .Y(new_n7056));
  nor_4  g06680(.A(new_n7053), .B(new_n7051), .Y(new_n7057));
  not_3  g06681(.A(new_n7057), .Y(new_n7058));
  nand_4 g06682(.A(new_n7058), .B(new_n7056), .Y(new_n7059));
  xnor_3 g06683(.A(new_n7059), .B(new_n7050), .Y(new_n7060));
  nand_4 g06684(.A(new_n7060), .B(new_n7048), .Y(new_n7061));
  nand_4 g06685(.A(new_n7061), .B(new_n7047), .Y(new_n7062));
  nand_4 g06686(.A(n4634), .B(n3172), .Y(new_n7063));
  nand_4 g06687(.A(n9195), .B(n1333), .Y(new_n7064));
  xor_3  g06688(.A(new_n7064), .B(new_n7063), .Y(new_n7065));
  xnor_3 g06689(.A(new_n7065), .B(new_n7062), .Y(new_n7066));
  nand_4 g06690(.A(n11757), .B(n10223), .Y(new_n7067));
  not_3  g06691(.A(new_n7067), .Y(new_n7068));
  nand_4 g06692(.A(n5240), .B(n2879), .Y(new_n7069));
  nand_4 g06693(.A(n11821), .B(n7265), .Y(new_n7070));
  xnor_3 g06694(.A(new_n7070), .B(new_n7069), .Y(new_n7071));
  not_3  g06695(.A(new_n7071), .Y(new_n7072));
  nor_4  g06696(.A(new_n7072), .B(new_n7068), .Y(new_n7073));
  nor_4  g06697(.A(new_n7071), .B(new_n7067), .Y(new_n7074));
  nor_4  g06698(.A(new_n7074), .B(new_n7073), .Y(new_n7075));
  nor_4  g06699(.A(new_n7057), .B(new_n7050), .Y(new_n7076));
  nor_4  g06700(.A(new_n7076), .B(new_n7055), .Y(new_n7077));
  not_3  g06701(.A(new_n7077), .Y(new_n7078));
  xor_3  g06702(.A(new_n7078), .B(new_n7075), .Y(new_n7079));
  xnor_3 g06703(.A(new_n7079), .B(new_n7066), .Y(new_n7080));
  not_3  g06704(.A(new_n7080), .Y(new_n7081));
  nand_4 g06705(.A(n9195), .B(n7862), .Y(new_n7082));
  xnor_3 g06706(.A(new_n7060), .B(new_n7048), .Y(new_n7083));
  nor_4  g06707(.A(new_n7083), .B(new_n7082), .Y(new_n7084));
  not_3  g06708(.A(new_n7084), .Y(new_n7085));
  not_3  g06709(.A(new_n6289), .Y(new_n7086));
  nand_4 g06710(.A(new_n6299), .B(new_n7086), .Y(new_n7087));
  xor_3  g06711(.A(new_n6299), .B(new_n7086), .Y(new_n7088));
  xor_3  g06712(.A(new_n6308), .B(new_n7044), .Y(new_n7089));
  nand_4 g06713(.A(new_n7089), .B(new_n7088), .Y(new_n7090));
  nand_4 g06714(.A(new_n7090), .B(new_n7087), .Y(new_n7091));
  not_3  g06715(.A(new_n7082), .Y(new_n7092));
  not_3  g06716(.A(new_n7083), .Y(new_n7093));
  nor_4  g06717(.A(new_n7093), .B(new_n7092), .Y(new_n7094));
  nor_4  g06718(.A(new_n7094), .B(new_n7084), .Y(new_n7095));
  nand_4 g06719(.A(new_n7095), .B(new_n7091), .Y(new_n7096));
  nand_4 g06720(.A(new_n7096), .B(new_n7085), .Y(new_n7097));
  nand_4 g06721(.A(new_n7097), .B(new_n7081), .Y(new_n7098));
  not_3  g06722(.A(new_n7075), .Y(new_n7099));
  nor_4  g06723(.A(new_n7077), .B(new_n7099), .Y(new_n7100));
  nor_4  g06724(.A(new_n7100), .B(new_n7073), .Y(new_n7101));
  nand_4 g06725(.A(n2253), .B(n1333), .Y(new_n7102));
  nand_4 g06726(.A(n9195), .B(n3172), .Y(new_n7103));
  nand_4 g06727(.A(n7862), .B(n3865), .Y(new_n7104));
  xor_3  g06728(.A(new_n7104), .B(new_n7103), .Y(new_n7105));
  xnor_3 g06729(.A(new_n7105), .B(new_n7102), .Y(new_n7106));
  xnor_3 g06730(.A(new_n7106), .B(new_n7101), .Y(new_n7107));
  nor_4  g06731(.A(new_n7070), .B(new_n7069), .Y(new_n7108));
  nand_4 g06732(.A(n11757), .B(n4634), .Y(new_n7109));
  not_3  g06733(.A(new_n7109), .Y(new_n7110));
  xor_3  g06734(.A(new_n7110), .B(new_n7108), .Y(new_n7111));
  nand_4 g06735(.A(n11821), .B(n2879), .Y(new_n7112));
  not_3  g06736(.A(new_n7112), .Y(new_n7113));
  nand_4 g06737(.A(n10223), .B(n5240), .Y(new_n7114));
  nand_4 g06738(.A(n9080), .B(n7265), .Y(new_n7115));
  xnor_3 g06739(.A(new_n7115), .B(new_n7114), .Y(new_n7116));
  and_4  g06740(.A(new_n7116), .B(new_n7113), .Y(new_n7117));
  nor_4  g06741(.A(new_n7116), .B(new_n7113), .Y(new_n7118));
  nor_4  g06742(.A(new_n7118), .B(new_n7117), .Y(new_n7119));
  xnor_3 g06743(.A(new_n7119), .B(new_n7111), .Y(new_n7120));
  not_3  g06744(.A(new_n7120), .Y(new_n7121));
  xnor_3 g06745(.A(new_n7121), .B(new_n7107), .Y(new_n7122));
  nand_4 g06746(.A(new_n7065), .B(new_n7062), .Y(new_n7123));
  nor_4  g06747(.A(new_n7064), .B(new_n7063), .Y(new_n7124));
  nor_4  g06748(.A(new_n7079), .B(new_n7066), .Y(new_n7125));
  xnor_3 g06749(.A(new_n7125), .B(new_n7124), .Y(new_n7126));
  nand_4 g06750(.A(new_n7126), .B(new_n7123), .Y(new_n7127));
  xnor_3 g06751(.A(new_n7127), .B(new_n7122), .Y(new_n7128));
  xnor_3 g06752(.A(new_n7128), .B(new_n7098), .Y(new_n7129));
  nand_4 g06753(.A(n7862), .B(n2253), .Y(new_n7130));
  not_3  g06754(.A(new_n7130), .Y(new_n7131));
  xnor_3 g06755(.A(new_n7097), .B(new_n7080), .Y(new_n7132));
  nand_4 g06756(.A(new_n7132), .B(new_n7131), .Y(new_n7133));
  not_3  g06757(.A(new_n6318), .Y(new_n7134));
  nor_4  g06758(.A(new_n7134), .B(new_n6310), .Y(new_n7135));
  not_3  g06759(.A(new_n7135), .Y(new_n7136));
  xnor_3 g06760(.A(new_n7095), .B(new_n7091), .Y(new_n7137));
  nor_4  g06761(.A(new_n7137), .B(new_n7136), .Y(new_n7138));
  xnor_3 g06762(.A(new_n7132), .B(new_n7130), .Y(new_n7139));
  nand_4 g06763(.A(new_n7139), .B(new_n7138), .Y(new_n7140));
  nand_4 g06764(.A(new_n7140), .B(new_n7133), .Y(new_n7141));
  xor_3  g06765(.A(new_n7141), .B(new_n7129), .Y(new_n7142));
  not_3  g06766(.A(new_n7142), .Y(new_n7143));
  not_3  g06767(.A(new_n7138), .Y(new_n7144));
  xnor_3 g06768(.A(new_n7139), .B(new_n7144), .Y(new_n7145));
  not_3  g06769(.A(new_n7145), .Y(new_n7146));
  not_3  g06770(.A(new_n7137), .Y(new_n7147));
  xor_3  g06771(.A(new_n7147), .B(new_n7136), .Y(new_n7148));
  not_3  g06772(.A(new_n6355), .Y(new_n7149));
  nand_4 g06773(.A(n12145), .B(n6877), .Y(new_n7150));
  nand_4 g06774(.A(n9400), .B(n2522), .Y(new_n7151));
  not_3  g06775(.A(new_n7151), .Y(new_n7152));
  nand_4 g06776(.A(n11311), .B(n2024), .Y(new_n7153));
  not_3  g06777(.A(new_n7153), .Y(new_n7154));
  nand_4 g06778(.A(n9189), .B(n2464), .Y(new_n7155));
  nand_4 g06779(.A(n7946), .B(n4187), .Y(new_n7156));
  xnor_3 g06780(.A(new_n7156), .B(new_n7155), .Y(new_n7157));
  xnor_3 g06781(.A(new_n7157), .B(new_n7154), .Y(new_n7158));
  xnor_3 g06782(.A(new_n7158), .B(new_n7152), .Y(new_n7159_1));
  and_4  g06783(.A(new_n6323), .B(new_n6322), .Y(new_n7160_1));
  nor_4  g06784(.A(new_n6328), .B(new_n7160_1), .Y(new_n7161));
  xnor_3 g06785(.A(new_n7161), .B(new_n7159_1), .Y(new_n7162));
  xnor_3 g06786(.A(new_n7162), .B(new_n7150), .Y(new_n7163));
  nor_4  g06787(.A(new_n6329), .B(new_n6320), .Y(new_n7164));
  nor_4  g06788(.A(new_n6342), .B(new_n7164), .Y(new_n7165));
  not_3  g06789(.A(new_n7165), .Y(new_n7166));
  xnor_3 g06790(.A(new_n7166), .B(new_n7163), .Y(new_n7167));
  nor_4  g06791(.A(new_n7167), .B(new_n7149), .Y(new_n7168));
  not_3  g06792(.A(new_n7167), .Y(new_n7169));
  nor_4  g06793(.A(new_n7169), .B(new_n6355), .Y(new_n7170));
  nor_4  g06794(.A(new_n7170), .B(new_n7168), .Y(new_n7171));
  not_3  g06795(.A(new_n6442), .Y(new_n7172));
  nand_4 g06796(.A(new_n6497), .B(new_n7172), .Y(new_n7173));
  xnor_3 g06797(.A(new_n7173), .B(new_n7171), .Y(new_n7174));
  not_3  g06798(.A(new_n6466), .Y(new_n7175));
  nand_4 g06799(.A(n11478), .B(n521), .Y(new_n7176));
  not_3  g06800(.A(new_n7176), .Y(new_n7177));
  not_3  g06801(.A(new_n6456), .Y(new_n7178));
  not_3  g06802(.A(new_n6457), .Y(new_n7179));
  nor_4  g06803(.A(new_n7179), .B(new_n7178), .Y(new_n7180));
  not_3  g06804(.A(new_n6455), .Y(new_n7181));
  nor_4  g06805(.A(new_n6457), .B(new_n6456), .Y(new_n7182));
  nor_4  g06806(.A(new_n7182), .B(new_n7181), .Y(new_n7183));
  nor_4  g06807(.A(new_n7183), .B(new_n7180), .Y(new_n7184));
  xnor_3 g06808(.A(new_n7184), .B(new_n7177), .Y(new_n7185));
  nand_4 g06809(.A(n2498), .B(n137), .Y(new_n7186));
  not_3  g06810(.A(new_n7186), .Y(new_n7187));
  nand_4 g06811(.A(n5579), .B(n5283), .Y(new_n7188));
  not_3  g06812(.A(new_n7188), .Y(new_n7189));
  nand_4 g06813(.A(n6294), .B(n2558), .Y(new_n7190));
  not_3  g06814(.A(new_n7190), .Y(new_n7191));
  nor_4  g06815(.A(new_n7191), .B(new_n7189), .Y(new_n7192));
  not_3  g06816(.A(new_n7192), .Y(new_n7193_1));
  nor_4  g06817(.A(new_n7190), .B(new_n7188), .Y(new_n7194));
  not_3  g06818(.A(new_n7194), .Y(new_n7195));
  nand_4 g06819(.A(new_n7195), .B(new_n7193_1), .Y(new_n7196));
  xnor_3 g06820(.A(new_n7196), .B(new_n7187), .Y(new_n7197));
  xnor_3 g06821(.A(new_n7197), .B(new_n7185), .Y(new_n7198));
  not_3  g06822(.A(new_n7198), .Y(new_n7199));
  nand_4 g06823(.A(n6016), .B(n4805), .Y(new_n7200));
  not_3  g06824(.A(new_n7200), .Y(new_n7201));
  not_3  g06825(.A(new_n6451), .Y(new_n7202));
  nand_4 g06826(.A(new_n6460), .B(new_n6454), .Y(new_n7203));
  nand_4 g06827(.A(new_n7203), .B(new_n7202), .Y(new_n7204));
  nor_4  g06828(.A(new_n7204), .B(new_n7201), .Y(new_n7205));
  not_3  g06829(.A(new_n7204), .Y(new_n7206));
  nor_4  g06830(.A(new_n7206), .B(new_n7200), .Y(new_n7207));
  nor_4  g06831(.A(new_n7207), .B(new_n7205), .Y(new_n7208));
  nand_4 g06832(.A(new_n7208), .B(new_n7199), .Y(new_n7209));
  not_3  g06833(.A(new_n7209), .Y(new_n7210));
  nor_4  g06834(.A(new_n7208), .B(new_n7199), .Y(new_n7211));
  nor_4  g06835(.A(new_n7211), .B(new_n7210), .Y(new_n7212));
  xnor_3 g06836(.A(new_n7212), .B(new_n7175), .Y(new_n7213));
  not_3  g06837(.A(new_n6490), .Y(new_n7214));
  nand_4 g06838(.A(n7270), .B(n7236), .Y(new_n7215));
  not_3  g06839(.A(new_n7215), .Y(new_n7216));
  not_3  g06840(.A(new_n6473), .Y(new_n7217));
  nand_4 g06841(.A(new_n6482), .B(new_n6476), .Y(new_n7218));
  nand_4 g06842(.A(new_n7218), .B(new_n7217), .Y(new_n7219));
  nor_4  g06843(.A(new_n7219), .B(new_n7216), .Y(new_n7220));
  not_3  g06844(.A(new_n7219), .Y(new_n7221));
  nor_4  g06845(.A(new_n7221), .B(new_n7215), .Y(new_n7222));
  nor_4  g06846(.A(new_n7222), .B(new_n7220), .Y(new_n7223));
  nand_4 g06847(.A(n3992), .B(n806), .Y(new_n7224));
  not_3  g06848(.A(new_n7224), .Y(new_n7225));
  not_3  g06849(.A(new_n6478), .Y(new_n7226));
  not_3  g06850(.A(new_n6479), .Y(new_n7227));
  nor_4  g06851(.A(new_n7227), .B(new_n7226), .Y(new_n7228));
  not_3  g06852(.A(new_n6477), .Y(new_n7229));
  nor_4  g06853(.A(new_n6479), .B(new_n6478), .Y(new_n7230));
  nor_4  g06854(.A(new_n7230), .B(new_n7229), .Y(new_n7231));
  nor_4  g06855(.A(new_n7231), .B(new_n7228), .Y(new_n7232));
  nand_4 g06856(.A(new_n7232), .B(new_n7225), .Y(new_n7233));
  not_3  g06857(.A(new_n7233), .Y(new_n7234));
  nor_4  g06858(.A(new_n7232), .B(new_n7225), .Y(new_n7235));
  nor_4  g06859(.A(new_n7235), .B(new_n7234), .Y(new_n7236_1));
  not_3  g06860(.A(new_n7236_1), .Y(new_n7237));
  nand_4 g06861(.A(n9111), .B(n6358), .Y(new_n7238));
  nand_4 g06862(.A(n8384), .B(n3342), .Y(new_n7239));
  nand_4 g06863(.A(n9763), .B(n5198), .Y(new_n7240));
  xnor_3 g06864(.A(new_n7240), .B(new_n7239), .Y(new_n7241));
  xnor_3 g06865(.A(new_n7241), .B(new_n7238), .Y(new_n7242));
  xnor_3 g06866(.A(new_n7242), .B(new_n7237), .Y(new_n7243));
  nand_4 g06867(.A(new_n7243), .B(new_n7223), .Y(new_n7244));
  not_3  g06868(.A(new_n7244), .Y(new_n7245));
  nor_4  g06869(.A(new_n7243), .B(new_n7223), .Y(new_n7246));
  nor_4  g06870(.A(new_n7246), .B(new_n7245), .Y(new_n7247));
  xnor_3 g06871(.A(new_n7247), .B(new_n7214), .Y(new_n7248));
  xnor_3 g06872(.A(new_n7248), .B(new_n7213), .Y(new_n7249));
  nor_4  g06873(.A(new_n6491), .B(new_n6467), .Y(new_n7250));
  nor_4  g06874(.A(new_n6494), .B(new_n6492), .Y(new_n7251));
  nor_4  g06875(.A(new_n7251), .B(new_n7250), .Y(new_n7252));
  xnor_3 g06876(.A(new_n7252), .B(new_n7249), .Y(new_n7253));
  xnor_3 g06877(.A(new_n7253), .B(new_n7174), .Y(new_n7254));
  not_3  g06878(.A(new_n7254), .Y(new_n7255));
  nand_4 g06879(.A(new_n7255), .B(new_n7148), .Y(new_n7256));
  xnor_3 g06880(.A(new_n7254), .B(new_n7148), .Y(new_n7257));
  nand_4 g06881(.A(new_n6526), .B(new_n6502), .Y(new_n7258));
  nand_4 g06882(.A(new_n7258), .B(new_n6501), .Y(new_n7259));
  nand_4 g06883(.A(new_n7259), .B(new_n7257), .Y(new_n7260));
  nand_4 g06884(.A(new_n7260), .B(new_n7256), .Y(new_n7261));
  nand_4 g06885(.A(new_n7261), .B(new_n7146), .Y(new_n7262));
  nor_4  g06886(.A(new_n7247), .B(new_n7214), .Y(new_n7263));
  not_3  g06887(.A(new_n7263), .Y(new_n7264));
  nand_4 g06888(.A(n7236), .B(n5153), .Y(new_n7265_1));
  nand_4 g06889(.A(n6358), .B(n3342), .Y(new_n7266));
  nand_4 g06890(.A(n9111), .B(n5198), .Y(new_n7267));
  nand_4 g06891(.A(n9763), .B(n1471), .Y(new_n7268));
  xnor_3 g06892(.A(new_n7268), .B(new_n7267), .Y(new_n7269));
  nor_4  g06893(.A(new_n7269), .B(new_n7266), .Y(new_n7270_1));
  not_3  g06894(.A(new_n7266), .Y(new_n7271));
  not_3  g06895(.A(new_n7269), .Y(new_n7272));
  nor_4  g06896(.A(new_n7272), .B(new_n7271), .Y(new_n7273));
  nor_4  g06897(.A(new_n7273), .B(new_n7270_1), .Y(new_n7274));
  and_4  g06898(.A(new_n7240), .B(new_n7239), .Y(new_n7275));
  not_3  g06899(.A(new_n7238), .Y(new_n7276));
  nor_4  g06900(.A(new_n7241), .B(new_n7276), .Y(new_n7277));
  nor_4  g06901(.A(new_n7277), .B(new_n7275), .Y(new_n7278));
  xnor_3 g06902(.A(new_n7278), .B(new_n7274), .Y(new_n7279));
  nand_4 g06903(.A(n7270), .B(n3992), .Y(new_n7280));
  nand_4 g06904(.A(n8384), .B(n806), .Y(new_n7281));
  not_3  g06905(.A(new_n7281), .Y(new_n7282));
  xor_3  g06906(.A(new_n7282), .B(new_n7280), .Y(new_n7283));
  xnor_3 g06907(.A(new_n7283), .B(new_n7279), .Y(new_n7284));
  nor_4  g06908(.A(new_n7242), .B(new_n7237), .Y(new_n7285));
  nor_4  g06909(.A(new_n7285), .B(new_n7234), .Y(new_n7286));
  xnor_3 g06910(.A(new_n7286), .B(new_n7284), .Y(new_n7287));
  not_3  g06911(.A(new_n7220), .Y(new_n7288));
  nand_4 g06912(.A(new_n7244), .B(new_n7288), .Y(new_n7289));
  xnor_3 g06913(.A(new_n7289), .B(new_n7287), .Y(new_n7290));
  xnor_3 g06914(.A(new_n7290), .B(new_n7265_1), .Y(new_n7291));
  xnor_3 g06915(.A(new_n7291), .B(new_n7264), .Y(new_n7292));
  nor_4  g06916(.A(new_n7212), .B(new_n7175), .Y(new_n7293));
  nand_4 g06917(.A(n5798), .B(n4805), .Y(new_n7294_1));
  nand_4 g06918(.A(n5579), .B(n137), .Y(new_n7295));
  nand_4 g06919(.A(n6797), .B(n2558), .Y(new_n7296));
  nand_4 g06920(.A(n6294), .B(n2498), .Y(new_n7297));
  xnor_3 g06921(.A(new_n7297), .B(new_n7296), .Y(new_n7298));
  nor_4  g06922(.A(new_n7298), .B(new_n7295), .Y(new_n7299));
  not_3  g06923(.A(new_n7295), .Y(new_n7300));
  not_3  g06924(.A(new_n7298), .Y(new_n7301));
  nor_4  g06925(.A(new_n7301), .B(new_n7300), .Y(new_n7302));
  nor_4  g06926(.A(new_n7302), .B(new_n7299), .Y(new_n7303));
  nor_4  g06927(.A(new_n7194), .B(new_n7187), .Y(new_n7304));
  nor_4  g06928(.A(new_n7304), .B(new_n7192), .Y(new_n7305));
  xnor_3 g06929(.A(new_n7305), .B(new_n7303), .Y(new_n7306));
  nand_4 g06930(.A(n11478), .B(n6016), .Y(new_n7307));
  nand_4 g06931(.A(n5283), .B(n521), .Y(new_n7308));
  xor_3  g06932(.A(new_n7308), .B(new_n7307), .Y(new_n7309));
  xnor_3 g06933(.A(new_n7309), .B(new_n7306), .Y(new_n7310));
  and_4  g06934(.A(new_n7184), .B(new_n7177), .Y(new_n7311));
  not_3  g06935(.A(new_n7197), .Y(new_n7312));
  nor_4  g06936(.A(new_n7312), .B(new_n7185), .Y(new_n7313));
  nor_4  g06937(.A(new_n7313), .B(new_n7311), .Y(new_n7314));
  xnor_3 g06938(.A(new_n7314), .B(new_n7310), .Y(new_n7315));
  not_3  g06939(.A(new_n7205), .Y(new_n7316));
  nand_4 g06940(.A(new_n7209), .B(new_n7316), .Y(new_n7317));
  xnor_3 g06941(.A(new_n7317), .B(new_n7315), .Y(new_n7318));
  not_3  g06942(.A(new_n7318), .Y(new_n7319));
  nand_4 g06943(.A(new_n7319), .B(new_n7294_1), .Y(new_n7320_1));
  not_3  g06944(.A(new_n7294_1), .Y(new_n7321));
  nand_4 g06945(.A(new_n7318), .B(new_n7321), .Y(new_n7322));
  nand_4 g06946(.A(new_n7322), .B(new_n7320_1), .Y(new_n7323));
  xnor_3 g06947(.A(new_n7323), .B(new_n7293), .Y(new_n7324));
  xnor_3 g06948(.A(new_n7324), .B(new_n7292), .Y(new_n7325));
  nand_4 g06949(.A(new_n7248), .B(new_n7213), .Y(new_n7326));
  not_3  g06950(.A(new_n7326), .Y(new_n7327));
  nor_4  g06951(.A(new_n7252), .B(new_n7249), .Y(new_n7328));
  nor_4  g06952(.A(new_n7328), .B(new_n7327), .Y(new_n7329));
  not_3  g06953(.A(new_n7329), .Y(new_n7330));
  nand_4 g06954(.A(new_n7330), .B(new_n7325), .Y(new_n7331));
  not_3  g06955(.A(new_n7331), .Y(new_n7332));
  nor_4  g06956(.A(new_n7330), .B(new_n7325), .Y(new_n7333));
  nor_4  g06957(.A(new_n7333), .B(new_n7332), .Y(new_n7334));
  nor_4  g06958(.A(new_n7173), .B(new_n7171), .Y(new_n7335));
  not_3  g06959(.A(new_n7335), .Y(new_n7336));
  not_3  g06960(.A(new_n7174), .Y(new_n7337));
  not_3  g06961(.A(new_n7253), .Y(new_n7338));
  nand_4 g06962(.A(new_n7338), .B(new_n7337), .Y(new_n7339));
  nand_4 g06963(.A(new_n7339), .B(new_n7336), .Y(new_n7340));
  not_3  g06964(.A(new_n7340), .Y(new_n7341));
  nand_4 g06965(.A(n12221), .B(n6877), .Y(new_n7342));
  not_3  g06966(.A(new_n7342), .Y(new_n7343));
  not_3  g06967(.A(new_n7150), .Y(new_n7344));
  nand_4 g06968(.A(new_n7162), .B(new_n7344), .Y(new_n7345));
  nand_4 g06969(.A(new_n7166), .B(new_n7163), .Y(new_n7346));
  nand_4 g06970(.A(new_n7346), .B(new_n7345), .Y(new_n7347));
  nor_4  g06971(.A(new_n7158), .B(new_n7152), .Y(new_n7348));
  nor_4  g06972(.A(new_n7161), .B(new_n7159_1), .Y(new_n7349));
  nor_4  g06973(.A(new_n7349), .B(new_n7348), .Y(new_n7350));
  not_3  g06974(.A(new_n7350), .Y(new_n7351));
  nand_4 g06975(.A(n11311), .B(n9189), .Y(new_n7352));
  not_3  g06976(.A(new_n7352), .Y(new_n7353));
  nand_4 g06977(.A(n4187), .B(n2024), .Y(new_n7354_1));
  nand_4 g06978(.A(n7946), .B(n4203), .Y(new_n7355));
  not_3  g06979(.A(new_n7355), .Y(new_n7356));
  xor_3  g06980(.A(new_n7356), .B(new_n7354_1), .Y(new_n7357));
  xnor_3 g06981(.A(new_n7357), .B(new_n7353), .Y(new_n7358));
  and_4  g06982(.A(new_n7156), .B(new_n7155), .Y(new_n7359));
  nor_4  g06983(.A(new_n7156), .B(new_n7155), .Y(new_n7360));
  nor_4  g06984(.A(new_n7360), .B(new_n7154), .Y(new_n7361));
  nor_4  g06985(.A(new_n7361), .B(new_n7359), .Y(new_n7362));
  not_3  g06986(.A(new_n7362), .Y(new_n7363));
  xnor_3 g06987(.A(new_n7363), .B(new_n7358), .Y(new_n7364));
  nand_4 g06988(.A(n12145), .B(n9400), .Y(new_n7365));
  nand_4 g06989(.A(n2522), .B(n2464), .Y(new_n7366));
  xor_3  g06990(.A(new_n7366), .B(new_n7365), .Y(new_n7367));
  xnor_3 g06991(.A(new_n7367), .B(new_n7364), .Y(new_n7368));
  xnor_3 g06992(.A(new_n7368), .B(new_n7351), .Y(new_n7369));
  xnor_3 g06993(.A(new_n7369), .B(new_n7347), .Y(new_n7370));
  xnor_3 g06994(.A(new_n7370), .B(new_n7343), .Y(new_n7371));
  xnor_3 g06995(.A(new_n7371), .B(new_n7168), .Y(new_n7372));
  xnor_3 g06996(.A(new_n7372), .B(new_n7341), .Y(new_n7373));
  xnor_3 g06997(.A(new_n7373), .B(new_n7334), .Y(new_n7374));
  xnor_3 g06998(.A(new_n7261), .B(new_n7145), .Y(new_n7375));
  nand_4 g06999(.A(new_n7375), .B(new_n7374), .Y(new_n7376));
  nand_4 g07000(.A(new_n7376), .B(new_n7262), .Y(new_n7377));
  nand_4 g07001(.A(new_n7377), .B(new_n7143), .Y(new_n7378));
  xnor_3 g07002(.A(new_n7377), .B(new_n7142), .Y(new_n7379));
  xnor_3 g07003(.A(new_n7368), .B(new_n7350), .Y(new_n7380));
  nand_4 g07004(.A(new_n7380), .B(new_n7347), .Y(new_n7381));
  nand_4 g07005(.A(new_n7357), .B(new_n7352), .Y(new_n7382));
  nand_4 g07006(.A(new_n7363), .B(new_n7358), .Y(new_n7383));
  nand_4 g07007(.A(new_n7383), .B(new_n7382), .Y(new_n7384));
  nand_4 g07008(.A(n12221), .B(n9400), .Y(new_n7385));
  not_3  g07009(.A(new_n7385), .Y(new_n7386));
  nand_4 g07010(.A(n12145), .B(n2464), .Y(new_n7387));
  nand_4 g07011(.A(n10217), .B(n6877), .Y(new_n7388_1));
  not_3  g07012(.A(new_n7388_1), .Y(new_n7389));
  xor_3  g07013(.A(new_n7389), .B(new_n7387), .Y(new_n7390));
  xnor_3 g07014(.A(new_n7390), .B(new_n7386), .Y(new_n7391));
  xnor_3 g07015(.A(new_n7391), .B(new_n7384), .Y(new_n7392));
  nor_4  g07016(.A(new_n7355), .B(new_n7354_1), .Y(new_n7393));
  nand_4 g07017(.A(n11311), .B(n2522), .Y(new_n7394));
  not_3  g07018(.A(new_n7394), .Y(new_n7395));
  xor_3  g07019(.A(new_n7395), .B(new_n7393), .Y(new_n7396));
  nand_4 g07020(.A(n4203), .B(n2024), .Y(new_n7397));
  nand_4 g07021(.A(n9189), .B(n4187), .Y(new_n7398));
  not_3  g07022(.A(new_n7398), .Y(new_n7399));
  nand_4 g07023(.A(n12753), .B(n7946), .Y(new_n7400));
  not_3  g07024(.A(new_n7400), .Y(new_n7401));
  nand_4 g07025(.A(new_n7401), .B(new_n7399), .Y(new_n7402));
  nand_4 g07026(.A(new_n7400), .B(new_n7398), .Y(new_n7403));
  nand_4 g07027(.A(new_n7403), .B(new_n7402), .Y(new_n7404));
  xor_3  g07028(.A(new_n7404), .B(new_n7397), .Y(new_n7405));
  xnor_3 g07029(.A(new_n7405), .B(new_n7396), .Y(new_n7406));
  xnor_3 g07030(.A(new_n7406), .B(new_n7392), .Y(new_n7407));
  nand_4 g07031(.A(new_n7367), .B(new_n7364), .Y(new_n7408));
  nor_4  g07032(.A(new_n7366), .B(new_n7365), .Y(new_n7409));
  nor_4  g07033(.A(new_n7367), .B(new_n7364), .Y(new_n7410));
  nor_4  g07034(.A(new_n7410), .B(new_n7351), .Y(new_n7411));
  xnor_3 g07035(.A(new_n7411), .B(new_n7409), .Y(new_n7412));
  nand_4 g07036(.A(new_n7412), .B(new_n7408), .Y(new_n7413));
  xnor_3 g07037(.A(new_n7413), .B(new_n7407), .Y(new_n7414));
  xnor_3 g07038(.A(new_n7414), .B(new_n7381), .Y(new_n7415));
  xnor_3 g07039(.A(new_n7380), .B(new_n7347), .Y(new_n7416));
  nor_4  g07040(.A(new_n7416), .B(new_n7342), .Y(new_n7417));
  not_3  g07041(.A(new_n7168), .Y(new_n7418));
  nor_4  g07042(.A(new_n7371), .B(new_n7418), .Y(new_n7419));
  nor_4  g07043(.A(new_n7419), .B(new_n7417), .Y(new_n7420));
  xnor_3 g07044(.A(new_n7420), .B(new_n7415), .Y(new_n7421));
  not_3  g07045(.A(new_n7317), .Y(new_n7422));
  nand_4 g07046(.A(new_n7422), .B(new_n7315), .Y(new_n7423));
  nand_4 g07047(.A(n4805), .B(n2347), .Y(new_n7424));
  nand_4 g07048(.A(n6016), .B(n5283), .Y(new_n7425));
  nand_4 g07049(.A(n11478), .B(n5798), .Y(new_n7426));
  not_3  g07050(.A(new_n7426), .Y(new_n7427));
  xor_3  g07051(.A(new_n7427), .B(new_n7425), .Y(new_n7428));
  xnor_3 g07052(.A(new_n7428), .B(new_n7424), .Y(new_n7429));
  nand_4 g07053(.A(new_n7305), .B(new_n7303), .Y(new_n7430));
  not_3  g07054(.A(new_n7430), .Y(new_n7431));
  nor_4  g07055(.A(new_n7431), .B(new_n7299), .Y(new_n7432));
  not_3  g07056(.A(new_n7432), .Y(new_n7433));
  xnor_3 g07057(.A(new_n7433), .B(new_n7429), .Y(new_n7434));
  nor_4  g07058(.A(new_n7297), .B(new_n7296), .Y(new_n7435));
  nand_4 g07059(.A(n521), .B(n137), .Y(new_n7436_1));
  xor_3  g07060(.A(new_n7436_1), .B(new_n7435), .Y(new_n7437));
  nand_4 g07061(.A(n6797), .B(n2498), .Y(new_n7438));
  nand_4 g07062(.A(n6294), .B(n5579), .Y(new_n7439));
  nand_4 g07063(.A(n3146), .B(n2558), .Y(new_n7440));
  not_3  g07064(.A(new_n7440), .Y(new_n7441));
  xor_3  g07065(.A(new_n7441), .B(new_n7439), .Y(new_n7442));
  xnor_3 g07066(.A(new_n7442), .B(new_n7438), .Y(new_n7443));
  xnor_3 g07067(.A(new_n7443), .B(new_n7437), .Y(new_n7444));
  xnor_3 g07068(.A(new_n7444), .B(new_n7434), .Y(new_n7445));
  not_3  g07069(.A(new_n7306), .Y(new_n7446));
  nand_4 g07070(.A(new_n7309), .B(new_n7446), .Y(new_n7447));
  nor_4  g07071(.A(new_n7308), .B(new_n7307), .Y(new_n7448));
  not_3  g07072(.A(new_n7310), .Y(new_n7449));
  nor_4  g07073(.A(new_n7314), .B(new_n7449), .Y(new_n7450));
  xnor_3 g07074(.A(new_n7450), .B(new_n7448), .Y(new_n7451));
  nand_4 g07075(.A(new_n7451), .B(new_n7447), .Y(new_n7452));
  xnor_3 g07076(.A(new_n7452), .B(new_n7445), .Y(new_n7453));
  xnor_3 g07077(.A(new_n7453), .B(new_n7423), .Y(new_n7454));
  nand_4 g07078(.A(new_n7320_1), .B(new_n7293), .Y(new_n7455));
  nand_4 g07079(.A(new_n7455), .B(new_n7322), .Y(new_n7456_1));
  xnor_3 g07080(.A(new_n7456_1), .B(new_n7454), .Y(new_n7457));
  nor_4  g07081(.A(new_n7289), .B(new_n7287), .Y(new_n7458));
  not_3  g07082(.A(new_n7458), .Y(new_n7459));
  not_3  g07083(.A(new_n7279), .Y(new_n7460));
  not_3  g07084(.A(new_n7283), .Y(new_n7461));
  nand_4 g07085(.A(new_n7461), .B(new_n7460), .Y(new_n7462));
  nor_4  g07086(.A(new_n7281), .B(new_n7280), .Y(new_n7463));
  nor_4  g07087(.A(new_n7286), .B(new_n7284), .Y(new_n7464));
  xnor_3 g07088(.A(new_n7464), .B(new_n7463), .Y(new_n7465));
  nand_4 g07089(.A(new_n7465), .B(new_n7462), .Y(new_n7466));
  nor_4  g07090(.A(new_n7268), .B(new_n7267), .Y(new_n7467));
  nand_4 g07091(.A(n6358), .B(n806), .Y(new_n7468));
  not_3  g07092(.A(new_n7468), .Y(new_n7469));
  xor_3  g07093(.A(new_n7469), .B(new_n7467), .Y(new_n7470));
  nand_4 g07094(.A(n9111), .B(n1471), .Y(new_n7471));
  nand_4 g07095(.A(n5198), .B(n3342), .Y(new_n7472));
  nand_4 g07096(.A(n9763), .B(n7646), .Y(new_n7473));
  nand_4 g07097(.A(new_n7473), .B(new_n7472), .Y(new_n7474));
  not_3  g07098(.A(new_n7472), .Y(new_n7475));
  not_3  g07099(.A(new_n7473), .Y(new_n7476));
  nand_4 g07100(.A(new_n7476), .B(new_n7475), .Y(new_n7477));
  nand_4 g07101(.A(new_n7477), .B(new_n7474), .Y(new_n7478));
  xor_3  g07102(.A(new_n7478), .B(new_n7471), .Y(new_n7479));
  xnor_3 g07103(.A(new_n7479), .B(new_n7470), .Y(new_n7480));
  not_3  g07104(.A(new_n7480), .Y(new_n7481));
  not_3  g07105(.A(new_n7270_1), .Y(new_n7482));
  nand_4 g07106(.A(new_n7278), .B(new_n7274), .Y(new_n7483));
  nand_4 g07107(.A(new_n7483), .B(new_n7482), .Y(new_n7484));
  nand_4 g07108(.A(n5153), .B(n3992), .Y(new_n7485));
  nand_4 g07109(.A(n8384), .B(n7270), .Y(new_n7486));
  nand_4 g07110(.A(n7236), .B(n2507), .Y(new_n7487));
  not_3  g07111(.A(new_n7487), .Y(new_n7488));
  xor_3  g07112(.A(new_n7488), .B(new_n7486), .Y(new_n7489));
  xnor_3 g07113(.A(new_n7489), .B(new_n7485), .Y(new_n7490));
  xnor_3 g07114(.A(new_n7490), .B(new_n7484), .Y(new_n7491));
  xnor_3 g07115(.A(new_n7491), .B(new_n7481), .Y(new_n7492));
  xnor_3 g07116(.A(new_n7492), .B(new_n7466), .Y(new_n7493));
  xnor_3 g07117(.A(new_n7493), .B(new_n7459), .Y(new_n7494));
  nor_4  g07118(.A(new_n7290), .B(new_n7265_1), .Y(new_n7495));
  not_3  g07119(.A(new_n7495), .Y(new_n7496));
  nand_4 g07120(.A(new_n7290), .B(new_n7265_1), .Y(new_n7497));
  nand_4 g07121(.A(new_n7497), .B(new_n7263), .Y(new_n7498));
  nand_4 g07122(.A(new_n7498), .B(new_n7496), .Y(new_n7499));
  xnor_3 g07123(.A(new_n7499), .B(new_n7494), .Y(new_n7500_1));
  xnor_3 g07124(.A(new_n7500_1), .B(new_n7457), .Y(new_n7501));
  not_3  g07125(.A(new_n7324), .Y(new_n7502));
  nand_4 g07126(.A(new_n7502), .B(new_n7292), .Y(new_n7503));
  nand_4 g07127(.A(new_n7331), .B(new_n7503), .Y(new_n7504));
  xnor_3 g07128(.A(new_n7504), .B(new_n7501), .Y(new_n7505));
  xnor_3 g07129(.A(new_n7505), .B(new_n7421), .Y(new_n7506));
  nand_4 g07130(.A(new_n7372), .B(new_n7341), .Y(new_n7507));
  not_3  g07131(.A(new_n7334), .Y(new_n7508));
  not_3  g07132(.A(new_n7373), .Y(new_n7509));
  nand_4 g07133(.A(new_n7509), .B(new_n7508), .Y(new_n7510));
  nand_4 g07134(.A(new_n7510), .B(new_n7507), .Y(new_n7511));
  xnor_3 g07135(.A(new_n7511), .B(new_n7506), .Y(new_n7512));
  nand_4 g07136(.A(new_n7512), .B(new_n7379), .Y(new_n7513));
  nand_4 g07137(.A(new_n7513), .B(new_n7378), .Y(new_n7514));
  not_3  g07138(.A(new_n7421), .Y(new_n7515));
  nand_4 g07139(.A(new_n7505), .B(new_n7515), .Y(new_n7516));
  nand_4 g07140(.A(new_n7511), .B(new_n7506), .Y(new_n7517));
  nand_4 g07141(.A(new_n7517), .B(new_n7516), .Y(new_n7518));
  nor_4  g07142(.A(new_n7453), .B(new_n7423), .Y(new_n7519));
  not_3  g07143(.A(new_n7456_1), .Y(new_n7520));
  nor_4  g07144(.A(new_n7520), .B(new_n7454), .Y(new_n7521));
  nor_4  g07145(.A(new_n7521), .B(new_n7519), .Y(new_n7522));
  xnor_3 g07146(.A(new_n7522), .B(new_n7518), .Y(new_n7523_1));
  not_3  g07147(.A(new_n7457), .Y(new_n7524));
  nand_4 g07148(.A(new_n7500_1), .B(new_n7524), .Y(new_n7525));
  nand_4 g07149(.A(new_n7504), .B(new_n7501), .Y(new_n7526));
  nand_4 g07150(.A(new_n7526), .B(new_n7525), .Y(new_n7527));
  nand_4 g07151(.A(new_n7432), .B(new_n7429), .Y(new_n7528));
  nand_4 g07152(.A(new_n7444), .B(new_n7434), .Y(new_n7529));
  nand_4 g07153(.A(new_n7529), .B(new_n7528), .Y(new_n7530));
  nand_4 g07154(.A(n11478), .B(n2347), .Y(new_n7531));
  not_3  g07155(.A(new_n7531), .Y(new_n7532));
  xnor_3 g07156(.A(new_n7532), .B(new_n7530), .Y(new_n7533));
  nand_4 g07157(.A(n3342), .B(n1471), .Y(new_n7534));
  not_3  g07158(.A(new_n7534), .Y(new_n7535));
  not_3  g07159(.A(new_n7435), .Y(new_n7536));
  nor_4  g07160(.A(new_n7436_1), .B(new_n7536), .Y(new_n7537));
  nor_4  g07161(.A(new_n7443), .B(new_n7437), .Y(new_n7538));
  nor_4  g07162(.A(new_n7538), .B(new_n7537), .Y(new_n7539));
  not_3  g07163(.A(new_n7387), .Y(new_n7540));
  nor_4  g07164(.A(new_n7389), .B(new_n7540), .Y(new_n7541));
  nor_4  g07165(.A(new_n7390), .B(new_n7386), .Y(new_n7542));
  nor_4  g07166(.A(new_n7542), .B(new_n7541), .Y(new_n7543));
  nand_4 g07167(.A(n7236), .B(n6431), .Y(new_n7544));
  not_3  g07168(.A(new_n7544), .Y(new_n7545));
  nand_4 g07169(.A(n9111), .B(n7646), .Y(new_n7546_1));
  nand_4 g07170(.A(n9763), .B(n4722), .Y(new_n7547));
  xor_3  g07171(.A(new_n7547), .B(new_n7546_1), .Y(new_n7548));
  xnor_3 g07172(.A(new_n7548), .B(new_n7545), .Y(new_n7549));
  xnor_3 g07173(.A(new_n7549), .B(new_n7543), .Y(new_n7550));
  xnor_3 g07174(.A(new_n7550), .B(new_n7539), .Y(new_n7551));
  xnor_3 g07175(.A(new_n7551), .B(new_n7535), .Y(new_n7552));
  not_3  g07176(.A(new_n7391), .Y(new_n7553));
  nand_4 g07177(.A(new_n7553), .B(new_n7384), .Y(new_n7554));
  nand_4 g07178(.A(new_n7406), .B(new_n7392), .Y(new_n7555));
  nand_4 g07179(.A(new_n7555), .B(new_n7554), .Y(new_n7556));
  nand_4 g07180(.A(new_n7395), .B(new_n7393), .Y(new_n7557));
  nand_4 g07181(.A(new_n7405), .B(new_n7396), .Y(new_n7558));
  nand_4 g07182(.A(new_n7558), .B(new_n7557), .Y(new_n7559));
  nand_4 g07183(.A(n10217), .B(n9400), .Y(new_n7560));
  not_3  g07184(.A(new_n7560), .Y(new_n7561));
  xnor_3 g07185(.A(new_n7561), .B(new_n7559), .Y(new_n7562));
  nand_4 g07186(.A(n9189), .B(n4203), .Y(new_n7563));
  not_3  g07187(.A(new_n7563), .Y(new_n7564));
  nand_4 g07188(.A(n4187), .B(n2522), .Y(new_n7565));
  nand_4 g07189(.A(n12145), .B(n11311), .Y(new_n7566));
  xor_3  g07190(.A(new_n7566), .B(new_n7565), .Y(new_n7567));
  xnor_3 g07191(.A(new_n7567), .B(new_n7564), .Y(new_n7568_1));
  nand_4 g07192(.A(n7823), .B(n6877), .Y(new_n7569));
  nand_4 g07193(.A(n12753), .B(n2024), .Y(new_n7570));
  not_3  g07194(.A(new_n7570), .Y(new_n7571));
  xor_3  g07195(.A(new_n7571), .B(new_n7569), .Y(new_n7572));
  xnor_3 g07196(.A(new_n7572), .B(new_n7568_1), .Y(new_n7573));
  not_3  g07197(.A(new_n7397), .Y(new_n7574));
  nand_4 g07198(.A(new_n7403), .B(new_n7574), .Y(new_n7575));
  and_4  g07199(.A(new_n7575), .B(new_n7402), .Y(new_n7576));
  nand_4 g07200(.A(n10174), .B(n7946), .Y(new_n7577));
  nand_4 g07201(.A(n12221), .B(n2464), .Y(new_n7578));
  xor_3  g07202(.A(new_n7578), .B(new_n7577), .Y(new_n7579));
  xnor_3 g07203(.A(new_n7579), .B(new_n7576), .Y(new_n7580));
  xnor_3 g07204(.A(new_n7580), .B(new_n7573), .Y(new_n7581));
  xnor_3 g07205(.A(new_n7581), .B(new_n7562), .Y(new_n7582));
  xnor_3 g07206(.A(new_n7582), .B(new_n7556), .Y(new_n7583));
  xnor_3 g07207(.A(new_n7583), .B(new_n7552), .Y(new_n7584));
  xnor_3 g07208(.A(new_n7584), .B(new_n7533), .Y(new_n7585));
  nand_4 g07209(.A(new_n7464), .B(new_n7463), .Y(new_n7586));
  not_3  g07210(.A(new_n7492), .Y(new_n7587));
  nand_4 g07211(.A(new_n7587), .B(new_n7466), .Y(new_n7588));
  nand_4 g07212(.A(new_n7588), .B(new_n7586), .Y(new_n7589));
  nand_4 g07213(.A(new_n7411), .B(new_n7409), .Y(new_n7590));
  nand_4 g07214(.A(new_n7413), .B(new_n7407), .Y(new_n7591));
  nand_4 g07215(.A(new_n7591), .B(new_n7590), .Y(new_n7592));
  xnor_3 g07216(.A(new_n7592), .B(new_n7589), .Y(new_n7593));
  xnor_3 g07217(.A(new_n7593), .B(new_n7585), .Y(new_n7594));
  not_3  g07218(.A(new_n7439), .Y(new_n7595));
  nor_4  g07219(.A(new_n7441), .B(new_n7595), .Y(new_n7596));
  not_3  g07220(.A(new_n7438), .Y(new_n7597));
  nor_4  g07221(.A(new_n7442), .B(new_n7597), .Y(new_n7598));
  or_4   g07222(.A(new_n7598), .B(new_n7596), .Y(new_n7599));
  nand_4 g07223(.A(new_n7493), .B(new_n7458), .Y(new_n7600));
  nand_4 g07224(.A(new_n7499), .B(new_n7494), .Y(new_n7601));
  nand_4 g07225(.A(new_n7601), .B(new_n7600), .Y(new_n7602));
  xnor_3 g07226(.A(new_n7602), .B(new_n7599), .Y(new_n7603));
  xnor_3 g07227(.A(new_n7603), .B(new_n7594), .Y(new_n7604));
  xnor_3 g07228(.A(new_n7604), .B(new_n7527), .Y(new_n7605));
  nor_4  g07229(.A(new_n7414), .B(new_n7381), .Y(new_n7606));
  nor_4  g07230(.A(new_n7420), .B(new_n7415), .Y(new_n7607));
  nor_4  g07231(.A(new_n7607), .B(new_n7606), .Y(new_n7608));
  not_3  g07232(.A(new_n7098), .Y(new_n7609));
  nand_4 g07233(.A(new_n7128), .B(new_n7609), .Y(new_n7610_1));
  nand_4 g07234(.A(new_n7141), .B(new_n7129), .Y(new_n7611));
  nand_4 g07235(.A(new_n7611), .B(new_n7610_1), .Y(new_n7612));
  nand_4 g07236(.A(new_n7125), .B(new_n7124), .Y(new_n7613));
  not_3  g07237(.A(new_n7122), .Y(new_n7614));
  nand_4 g07238(.A(new_n7127), .B(new_n7614), .Y(new_n7615));
  nand_4 g07239(.A(new_n7615), .B(new_n7613), .Y(new_n7616));
  not_3  g07240(.A(new_n7425), .Y(new_n7617));
  nor_4  g07241(.A(new_n7427), .B(new_n7617), .Y(new_n7618));
  not_3  g07242(.A(new_n7424), .Y(new_n7619));
  nor_4  g07243(.A(new_n7428), .B(new_n7619), .Y(new_n7620));
  nor_4  g07244(.A(new_n7620), .B(new_n7618), .Y(new_n7621));
  nor_4  g07245(.A(new_n7106), .B(new_n7101), .Y(new_n7622));
  nor_4  g07246(.A(new_n7120), .B(new_n7107), .Y(new_n7623));
  nor_4  g07247(.A(new_n7623), .B(new_n7622), .Y(new_n7624));
  nand_4 g07248(.A(n7862), .B(n2512), .Y(new_n7625));
  not_3  g07249(.A(new_n7108), .Y(new_n7626));
  nand_4 g07250(.A(new_n7109), .B(new_n7626), .Y(new_n7627));
  nand_4 g07251(.A(new_n7119), .B(new_n7111), .Y(new_n7628));
  nand_4 g07252(.A(new_n7628), .B(new_n7627), .Y(new_n7629));
  xnor_3 g07253(.A(new_n7629), .B(new_n7625), .Y(new_n7630));
  nor_4  g07254(.A(new_n7104), .B(new_n7103), .Y(new_n7631));
  not_3  g07255(.A(new_n7102), .Y(new_n7632));
  nand_4 g07256(.A(new_n7104), .B(new_n7103), .Y(new_n7633));
  nand_4 g07257(.A(new_n7633), .B(new_n7632), .Y(new_n7634));
  not_3  g07258(.A(new_n7634), .Y(new_n7635));
  nor_4  g07259(.A(new_n7635), .B(new_n7631), .Y(new_n7636));
  nand_4 g07260(.A(n11821), .B(n10223), .Y(new_n7637));
  nand_4 g07261(.A(n5240), .B(n4634), .Y(new_n7638));
  nand_4 g07262(.A(n9080), .B(n2879), .Y(new_n7639));
  xnor_3 g07263(.A(new_n7639), .B(new_n7638), .Y(new_n7640));
  and_4  g07264(.A(new_n7640), .B(new_n7637), .Y(new_n7641));
  nor_4  g07265(.A(new_n7640), .B(new_n7637), .Y(new_n7642));
  nor_4  g07266(.A(new_n7642), .B(new_n7641), .Y(new_n7643));
  xnor_3 g07267(.A(new_n7643), .B(new_n7636), .Y(new_n7644));
  and_4  g07268(.A(new_n7115), .B(new_n7114), .Y(new_n7645));
  nor_4  g07269(.A(new_n7118), .B(new_n7645), .Y(new_n7646_1));
  nand_4 g07270(.A(n11757), .B(n9195), .Y(new_n7647));
  not_3  g07271(.A(new_n7647), .Y(new_n7648));
  nand_4 g07272(.A(n3172), .B(n2253), .Y(new_n7649));
  nand_4 g07273(.A(n3865), .B(n1333), .Y(new_n7650));
  xnor_3 g07274(.A(new_n7650), .B(new_n7649), .Y(new_n7651));
  xnor_3 g07275(.A(new_n7651), .B(new_n7648), .Y(new_n7652));
  xnor_3 g07276(.A(new_n7652), .B(new_n7646_1), .Y(new_n7653));
  xnor_3 g07277(.A(new_n7653), .B(new_n7644), .Y(new_n7654));
  xnor_3 g07278(.A(new_n7654), .B(new_n7630), .Y(new_n7655));
  xnor_3 g07279(.A(new_n7655), .B(new_n7624), .Y(new_n7656));
  xnor_3 g07280(.A(new_n7656), .B(new_n7621), .Y(new_n7657));
  not_3  g07281(.A(new_n7484), .Y(new_n7658));
  nand_4 g07282(.A(new_n7490), .B(new_n7658), .Y(new_n7659));
  nand_4 g07283(.A(new_n7491), .B(new_n7480), .Y(new_n7660));
  nand_4 g07284(.A(new_n7660), .B(new_n7659), .Y(new_n7661));
  nand_4 g07285(.A(n5798), .B(n5283), .Y(new_n7662));
  nand_4 g07286(.A(n7265), .B(n6826), .Y(new_n7663));
  nand_4 g07287(.A(n6294), .B(n521), .Y(new_n7664));
  xor_3  g07288(.A(new_n7664), .B(new_n7663), .Y(new_n7665));
  xor_3  g07289(.A(new_n7665), .B(new_n7662), .Y(new_n7666));
  xnor_3 g07290(.A(new_n7666), .B(new_n7661), .Y(new_n7667));
  xnor_3 g07291(.A(new_n7667), .B(new_n7657), .Y(new_n7668));
  xnor_3 g07292(.A(new_n7668), .B(new_n7616), .Y(new_n7669));
  xnor_3 g07293(.A(new_n7669), .B(new_n7612), .Y(new_n7670));
  xnor_3 g07294(.A(new_n7670), .B(new_n7608), .Y(new_n7671));
  nand_4 g07295(.A(new_n7450), .B(new_n7448), .Y(new_n7672));
  nand_4 g07296(.A(new_n7452), .B(new_n7445), .Y(new_n7673));
  nand_4 g07297(.A(new_n7673), .B(new_n7672), .Y(new_n7674));
  nand_4 g07298(.A(n6797), .B(n5579), .Y(new_n7675));
  not_3  g07299(.A(new_n7675), .Y(new_n7676_1));
  nand_4 g07300(.A(new_n7469), .B(new_n7467), .Y(new_n7677));
  nand_4 g07301(.A(new_n7479), .B(new_n7470), .Y(new_n7678));
  nand_4 g07302(.A(new_n7678), .B(new_n7677), .Y(new_n7679));
  xor_3  g07303(.A(new_n7679), .B(new_n7676_1), .Y(new_n7680));
  nand_4 g07304(.A(n4805), .B(n1576), .Y(new_n7681));
  nand_4 g07305(.A(n3992), .B(n2507), .Y(new_n7682));
  xor_3  g07306(.A(new_n7682), .B(new_n7681), .Y(new_n7683));
  nand_4 g07307(.A(n3146), .B(n2498), .Y(new_n7684));
  nand_4 g07308(.A(n6016), .B(n137), .Y(new_n7685));
  xor_3  g07309(.A(new_n7685), .B(new_n7684), .Y(new_n7686));
  xor_3  g07310(.A(new_n7686), .B(new_n7683), .Y(new_n7687));
  nand_4 g07311(.A(n8384), .B(n5153), .Y(new_n7688));
  nand_4 g07312(.A(n7270), .B(n6358), .Y(new_n7689));
  xor_3  g07313(.A(new_n7689), .B(new_n7688), .Y(new_n7690_1));
  not_3  g07314(.A(new_n7471), .Y(new_n7691));
  nand_4 g07315(.A(new_n7474), .B(new_n7691), .Y(new_n7692));
  and_4  g07316(.A(new_n7692), .B(new_n7477), .Y(new_n7693));
  xor_3  g07317(.A(new_n7693), .B(new_n7690_1), .Y(new_n7694));
  xnor_3 g07318(.A(new_n7694), .B(new_n7687), .Y(new_n7695));
  not_3  g07319(.A(new_n7486), .Y(new_n7696));
  nor_4  g07320(.A(new_n7488), .B(new_n7696), .Y(new_n7697));
  not_3  g07321(.A(new_n7485), .Y(new_n7698));
  nor_4  g07322(.A(new_n7489), .B(new_n7698), .Y(new_n7699));
  nor_4  g07323(.A(new_n7699), .B(new_n7697), .Y(new_n7700));
  nand_4 g07324(.A(n4938), .B(n2558), .Y(new_n7701));
  nand_4 g07325(.A(n5198), .B(n806), .Y(new_n7702));
  xor_3  g07326(.A(new_n7702), .B(new_n7701), .Y(new_n7703));
  xor_3  g07327(.A(new_n7703), .B(new_n7700), .Y(new_n7704));
  xnor_3 g07328(.A(new_n7704), .B(new_n7695), .Y(new_n7705));
  xnor_3 g07329(.A(new_n7705), .B(new_n7680), .Y(new_n7706));
  xnor_3 g07330(.A(new_n7706), .B(new_n7674), .Y(new_n7707));
  xnor_3 g07331(.A(new_n7707), .B(new_n7671), .Y(new_n7708));
  xnor_3 g07332(.A(new_n7708), .B(new_n7605), .Y(new_n7709));
  xnor_3 g07333(.A(new_n7709), .B(new_n7523_1), .Y(new_n7710));
  xnor_3 g07334(.A(new_n7710), .B(new_n7514), .Y(n2383));
  not_3  g07335(.A(new_n6272), .Y(new_n7712));
  xor_3  g07336(.A(new_n6282), .B(new_n7712), .Y(n2425));
  not_3  g07337(.A(new_n3043), .Y(new_n7714));
  nor_4  g07338(.A(new_n7714), .B(new_n3041), .Y(new_n7715));
  xnor_3 g07339(.A(new_n7715), .B(new_n3093), .Y(n2431));
  xnor_3 g07340(.A(new_n2187), .B(new_n2186), .Y(n2434));
  not_3  g07341(.A(new_n5266), .Y(new_n7718));
  xor_3  g07342(.A(new_n5267), .B(new_n7718), .Y(n2581));
  nand_4 g07343(.A(new_n7026), .B(new_n7025), .Y(new_n7720));
  xnor_3 g07344(.A(new_n7720), .B(new_n7037), .Y(n2624));
  nand_4 g07345(.A(n6126), .B(n2226), .Y(new_n7722));
  nand_4 g07346(.A(n3602), .B(n1094), .Y(new_n7723));
  nand_4 g07347(.A(n10678), .B(n3719), .Y(new_n7724));
  not_3  g07348(.A(new_n7724), .Y(new_n7725));
  xor_3  g07349(.A(new_n7725), .B(new_n7723), .Y(new_n7726));
  xnor_3 g07350(.A(new_n7726), .B(new_n7722), .Y(new_n7727));
  and_4  g07351(.A(new_n4487), .B(new_n4486), .Y(new_n7728));
  nor_4  g07352(.A(new_n4488), .B(new_n4485), .Y(new_n7729));
  nor_4  g07353(.A(new_n7729), .B(new_n7728), .Y(new_n7730_1));
  xnor_3 g07354(.A(new_n7730_1), .B(new_n7727), .Y(new_n7731));
  nand_4 g07355(.A(n10928), .B(n10439), .Y(new_n7732));
  nand_4 g07356(.A(n8595), .B(n6986), .Y(new_n7733_1));
  xor_3  g07357(.A(new_n7733_1), .B(new_n7732), .Y(new_n7734));
  xnor_3 g07358(.A(new_n7734), .B(new_n7731), .Y(new_n7735));
  and_4  g07359(.A(new_n4481), .B(new_n4476), .Y(new_n7736));
  nor_4  g07360(.A(new_n4489), .B(new_n4483), .Y(new_n7737));
  nor_4  g07361(.A(new_n7737), .B(new_n7736), .Y(new_n7738));
  xnor_3 g07362(.A(new_n7738), .B(new_n7735), .Y(new_n7739));
  nand_4 g07363(.A(new_n4473), .B(new_n4472), .Y(new_n7740));
  nand_4 g07364(.A(new_n4494), .B(new_n4493), .Y(new_n7741));
  nand_4 g07365(.A(new_n7741), .B(new_n7740), .Y(new_n7742));
  not_3  g07366(.A(new_n7742), .Y(new_n7743));
  nor_4  g07367(.A(new_n7743), .B(new_n7739), .Y(new_n7744));
  not_3  g07368(.A(new_n7722), .Y(new_n7745));
  not_3  g07369(.A(new_n7726), .Y(new_n7746));
  nor_4  g07370(.A(new_n7746), .B(new_n7745), .Y(new_n7747));
  nor_4  g07371(.A(new_n7730_1), .B(new_n7727), .Y(new_n7748));
  nor_4  g07372(.A(new_n7748), .B(new_n7747), .Y(new_n7749));
  nand_4 g07373(.A(n10928), .B(n8065), .Y(new_n7750));
  nand_4 g07374(.A(n10439), .B(n6986), .Y(new_n7751));
  nand_4 g07375(.A(n10391), .B(n8336), .Y(new_n7752));
  not_3  g07376(.A(new_n7752), .Y(new_n7753));
  xor_3  g07377(.A(new_n7753), .B(new_n7751), .Y(new_n7754));
  xnor_3 g07378(.A(new_n7754), .B(new_n7750), .Y(new_n7755));
  xnor_3 g07379(.A(new_n7755), .B(new_n7749), .Y(new_n7756));
  nor_4  g07380(.A(new_n7724), .B(new_n7723), .Y(new_n7757));
  nand_4 g07381(.A(n8595), .B(n2226), .Y(new_n7758));
  not_3  g07382(.A(new_n7758), .Y(new_n7759));
  xor_3  g07383(.A(new_n7759), .B(new_n7757), .Y(new_n7760));
  not_3  g07384(.A(new_n7760), .Y(new_n7761));
  nand_4 g07385(.A(n10678), .B(n3602), .Y(new_n7762));
  nand_4 g07386(.A(n6126), .B(n1094), .Y(new_n7763));
  nand_4 g07387(.A(n7320), .B(n3719), .Y(new_n7764));
  not_3  g07388(.A(new_n7764), .Y(new_n7765));
  xor_3  g07389(.A(new_n7765), .B(new_n7763), .Y(new_n7766));
  xnor_3 g07390(.A(new_n7766), .B(new_n7762), .Y(new_n7767));
  not_3  g07391(.A(new_n7767), .Y(new_n7768));
  xor_3  g07392(.A(new_n7768), .B(new_n7761), .Y(new_n7769));
  xnor_3 g07393(.A(new_n7769), .B(new_n7756), .Y(new_n7770));
  not_3  g07394(.A(new_n7770), .Y(new_n7771));
  nand_4 g07395(.A(new_n7734), .B(new_n7731), .Y(new_n7772));
  nor_4  g07396(.A(new_n7733_1), .B(new_n7732), .Y(new_n7773));
  not_3  g07397(.A(new_n7773), .Y(new_n7774));
  not_3  g07398(.A(new_n7734), .Y(new_n7775));
  xnor_3 g07399(.A(new_n7775), .B(new_n7731), .Y(new_n7776));
  not_3  g07400(.A(new_n7738), .Y(new_n7777));
  nand_4 g07401(.A(new_n7777), .B(new_n7776), .Y(new_n7778));
  xnor_3 g07402(.A(new_n7778), .B(new_n7774), .Y(new_n7779));
  nand_4 g07403(.A(new_n7779), .B(new_n7772), .Y(new_n7780));
  xnor_3 g07404(.A(new_n7780), .B(new_n7771), .Y(new_n7781));
  xnor_3 g07405(.A(new_n7781), .B(new_n7744), .Y(new_n7782));
  nand_4 g07406(.A(n8336), .B(n8065), .Y(new_n7783));
  xnor_3 g07407(.A(new_n7743), .B(new_n7739), .Y(new_n7784));
  nand_4 g07408(.A(new_n7784), .B(new_n7783), .Y(new_n7785));
  nand_4 g07409(.A(new_n4496), .B(new_n4470), .Y(new_n7786));
  xnor_3 g07410(.A(new_n7742), .B(new_n7739), .Y(new_n7787));
  xnor_3 g07411(.A(new_n7787), .B(new_n7783), .Y(new_n7788));
  nand_4 g07412(.A(new_n7788), .B(new_n7786), .Y(new_n7789));
  nand_4 g07413(.A(new_n7789), .B(new_n7785), .Y(new_n7790));
  xnor_3 g07414(.A(new_n7790), .B(new_n7782), .Y(new_n7791));
  nand_4 g07415(.A(n7160), .B(n4826), .Y(new_n7792));
  nand_4 g07416(.A(n7733), .B(n4828), .Y(new_n7793));
  nand_4 g07417(.A(n12925), .B(n2515), .Y(new_n7794));
  xnor_3 g07418(.A(new_n7794), .B(new_n7793), .Y(new_n7795));
  nor_4  g07419(.A(new_n7795), .B(new_n7792), .Y(new_n7796));
  not_3  g07420(.A(new_n7792), .Y(new_n7797));
  not_3  g07421(.A(new_n7795), .Y(new_n7798));
  nor_4  g07422(.A(new_n7798), .B(new_n7797), .Y(new_n7799));
  nor_4  g07423(.A(new_n7799), .B(new_n7796), .Y(new_n7800));
  not_3  g07424(.A(new_n4540), .Y(new_n7801));
  not_3  g07425(.A(new_n4541), .Y(new_n7802));
  nor_4  g07426(.A(new_n7802), .B(new_n7801), .Y(new_n7803));
  not_3  g07427(.A(new_n4539), .Y(new_n7804));
  nor_4  g07428(.A(new_n4542), .B(new_n7804), .Y(new_n7805));
  nor_4  g07429(.A(new_n7805), .B(new_n7803), .Y(new_n7806));
  xnor_3 g07430(.A(new_n7806), .B(new_n7800), .Y(new_n7807));
  not_3  g07431(.A(new_n7807), .Y(new_n7808));
  nand_4 g07432(.A(n12391), .B(n4970), .Y(new_n7809));
  nand_4 g07433(.A(n7891), .B(n7610), .Y(new_n7810));
  xor_3  g07434(.A(new_n7810), .B(new_n7809), .Y(new_n7811));
  xnor_3 g07435(.A(new_n7811), .B(new_n7808), .Y(new_n7812));
  nand_4 g07436(.A(new_n4537), .B(new_n4535), .Y(new_n7813));
  not_3  g07437(.A(new_n7813), .Y(new_n7814));
  nor_4  g07438(.A(new_n4543), .B(new_n4538), .Y(new_n7815));
  nor_4  g07439(.A(new_n7815), .B(new_n7814), .Y(new_n7816));
  xnor_3 g07440(.A(new_n7816), .B(new_n7812), .Y(new_n7817));
  nor_4  g07441(.A(new_n4544), .B(new_n4533), .Y(new_n7818));
  nor_4  g07442(.A(new_n4548), .B(new_n4545), .Y(new_n7819));
  nor_4  g07443(.A(new_n7819), .B(new_n7818), .Y(new_n7820));
  nor_4  g07444(.A(new_n7820), .B(new_n7817), .Y(new_n7821));
  not_3  g07445(.A(new_n7821), .Y(new_n7822));
  not_3  g07446(.A(new_n7796), .Y(new_n7823_1));
  nand_4 g07447(.A(new_n7806), .B(new_n7800), .Y(new_n7824));
  nand_4 g07448(.A(new_n7824), .B(new_n7823_1), .Y(new_n7825));
  nand_4 g07449(.A(n12391), .B(n503), .Y(new_n7826));
  not_3  g07450(.A(new_n7826), .Y(new_n7827));
  nand_4 g07451(.A(n7891), .B(n4970), .Y(new_n7828));
  nand_4 g07452(.A(n12069), .B(n10965), .Y(new_n7829));
  xnor_3 g07453(.A(new_n7829), .B(new_n7828), .Y(new_n7830));
  xor_3  g07454(.A(new_n7830), .B(new_n7827), .Y(new_n7831));
  xnor_3 g07455(.A(new_n7831), .B(new_n7825), .Y(new_n7832));
  nor_4  g07456(.A(new_n7794), .B(new_n7793), .Y(new_n7833));
  not_3  g07457(.A(new_n7833), .Y(new_n7834));
  nand_4 g07458(.A(n7610), .B(n7160), .Y(new_n7835));
  xor_3  g07459(.A(new_n7835), .B(new_n7834), .Y(new_n7836));
  nand_4 g07460(.A(n7733), .B(n2515), .Y(new_n7837));
  not_3  g07461(.A(new_n7837), .Y(new_n7838));
  nand_4 g07462(.A(n4828), .B(n4826), .Y(new_n7839));
  nand_4 g07463(.A(n12925), .B(n1199), .Y(new_n7840));
  xnor_3 g07464(.A(new_n7840), .B(new_n7839), .Y(new_n7841));
  xor_3  g07465(.A(new_n7841), .B(new_n7838), .Y(new_n7842));
  xnor_3 g07466(.A(new_n7842), .B(new_n7836), .Y(new_n7843));
  xnor_3 g07467(.A(new_n7843), .B(new_n7832), .Y(new_n7844));
  nand_4 g07468(.A(new_n7811), .B(new_n7808), .Y(new_n7845));
  nor_4  g07469(.A(new_n7810), .B(new_n7809), .Y(new_n7846));
  xnor_3 g07470(.A(new_n7811), .B(new_n7807), .Y(new_n7847));
  not_3  g07471(.A(new_n7816), .Y(new_n7848));
  nand_4 g07472(.A(new_n7848), .B(new_n7847), .Y(new_n7849));
  not_3  g07473(.A(new_n7849), .Y(new_n7850));
  xnor_3 g07474(.A(new_n7850), .B(new_n7846), .Y(new_n7851));
  nand_4 g07475(.A(new_n7851), .B(new_n7845), .Y(new_n7852));
  xnor_3 g07476(.A(new_n7852), .B(new_n7844), .Y(new_n7853));
  xnor_3 g07477(.A(new_n7853), .B(new_n7822), .Y(new_n7854));
  nand_4 g07478(.A(n12069), .B(n503), .Y(new_n7855));
  not_3  g07479(.A(new_n7855), .Y(new_n7856));
  not_3  g07480(.A(new_n7817), .Y(new_n7857));
  xnor_3 g07481(.A(new_n7820), .B(new_n7857), .Y(new_n7858));
  nand_4 g07482(.A(new_n7858), .B(new_n7856), .Y(new_n7859));
  nor_4  g07483(.A(new_n4549), .B(new_n4532), .Y(new_n7860));
  xnor_3 g07484(.A(new_n7858), .B(new_n7855), .Y(new_n7861));
  nand_4 g07485(.A(new_n7861), .B(new_n7860), .Y(new_n7862_1));
  nand_4 g07486(.A(new_n7862_1), .B(new_n7859), .Y(new_n7863));
  xnor_3 g07487(.A(new_n7863), .B(new_n7854), .Y(new_n7864));
  nand_4 g07488(.A(n11222), .B(n6359), .Y(new_n7865));
  not_3  g07489(.A(new_n7865), .Y(new_n7866));
  nand_4 g07490(.A(n4086), .B(n996), .Y(new_n7867));
  nand_4 g07491(.A(n5767), .B(n405), .Y(new_n7868));
  nand_4 g07492(.A(n8433), .B(n5319), .Y(new_n7869));
  xnor_3 g07493(.A(new_n7869), .B(new_n7868), .Y(new_n7870));
  nor_4  g07494(.A(new_n7870), .B(new_n7867), .Y(new_n7871));
  not_3  g07495(.A(new_n7867), .Y(new_n7872));
  not_3  g07496(.A(new_n7870), .Y(new_n7873));
  nor_4  g07497(.A(new_n7873), .B(new_n7872), .Y(new_n7874));
  nor_4  g07498(.A(new_n7874), .B(new_n7871), .Y(new_n7875));
  not_3  g07499(.A(new_n4502), .Y(new_n7876));
  nor_4  g07500(.A(new_n4508), .B(new_n7876), .Y(new_n7877));
  nor_4  g07501(.A(new_n7877), .B(new_n4507), .Y(new_n7878));
  xnor_3 g07502(.A(new_n7878), .B(new_n7875), .Y(new_n7879));
  nand_4 g07503(.A(n11153), .B(n6611), .Y(new_n7880));
  nand_4 g07504(.A(n5314), .B(n217), .Y(new_n7881));
  xor_3  g07505(.A(new_n7881), .B(new_n7880), .Y(new_n7882));
  xnor_3 g07506(.A(new_n7882), .B(new_n7879), .Y(new_n7883));
  not_3  g07507(.A(new_n4501), .Y(new_n7884));
  nand_4 g07508(.A(new_n4510), .B(new_n7884), .Y(new_n7885));
  nand_4 g07509(.A(new_n4517), .B(new_n4511), .Y(new_n7886));
  nand_4 g07510(.A(new_n7886), .B(new_n7885), .Y(new_n7887));
  xnor_3 g07511(.A(new_n7887), .B(new_n7883), .Y(new_n7888));
  not_3  g07512(.A(new_n4526), .Y(new_n7889));
  nand_4 g07513(.A(new_n7889), .B(new_n4521), .Y(new_n7890));
  nand_4 g07514(.A(new_n7890), .B(new_n4519), .Y(new_n7891_1));
  not_3  g07515(.A(new_n7891_1), .Y(new_n7892));
  nor_4  g07516(.A(new_n7892), .B(new_n7888), .Y(new_n7893));
  not_3  g07517(.A(new_n7888), .Y(new_n7894));
  nor_4  g07518(.A(new_n7891_1), .B(new_n7894), .Y(new_n7895));
  nor_4  g07519(.A(new_n7895), .B(new_n7893), .Y(new_n7896));
  nand_4 g07520(.A(new_n7896), .B(new_n7866), .Y(new_n7897));
  xnor_3 g07521(.A(new_n7896), .B(new_n7865), .Y(new_n7898));
  nand_4 g07522(.A(new_n7898), .B(new_n4528), .Y(new_n7899));
  nand_4 g07523(.A(new_n7899), .B(new_n7897), .Y(new_n7900));
  nor_4  g07524(.A(new_n7869), .B(new_n7868), .Y(new_n7901));
  nand_4 g07525(.A(n996), .B(n217), .Y(new_n7902));
  not_3  g07526(.A(new_n7902), .Y(new_n7903));
  xor_3  g07527(.A(new_n7903), .B(new_n7901), .Y(new_n7904));
  not_3  g07528(.A(new_n7904), .Y(new_n7905));
  nand_4 g07529(.A(n5319), .B(n405), .Y(new_n7906));
  not_3  g07530(.A(new_n7906), .Y(new_n7907));
  nand_4 g07531(.A(n5767), .B(n4086), .Y(new_n7908));
  nand_4 g07532(.A(n9457), .B(n8433), .Y(new_n7909));
  xnor_3 g07533(.A(new_n7909), .B(new_n7908), .Y(new_n7910));
  xor_3  g07534(.A(new_n7910), .B(new_n7907), .Y(new_n7911));
  nor_4  g07535(.A(new_n7911), .B(new_n7905), .Y(new_n7912));
  not_3  g07536(.A(new_n7911), .Y(new_n7913));
  nor_4  g07537(.A(new_n7913), .B(new_n7904), .Y(new_n7914));
  nor_4  g07538(.A(new_n7914), .B(new_n7912), .Y(new_n7915));
  nand_4 g07539(.A(new_n7878), .B(new_n7875), .Y(new_n7916));
  not_3  g07540(.A(new_n7916), .Y(new_n7917));
  nor_4  g07541(.A(new_n7917), .B(new_n7871), .Y(new_n7918));
  not_3  g07542(.A(new_n7918), .Y(new_n7919));
  nand_4 g07543(.A(n11153), .B(n6359), .Y(new_n7920));
  not_3  g07544(.A(new_n7920), .Y(new_n7921));
  nand_4 g07545(.A(n6611), .B(n5314), .Y(new_n7922));
  nand_4 g07546(.A(n11296), .B(n11222), .Y(new_n7923));
  nand_4 g07547(.A(new_n7923), .B(new_n7922), .Y(new_n7924));
  not_3  g07548(.A(new_n7922), .Y(new_n7925));
  not_3  g07549(.A(new_n7923), .Y(new_n7926));
  nand_4 g07550(.A(new_n7926), .B(new_n7925), .Y(new_n7927));
  nand_4 g07551(.A(new_n7927), .B(new_n7924), .Y(new_n7928));
  xor_3  g07552(.A(new_n7928), .B(new_n7921), .Y(new_n7929));
  xnor_3 g07553(.A(new_n7929), .B(new_n7919), .Y(new_n7930));
  xnor_3 g07554(.A(new_n7930), .B(new_n7915), .Y(new_n7931));
  not_3  g07555(.A(new_n7879), .Y(new_n7932));
  nand_4 g07556(.A(new_n7882), .B(new_n7932), .Y(new_n7933));
  nor_4  g07557(.A(new_n7881), .B(new_n7880), .Y(new_n7934));
  nand_4 g07558(.A(new_n7887), .B(new_n7883), .Y(new_n7935));
  not_3  g07559(.A(new_n7935), .Y(new_n7936));
  xnor_3 g07560(.A(new_n7936), .B(new_n7934), .Y(new_n7937));
  nand_4 g07561(.A(new_n7937), .B(new_n7933), .Y(new_n7938));
  xnor_3 g07562(.A(new_n7938), .B(new_n7931), .Y(new_n7939));
  xnor_3 g07563(.A(new_n7939), .B(new_n7893), .Y(new_n7940));
  xnor_3 g07564(.A(new_n7940), .B(new_n7900), .Y(new_n7941));
  xnor_3 g07565(.A(new_n7941), .B(new_n7864), .Y(new_n7942));
  xnor_3 g07566(.A(new_n7861), .B(new_n7860), .Y(new_n7943));
  not_3  g07567(.A(new_n7943), .Y(new_n7944));
  not_3  g07568(.A(new_n4528), .Y(new_n7945));
  xnor_3 g07569(.A(new_n7898), .B(new_n7945), .Y(new_n7946_1));
  nor_4  g07570(.A(new_n7946_1), .B(new_n7944), .Y(new_n7947));
  not_3  g07571(.A(new_n4550), .Y(new_n7948));
  not_3  g07572(.A(new_n4554), .Y(new_n7949));
  nor_4  g07573(.A(new_n7949), .B(new_n7948), .Y(new_n7950));
  nor_4  g07574(.A(new_n4555), .B(new_n4531), .Y(new_n7951));
  nor_4  g07575(.A(new_n7951), .B(new_n7950), .Y(new_n7952));
  xnor_3 g07576(.A(new_n7946_1), .B(new_n7944), .Y(new_n7953));
  nor_4  g07577(.A(new_n7953), .B(new_n7952), .Y(new_n7954));
  nor_4  g07578(.A(new_n7954), .B(new_n7947), .Y(new_n7955));
  xnor_3 g07579(.A(new_n7955), .B(new_n7942), .Y(new_n7956));
  nand_4 g07580(.A(new_n7956), .B(new_n7791), .Y(new_n7957));
  xnor_3 g07581(.A(new_n7956), .B(new_n7791), .Y(new_n7958));
  not_3  g07582(.A(new_n7958), .Y(new_n7959));
  not_3  g07583(.A(new_n7783), .Y(new_n7960));
  nand_4 g07584(.A(new_n7787), .B(new_n7960), .Y(new_n7961));
  nand_4 g07585(.A(new_n7961), .B(new_n7785), .Y(new_n7962));
  xnor_3 g07586(.A(new_n7962), .B(new_n7786), .Y(new_n7963));
  xnor_3 g07587(.A(new_n7953), .B(new_n7952), .Y(new_n7964));
  not_3  g07588(.A(new_n7964), .Y(new_n7965_1));
  nand_4 g07589(.A(new_n7965_1), .B(new_n7963), .Y(new_n7966_1));
  xnor_3 g07590(.A(new_n7964), .B(new_n7963), .Y(new_n7967));
  nor_4  g07591(.A(new_n4557), .B(new_n4497), .Y(new_n7968));
  not_3  g07592(.A(new_n4563), .Y(new_n7969));
  nor_4  g07593(.A(new_n7969), .B(new_n4558), .Y(new_n7970));
  nor_4  g07594(.A(new_n7970), .B(new_n7968), .Y(new_n7971));
  nand_4 g07595(.A(new_n7971), .B(new_n7967), .Y(new_n7972));
  nand_4 g07596(.A(new_n7972), .B(new_n7966_1), .Y(new_n7973));
  nand_4 g07597(.A(new_n7973), .B(new_n7959), .Y(new_n7974));
  nand_4 g07598(.A(new_n7974), .B(new_n7957), .Y(new_n7975));
  nand_4 g07599(.A(new_n7781), .B(new_n7744), .Y(new_n7976));
  not_3  g07600(.A(new_n7976), .Y(new_n7977));
  nor_4  g07601(.A(new_n7790), .B(new_n7782), .Y(new_n7978));
  nor_4  g07602(.A(new_n7978), .B(new_n7977), .Y(new_n7979));
  xnor_3 g07603(.A(new_n7979), .B(new_n7975), .Y(new_n7980));
  not_3  g07604(.A(new_n7941), .Y(new_n7981_1));
  nand_4 g07605(.A(new_n7981_1), .B(new_n7864), .Y(new_n7982));
  not_3  g07606(.A(new_n7947), .Y(new_n7983));
  not_3  g07607(.A(new_n7952), .Y(new_n7984));
  xnor_3 g07608(.A(new_n7946_1), .B(new_n7943), .Y(new_n7985));
  nand_4 g07609(.A(new_n7985), .B(new_n7984), .Y(new_n7986));
  nand_4 g07610(.A(new_n7986), .B(new_n7983), .Y(new_n7987));
  nand_4 g07611(.A(new_n7987), .B(new_n7942), .Y(new_n7988));
  nand_4 g07612(.A(new_n7988), .B(new_n7982), .Y(new_n7989));
  nand_4 g07613(.A(new_n7853), .B(new_n7821), .Y(new_n7990));
  nand_4 g07614(.A(new_n7863), .B(new_n7854), .Y(new_n7991));
  nand_4 g07615(.A(new_n7991), .B(new_n7990), .Y(new_n7992));
  and_4  g07616(.A(new_n7909), .B(new_n7908), .Y(new_n7993));
  nor_4  g07617(.A(new_n7910), .B(new_n7907), .Y(new_n7994));
  nor_4  g07618(.A(new_n7994), .B(new_n7993), .Y(new_n7995));
  nand_4 g07619(.A(n11296), .B(n11153), .Y(new_n7996));
  xor_3  g07620(.A(new_n7996), .B(new_n7995), .Y(new_n7997));
  not_3  g07621(.A(new_n7751), .Y(new_n7998));
  nor_4  g07622(.A(new_n7753), .B(new_n7998), .Y(new_n7999));
  not_3  g07623(.A(new_n7750), .Y(new_n8000));
  nor_4  g07624(.A(new_n7754), .B(new_n8000), .Y(new_n8001));
  nor_4  g07625(.A(new_n8001), .B(new_n7999), .Y(new_n8002));
  nand_4 g07626(.A(n6611), .B(n996), .Y(new_n8003));
  nand_4 g07627(.A(n6359), .B(n5314), .Y(new_n8004));
  xor_3  g07628(.A(new_n8004), .B(new_n8003), .Y(new_n8005));
  nand_4 g07629(.A(n12069), .B(n7546), .Y(new_n8006));
  nand_4 g07630(.A(n12925), .B(n6578), .Y(new_n8007));
  xor_3  g07631(.A(new_n8007), .B(new_n8006), .Y(new_n8008));
  xnor_3 g07632(.A(new_n8008), .B(new_n8005), .Y(new_n8009));
  nand_4 g07633(.A(n7733), .B(n1199), .Y(new_n8010));
  nand_4 g07634(.A(n7160), .B(n4970), .Y(new_n8011));
  not_3  g07635(.A(new_n8011), .Y(new_n8012));
  xor_3  g07636(.A(new_n8012), .B(new_n8010), .Y(new_n8013));
  xnor_3 g07637(.A(new_n8013), .B(new_n8009), .Y(new_n8014));
  xnor_3 g07638(.A(new_n8014), .B(new_n8002), .Y(new_n8015));
  nand_4 g07639(.A(new_n7903), .B(new_n7901), .Y(new_n8016));
  nand_4 g07640(.A(new_n7913), .B(new_n7904), .Y(new_n8017));
  nand_4 g07641(.A(new_n8017), .B(new_n8016), .Y(new_n8018));
  nand_4 g07642(.A(n5767), .B(n217), .Y(new_n8019));
  nand_4 g07643(.A(new_n7924), .B(new_n7921), .Y(new_n8020));
  nand_4 g07644(.A(new_n8020), .B(new_n7927), .Y(new_n8021));
  xor_3  g07645(.A(new_n8021), .B(new_n8019), .Y(new_n8022));
  xor_3  g07646(.A(new_n8022), .B(new_n8018), .Y(new_n8023));
  xnor_3 g07647(.A(new_n8023), .B(new_n8015), .Y(new_n8024));
  xnor_3 g07648(.A(new_n8024), .B(new_n7997), .Y(new_n8025));
  nand_4 g07649(.A(new_n7929), .B(new_n7918), .Y(new_n8026));
  not_3  g07650(.A(new_n7915), .Y(new_n8027));
  nand_4 g07651(.A(new_n7930), .B(new_n8027), .Y(new_n8028_1));
  nand_4 g07652(.A(new_n8028_1), .B(new_n8026), .Y(new_n8029));
  nand_4 g07653(.A(n7610), .B(n4828), .Y(new_n8030));
  nand_4 g07654(.A(n4826), .B(n2515), .Y(new_n8031));
  not_3  g07655(.A(new_n8031), .Y(new_n8032));
  xor_3  g07656(.A(new_n8032), .B(new_n8030), .Y(new_n8033));
  xnor_3 g07657(.A(new_n8033), .B(new_n8029), .Y(new_n8034));
  nand_4 g07658(.A(n4921), .B(n4516), .Y(new_n8035));
  nand_4 g07659(.A(n2564), .B(n1835), .Y(new_n8036));
  xor_3  g07660(.A(new_n8036), .B(new_n8035), .Y(new_n8037));
  xnor_3 g07661(.A(new_n8037), .B(new_n8034), .Y(new_n8038));
  xnor_3 g07662(.A(new_n8038), .B(new_n8025), .Y(new_n8039));
  xnor_3 g07663(.A(new_n8039), .B(new_n7992), .Y(new_n8040));
  xnor_3 g07664(.A(new_n8040), .B(new_n7989), .Y(new_n8041));
  nand_4 g07665(.A(new_n7939), .B(new_n7893), .Y(new_n8042));
  not_3  g07666(.A(new_n7940), .Y(new_n8043));
  nand_4 g07667(.A(new_n8043), .B(new_n7900), .Y(new_n8044));
  nand_4 g07668(.A(new_n8044), .B(new_n8042), .Y(new_n8045));
  nand_4 g07669(.A(new_n7850), .B(new_n7846), .Y(new_n8046));
  not_3  g07670(.A(new_n7844), .Y(new_n8047));
  nand_4 g07671(.A(new_n7852), .B(new_n8047), .Y(new_n8048));
  nand_4 g07672(.A(new_n8048), .B(new_n8046), .Y(new_n8049));
  nand_4 g07673(.A(n4189), .B(n2577), .Y(new_n8050));
  not_3  g07674(.A(new_n8050), .Y(new_n8051));
  nand_4 g07675(.A(n6687), .B(n1835), .Y(new_n8052));
  not_3  g07676(.A(new_n8052), .Y(new_n8053));
  nor_4  g07677(.A(new_n8053), .B(new_n8051), .Y(new_n8054));
  nand_4 g07678(.A(n9637), .B(n2564), .Y(new_n8055));
  not_3  g07679(.A(new_n8055), .Y(new_n8056));
  xor_3  g07680(.A(new_n8053), .B(new_n8050), .Y(new_n8057));
  nor_4  g07681(.A(new_n8057), .B(new_n8056), .Y(new_n8058));
  nor_4  g07682(.A(new_n8058), .B(new_n8054), .Y(new_n8059));
  xnor_3 g07683(.A(new_n8059), .B(new_n8049), .Y(new_n8060));
  nand_4 g07684(.A(n11917), .B(n6770), .Y(new_n8061));
  not_3  g07685(.A(new_n8061), .Y(new_n8062));
  nand_4 g07686(.A(n9920), .B(n4921), .Y(new_n8063));
  nand_4 g07687(.A(n9956), .B(n3627), .Y(new_n8064));
  not_3  g07688(.A(new_n8064), .Y(new_n8065_1));
  xor_3  g07689(.A(new_n8065_1), .B(new_n8063), .Y(new_n8066));
  not_3  g07690(.A(new_n8066), .Y(new_n8067));
  nor_4  g07691(.A(new_n8067), .B(new_n8062), .Y(new_n8068));
  xor_3  g07692(.A(new_n8067), .B(new_n8062), .Y(new_n8069));
  not_3  g07693(.A(new_n8069), .Y(new_n8070));
  not_3  g07694(.A(new_n4263), .Y(new_n8071));
  nor_4  g07695(.A(new_n4265), .B(new_n8071), .Y(new_n8072));
  not_3  g07696(.A(new_n4262), .Y(new_n8073));
  nor_4  g07697(.A(new_n4266), .B(new_n8073), .Y(new_n8074));
  nor_4  g07698(.A(new_n8074), .B(new_n8072), .Y(new_n8075));
  nor_4  g07699(.A(new_n8075), .B(new_n8070), .Y(new_n8076));
  nor_4  g07700(.A(new_n8076), .B(new_n8068), .Y(new_n8077));
  xnor_3 g07701(.A(new_n8057), .B(new_n8055), .Y(new_n8078));
  not_3  g07702(.A(new_n8078), .Y(new_n8079));
  nand_4 g07703(.A(new_n8079), .B(new_n8077), .Y(new_n8080));
  nor_4  g07704(.A(new_n8064), .B(new_n8063), .Y(new_n8081));
  nand_4 g07705(.A(n6770), .B(n3842), .Y(new_n8082));
  xor_3  g07706(.A(new_n8082), .B(new_n8081), .Y(new_n8083));
  nand_4 g07707(.A(n4921), .B(n3627), .Y(new_n8084));
  nand_4 g07708(.A(n11917), .B(n9920), .Y(new_n8085));
  nand_4 g07709(.A(n9956), .B(n4516), .Y(new_n8086));
  not_3  g07710(.A(new_n8086), .Y(new_n8087));
  xor_3  g07711(.A(new_n8087), .B(new_n8085), .Y(new_n8088));
  xnor_3 g07712(.A(new_n8088), .B(new_n8084), .Y(new_n8089));
  not_3  g07713(.A(new_n8089), .Y(new_n8090));
  xor_3  g07714(.A(new_n8090), .B(new_n8083), .Y(new_n8091));
  not_3  g07715(.A(new_n8091), .Y(new_n8092));
  xnor_3 g07716(.A(new_n8078), .B(new_n8077), .Y(new_n8093));
  nand_4 g07717(.A(new_n8093), .B(new_n8092), .Y(new_n8094));
  nand_4 g07718(.A(new_n8094), .B(new_n8080), .Y(new_n8095));
  nand_4 g07719(.A(n9920), .B(n3842), .Y(new_n8096));
  xnor_3 g07720(.A(new_n8096), .B(new_n8095), .Y(new_n8097));
  xnor_3 g07721(.A(new_n8097), .B(new_n8060), .Y(new_n8098));
  xnor_3 g07722(.A(new_n8098), .B(new_n8045), .Y(new_n8099));
  nand_4 g07723(.A(new_n7936), .B(new_n7934), .Y(new_n8100_1));
  not_3  g07724(.A(new_n7931), .Y(new_n8101));
  nand_4 g07725(.A(new_n7938), .B(new_n8101), .Y(new_n8102));
  nand_4 g07726(.A(new_n8102), .B(new_n8100_1), .Y(new_n8103));
  nand_4 g07727(.A(new_n7759), .B(new_n7757), .Y(new_n8104));
  nand_4 g07728(.A(new_n7768), .B(new_n7760), .Y(new_n8105));
  nand_4 g07729(.A(new_n8105), .B(new_n8104), .Y(new_n8106));
  nand_4 g07730(.A(n10439), .B(n2226), .Y(new_n8107));
  nand_4 g07731(.A(n10678), .B(n6126), .Y(new_n8108));
  xor_3  g07732(.A(new_n8108), .B(new_n8107), .Y(new_n8109));
  nand_4 g07733(.A(n11222), .B(n1357), .Y(new_n8110));
  nand_4 g07734(.A(n8433), .B(n4817), .Y(new_n8111));
  xor_3  g07735(.A(new_n8111), .B(new_n8110), .Y(new_n8112));
  nand_4 g07736(.A(n10928), .B(n10391), .Y(new_n8113));
  nand_4 g07737(.A(n8595), .B(n1094), .Y(new_n8114));
  not_3  g07738(.A(new_n8114), .Y(new_n8115));
  xor_3  g07739(.A(new_n8115), .B(new_n8113), .Y(new_n8116));
  xor_3  g07740(.A(new_n8116), .B(new_n8112), .Y(new_n8117));
  xnor_3 g07741(.A(new_n8117), .B(new_n8109), .Y(new_n8118));
  xnor_3 g07742(.A(new_n8118), .B(new_n8106), .Y(new_n8119));
  not_3  g07743(.A(new_n7763), .Y(new_n8120));
  nor_4  g07744(.A(new_n7765), .B(new_n8120), .Y(new_n8121));
  not_3  g07745(.A(new_n7762), .Y(new_n8122));
  nor_4  g07746(.A(new_n7766), .B(new_n8122), .Y(new_n8123));
  nor_4  g07747(.A(new_n8123), .B(new_n8121), .Y(new_n8124));
  nand_4 g07748(.A(n9457), .B(n405), .Y(new_n8125));
  not_3  g07749(.A(new_n8125), .Y(new_n8126));
  xnor_3 g07750(.A(new_n8126), .B(new_n8124), .Y(new_n8127));
  nand_4 g07751(.A(n8065), .B(n6986), .Y(new_n8128));
  nand_4 g07752(.A(n8336), .B(n4190), .Y(new_n8129));
  not_3  g07753(.A(new_n8129), .Y(new_n8130));
  xor_3  g07754(.A(new_n8130), .B(new_n8128), .Y(new_n8131));
  nand_4 g07755(.A(n7523), .B(n3719), .Y(new_n8132));
  nand_4 g07756(.A(n7320), .B(n3602), .Y(new_n8133));
  xor_3  g07757(.A(new_n8133), .B(new_n8132), .Y(new_n8134));
  xor_3  g07758(.A(new_n8134), .B(new_n8131), .Y(new_n8135));
  xnor_3 g07759(.A(new_n8135), .B(new_n8127), .Y(new_n8136));
  nand_4 g07760(.A(n11536), .B(n6687), .Y(new_n8137));
  and_4  g07761(.A(new_n7829), .B(new_n7828), .Y(new_n8138_1));
  nor_4  g07762(.A(new_n7830), .B(new_n7827), .Y(new_n8139));
  nor_4  g07763(.A(new_n8139), .B(new_n8138_1), .Y(new_n8140));
  xor_3  g07764(.A(new_n8140), .B(new_n8137), .Y(new_n8141));
  xnor_3 g07765(.A(new_n8141), .B(new_n8136), .Y(new_n8142));
  xnor_3 g07766(.A(new_n8142), .B(new_n8119), .Y(new_n8143));
  xnor_3 g07767(.A(new_n8143), .B(new_n8103), .Y(new_n8144));
  not_3  g07768(.A(new_n7749), .Y(new_n8145));
  nand_4 g07769(.A(new_n7755), .B(new_n8145), .Y(new_n8146));
  nand_4 g07770(.A(new_n7769), .B(new_n7756), .Y(new_n8147));
  nand_4 g07771(.A(new_n8147), .B(new_n8146), .Y(new_n8148));
  not_3  g07772(.A(new_n8082), .Y(new_n8149));
  nor_4  g07773(.A(new_n8149), .B(new_n8081), .Y(new_n8150));
  nor_4  g07774(.A(new_n8090), .B(new_n8083), .Y(new_n8151));
  nor_4  g07775(.A(new_n8151), .B(new_n8150), .Y(new_n8152));
  nand_4 g07776(.A(n9637), .B(n4189), .Y(new_n8153));
  not_3  g07777(.A(new_n8085), .Y(new_n8154));
  nor_4  g07778(.A(new_n8087), .B(new_n8154), .Y(new_n8155));
  not_3  g07779(.A(new_n8084), .Y(new_n8156));
  nor_4  g07780(.A(new_n8088), .B(new_n8156), .Y(new_n8157));
  nor_4  g07781(.A(new_n8157), .B(new_n8155), .Y(new_n8158));
  nand_4 g07782(.A(n5319), .B(n4086), .Y(new_n8159));
  not_3  g07783(.A(new_n8159), .Y(new_n8160));
  nand_4 g07784(.A(n6770), .B(n2577), .Y(new_n8161));
  nand_4 g07785(.A(n11917), .B(n3627), .Y(new_n8162));
  xor_3  g07786(.A(new_n8162), .B(new_n8161), .Y(new_n8163));
  xnor_3 g07787(.A(new_n8163), .B(new_n8160), .Y(new_n8164));
  xnor_3 g07788(.A(new_n8164), .B(new_n8158), .Y(new_n8165));
  xnor_3 g07789(.A(new_n8165), .B(new_n8153), .Y(new_n8166));
  xnor_3 g07790(.A(new_n8166), .B(new_n8152), .Y(new_n8167));
  nand_4 g07791(.A(n9956), .B(n2087), .Y(new_n8168));
  nor_4  g07792(.A(new_n7835), .B(new_n7834), .Y(new_n8169));
  not_3  g07793(.A(new_n7836), .Y(new_n8170));
  nor_4  g07794(.A(new_n7842), .B(new_n8170), .Y(new_n8171));
  nor_4  g07795(.A(new_n8171), .B(new_n8169), .Y(new_n8172));
  and_4  g07796(.A(new_n7840), .B(new_n7839), .Y(new_n8173));
  nor_4  g07797(.A(new_n7841), .B(new_n7838), .Y(new_n8174));
  nor_4  g07798(.A(new_n8174), .B(new_n8173), .Y(new_n8175));
  nand_4 g07799(.A(n12391), .B(n10965), .Y(new_n8176));
  nand_4 g07800(.A(n7891), .B(n503), .Y(new_n8177));
  xor_3  g07801(.A(new_n8177), .B(new_n8176), .Y(new_n8178));
  xnor_3 g07802(.A(new_n8178), .B(new_n8175), .Y(new_n8179));
  xnor_3 g07803(.A(new_n8179), .B(new_n8172), .Y(new_n8180));
  xnor_3 g07804(.A(new_n8180), .B(new_n8168), .Y(new_n8181));
  xnor_3 g07805(.A(new_n8181), .B(new_n8167), .Y(new_n8182));
  xnor_3 g07806(.A(new_n8182), .B(new_n8148), .Y(new_n8183));
  not_3  g07807(.A(new_n7778), .Y(new_n8184));
  nand_4 g07808(.A(new_n8184), .B(new_n7773), .Y(new_n8185));
  nand_4 g07809(.A(new_n7780), .B(new_n7770), .Y(new_n8186));
  nand_4 g07810(.A(new_n8186), .B(new_n8185), .Y(new_n8187));
  nand_4 g07811(.A(n2577), .B(n2564), .Y(new_n8188));
  nand_4 g07812(.A(n4189), .B(n3842), .Y(new_n8189));
  nor_4  g07813(.A(new_n8189), .B(new_n8188), .Y(new_n8190));
  xnor_3 g07814(.A(new_n8075), .B(new_n8069), .Y(new_n8191));
  not_3  g07815(.A(new_n8191), .Y(new_n8192));
  xor_3  g07816(.A(new_n8189), .B(new_n8188), .Y(new_n8193));
  xnor_3 g07817(.A(new_n8193), .B(new_n8192), .Y(new_n8194));
  not_3  g07818(.A(new_n4257), .Y(new_n8195));
  and_4  g07819(.A(new_n4259), .B(new_n8195), .Y(new_n8196));
  nor_4  g07820(.A(new_n4267), .B(new_n4260), .Y(new_n8197));
  nor_4  g07821(.A(new_n8197), .B(new_n8196), .Y(new_n8198));
  nor_4  g07822(.A(new_n8198), .B(new_n8194), .Y(new_n8199));
  nand_4 g07823(.A(new_n8199), .B(new_n8190), .Y(new_n8200));
  xnor_3 g07824(.A(new_n8093), .B(new_n8091), .Y(new_n8201));
  nand_4 g07825(.A(new_n8193), .B(new_n8192), .Y(new_n8202_1));
  xnor_3 g07826(.A(new_n8199), .B(new_n8190), .Y(new_n8203));
  nand_4 g07827(.A(new_n8203), .B(new_n8202_1), .Y(new_n8204));
  nand_4 g07828(.A(new_n8204), .B(new_n8201), .Y(new_n8205));
  nand_4 g07829(.A(new_n8205), .B(new_n8200), .Y(new_n8206));
  xnor_3 g07830(.A(new_n8206), .B(new_n8187), .Y(new_n8207));
  xnor_3 g07831(.A(new_n8207), .B(new_n8183), .Y(new_n8208));
  xnor_3 g07832(.A(new_n8208), .B(new_n8144), .Y(new_n8209));
  xnor_3 g07833(.A(new_n8209), .B(new_n8099), .Y(new_n8210));
  xnor_3 g07834(.A(new_n8210), .B(new_n8041), .Y(new_n8211));
  xnor_3 g07835(.A(new_n8211), .B(new_n7980), .Y(new_n8212));
  xnor_3 g07836(.A(new_n8198), .B(new_n8194), .Y(new_n8213));
  not_3  g07837(.A(new_n4250), .Y(new_n8214));
  nand_4 g07838(.A(new_n4254), .B(new_n8214), .Y(new_n8215));
  nand_4 g07839(.A(new_n4269), .B(new_n4256), .Y(new_n8216));
  nand_4 g07840(.A(new_n8216), .B(new_n8215), .Y(new_n8217));
  not_3  g07841(.A(new_n8217), .Y(new_n8218));
  nor_4  g07842(.A(new_n8218), .B(new_n8213), .Y(new_n8219));
  xnor_3 g07843(.A(new_n8204), .B(new_n8201), .Y(new_n8220));
  xnor_3 g07844(.A(new_n8220), .B(new_n8219), .Y(new_n8221));
  nand_4 g07845(.A(n9637), .B(n6687), .Y(new_n8222));
  not_3  g07846(.A(new_n8222), .Y(new_n8223));
  not_3  g07847(.A(new_n8213), .Y(new_n8224));
  nor_4  g07848(.A(new_n8217), .B(new_n8224), .Y(new_n8225));
  nor_4  g07849(.A(new_n8225), .B(new_n8219), .Y(new_n8226));
  nand_4 g07850(.A(new_n8226), .B(new_n8223), .Y(new_n8227));
  nor_4  g07851(.A(new_n4270), .B(new_n4249), .Y(new_n8228));
  xnor_3 g07852(.A(new_n8226), .B(new_n8222), .Y(new_n8229));
  nand_4 g07853(.A(new_n8229), .B(new_n8228), .Y(new_n8230));
  nand_4 g07854(.A(new_n8230), .B(new_n8227), .Y(new_n8231));
  xnor_3 g07855(.A(new_n8231), .B(new_n8221), .Y(new_n8232));
  not_3  g07856(.A(new_n8232), .Y(new_n8233));
  xnor_3 g07857(.A(new_n7973), .B(new_n7958), .Y(new_n8234));
  not_3  g07858(.A(new_n8234), .Y(new_n8235));
  nand_4 g07859(.A(new_n8235), .B(new_n8233), .Y(new_n8236_1));
  nand_4 g07860(.A(new_n8234), .B(new_n8232), .Y(new_n8237));
  not_3  g07861(.A(new_n8229), .Y(new_n8238));
  xnor_3 g07862(.A(new_n8238), .B(new_n8228), .Y(new_n8239));
  not_3  g07863(.A(new_n4271), .Y(new_n8240));
  nand_4 g07864(.A(new_n4467), .B(new_n8240), .Y(new_n8241));
  nand_4 g07865(.A(new_n4564), .B(new_n4468), .Y(new_n8242));
  nand_4 g07866(.A(new_n8242), .B(new_n8241), .Y(new_n8243));
  nor_4  g07867(.A(new_n8243), .B(new_n8239), .Y(new_n8244));
  xnor_3 g07868(.A(new_n7971), .B(new_n7967), .Y(new_n8245));
  xnor_3 g07869(.A(new_n8243), .B(new_n8239), .Y(new_n8246));
  nor_4  g07870(.A(new_n8246), .B(new_n8245), .Y(new_n8247));
  nor_4  g07871(.A(new_n8247), .B(new_n8244), .Y(new_n8248));
  nand_4 g07872(.A(new_n8248), .B(new_n8237), .Y(new_n8249));
  nand_4 g07873(.A(new_n8249), .B(new_n8236_1), .Y(new_n8250));
  not_3  g07874(.A(new_n8220), .Y(new_n8251));
  nand_4 g07875(.A(new_n8251), .B(new_n8219), .Y(new_n8252));
  nand_4 g07876(.A(new_n8231), .B(new_n8221), .Y(new_n8253));
  nand_4 g07877(.A(new_n8253), .B(new_n8252), .Y(new_n8254));
  not_3  g07878(.A(new_n7831), .Y(new_n8255));
  nor_4  g07879(.A(new_n8255), .B(new_n7825), .Y(new_n8256));
  not_3  g07880(.A(new_n7832), .Y(new_n8257));
  nor_4  g07881(.A(new_n7843), .B(new_n8257), .Y(new_n8258));
  nor_4  g07882(.A(new_n8258), .B(new_n8256), .Y(new_n8259));
  xnor_3 g07883(.A(new_n8259), .B(new_n8254), .Y(new_n8260));
  xnor_3 g07884(.A(new_n8260), .B(new_n8250), .Y(new_n8261));
  xnor_3 g07885(.A(new_n8261), .B(new_n8212), .Y(n2679));
  not_3  g07886(.A(new_n6000), .Y(new_n8263));
  nor_4  g07887(.A(new_n8263), .B(new_n5972), .Y(new_n8264));
  nand_4 g07888(.A(n6687), .B(n2253), .Y(new_n8265));
  not_3  g07889(.A(new_n8265), .Y(new_n8266));
  nand_4 g07890(.A(n10223), .B(n6770), .Y(new_n8267));
  not_3  g07891(.A(new_n8267), .Y(new_n8268));
  nand_4 g07892(.A(n9920), .B(n2879), .Y(new_n8269));
  nand_4 g07893(.A(n7265), .B(n3627), .Y(new_n8270));
  xnor_3 g07894(.A(new_n8270), .B(new_n8269), .Y(new_n8271));
  xnor_3 g07895(.A(new_n8271), .B(new_n8268), .Y(new_n8272));
  not_3  g07896(.A(new_n5977), .Y(new_n8273));
  not_3  g07897(.A(new_n5978), .Y(new_n8274));
  nor_4  g07898(.A(new_n8274), .B(new_n8273), .Y(new_n8275));
  not_3  g07899(.A(new_n5976), .Y(new_n8276_1));
  nor_4  g07900(.A(new_n5979), .B(new_n8276_1), .Y(new_n8277));
  nor_4  g07901(.A(new_n8277), .B(new_n8275), .Y(new_n8278));
  xnor_3 g07902(.A(new_n8278), .B(new_n8272), .Y(new_n8279));
  not_3  g07903(.A(new_n8279), .Y(new_n8280));
  nand_4 g07904(.A(n9195), .B(n2564), .Y(new_n8281));
  nand_4 g07905(.A(n4634), .B(n4189), .Y(new_n8282));
  xor_3  g07906(.A(new_n8282), .B(new_n8281), .Y(new_n8283));
  not_3  g07907(.A(new_n8283), .Y(new_n8284));
  xor_3  g07908(.A(new_n8284), .B(new_n8280), .Y(new_n8285));
  nor_4  g07909(.A(new_n5980), .B(new_n5975), .Y(new_n8286));
  not_3  g07910(.A(new_n5986), .Y(new_n8287));
  nor_4  g07911(.A(new_n8287), .B(new_n5981), .Y(new_n8288));
  nor_4  g07912(.A(new_n8288), .B(new_n8286), .Y(new_n8289));
  xnor_3 g07913(.A(new_n8289), .B(new_n8285), .Y(new_n8290));
  not_3  g07914(.A(new_n5989), .Y(new_n8291));
  nand_4 g07915(.A(new_n5997), .B(new_n8291), .Y(new_n8292));
  xnor_3 g07916(.A(new_n8292), .B(new_n8290), .Y(new_n8293));
  xnor_3 g07917(.A(new_n8293), .B(new_n8266), .Y(new_n8294));
  xor_3  g07918(.A(new_n8294), .B(new_n8264), .Y(new_n8295));
  not_3  g07919(.A(new_n6001), .Y(new_n8296));
  nand_4 g07920(.A(new_n6254_1), .B(new_n8296), .Y(new_n8297));
  nand_4 g07921(.A(new_n6287), .B(new_n6255), .Y(new_n8298));
  nand_4 g07922(.A(new_n8298), .B(new_n8297), .Y(new_n8299));
  xnor_3 g07923(.A(new_n8299), .B(new_n8295), .Y(new_n8300));
  nor_4  g07924(.A(new_n6054), .B(new_n6031), .Y(new_n8301));
  nand_4 g07925(.A(n12221), .B(n8336), .Y(new_n8302));
  not_3  g07926(.A(new_n8302), .Y(new_n8303_1));
  nand_4 g07927(.A(n9189), .B(n2226), .Y(new_n8304));
  nand_4 g07928(.A(n2024), .B(n1094), .Y(new_n8305));
  nand_4 g07929(.A(n10678), .B(n7946), .Y(new_n8306));
  xnor_3 g07930(.A(new_n8306), .B(new_n8305), .Y(new_n8307));
  nor_4  g07931(.A(new_n8307), .B(new_n8304), .Y(new_n8308));
  not_3  g07932(.A(new_n8304), .Y(new_n8309));
  not_3  g07933(.A(new_n8307), .Y(new_n8310));
  nor_4  g07934(.A(new_n8310), .B(new_n8309), .Y(new_n8311));
  nor_4  g07935(.A(new_n8311), .B(new_n8308), .Y(new_n8312));
  not_3  g07936(.A(new_n6041), .Y(new_n8313));
  not_3  g07937(.A(new_n6042), .Y(new_n8314));
  nor_4  g07938(.A(new_n8314), .B(new_n8313), .Y(new_n8315));
  nor_4  g07939(.A(new_n6043), .B(new_n6040), .Y(new_n8316));
  nor_4  g07940(.A(new_n8316), .B(new_n8315), .Y(new_n8317));
  xnor_3 g07941(.A(new_n8317), .B(new_n8312), .Y(new_n8318));
  not_3  g07942(.A(new_n8318), .Y(new_n8319));
  nand_4 g07943(.A(n12145), .B(n10928), .Y(new_n8320));
  nand_4 g07944(.A(n6986), .B(n2522), .Y(new_n8321));
  xor_3  g07945(.A(new_n8321), .B(new_n8320), .Y(new_n8322));
  not_3  g07946(.A(new_n8322), .Y(new_n8323));
  xor_3  g07947(.A(new_n8323), .B(new_n8319), .Y(new_n8324));
  not_3  g07948(.A(new_n6034), .Y(new_n8325));
  and_4  g07949(.A(new_n6037), .B(new_n8325), .Y(new_n8326));
  nor_4  g07950(.A(new_n6044), .B(new_n6038_1), .Y(new_n8327));
  nor_4  g07951(.A(new_n8327), .B(new_n8326), .Y(new_n8328));
  xnor_3 g07952(.A(new_n8328), .B(new_n8324), .Y(new_n8329));
  nand_4 g07953(.A(new_n6046), .B(new_n6033), .Y(new_n8330));
  nand_4 g07954(.A(new_n6053), .B(new_n6047), .Y(new_n8331));
  nand_4 g07955(.A(new_n8331), .B(new_n8330), .Y(new_n8332));
  not_3  g07956(.A(new_n8332), .Y(new_n8333));
  nor_4  g07957(.A(new_n8333), .B(new_n8329), .Y(new_n8334));
  not_3  g07958(.A(new_n8329), .Y(new_n8335));
  nor_4  g07959(.A(new_n8332), .B(new_n8335), .Y(new_n8336_1));
  nor_4  g07960(.A(new_n8336_1), .B(new_n8334), .Y(new_n8337));
  xnor_3 g07961(.A(new_n8337), .B(new_n8303_1), .Y(new_n8338));
  xnor_3 g07962(.A(new_n8338), .B(new_n8301), .Y(new_n8339));
  not_3  g07963(.A(new_n6190), .Y(new_n8340));
  nor_4  g07964(.A(new_n8340), .B(new_n6055), .Y(new_n8341));
  not_3  g07965(.A(new_n8341), .Y(new_n8342));
  nand_4 g07966(.A(new_n6253), .B(new_n6191), .Y(new_n8343));
  nand_4 g07967(.A(new_n8343), .B(new_n8342), .Y(new_n8344));
  xnor_3 g07968(.A(new_n8344), .B(new_n8339), .Y(new_n8345));
  not_3  g07969(.A(new_n6091), .Y(new_n8346));
  nor_4  g07970(.A(new_n6212), .B(new_n8346), .Y(new_n8347));
  not_3  g07971(.A(new_n8347), .Y(new_n8348));
  nand_4 g07972(.A(n12069), .B(n5798), .Y(new_n8349));
  nand_4 g07973(.A(n7160), .B(n5579), .Y(new_n8350));
  not_3  g07974(.A(new_n8350), .Y(new_n8351));
  nor_4  g07975(.A(new_n6205), .B(new_n6200), .Y(new_n8352));
  nor_4  g07976(.A(new_n8352), .B(new_n8351), .Y(new_n8353));
  nor_4  g07977(.A(new_n8352), .B(new_n6081), .Y(new_n8354));
  nor_4  g07978(.A(new_n8354), .B(new_n8350), .Y(new_n8355));
  nor_4  g07979(.A(new_n8355), .B(new_n8353), .Y(new_n8356));
  nand_4 g07980(.A(n4828), .B(n2498), .Y(new_n8357));
  nand_4 g07981(.A(n2558), .B(n2515), .Y(new_n8358));
  xor_3  g07982(.A(new_n8358), .B(new_n8357), .Y(new_n8359));
  xnor_3 g07983(.A(new_n8359), .B(new_n8356), .Y(new_n8360));
  nand_4 g07984(.A(n12391), .B(n6016), .Y(new_n8361));
  nand_4 g07985(.A(n7891), .B(n521), .Y(new_n8362));
  not_3  g07986(.A(new_n8362), .Y(new_n8363));
  xor_3  g07987(.A(new_n8363), .B(new_n8361), .Y(new_n8364));
  xnor_3 g07988(.A(new_n8364), .B(new_n8360), .Y(new_n8365));
  and_4  g07989(.A(new_n6196), .B(new_n6194), .Y(new_n8366));
  nor_4  g07990(.A(new_n6206), .B(new_n6197), .Y(new_n8367));
  nor_4  g07991(.A(new_n8367), .B(new_n8366), .Y(new_n8368));
  xnor_3 g07992(.A(new_n8368), .B(new_n8365), .Y(new_n8369));
  nor_4  g07993(.A(new_n6207), .B(new_n6192_1), .Y(new_n8370));
  nor_4  g07994(.A(new_n6211), .B(new_n6208), .Y(new_n8371));
  nor_4  g07995(.A(new_n8371), .B(new_n8370), .Y(new_n8372));
  xnor_3 g07996(.A(new_n8372), .B(new_n8369), .Y(new_n8373));
  xnor_3 g07997(.A(new_n8373), .B(new_n8349), .Y(new_n8374));
  xnor_3 g07998(.A(new_n8374), .B(new_n8348), .Y(new_n8375));
  not_3  g07999(.A(new_n6248), .Y(new_n8376));
  nand_4 g08000(.A(n11222), .B(n5153), .Y(new_n8377));
  nand_4 g08001(.A(n3342), .B(n996), .Y(new_n8378));
  nand_4 g08002(.A(n9111), .B(n5767), .Y(new_n8379));
  nand_4 g08003(.A(n9763), .B(n5319), .Y(new_n8380));
  xnor_3 g08004(.A(new_n8380), .B(new_n8379), .Y(new_n8381));
  nor_4  g08005(.A(new_n8381), .B(new_n8378), .Y(new_n8382));
  not_3  g08006(.A(new_n8378), .Y(new_n8383));
  not_3  g08007(.A(new_n8381), .Y(new_n8384_1));
  nor_4  g08008(.A(new_n8384_1), .B(new_n8383), .Y(new_n8385));
  nor_4  g08009(.A(new_n8385), .B(new_n8382), .Y(new_n8386));
  nor_4  g08010(.A(new_n6233), .B(new_n6227), .Y(new_n8387));
  nor_4  g08011(.A(new_n8387), .B(new_n6232), .Y(new_n8388));
  xnor_3 g08012(.A(new_n8388), .B(new_n8386), .Y(new_n8389));
  not_3  g08013(.A(new_n8389), .Y(new_n8390));
  nand_4 g08014(.A(n11153), .B(n7270), .Y(new_n8391));
  nand_4 g08015(.A(n5314), .B(n806), .Y(new_n8392));
  xor_3  g08016(.A(new_n8392), .B(new_n8391), .Y(new_n8393));
  xnor_3 g08017(.A(new_n8393), .B(new_n8390), .Y(new_n8394));
  and_4  g08018(.A(new_n6224), .B(new_n6217), .Y(new_n8395));
  nor_4  g08019(.A(new_n6235), .B(new_n6225), .Y(new_n8396));
  nor_4  g08020(.A(new_n8396), .B(new_n8395), .Y(new_n8397));
  xnor_3 g08021(.A(new_n8397), .B(new_n8394), .Y(new_n8398_1));
  not_3  g08022(.A(new_n6237), .Y(new_n8399));
  nand_4 g08023(.A(new_n6243), .B(new_n6241), .Y(new_n8400));
  nand_4 g08024(.A(new_n8400), .B(new_n8399), .Y(new_n8401));
  not_3  g08025(.A(new_n8401), .Y(new_n8402));
  xnor_3 g08026(.A(new_n8402), .B(new_n8398_1), .Y(new_n8403));
  xnor_3 g08027(.A(new_n8403), .B(new_n8377), .Y(new_n8404));
  not_3  g08028(.A(new_n8404), .Y(new_n8405));
  nor_4  g08029(.A(new_n8405), .B(new_n8376), .Y(new_n8406));
  nor_4  g08030(.A(new_n8404), .B(new_n6248), .Y(new_n8407));
  nor_4  g08031(.A(new_n8407), .B(new_n8406), .Y(new_n8408));
  nand_4 g08032(.A(new_n8408), .B(new_n8375), .Y(new_n8409));
  not_3  g08033(.A(new_n8375), .Y(new_n8410));
  not_3  g08034(.A(new_n8408), .Y(new_n8411));
  nand_4 g08035(.A(new_n8411), .B(new_n8410), .Y(new_n8412));
  nand_4 g08036(.A(new_n8412), .B(new_n8409), .Y(new_n8413));
  nor_4  g08037(.A(new_n6249), .B(new_n6214), .Y(new_n8414));
  nor_4  g08038(.A(new_n6252), .B(new_n6250), .Y(new_n8415));
  nor_4  g08039(.A(new_n8415), .B(new_n8414), .Y(new_n8416));
  xnor_3 g08040(.A(new_n8416), .B(new_n8413), .Y(new_n8417));
  not_3  g08041(.A(new_n8417), .Y(new_n8418));
  xnor_3 g08042(.A(new_n8418), .B(new_n8345), .Y(new_n8419));
  nor_4  g08043(.A(new_n8419), .B(new_n8300), .Y(new_n8420));
  not_3  g08044(.A(new_n8300), .Y(new_n8421));
  not_3  g08045(.A(new_n8419), .Y(new_n8422));
  nor_4  g08046(.A(new_n8422), .B(new_n8421), .Y(new_n8423));
  nor_4  g08047(.A(new_n8423), .B(new_n8420), .Y(n2708));
  xor_3  g08048(.A(new_n1050), .B(new_n1049), .Y(n2818));
  xnor_3 g08049(.A(new_n2189), .B(new_n2164), .Y(n2902));
  nand_4 g08050(.A(n11407), .B(n5305), .Y(new_n8427));
  not_3  g08051(.A(new_n8427), .Y(new_n8428));
  nand_4 g08052(.A(n12709), .B(n8759), .Y(new_n8429));
  not_3  g08053(.A(new_n8429), .Y(new_n8430));
  nand_4 g08054(.A(n12489), .B(n5331), .Y(new_n8431));
  nand_4 g08055(.A(n10990), .B(n7965), .Y(new_n8432));
  not_3  g08056(.A(new_n8432), .Y(new_n8433_1));
  xor_3  g08057(.A(new_n8433_1), .B(new_n8431), .Y(new_n8434));
  not_3  g08058(.A(new_n8434), .Y(new_n8435));
  xor_3  g08059(.A(new_n8435), .B(new_n8430), .Y(new_n8436));
  xor_3  g08060(.A(new_n8436), .B(new_n8428), .Y(n3071));
  not_3  g08061(.A(new_n3084), .Y(new_n8438));
  xor_3  g08062(.A(new_n3087), .B(new_n8438), .Y(n3124));
  nand_4 g08063(.A(new_n8436), .B(new_n8428), .Y(new_n8440));
  nand_4 g08064(.A(n11407), .B(n5964), .Y(new_n8441));
  nand_4 g08065(.A(n5305), .B(n5212), .Y(new_n8442));
  xor_3  g08066(.A(new_n8442), .B(new_n8441), .Y(new_n8443));
  not_3  g08067(.A(new_n8443), .Y(new_n8444));
  nand_4 g08068(.A(new_n8444), .B(new_n8440), .Y(new_n8445));
  nor_4  g08069(.A(new_n8434), .B(new_n8429), .Y(new_n8446));
  nand_4 g08070(.A(n11728), .B(n8759), .Y(new_n8447));
  nand_4 g08071(.A(n12709), .B(n6776), .Y(new_n8448));
  not_3  g08072(.A(new_n8448), .Y(new_n8449));
  xor_3  g08073(.A(new_n8449), .B(new_n8447), .Y(new_n8450));
  not_3  g08074(.A(new_n8450), .Y(new_n8451));
  nand_4 g08075(.A(new_n8451), .B(new_n8446), .Y(new_n8452));
  not_3  g08076(.A(new_n8452), .Y(new_n8453));
  nor_4  g08077(.A(new_n8451), .B(new_n8446), .Y(new_n8454));
  nor_4  g08078(.A(new_n8454), .B(new_n8453), .Y(new_n8455));
  not_3  g08079(.A(new_n8455), .Y(new_n8456));
  nor_4  g08080(.A(new_n8432), .B(new_n8431), .Y(new_n8457));
  nand_4 g08081(.A(n7159), .B(n5331), .Y(new_n8458));
  nand_4 g08082(.A(n12489), .B(n8476), .Y(new_n8459));
  not_3  g08083(.A(new_n8459), .Y(new_n8460));
  xor_3  g08084(.A(new_n8460), .B(new_n8458), .Y(new_n8461));
  not_3  g08085(.A(new_n8461), .Y(new_n8462));
  xor_3  g08086(.A(new_n8462), .B(new_n8457), .Y(new_n8463));
  nand_4 g08087(.A(n7965), .B(n5760), .Y(new_n8464));
  nand_4 g08088(.A(n10990), .B(n7388), .Y(new_n8465));
  xor_3  g08089(.A(new_n8465), .B(new_n8464), .Y(new_n8466));
  not_3  g08090(.A(new_n8466), .Y(new_n8467));
  nor_4  g08091(.A(new_n8467), .B(new_n8463), .Y(new_n8468));
  not_3  g08092(.A(new_n8463), .Y(new_n8469));
  nor_4  g08093(.A(new_n8466), .B(new_n8469), .Y(new_n8470));
  nor_4  g08094(.A(new_n8470), .B(new_n8468), .Y(new_n8471));
  xnor_3 g08095(.A(new_n8471), .B(new_n8456), .Y(new_n8472));
  not_3  g08096(.A(new_n8445), .Y(new_n8473));
  nor_4  g08097(.A(new_n8444), .B(new_n8440), .Y(new_n8474));
  nor_4  g08098(.A(new_n8474), .B(new_n8473), .Y(new_n8475));
  nand_4 g08099(.A(new_n8475), .B(new_n8472), .Y(new_n8476_1));
  nand_4 g08100(.A(new_n8476_1), .B(new_n8445), .Y(new_n8477));
  nand_4 g08101(.A(n5964), .B(n5212), .Y(new_n8478));
  nor_4  g08102(.A(new_n8478), .B(new_n8428), .Y(new_n8479));
  nand_4 g08103(.A(n11407), .B(n1097), .Y(new_n8480));
  nand_4 g08104(.A(n11877), .B(n5305), .Y(new_n8481));
  nand_4 g08105(.A(new_n8481), .B(new_n8480), .Y(new_n8482));
  nor_4  g08106(.A(new_n8482), .B(new_n8479), .Y(new_n8483));
  nor_4  g08107(.A(new_n8481), .B(new_n8480), .Y(new_n8484));
  nor_4  g08108(.A(new_n8484), .B(new_n8483), .Y(new_n8485));
  not_3  g08109(.A(new_n8485), .Y(new_n8486));
  not_3  g08110(.A(new_n8479), .Y(new_n8487));
  not_3  g08111(.A(new_n8482), .Y(new_n8488));
  nor_4  g08112(.A(new_n8488), .B(new_n8487), .Y(new_n8489));
  nor_4  g08113(.A(new_n8489), .B(new_n8486), .Y(new_n8490));
  not_3  g08114(.A(new_n8490), .Y(new_n8491));
  nor_4  g08115(.A(new_n8491), .B(new_n8477), .Y(new_n8492));
  not_3  g08116(.A(new_n8477), .Y(new_n8493));
  nor_4  g08117(.A(new_n8490), .B(new_n8493), .Y(new_n8494));
  nor_4  g08118(.A(new_n8494), .B(new_n8492), .Y(new_n8495));
  nor_4  g08119(.A(new_n8471), .B(new_n8456), .Y(new_n8496));
  nor_4  g08120(.A(new_n8496), .B(new_n8453), .Y(new_n8497));
  nand_4 g08121(.A(n11728), .B(n6776), .Y(new_n8498));
  nor_4  g08122(.A(new_n8498), .B(new_n8430), .Y(new_n8499));
  nand_4 g08123(.A(n12709), .B(n12299), .Y(new_n8500));
  not_3  g08124(.A(new_n8500), .Y(new_n8501));
  nand_4 g08125(.A(n8759), .B(n6429), .Y(new_n8502));
  not_3  g08126(.A(new_n8502), .Y(new_n8503));
  nand_4 g08127(.A(new_n8503), .B(new_n8501), .Y(new_n8504));
  nand_4 g08128(.A(new_n8502), .B(new_n8500), .Y(new_n8505));
  and_4  g08129(.A(new_n8505), .B(new_n8504), .Y(new_n8506));
  nor_4  g08130(.A(new_n8506), .B(new_n8499), .Y(new_n8507));
  not_3  g08131(.A(new_n8498), .Y(new_n8508));
  nand_4 g08132(.A(new_n8505), .B(new_n8508), .Y(new_n8509));
  nor_4  g08133(.A(new_n8509), .B(new_n8430), .Y(new_n8510));
  nor_4  g08134(.A(new_n8510), .B(new_n8507), .Y(new_n8511));
  xnor_3 g08135(.A(new_n8511), .B(new_n8497), .Y(new_n8512));
  not_3  g08136(.A(new_n8431), .Y(new_n8513));
  nand_4 g08137(.A(n8476), .B(n7159), .Y(new_n8514));
  nor_4  g08138(.A(new_n8514), .B(new_n8513), .Y(new_n8515));
  nand_4 g08139(.A(n12489), .B(n2530), .Y(new_n8516));
  not_3  g08140(.A(new_n8516), .Y(new_n8517));
  nand_4 g08141(.A(n12777), .B(n5331), .Y(new_n8518));
  not_3  g08142(.A(new_n8518), .Y(new_n8519));
  nor_4  g08143(.A(new_n8519), .B(new_n8517), .Y(new_n8520));
  nor_4  g08144(.A(new_n8518), .B(new_n8516), .Y(new_n8521));
  nor_4  g08145(.A(new_n8521), .B(new_n8520), .Y(new_n8522));
  nor_4  g08146(.A(new_n8522), .B(new_n8515), .Y(new_n8523));
  not_3  g08147(.A(new_n8523), .Y(new_n8524));
  not_3  g08148(.A(new_n8520), .Y(new_n8525));
  nand_4 g08149(.A(new_n8525), .B(new_n8515), .Y(new_n8526));
  nand_4 g08150(.A(new_n8526), .B(new_n8524), .Y(new_n8527));
  nand_4 g08151(.A(n7388), .B(n5760), .Y(new_n8528));
  nor_4  g08152(.A(new_n8528), .B(new_n8433_1), .Y(new_n8529));
  nand_4 g08153(.A(n11892), .B(n10990), .Y(new_n8530));
  not_3  g08154(.A(new_n8530), .Y(new_n8531));
  nand_4 g08155(.A(n7965), .B(n1478), .Y(new_n8532));
  not_3  g08156(.A(new_n8532), .Y(new_n8533));
  nor_4  g08157(.A(new_n8533), .B(new_n8531), .Y(new_n8534));
  nor_4  g08158(.A(new_n8532), .B(new_n8530), .Y(new_n8535));
  nor_4  g08159(.A(new_n8535), .B(new_n8534), .Y(new_n8536));
  nor_4  g08160(.A(new_n8536), .B(new_n8529), .Y(new_n8537));
  not_3  g08161(.A(new_n8537), .Y(new_n8538));
  not_3  g08162(.A(new_n8534), .Y(new_n8539));
  nand_4 g08163(.A(new_n8539), .B(new_n8529), .Y(new_n8540));
  nand_4 g08164(.A(new_n8540), .B(new_n8538), .Y(new_n8541));
  xor_3  g08165(.A(new_n8541), .B(new_n8527), .Y(new_n8542));
  nor_4  g08166(.A(new_n8462), .B(new_n8457), .Y(new_n8543));
  nor_4  g08167(.A(new_n8470), .B(new_n8543), .Y(new_n8544));
  nand_4 g08168(.A(new_n8544), .B(new_n8542), .Y(new_n8545));
  not_3  g08169(.A(new_n8545), .Y(new_n8546));
  nor_4  g08170(.A(new_n8544), .B(new_n8542), .Y(new_n8547));
  nor_4  g08171(.A(new_n8547), .B(new_n8546), .Y(new_n8548));
  nand_4 g08172(.A(new_n8548), .B(new_n8512), .Y(new_n8549));
  not_3  g08173(.A(new_n8549), .Y(new_n8550));
  nor_4  g08174(.A(new_n8548), .B(new_n8512), .Y(new_n8551));
  nor_4  g08175(.A(new_n8551), .B(new_n8550), .Y(new_n8552));
  xor_3  g08176(.A(new_n8552), .B(new_n8495), .Y(n3214));
  not_3  g08177(.A(new_n5802), .Y(new_n8554));
  nor_4  g08178(.A(new_n5798_1), .B(new_n5796), .Y(new_n8555));
  xor_3  g08179(.A(new_n8555), .B(new_n8554), .Y(n3230));
  not_3  g08180(.A(new_n5279), .Y(new_n8557));
  nand_4 g08181(.A(new_n5225), .B(new_n5223), .Y(new_n8558));
  xnor_3 g08182(.A(new_n8558), .B(new_n8557), .Y(n3272));
  nand_4 g08183(.A(n5964), .B(n4370), .Y(new_n8560));
  not_3  g08184(.A(new_n8560), .Y(new_n8561));
  nand_4 g08185(.A(n11407), .B(n4312), .Y(new_n8562));
  not_3  g08186(.A(new_n8562), .Y(new_n8563));
  nand_4 g08187(.A(n11877), .B(n5964), .Y(new_n8564));
  not_3  g08188(.A(new_n8564), .Y(new_n8565));
  nor_4  g08189(.A(new_n8565), .B(new_n8563), .Y(new_n8566));
  nor_4  g08190(.A(new_n8564), .B(new_n8562), .Y(new_n8567));
  nand_4 g08191(.A(n5212), .B(n1097), .Y(new_n8568));
  not_3  g08192(.A(new_n8568), .Y(new_n8569));
  nor_4  g08193(.A(new_n8569), .B(new_n8567), .Y(new_n8570));
  nor_4  g08194(.A(new_n8570), .B(new_n8566), .Y(new_n8571));
  nand_4 g08195(.A(new_n8571), .B(new_n8561), .Y(new_n8572));
  xor_3  g08196(.A(new_n8571), .B(new_n8561), .Y(new_n8573));
  nand_4 g08197(.A(n5212), .B(n4312), .Y(new_n8574));
  not_3  g08198(.A(new_n8574), .Y(new_n8575));
  nand_4 g08199(.A(n11877), .B(n1097), .Y(new_n8576));
  not_3  g08200(.A(new_n8576), .Y(new_n8577));
  nand_4 g08201(.A(n12705), .B(n11407), .Y(new_n8578));
  not_3  g08202(.A(new_n8578), .Y(new_n8579));
  nor_4  g08203(.A(new_n8579), .B(new_n8577), .Y(new_n8580));
  nor_4  g08204(.A(new_n8578), .B(new_n8576), .Y(new_n8581));
  nor_4  g08205(.A(new_n8581), .B(new_n8580), .Y(new_n8582));
  xor_3  g08206(.A(new_n8582), .B(new_n8575), .Y(new_n8583));
  nand_4 g08207(.A(new_n8583), .B(new_n8573), .Y(new_n8584));
  nand_4 g08208(.A(new_n8584), .B(new_n8572), .Y(new_n8585));
  not_3  g08209(.A(new_n8585), .Y(new_n8586));
  nand_4 g08210(.A(n5964), .B(n5320), .Y(new_n8587));
  nand_4 g08211(.A(n4370), .B(n1097), .Y(new_n8588));
  xor_3  g08212(.A(new_n8588), .B(new_n8587), .Y(new_n8589));
  not_3  g08213(.A(new_n8589), .Y(new_n8590));
  xor_3  g08214(.A(new_n8590), .B(new_n8586), .Y(new_n8591));
  nand_4 g08215(.A(n11877), .B(n4312), .Y(new_n8592));
  not_3  g08216(.A(new_n8592), .Y(new_n8593));
  nand_4 g08217(.A(n12705), .B(n5212), .Y(new_n8594));
  nand_4 g08218(.A(n12025), .B(n11407), .Y(new_n8595_1));
  xnor_3 g08219(.A(new_n8595_1), .B(new_n8594), .Y(new_n8596));
  xnor_3 g08220(.A(new_n8596), .B(new_n8593), .Y(new_n8597));
  nor_4  g08221(.A(new_n8581), .B(new_n8575), .Y(new_n8598));
  nor_4  g08222(.A(new_n8598), .B(new_n8580), .Y(new_n8599));
  xor_3  g08223(.A(new_n8599), .B(new_n8597), .Y(new_n8600));
  xnor_3 g08224(.A(new_n8600), .B(new_n8591), .Y(new_n8601));
  nand_4 g08225(.A(n5320), .B(n5305), .Y(new_n8602));
  xnor_3 g08226(.A(new_n8583), .B(new_n8573), .Y(new_n8603));
  nand_4 g08227(.A(new_n8603), .B(new_n8602), .Y(new_n8604));
  not_3  g08228(.A(new_n8602), .Y(new_n8605));
  not_3  g08229(.A(new_n8603), .Y(new_n8606));
  xor_3  g08230(.A(new_n8606), .B(new_n8605), .Y(new_n8607));
  nand_4 g08231(.A(n5305), .B(n4370), .Y(new_n8608));
  not_3  g08232(.A(new_n8608), .Y(new_n8609));
  not_3  g08233(.A(new_n8478), .Y(new_n8610));
  nor_4  g08234(.A(new_n8484), .B(new_n8610), .Y(new_n8611));
  nor_4  g08235(.A(new_n8611), .B(new_n8488), .Y(new_n8612));
  and_4  g08236(.A(new_n8612), .B(new_n8609), .Y(new_n8613));
  xor_3  g08237(.A(new_n8612), .B(new_n8608), .Y(new_n8614));
  nor_4  g08238(.A(new_n8567), .B(new_n8566), .Y(new_n8615));
  xor_3  g08239(.A(new_n8615), .B(new_n8568), .Y(new_n8616));
  nor_4  g08240(.A(new_n8616), .B(new_n8614), .Y(new_n8617));
  nor_4  g08241(.A(new_n8617), .B(new_n8613), .Y(new_n8618));
  nand_4 g08242(.A(new_n8618), .B(new_n8607), .Y(new_n8619));
  nand_4 g08243(.A(new_n8619), .B(new_n8604), .Y(new_n8620));
  nor_4  g08244(.A(new_n8620), .B(new_n8601), .Y(new_n8621));
  not_3  g08245(.A(new_n8621), .Y(new_n8622));
  nand_4 g08246(.A(new_n8596), .B(new_n8592), .Y(new_n8623));
  not_3  g08247(.A(new_n8599), .Y(new_n8624));
  nand_4 g08248(.A(new_n8624), .B(new_n8597), .Y(new_n8625));
  and_4  g08249(.A(new_n8625), .B(new_n8623), .Y(new_n8626));
  nand_4 g08250(.A(n12000), .B(n5964), .Y(new_n8627));
  nand_4 g08251(.A(n5320), .B(n1097), .Y(new_n8628));
  nand_4 g08252(.A(n9725), .B(n5305), .Y(new_n8629));
  not_3  g08253(.A(new_n8629), .Y(new_n8630));
  xor_3  g08254(.A(new_n8630), .B(new_n8628), .Y(new_n8631));
  xnor_3 g08255(.A(new_n8631), .B(new_n8627), .Y(new_n8632));
  xnor_3 g08256(.A(new_n8632), .B(new_n8626), .Y(new_n8633));
  not_3  g08257(.A(new_n8633), .Y(new_n8634));
  nor_4  g08258(.A(new_n8595_1), .B(new_n8594), .Y(new_n8635));
  nand_4 g08259(.A(n4370), .B(n4312), .Y(new_n8636));
  xor_3  g08260(.A(new_n8636), .B(new_n8635), .Y(new_n8637));
  nand_4 g08261(.A(n12025), .B(n5212), .Y(new_n8638));
  nand_4 g08262(.A(n12705), .B(n11877), .Y(new_n8639));
  nand_4 g08263(.A(n11407), .B(n11257), .Y(new_n8640));
  not_3  g08264(.A(new_n8640), .Y(new_n8641));
  xor_3  g08265(.A(new_n8641), .B(new_n8639), .Y(new_n8642));
  xnor_3 g08266(.A(new_n8642), .B(new_n8638), .Y(new_n8643));
  xnor_3 g08267(.A(new_n8643), .B(new_n8637), .Y(new_n8644));
  xnor_3 g08268(.A(new_n8644), .B(new_n8634), .Y(new_n8645));
  nor_4  g08269(.A(new_n8590), .B(new_n8586), .Y(new_n8646));
  nor_4  g08270(.A(new_n8588), .B(new_n8587), .Y(new_n8647));
  nand_4 g08271(.A(new_n8600), .B(new_n8591), .Y(new_n8648));
  xnor_3 g08272(.A(new_n8648), .B(new_n8647), .Y(new_n8649));
  nor_4  g08273(.A(new_n8649), .B(new_n8646), .Y(new_n8650));
  not_3  g08274(.A(new_n8650), .Y(new_n8651));
  xnor_3 g08275(.A(new_n8651), .B(new_n8645), .Y(new_n8652));
  xnor_3 g08276(.A(new_n8652), .B(new_n8622), .Y(new_n8653));
  nand_4 g08277(.A(n12000), .B(n5305), .Y(new_n8654));
  xnor_3 g08278(.A(new_n8620), .B(new_n8601), .Y(new_n8655));
  nor_4  g08279(.A(new_n8655), .B(new_n8654), .Y(new_n8656));
  not_3  g08280(.A(new_n8656), .Y(new_n8657));
  xor_3  g08281(.A(new_n8616), .B(new_n8614), .Y(new_n8658));
  nor_4  g08282(.A(new_n8485), .B(new_n8478), .Y(new_n8659));
  nand_4 g08283(.A(new_n8659), .B(new_n8658), .Y(new_n8660));
  not_3  g08284(.A(new_n8619), .Y(new_n8661));
  nor_4  g08285(.A(new_n8618), .B(new_n8607), .Y(new_n8662));
  nor_4  g08286(.A(new_n8662), .B(new_n8661), .Y(new_n8663));
  nor_4  g08287(.A(new_n8663), .B(new_n8660), .Y(new_n8664));
  not_3  g08288(.A(new_n8654), .Y(new_n8665_1));
  not_3  g08289(.A(new_n8655), .Y(new_n8666));
  nor_4  g08290(.A(new_n8666), .B(new_n8665_1), .Y(new_n8667));
  nor_4  g08291(.A(new_n8667), .B(new_n8656), .Y(new_n8668));
  nand_4 g08292(.A(new_n8668), .B(new_n8664), .Y(new_n8669));
  nand_4 g08293(.A(new_n8669), .B(new_n8657), .Y(new_n8670));
  xnor_3 g08294(.A(new_n8670), .B(new_n8653), .Y(new_n8671));
  not_3  g08295(.A(new_n8671), .Y(new_n8672));
  nand_4 g08296(.A(n8759), .B(n8717), .Y(new_n8673));
  not_3  g08297(.A(new_n8673), .Y(new_n8674));
  nand_4 g08298(.A(n7436), .B(n6429), .Y(new_n8675));
  not_3  g08299(.A(new_n8675), .Y(new_n8676));
  nand_4 g08300(.A(n12709), .B(n9241), .Y(new_n8677));
  nand_4 g08301(.A(n11728), .B(n8276), .Y(new_n8678));
  xnor_3 g08302(.A(new_n8678), .B(new_n8677), .Y(new_n8679));
  xnor_3 g08303(.A(new_n8679), .B(new_n8676), .Y(new_n8680));
  nand_4 g08304(.A(n12299), .B(n6429), .Y(new_n8681));
  not_3  g08305(.A(new_n8681), .Y(new_n8682));
  nand_4 g08306(.A(n12709), .B(n8276), .Y(new_n8683));
  not_3  g08307(.A(new_n8683), .Y(new_n8684));
  nor_4  g08308(.A(new_n8684), .B(new_n8682), .Y(new_n8685));
  nor_4  g08309(.A(new_n8683), .B(new_n8681), .Y(new_n8686));
  nand_4 g08310(.A(n11728), .B(n7436), .Y(new_n8687));
  not_3  g08311(.A(new_n8687), .Y(new_n8688));
  nor_4  g08312(.A(new_n8688), .B(new_n8686), .Y(new_n8689));
  nor_4  g08313(.A(new_n8689), .B(new_n8685), .Y(new_n8690));
  xor_3  g08314(.A(new_n8690), .B(new_n8680), .Y(new_n8691));
  nand_4 g08315(.A(n6776), .B(n2433), .Y(new_n8692));
  nand_4 g08316(.A(n12299), .B(n8819), .Y(new_n8693));
  xor_3  g08317(.A(new_n8693), .B(new_n8692), .Y(new_n8694));
  xnor_3 g08318(.A(new_n8694), .B(new_n8691), .Y(new_n8695));
  not_3  g08319(.A(new_n8695), .Y(new_n8696));
  nand_4 g08320(.A(n8819), .B(n6776), .Y(new_n8697));
  not_3  g08321(.A(new_n8697), .Y(new_n8698));
  nand_4 g08322(.A(n12709), .B(n7436), .Y(new_n8699));
  not_3  g08323(.A(new_n8699), .Y(new_n8700));
  nand_4 g08324(.A(n6776), .B(n6429), .Y(new_n8701));
  not_3  g08325(.A(new_n8701), .Y(new_n8702));
  nor_4  g08326(.A(new_n8702), .B(new_n8700), .Y(new_n8703));
  nor_4  g08327(.A(new_n8701), .B(new_n8699), .Y(new_n8704));
  nand_4 g08328(.A(n12299), .B(n11728), .Y(new_n8705));
  not_3  g08329(.A(new_n8705), .Y(new_n8706));
  nor_4  g08330(.A(new_n8706), .B(new_n8704), .Y(new_n8707));
  nor_4  g08331(.A(new_n8707), .B(new_n8703), .Y(new_n8708));
  and_4  g08332(.A(new_n8708), .B(new_n8698), .Y(new_n8709));
  xor_3  g08333(.A(new_n8708), .B(new_n8697), .Y(new_n8710));
  nor_4  g08334(.A(new_n8686), .B(new_n8685), .Y(new_n8711));
  xor_3  g08335(.A(new_n8711), .B(new_n8687), .Y(new_n8712));
  nor_4  g08336(.A(new_n8712), .B(new_n8710), .Y(new_n8713));
  nor_4  g08337(.A(new_n8713), .B(new_n8709), .Y(new_n8714));
  xnor_3 g08338(.A(new_n8714), .B(new_n8696), .Y(new_n8715));
  nand_4 g08339(.A(n8759), .B(n2433), .Y(new_n8716));
  xnor_3 g08340(.A(new_n8712), .B(new_n8710), .Y(new_n8717_1));
  nand_4 g08341(.A(new_n8717_1), .B(new_n8716), .Y(new_n8718));
  not_3  g08342(.A(new_n8716), .Y(new_n8719));
  not_3  g08343(.A(new_n8717_1), .Y(new_n8720));
  xor_3  g08344(.A(new_n8720), .B(new_n8719), .Y(new_n8721));
  nand_4 g08345(.A(n8819), .B(n8759), .Y(new_n8722));
  nand_4 g08346(.A(new_n8509), .B(new_n8504), .Y(new_n8723));
  not_3  g08347(.A(new_n8723), .Y(new_n8724));
  nor_4  g08348(.A(new_n8724), .B(new_n8722), .Y(new_n8725));
  xor_3  g08349(.A(new_n8723), .B(new_n8722), .Y(new_n8726));
  nor_4  g08350(.A(new_n8704), .B(new_n8703), .Y(new_n8727));
  xor_3  g08351(.A(new_n8727), .B(new_n8705), .Y(new_n8728));
  nor_4  g08352(.A(new_n8728), .B(new_n8726), .Y(new_n8729));
  nor_4  g08353(.A(new_n8729), .B(new_n8725), .Y(new_n8730));
  nand_4 g08354(.A(new_n8730), .B(new_n8721), .Y(new_n8731));
  nand_4 g08355(.A(new_n8731), .B(new_n8718), .Y(new_n8732));
  xnor_3 g08356(.A(new_n8732), .B(new_n8715), .Y(new_n8733));
  nand_4 g08357(.A(new_n8733), .B(new_n8674), .Y(new_n8734));
  not_3  g08358(.A(new_n8726), .Y(new_n8735));
  not_3  g08359(.A(new_n8728), .Y(new_n8736));
  xor_3  g08360(.A(new_n8736), .B(new_n8735), .Y(new_n8737));
  not_3  g08361(.A(new_n8737), .Y(new_n8738));
  not_3  g08362(.A(new_n8507), .Y(new_n8739));
  nor_4  g08363(.A(new_n8739), .B(new_n8498), .Y(new_n8740));
  not_3  g08364(.A(new_n8740), .Y(new_n8741));
  nor_4  g08365(.A(new_n8741), .B(new_n8738), .Y(new_n8742));
  xnor_3 g08366(.A(new_n8730), .B(new_n8721), .Y(new_n8743));
  nand_4 g08367(.A(new_n8743), .B(new_n8742), .Y(new_n8744));
  not_3  g08368(.A(new_n8744), .Y(new_n8745));
  xnor_3 g08369(.A(new_n8733), .B(new_n8673), .Y(new_n8746));
  nand_4 g08370(.A(new_n8746), .B(new_n8745), .Y(new_n8747));
  nand_4 g08371(.A(new_n8747), .B(new_n8734), .Y(new_n8748));
  not_3  g08372(.A(new_n8715), .Y(new_n8749));
  nor_4  g08373(.A(new_n8732), .B(new_n8749), .Y(new_n8750));
  nand_4 g08374(.A(new_n8679), .B(new_n8675), .Y(new_n8751));
  not_3  g08375(.A(new_n8690), .Y(new_n8752));
  nand_4 g08376(.A(new_n8752), .B(new_n8680), .Y(new_n8753));
  and_4  g08377(.A(new_n8753), .B(new_n8751), .Y(new_n8754));
  nand_4 g08378(.A(n8717), .B(n6776), .Y(new_n8755));
  not_3  g08379(.A(new_n8755), .Y(new_n8756));
  nand_4 g08380(.A(n12299), .B(n2433), .Y(new_n8757));
  nand_4 g08381(.A(n8759), .B(n7730), .Y(new_n8758));
  nor_4  g08382(.A(new_n8758), .B(new_n8757), .Y(new_n8759_1));
  not_3  g08383(.A(new_n8757), .Y(new_n8760));
  not_3  g08384(.A(new_n8758), .Y(new_n8761));
  nor_4  g08385(.A(new_n8761), .B(new_n8760), .Y(new_n8762));
  nor_4  g08386(.A(new_n8762), .B(new_n8759_1), .Y(new_n8763));
  xnor_3 g08387(.A(new_n8763), .B(new_n8756), .Y(new_n8764));
  xnor_3 g08388(.A(new_n8764), .B(new_n8754), .Y(new_n8765));
  not_3  g08389(.A(new_n8765), .Y(new_n8766));
  nor_4  g08390(.A(new_n8678), .B(new_n8677), .Y(new_n8767));
  nand_4 g08391(.A(n8819), .B(n7436), .Y(new_n8768));
  xor_3  g08392(.A(new_n8768), .B(new_n8767), .Y(new_n8769));
  nand_4 g08393(.A(n11728), .B(n9241), .Y(new_n8770));
  nand_4 g08394(.A(n8276), .B(n6429), .Y(new_n8771));
  nand_4 g08395(.A(n12709), .B(n10510), .Y(new_n8772));
  not_3  g08396(.A(new_n8772), .Y(new_n8773));
  xor_3  g08397(.A(new_n8773), .B(new_n8771), .Y(new_n8774));
  xnor_3 g08398(.A(new_n8774), .B(new_n8770), .Y(new_n8775));
  xnor_3 g08399(.A(new_n8775), .B(new_n8769), .Y(new_n8776));
  not_3  g08400(.A(new_n8776), .Y(new_n8777));
  xor_3  g08401(.A(new_n8777), .B(new_n8766), .Y(new_n8778));
  nand_4 g08402(.A(new_n8694), .B(new_n8691), .Y(new_n8779));
  nor_4  g08403(.A(new_n8693), .B(new_n8692), .Y(new_n8780));
  nor_4  g08404(.A(new_n8714), .B(new_n8695), .Y(new_n8781));
  xnor_3 g08405(.A(new_n8781), .B(new_n8780), .Y(new_n8782));
  nand_4 g08406(.A(new_n8782), .B(new_n8779), .Y(new_n8783));
  xnor_3 g08407(.A(new_n8783), .B(new_n8778), .Y(new_n8784));
  xnor_3 g08408(.A(new_n8784), .B(new_n8750), .Y(new_n8785));
  xnor_3 g08409(.A(new_n8785), .B(new_n8748), .Y(new_n8786));
  nand_4 g08410(.A(n2393), .B(n1478), .Y(new_n8787));
  nand_4 g08411(.A(n5860), .B(n5760), .Y(new_n8788));
  nand_4 g08412(.A(n10990), .B(n3986), .Y(new_n8789));
  xnor_3 g08413(.A(new_n8789), .B(new_n8788), .Y(new_n8790));
  nor_4  g08414(.A(new_n8790), .B(new_n8787), .Y(new_n8791));
  not_3  g08415(.A(new_n8787), .Y(new_n8792));
  not_3  g08416(.A(new_n8790), .Y(new_n8793));
  nor_4  g08417(.A(new_n8793), .B(new_n8792), .Y(new_n8794));
  nor_4  g08418(.A(new_n8794), .B(new_n8791), .Y(new_n8795));
  nand_4 g08419(.A(n11892), .B(n1478), .Y(new_n8796));
  not_3  g08420(.A(new_n8796), .Y(new_n8797));
  nand_4 g08421(.A(n10990), .B(n5860), .Y(new_n8798));
  not_3  g08422(.A(new_n8798), .Y(new_n8799));
  nor_4  g08423(.A(new_n8799), .B(new_n8797), .Y(new_n8800));
  nor_4  g08424(.A(new_n8798), .B(new_n8796), .Y(new_n8801));
  nand_4 g08425(.A(n5760), .B(n2393), .Y(new_n8802));
  not_3  g08426(.A(new_n8802), .Y(new_n8803));
  nor_4  g08427(.A(new_n8803), .B(new_n8801), .Y(new_n8804));
  nor_4  g08428(.A(new_n8804), .B(new_n8800), .Y(new_n8805));
  xnor_3 g08429(.A(new_n8805), .B(new_n8795), .Y(new_n8806));
  not_3  g08430(.A(new_n8806), .Y(new_n8807));
  nand_4 g08431(.A(n12947), .B(n7388), .Y(new_n8808));
  nand_4 g08432(.A(n11892), .B(n11791), .Y(new_n8809));
  xor_3  g08433(.A(new_n8809), .B(new_n8808), .Y(new_n8810));
  xnor_3 g08434(.A(new_n8810), .B(new_n8807), .Y(new_n8811));
  nand_4 g08435(.A(n11791), .B(n7388), .Y(new_n8812));
  not_3  g08436(.A(new_n8812), .Y(new_n8813));
  nand_4 g08437(.A(n10990), .B(n2393), .Y(new_n8814));
  not_3  g08438(.A(new_n8814), .Y(new_n8815));
  nand_4 g08439(.A(n7388), .B(n1478), .Y(new_n8816));
  not_3  g08440(.A(new_n8816), .Y(new_n8817));
  nor_4  g08441(.A(new_n8817), .B(new_n8815), .Y(new_n8818));
  nor_4  g08442(.A(new_n8816), .B(new_n8814), .Y(new_n8819_1));
  nand_4 g08443(.A(n11892), .B(n5760), .Y(new_n8820));
  not_3  g08444(.A(new_n8820), .Y(new_n8821));
  nor_4  g08445(.A(new_n8821), .B(new_n8819_1), .Y(new_n8822));
  nor_4  g08446(.A(new_n8822), .B(new_n8818), .Y(new_n8823));
  and_4  g08447(.A(new_n8823), .B(new_n8813), .Y(new_n8824));
  xnor_3 g08448(.A(new_n8823), .B(new_n8813), .Y(new_n8825));
  nor_4  g08449(.A(new_n8801), .B(new_n8800), .Y(new_n8826));
  xnor_3 g08450(.A(new_n8826), .B(new_n8803), .Y(new_n8827));
  nor_4  g08451(.A(new_n8827), .B(new_n8825), .Y(new_n8828));
  nor_4  g08452(.A(new_n8828), .B(new_n8824), .Y(new_n8829));
  xnor_3 g08453(.A(new_n8829), .B(new_n8811), .Y(new_n8830));
  nand_4 g08454(.A(n12947), .B(n7965), .Y(new_n8831));
  not_3  g08455(.A(new_n8831), .Y(new_n8832));
  nand_4 g08456(.A(n11791), .B(n7965), .Y(new_n8833));
  not_3  g08457(.A(new_n8833), .Y(new_n8834));
  not_3  g08458(.A(new_n8528), .Y(new_n8835));
  nor_4  g08459(.A(new_n8535), .B(new_n8835), .Y(new_n8836));
  nor_4  g08460(.A(new_n8836), .B(new_n8534), .Y(new_n8837));
  nand_4 g08461(.A(new_n8837), .B(new_n8834), .Y(new_n8838));
  xnor_3 g08462(.A(new_n8837), .B(new_n8833), .Y(new_n8839));
  xnor_3 g08463(.A(new_n8816), .B(new_n8814), .Y(new_n8840));
  xnor_3 g08464(.A(new_n8840), .B(new_n8820), .Y(new_n8841));
  not_3  g08465(.A(new_n8841), .Y(new_n8842));
  nand_4 g08466(.A(new_n8842), .B(new_n8839), .Y(new_n8843));
  nand_4 g08467(.A(new_n8843), .B(new_n8838), .Y(new_n8844));
  nor_4  g08468(.A(new_n8844), .B(new_n8832), .Y(new_n8845));
  not_3  g08469(.A(new_n8845), .Y(new_n8846));
  xnor_3 g08470(.A(new_n8827), .B(new_n8825), .Y(new_n8847));
  not_3  g08471(.A(new_n8844), .Y(new_n8848));
  nor_4  g08472(.A(new_n8848), .B(new_n8831), .Y(new_n8849));
  nor_4  g08473(.A(new_n8849), .B(new_n8845), .Y(new_n8850));
  nand_4 g08474(.A(new_n8850), .B(new_n8847), .Y(new_n8851));
  nand_4 g08475(.A(new_n8851), .B(new_n8846), .Y(new_n8852));
  nor_4  g08476(.A(new_n8852), .B(new_n8830), .Y(new_n8853));
  nor_4  g08477(.A(new_n8789), .B(new_n8788), .Y(new_n8854));
  nand_4 g08478(.A(n11791), .B(n2393), .Y(new_n8855));
  not_3  g08479(.A(new_n8855), .Y(new_n8856));
  xor_3  g08480(.A(new_n8856), .B(new_n8854), .Y(new_n8857));
  not_3  g08481(.A(new_n8857), .Y(new_n8858));
  nand_4 g08482(.A(n5760), .B(n3986), .Y(new_n8859));
  nand_4 g08483(.A(n5860), .B(n1478), .Y(new_n8860));
  nand_4 g08484(.A(n10990), .B(n5857), .Y(new_n8861));
  nand_4 g08485(.A(new_n8861), .B(new_n8860), .Y(new_n8862));
  not_3  g08486(.A(new_n8860), .Y(new_n8863));
  not_3  g08487(.A(new_n8861), .Y(new_n8864));
  nand_4 g08488(.A(new_n8864), .B(new_n8863), .Y(new_n8865));
  nand_4 g08489(.A(new_n8865), .B(new_n8862), .Y(new_n8866));
  xor_3  g08490(.A(new_n8866), .B(new_n8859), .Y(new_n8867));
  xnor_3 g08491(.A(new_n8867), .B(new_n8858), .Y(new_n8868));
  nand_4 g08492(.A(new_n8805), .B(new_n8795), .Y(new_n8869));
  not_3  g08493(.A(new_n8869), .Y(new_n8870));
  nor_4  g08494(.A(new_n8870), .B(new_n8791), .Y(new_n8871));
  nand_4 g08495(.A(n7388), .B(n6441), .Y(new_n8872));
  nand_4 g08496(.A(n12947), .B(n11892), .Y(new_n8873));
  nand_4 g08497(.A(n11999), .B(n7965), .Y(new_n8874));
  xor_3  g08498(.A(new_n8874), .B(new_n8873), .Y(new_n8875));
  xnor_3 g08499(.A(new_n8875), .B(new_n8872), .Y(new_n8876));
  xnor_3 g08500(.A(new_n8876), .B(new_n8871), .Y(new_n8877));
  not_3  g08501(.A(new_n8877), .Y(new_n8878));
  nor_4  g08502(.A(new_n8878), .B(new_n8868), .Y(new_n8879));
  xnor_3 g08503(.A(new_n8867), .B(new_n8857), .Y(new_n8880));
  nor_4  g08504(.A(new_n8877), .B(new_n8880), .Y(new_n8881));
  nor_4  g08505(.A(new_n8881), .B(new_n8879), .Y(new_n8882));
  nand_4 g08506(.A(new_n8810), .B(new_n8807), .Y(new_n8883));
  nor_4  g08507(.A(new_n8809), .B(new_n8808), .Y(new_n8884));
  nor_4  g08508(.A(new_n8829), .B(new_n8811), .Y(new_n8885));
  xnor_3 g08509(.A(new_n8885), .B(new_n8884), .Y(new_n8886));
  nand_4 g08510(.A(new_n8886), .B(new_n8883), .Y(new_n8887));
  xnor_3 g08511(.A(new_n8887), .B(new_n8882), .Y(new_n8888));
  xnor_3 g08512(.A(new_n8888), .B(new_n8853), .Y(new_n8889));
  nand_4 g08513(.A(n7965), .B(n6441), .Y(new_n8890));
  not_3  g08514(.A(new_n8890), .Y(new_n8891));
  xnor_3 g08515(.A(new_n8852), .B(new_n8830), .Y(new_n8892));
  not_3  g08516(.A(new_n8892), .Y(new_n8893));
  nand_4 g08517(.A(new_n8893), .B(new_n8891), .Y(new_n8894));
  nand_4 g08518(.A(new_n8892), .B(new_n8890), .Y(new_n8895));
  xor_3  g08519(.A(new_n8841), .B(new_n8839), .Y(new_n8896));
  not_3  g08520(.A(new_n8896), .Y(new_n8897));
  nand_4 g08521(.A(new_n8537), .B(new_n8835), .Y(new_n8898));
  not_3  g08522(.A(new_n8898), .Y(new_n8899));
  nand_4 g08523(.A(new_n8899), .B(new_n8897), .Y(new_n8900));
  xnor_3 g08524(.A(new_n8850), .B(new_n8847), .Y(new_n8901));
  not_3  g08525(.A(new_n8901), .Y(new_n8902));
  nor_4  g08526(.A(new_n8902), .B(new_n8900), .Y(new_n8903));
  nand_4 g08527(.A(new_n8903), .B(new_n8895), .Y(new_n8904));
  nand_4 g08528(.A(new_n8904), .B(new_n8894), .Y(new_n8905));
  xnor_3 g08529(.A(new_n8905), .B(new_n8889), .Y(new_n8906));
  nand_4 g08530(.A(n12777), .B(n12648), .Y(new_n8907));
  nand_4 g08531(.A(n10545), .B(n7159), .Y(new_n8908));
  nand_4 g08532(.A(n12489), .B(n7690), .Y(new_n8909));
  xnor_3 g08533(.A(new_n8909), .B(new_n8908), .Y(new_n8910));
  nor_4  g08534(.A(new_n8910), .B(new_n8907), .Y(new_n8911));
  not_3  g08535(.A(new_n8907), .Y(new_n8912));
  not_3  g08536(.A(new_n8910), .Y(new_n8913));
  nor_4  g08537(.A(new_n8913), .B(new_n8912), .Y(new_n8914));
  nor_4  g08538(.A(new_n8914), .B(new_n8911), .Y(new_n8915));
  nand_4 g08539(.A(n12777), .B(n2530), .Y(new_n8916));
  not_3  g08540(.A(new_n8916), .Y(new_n8917));
  nand_4 g08541(.A(n12489), .B(n10545), .Y(new_n8918));
  not_3  g08542(.A(new_n8918), .Y(new_n8919));
  nor_4  g08543(.A(new_n8919), .B(new_n8917), .Y(new_n8920));
  nor_4  g08544(.A(new_n8918), .B(new_n8916), .Y(new_n8921));
  nand_4 g08545(.A(n12648), .B(n7159), .Y(new_n8922));
  not_3  g08546(.A(new_n8922), .Y(new_n8923));
  nor_4  g08547(.A(new_n8923), .B(new_n8921), .Y(new_n8924));
  nor_4  g08548(.A(new_n8924), .B(new_n8920), .Y(new_n8925));
  xnor_3 g08549(.A(new_n8925), .B(new_n8915), .Y(new_n8926));
  not_3  g08550(.A(new_n8926), .Y(new_n8927));
  nand_4 g08551(.A(n11967), .B(n8476), .Y(new_n8928));
  nand_4 g08552(.A(n6254), .B(n2530), .Y(new_n8929));
  xor_3  g08553(.A(new_n8929), .B(new_n8928), .Y(new_n8930));
  xnor_3 g08554(.A(new_n8930), .B(new_n8927), .Y(new_n8931));
  nand_4 g08555(.A(n8476), .B(n6254), .Y(new_n8932));
  not_3  g08556(.A(new_n8932), .Y(new_n8933));
  nand_4 g08557(.A(n12648), .B(n12489), .Y(new_n8934));
  not_3  g08558(.A(new_n8934), .Y(new_n8935));
  nand_4 g08559(.A(n12777), .B(n8476), .Y(new_n8936));
  not_3  g08560(.A(new_n8936), .Y(new_n8937));
  nor_4  g08561(.A(new_n8937), .B(new_n8935), .Y(new_n8938));
  nor_4  g08562(.A(new_n8936), .B(new_n8934), .Y(new_n8939));
  nand_4 g08563(.A(n7159), .B(n2530), .Y(new_n8940));
  not_3  g08564(.A(new_n8940), .Y(new_n8941));
  nor_4  g08565(.A(new_n8941), .B(new_n8939), .Y(new_n8942));
  nor_4  g08566(.A(new_n8942), .B(new_n8938), .Y(new_n8943));
  and_4  g08567(.A(new_n8943), .B(new_n8933), .Y(new_n8944));
  xnor_3 g08568(.A(new_n8943), .B(new_n8933), .Y(new_n8945));
  nor_4  g08569(.A(new_n8921), .B(new_n8920), .Y(new_n8946));
  xnor_3 g08570(.A(new_n8946), .B(new_n8923), .Y(new_n8947));
  nor_4  g08571(.A(new_n8947), .B(new_n8945), .Y(new_n8948));
  nor_4  g08572(.A(new_n8948), .B(new_n8944), .Y(new_n8949));
  xnor_3 g08573(.A(new_n8949), .B(new_n8931), .Y(new_n8950));
  nand_4 g08574(.A(n11967), .B(n5331), .Y(new_n8951));
  not_3  g08575(.A(new_n8951), .Y(new_n8952));
  xnor_3 g08576(.A(new_n8947), .B(new_n8945), .Y(new_n8953));
  not_3  g08577(.A(new_n8953), .Y(new_n8954));
  nor_4  g08578(.A(new_n8954), .B(new_n8952), .Y(new_n8955));
  not_3  g08579(.A(new_n8955), .Y(new_n8956));
  nor_4  g08580(.A(new_n8953), .B(new_n8951), .Y(new_n8957));
  nor_4  g08581(.A(new_n8957), .B(new_n8955), .Y(new_n8958));
  nand_4 g08582(.A(n6254), .B(n5331), .Y(new_n8959));
  not_3  g08583(.A(new_n8959), .Y(new_n8960));
  not_3  g08584(.A(new_n8514), .Y(new_n8961));
  nor_4  g08585(.A(new_n8521), .B(new_n8961), .Y(new_n8962));
  nor_4  g08586(.A(new_n8962), .B(new_n8520), .Y(new_n8963));
  nand_4 g08587(.A(new_n8963), .B(new_n8960), .Y(new_n8964));
  not_3  g08588(.A(new_n8964), .Y(new_n8965));
  xnor_3 g08589(.A(new_n8963), .B(new_n8960), .Y(new_n8966));
  nor_4  g08590(.A(new_n8939), .B(new_n8938), .Y(new_n8967));
  xnor_3 g08591(.A(new_n8967), .B(new_n8941), .Y(new_n8968));
  nor_4  g08592(.A(new_n8968), .B(new_n8966), .Y(new_n8969));
  nor_4  g08593(.A(new_n8969), .B(new_n8965), .Y(new_n8970));
  nand_4 g08594(.A(new_n8970), .B(new_n8958), .Y(new_n8971));
  nand_4 g08595(.A(new_n8971), .B(new_n8956), .Y(new_n8972));
  nor_4  g08596(.A(new_n8972), .B(new_n8950), .Y(new_n8973));
  not_3  g08597(.A(new_n8973), .Y(new_n8974));
  nand_4 g08598(.A(n5331), .B(n1353), .Y(new_n8975));
  nand_4 g08599(.A(n11967), .B(n2530), .Y(new_n8976));
  nand_4 g08600(.A(n8476), .B(n447), .Y(new_n8977));
  not_3  g08601(.A(new_n8977), .Y(new_n8978));
  xor_3  g08602(.A(new_n8978), .B(new_n8976), .Y(new_n8979));
  xnor_3 g08603(.A(new_n8979), .B(new_n8975), .Y(new_n8980));
  nand_4 g08604(.A(new_n8925), .B(new_n8915), .Y(new_n8981));
  not_3  g08605(.A(new_n8981), .Y(new_n8982));
  nor_4  g08606(.A(new_n8982), .B(new_n8911), .Y(new_n8983));
  not_3  g08607(.A(new_n8983), .Y(new_n8984));
  xnor_3 g08608(.A(new_n8984), .B(new_n8980), .Y(new_n8985));
  nor_4  g08609(.A(new_n8909), .B(new_n8908), .Y(new_n8986));
  nand_4 g08610(.A(n12648), .B(n6254), .Y(new_n8987));
  not_3  g08611(.A(new_n8987), .Y(new_n8988));
  xor_3  g08612(.A(new_n8988), .B(new_n8986), .Y(new_n8989));
  not_3  g08613(.A(new_n8989), .Y(new_n8990));
  nand_4 g08614(.A(n7690), .B(n7159), .Y(new_n8991));
  not_3  g08615(.A(new_n8991), .Y(new_n8992));
  nand_4 g08616(.A(n12777), .B(n10545), .Y(new_n8993));
  nand_4 g08617(.A(n12489), .B(n3616), .Y(new_n8994));
  not_3  g08618(.A(new_n8994), .Y(new_n8995));
  xor_3  g08619(.A(new_n8995), .B(new_n8993), .Y(new_n8996));
  xnor_3 g08620(.A(new_n8996), .B(new_n8992), .Y(new_n8997));
  xnor_3 g08621(.A(new_n8997), .B(new_n8990), .Y(new_n8998));
  xnor_3 g08622(.A(new_n8998), .B(new_n8985), .Y(new_n8999));
  nand_4 g08623(.A(new_n8930), .B(new_n8927), .Y(new_n9000));
  nor_4  g08624(.A(new_n8929), .B(new_n8928), .Y(new_n9001));
  nor_4  g08625(.A(new_n8949), .B(new_n8931), .Y(new_n9002));
  xnor_3 g08626(.A(new_n9002), .B(new_n9001), .Y(new_n9003));
  nand_4 g08627(.A(new_n9003), .B(new_n9000), .Y(new_n9004));
  xnor_3 g08628(.A(new_n9004), .B(new_n8999), .Y(new_n9005));
  xnor_3 g08629(.A(new_n9005), .B(new_n8974), .Y(new_n9006));
  nand_4 g08630(.A(n5331), .B(n447), .Y(new_n9007));
  not_3  g08631(.A(new_n9007), .Y(new_n9008));
  xnor_3 g08632(.A(new_n8972), .B(new_n8950), .Y(new_n9009));
  not_3  g08633(.A(new_n9009), .Y(new_n9010));
  nand_4 g08634(.A(new_n9010), .B(new_n9008), .Y(new_n9011));
  nand_4 g08635(.A(new_n9009), .B(new_n9007), .Y(new_n9012));
  not_3  g08636(.A(new_n8966), .Y(new_n9013));
  xor_3  g08637(.A(new_n8968), .B(new_n9013), .Y(new_n9014));
  nand_4 g08638(.A(new_n8523), .B(new_n8961), .Y(new_n9015));
  nor_4  g08639(.A(new_n9015), .B(new_n9014), .Y(new_n9016));
  xnor_3 g08640(.A(new_n8970), .B(new_n8958), .Y(new_n9017));
  nand_4 g08641(.A(new_n9017), .B(new_n9016), .Y(new_n9018));
  not_3  g08642(.A(new_n9018), .Y(new_n9019));
  nand_4 g08643(.A(new_n9019), .B(new_n9012), .Y(new_n9020));
  nand_4 g08644(.A(new_n9020), .B(new_n9011), .Y(new_n9021));
  xnor_3 g08645(.A(new_n9021), .B(new_n9006), .Y(new_n9022));
  xnor_3 g08646(.A(new_n9022), .B(new_n8906), .Y(new_n9023));
  nand_4 g08647(.A(new_n8895), .B(new_n8894), .Y(new_n9024));
  xnor_3 g08648(.A(new_n9024), .B(new_n8903), .Y(new_n9025));
  not_3  g08649(.A(new_n9025), .Y(new_n9026));
  nand_4 g08650(.A(new_n9012), .B(new_n9011), .Y(new_n9027));
  xnor_3 g08651(.A(new_n9027), .B(new_n9019), .Y(new_n9028));
  not_3  g08652(.A(new_n9028), .Y(new_n9029));
  nand_4 g08653(.A(new_n9029), .B(new_n9026), .Y(new_n9030));
  nand_4 g08654(.A(new_n9028), .B(new_n9025), .Y(new_n9031));
  xnor_3 g08655(.A(new_n9017), .B(new_n9016), .Y(new_n9032));
  xnor_3 g08656(.A(new_n8902), .B(new_n8900), .Y(new_n9033));
  nand_4 g08657(.A(new_n9033), .B(new_n9032), .Y(new_n9034));
  xnor_3 g08658(.A(new_n9033), .B(new_n9032), .Y(new_n9035));
  not_3  g08659(.A(new_n9035), .Y(new_n9036));
  xnor_3 g08660(.A(new_n9015), .B(new_n9014), .Y(new_n9037));
  xor_3  g08661(.A(new_n8898), .B(new_n8897), .Y(new_n9038));
  nor_4  g08662(.A(new_n9038), .B(new_n9037), .Y(new_n9039));
  nor_4  g08663(.A(new_n8541), .B(new_n8527), .Y(new_n9040));
  nor_4  g08664(.A(new_n8546), .B(new_n9040), .Y(new_n9041));
  xnor_3 g08665(.A(new_n9038), .B(new_n9037), .Y(new_n9042));
  nor_4  g08666(.A(new_n9042), .B(new_n9041), .Y(new_n9043));
  nor_4  g08667(.A(new_n9043), .B(new_n9039), .Y(new_n9044));
  nand_4 g08668(.A(new_n9044), .B(new_n9036), .Y(new_n9045));
  nand_4 g08669(.A(new_n9045), .B(new_n9034), .Y(new_n9046));
  nand_4 g08670(.A(new_n9046), .B(new_n9031), .Y(new_n9047));
  nand_4 g08671(.A(new_n9047), .B(new_n9030), .Y(new_n9048));
  xnor_3 g08672(.A(new_n9048), .B(new_n9023), .Y(new_n9049));
  xnor_3 g08673(.A(new_n9049), .B(new_n8786), .Y(new_n9050));
  not_3  g08674(.A(new_n8747), .Y(new_n9051));
  nor_4  g08675(.A(new_n8746), .B(new_n8745), .Y(new_n9052));
  nor_4  g08676(.A(new_n9052), .B(new_n9051), .Y(new_n9053));
  not_3  g08677(.A(new_n9034), .Y(new_n9054));
  not_3  g08678(.A(new_n9014), .Y(new_n9055));
  not_3  g08679(.A(new_n9015), .Y(new_n9056));
  nor_4  g08680(.A(new_n9056), .B(new_n9055), .Y(new_n9057));
  nor_4  g08681(.A(new_n9057), .B(new_n9016), .Y(new_n9058));
  xor_3  g08682(.A(new_n8899), .B(new_n8897), .Y(new_n9059));
  nand_4 g08683(.A(new_n9059), .B(new_n9058), .Y(new_n9060));
  not_3  g08684(.A(new_n9041), .Y(new_n9061));
  nor_4  g08685(.A(new_n9059), .B(new_n9058), .Y(new_n9062));
  nor_4  g08686(.A(new_n9062), .B(new_n9039), .Y(new_n9063));
  nand_4 g08687(.A(new_n9063), .B(new_n9061), .Y(new_n9064));
  nand_4 g08688(.A(new_n9064), .B(new_n9060), .Y(new_n9065));
  nor_4  g08689(.A(new_n9065), .B(new_n9035), .Y(new_n9066));
  nor_4  g08690(.A(new_n9066), .B(new_n9054), .Y(new_n9067));
  nand_4 g08691(.A(new_n9031), .B(new_n9030), .Y(new_n9068));
  xnor_3 g08692(.A(new_n9068), .B(new_n9067), .Y(new_n9069));
  nand_4 g08693(.A(new_n9069), .B(new_n9053), .Y(new_n9070));
  not_3  g08694(.A(new_n9053), .Y(new_n9071));
  xnor_3 g08695(.A(new_n9068), .B(new_n9046), .Y(new_n9072));
  nand_4 g08696(.A(new_n9072), .B(new_n9071), .Y(new_n9073));
  xnor_3 g08697(.A(new_n8743), .B(new_n8742), .Y(new_n9074));
  not_3  g08698(.A(new_n9074), .Y(new_n9075));
  xnor_3 g08699(.A(new_n9065), .B(new_n9035), .Y(new_n9076));
  nand_4 g08700(.A(new_n9076), .B(new_n9075), .Y(new_n9077));
  nor_4  g08701(.A(new_n8740), .B(new_n8737), .Y(new_n9078));
  nor_4  g08702(.A(new_n9078), .B(new_n8742), .Y(new_n9079));
  xnor_3 g08703(.A(new_n9042), .B(new_n9061), .Y(new_n9080_1));
  nand_4 g08704(.A(new_n9080_1), .B(new_n9079), .Y(new_n9081));
  not_3  g08705(.A(new_n9079), .Y(new_n9082));
  xnor_3 g08706(.A(new_n9042), .B(new_n9041), .Y(new_n9083));
  nor_4  g08707(.A(new_n9083), .B(new_n9082), .Y(new_n9084));
  nor_4  g08708(.A(new_n9080_1), .B(new_n9079), .Y(new_n9085));
  nor_4  g08709(.A(new_n9085), .B(new_n9084), .Y(new_n9086));
  not_3  g08710(.A(new_n8511), .Y(new_n9087));
  nor_4  g08711(.A(new_n9087), .B(new_n8497), .Y(new_n9088));
  not_3  g08712(.A(new_n9088), .Y(new_n9089));
  nand_4 g08713(.A(new_n8549), .B(new_n9089), .Y(new_n9090));
  nand_4 g08714(.A(new_n9090), .B(new_n9086), .Y(new_n9091));
  nand_4 g08715(.A(new_n9091), .B(new_n9081), .Y(new_n9092));
  xnor_3 g08716(.A(new_n9076), .B(new_n9074), .Y(new_n9093));
  nand_4 g08717(.A(new_n9093), .B(new_n9092), .Y(new_n9094));
  nand_4 g08718(.A(new_n9094), .B(new_n9077), .Y(new_n9095));
  nand_4 g08719(.A(new_n9095), .B(new_n9073), .Y(new_n9096));
  nand_4 g08720(.A(new_n9096), .B(new_n9070), .Y(new_n9097));
  xnor_3 g08721(.A(new_n9097), .B(new_n9050), .Y(new_n9098));
  nand_4 g08722(.A(new_n9098), .B(new_n8672), .Y(new_n9099));
  xnor_3 g08723(.A(new_n9098), .B(new_n8671), .Y(new_n9100));
  xnor_3 g08724(.A(new_n8668), .B(new_n8664), .Y(new_n9101));
  not_3  g08725(.A(new_n9077), .Y(new_n9102));
  xnor_3 g08726(.A(new_n9083), .B(new_n9082), .Y(new_n9103));
  not_3  g08727(.A(new_n9090), .Y(new_n9104));
  nor_4  g08728(.A(new_n9104), .B(new_n9103), .Y(new_n9105));
  nor_4  g08729(.A(new_n9105), .B(new_n9084), .Y(new_n9106));
  xnor_3 g08730(.A(new_n9076), .B(new_n9075), .Y(new_n9107));
  nor_4  g08731(.A(new_n9107), .B(new_n9106), .Y(new_n9108));
  nor_4  g08732(.A(new_n9108), .B(new_n9102), .Y(new_n9109));
  nand_4 g08733(.A(new_n9073), .B(new_n9070), .Y(new_n9110));
  xnor_3 g08734(.A(new_n9110), .B(new_n9109), .Y(new_n9111_1));
  nand_4 g08735(.A(new_n9111_1), .B(new_n9101), .Y(new_n9112));
  not_3  g08736(.A(new_n9112), .Y(new_n9113));
  not_3  g08737(.A(new_n9101), .Y(new_n9114));
  xnor_3 g08738(.A(new_n9110), .B(new_n9095), .Y(new_n9115));
  nand_4 g08739(.A(new_n9115), .B(new_n9114), .Y(new_n9116));
  nand_4 g08740(.A(new_n9116), .B(new_n9112), .Y(new_n9117));
  not_3  g08741(.A(new_n8660), .Y(new_n9118));
  not_3  g08742(.A(new_n8663), .Y(new_n9119));
  nor_4  g08743(.A(new_n9119), .B(new_n9118), .Y(new_n9120));
  nor_4  g08744(.A(new_n9120), .B(new_n8664), .Y(new_n9121));
  not_3  g08745(.A(new_n9121), .Y(new_n9122));
  xnor_3 g08746(.A(new_n9107), .B(new_n9106), .Y(new_n9123));
  nand_4 g08747(.A(new_n9123), .B(new_n9122), .Y(new_n9124));
  not_3  g08748(.A(new_n9124), .Y(new_n9125));
  nor_4  g08749(.A(new_n9093), .B(new_n9092), .Y(new_n9126));
  nor_4  g08750(.A(new_n9126), .B(new_n9108), .Y(new_n9127));
  nand_4 g08751(.A(new_n9127), .B(new_n9121), .Y(new_n9128));
  nand_4 g08752(.A(new_n9128), .B(new_n9124), .Y(new_n9129));
  nor_4  g08753(.A(new_n8659), .B(new_n8658), .Y(new_n9130));
  nor_4  g08754(.A(new_n9130), .B(new_n9118), .Y(new_n9131));
  xnor_3 g08755(.A(new_n9090), .B(new_n9103), .Y(new_n9132));
  nor_4  g08756(.A(new_n9132), .B(new_n9131), .Y(new_n9133));
  not_3  g08757(.A(new_n8492), .Y(new_n9134));
  nand_4 g08758(.A(new_n8552), .B(new_n8495), .Y(new_n9135));
  nand_4 g08759(.A(new_n9135), .B(new_n9134), .Y(new_n9136));
  xnor_3 g08760(.A(new_n9132), .B(new_n9131), .Y(new_n9137_1));
  nor_4  g08761(.A(new_n9137_1), .B(new_n9136), .Y(new_n9138));
  nor_4  g08762(.A(new_n9138), .B(new_n9133), .Y(new_n9139));
  nor_4  g08763(.A(new_n9139), .B(new_n9129), .Y(new_n9140));
  nor_4  g08764(.A(new_n9140), .B(new_n9125), .Y(new_n9141));
  nor_4  g08765(.A(new_n9141), .B(new_n9117), .Y(new_n9142));
  nor_4  g08766(.A(new_n9142), .B(new_n9113), .Y(new_n9143));
  nand_4 g08767(.A(new_n9143), .B(new_n9100), .Y(new_n9144));
  nand_4 g08768(.A(new_n9144), .B(new_n9099), .Y(new_n9145));
  nor_4  g08769(.A(new_n9049), .B(new_n8786), .Y(new_n9146));
  nor_4  g08770(.A(new_n9097), .B(new_n9050), .Y(new_n9147));
  nor_4  g08771(.A(new_n9147), .B(new_n9146), .Y(new_n9148));
  not_3  g08772(.A(new_n8906), .Y(new_n9149));
  nand_4 g08773(.A(new_n9022), .B(new_n9149), .Y(new_n9150));
  nand_4 g08774(.A(new_n9048), .B(new_n9023), .Y(new_n9151));
  nand_4 g08775(.A(new_n9151), .B(new_n9150), .Y(new_n9152));
  nand_4 g08776(.A(new_n8888), .B(new_n8853), .Y(new_n9153));
  not_3  g08777(.A(new_n8889), .Y(new_n9154));
  nand_4 g08778(.A(new_n8905), .B(new_n9154), .Y(new_n9155));
  nand_4 g08779(.A(new_n9155), .B(new_n9153), .Y(new_n9156));
  nand_4 g08780(.A(new_n8885), .B(new_n8884), .Y(new_n9157));
  not_3  g08781(.A(new_n8882), .Y(new_n9158));
  nand_4 g08782(.A(new_n8887), .B(new_n9158), .Y(new_n9159));
  nand_4 g08783(.A(new_n9159), .B(new_n9157), .Y(new_n9160));
  not_3  g08784(.A(new_n8767), .Y(new_n9161));
  nor_4  g08785(.A(new_n8768), .B(new_n9161), .Y(new_n9162));
  nor_4  g08786(.A(new_n8775), .B(new_n8769), .Y(new_n9163));
  nor_4  g08787(.A(new_n9163), .B(new_n9162), .Y(new_n9164));
  nand_4 g08788(.A(n9241), .B(n6429), .Y(new_n9165));
  nand_4 g08789(.A(n12299), .B(n8717), .Y(new_n9166));
  xor_3  g08790(.A(new_n9166), .B(new_n9165), .Y(new_n9167));
  nand_4 g08791(.A(n7730), .B(n6776), .Y(new_n9168));
  nand_4 g08792(.A(n8819), .B(n8276), .Y(new_n9169));
  xor_3  g08793(.A(new_n9169), .B(new_n9168), .Y(new_n9170));
  xor_3  g08794(.A(new_n9170), .B(new_n9167), .Y(new_n9171));
  not_3  g08795(.A(new_n8771), .Y(new_n9172));
  nor_4  g08796(.A(new_n8773), .B(new_n9172), .Y(new_n9173));
  not_3  g08797(.A(new_n8770), .Y(new_n9174));
  nor_4  g08798(.A(new_n8774), .B(new_n9174), .Y(new_n9175));
  nor_4  g08799(.A(new_n9175), .B(new_n9173), .Y(new_n9176));
  nand_4 g08800(.A(n7436), .B(n2433), .Y(new_n9177));
  xnor_3 g08801(.A(new_n9177), .B(new_n9176), .Y(new_n9178));
  xnor_3 g08802(.A(new_n9178), .B(new_n9171), .Y(new_n9179));
  xnor_3 g08803(.A(new_n9179), .B(new_n9164), .Y(new_n9180));
  or_4   g08804(.A(new_n8762), .B(new_n8755), .Y(new_n9181));
  not_3  g08805(.A(new_n9181), .Y(new_n9182));
  nor_4  g08806(.A(new_n9182), .B(new_n8759_1), .Y(new_n9183));
  nand_4 g08807(.A(n12777), .B(n7690), .Y(new_n9184));
  nand_4 g08808(.A(n7159), .B(n3616), .Y(new_n9185));
  xor_3  g08809(.A(new_n9185), .B(new_n9184), .Y(new_n9186));
  nand_4 g08810(.A(n11999), .B(n7388), .Y(new_n9187));
  nand_4 g08811(.A(n11892), .B(n6441), .Y(new_n9188));
  xor_3  g08812(.A(new_n9188), .B(new_n9187), .Y(new_n9189_1));
  xnor_3 g08813(.A(new_n9189_1), .B(new_n9186), .Y(new_n9190));
  nand_4 g08814(.A(n10022), .B(n7965), .Y(new_n9191));
  nand_4 g08815(.A(n10990), .B(n45), .Y(new_n9192));
  xor_3  g08816(.A(new_n9192), .B(new_n9191), .Y(new_n9193));
  nand_4 g08817(.A(n3986), .B(n1478), .Y(new_n9194));
  nand_4 g08818(.A(n5857), .B(n5760), .Y(new_n9195_1));
  xor_3  g08819(.A(new_n9195_1), .B(new_n9194), .Y(new_n9196));
  xnor_3 g08820(.A(new_n9196), .B(new_n9193), .Y(new_n9197));
  xnor_3 g08821(.A(new_n9197), .B(new_n9190), .Y(new_n9198));
  not_3  g08822(.A(new_n8993), .Y(new_n9199));
  nor_4  g08823(.A(new_n8995), .B(new_n9199), .Y(new_n9200));
  nor_4  g08824(.A(new_n8996), .B(new_n8992), .Y(new_n9201));
  nor_4  g08825(.A(new_n9201), .B(new_n9200), .Y(new_n9202));
  nand_4 g08826(.A(n8476), .B(n1353), .Y(new_n9203));
  not_3  g08827(.A(new_n9203), .Y(new_n9204));
  xnor_3 g08828(.A(new_n9204), .B(new_n9202), .Y(new_n9205));
  xnor_3 g08829(.A(new_n9205), .B(new_n9198), .Y(new_n9206));
  xnor_3 g08830(.A(new_n9206), .B(new_n9183), .Y(new_n9207));
  xnor_3 g08831(.A(new_n9207), .B(new_n9180), .Y(new_n9208));
  xnor_3 g08832(.A(new_n9208), .B(new_n9160), .Y(new_n9209));
  xnor_3 g08833(.A(new_n9209), .B(new_n9156), .Y(new_n9210));
  xnor_3 g08834(.A(new_n9210), .B(new_n9152), .Y(new_n9211));
  xnor_3 g08835(.A(new_n9211), .B(new_n9148), .Y(new_n9212));
  nand_4 g08836(.A(new_n8784), .B(new_n8750), .Y(new_n9213));
  not_3  g08837(.A(new_n8785), .Y(new_n9214));
  nand_4 g08838(.A(new_n9214), .B(new_n8748), .Y(new_n9215));
  nand_4 g08839(.A(new_n9215), .B(new_n9213), .Y(new_n9216));
  nand_4 g08840(.A(n2530), .B(n447), .Y(new_n9217));
  xnor_3 g08841(.A(new_n9217), .B(new_n9216), .Y(new_n9218));
  nand_4 g08842(.A(new_n8781), .B(new_n8780), .Y(new_n9219));
  not_3  g08843(.A(new_n8778), .Y(new_n9220));
  nand_4 g08844(.A(new_n8783), .B(new_n9220), .Y(new_n9221));
  nand_4 g08845(.A(new_n9221), .B(new_n9219), .Y(new_n9222));
  nand_4 g08846(.A(n12648), .B(n11967), .Y(new_n9223));
  nand_4 g08847(.A(n11791), .B(n5860), .Y(new_n9224));
  xor_3  g08848(.A(new_n9224), .B(new_n9223), .Y(new_n9225));
  nand_4 g08849(.A(n5331), .B(n4436), .Y(new_n9226));
  nand_4 g08850(.A(n12489), .B(n4499), .Y(new_n9227));
  xor_3  g08851(.A(new_n9227), .B(new_n9226), .Y(new_n9228));
  xor_3  g08852(.A(new_n9228), .B(new_n9225), .Y(new_n9229));
  not_3  g08853(.A(new_n8859), .Y(new_n9230));
  nand_4 g08854(.A(new_n8862), .B(new_n9230), .Y(new_n9231));
  nand_4 g08855(.A(new_n9231), .B(new_n8865), .Y(new_n9232));
  nor_4  g08856(.A(new_n8874), .B(new_n8873), .Y(new_n9233));
  not_3  g08857(.A(new_n8872), .Y(new_n9234));
  nand_4 g08858(.A(new_n8874), .B(new_n8873), .Y(new_n9235));
  nand_4 g08859(.A(new_n9235), .B(new_n9234), .Y(new_n9236));
  not_3  g08860(.A(new_n9236), .Y(new_n9237));
  nor_4  g08861(.A(new_n9237), .B(new_n9233), .Y(new_n9238));
  xor_3  g08862(.A(new_n9238), .B(new_n9232), .Y(new_n9239));
  xnor_3 g08863(.A(new_n9239), .B(new_n9229), .Y(new_n9240));
  xnor_3 g08864(.A(new_n9240), .B(new_n9222), .Y(new_n9241_1));
  not_3  g08865(.A(new_n8647), .Y(new_n9242));
  nor_4  g08866(.A(new_n8648), .B(new_n9242), .Y(new_n9243));
  nor_4  g08867(.A(new_n8650), .B(new_n8645), .Y(new_n9244));
  nor_4  g08868(.A(new_n9244), .B(new_n9243), .Y(new_n9245));
  nand_4 g08869(.A(n11257), .B(n5212), .Y(new_n9246));
  not_3  g08870(.A(new_n8754), .Y(new_n9247));
  nand_4 g08871(.A(new_n8764), .B(new_n9247), .Y(new_n9248));
  nand_4 g08872(.A(new_n8776), .B(new_n8765), .Y(new_n9249));
  nand_4 g08873(.A(new_n9249), .B(new_n9248), .Y(new_n9250));
  nand_4 g08874(.A(n12709), .B(n10644), .Y(new_n9251));
  not_3  g08875(.A(new_n9251), .Y(new_n9252));
  xnor_3 g08876(.A(new_n9252), .B(new_n9250), .Y(new_n9253));
  nand_4 g08877(.A(n11728), .B(n10510), .Y(new_n9254));
  not_3  g08878(.A(new_n8626), .Y(new_n9255));
  nand_4 g08879(.A(new_n8632), .B(new_n9255), .Y(new_n9256));
  nand_4 g08880(.A(new_n8644), .B(new_n8633), .Y(new_n9257));
  nand_4 g08881(.A(new_n9257), .B(new_n9256), .Y(new_n9258));
  xnor_3 g08882(.A(new_n9258), .B(new_n9254), .Y(new_n9259));
  xnor_3 g08883(.A(new_n9259), .B(new_n9253), .Y(new_n9260));
  xnor_3 g08884(.A(new_n9260), .B(new_n9246), .Y(new_n9261));
  xnor_3 g08885(.A(new_n9261), .B(new_n9245), .Y(new_n9262));
  xnor_3 g08886(.A(new_n9262), .B(new_n9241_1), .Y(new_n9263));
  nand_4 g08887(.A(new_n9005), .B(new_n8973), .Y(new_n9264));
  nand_4 g08888(.A(new_n9021), .B(new_n9006), .Y(new_n9265));
  nand_4 g08889(.A(new_n9265), .B(new_n9264), .Y(new_n9266));
  nand_4 g08890(.A(n12947), .B(n2393), .Y(new_n9267));
  not_3  g08891(.A(new_n9267), .Y(new_n9268));
  nand_4 g08892(.A(new_n8856), .B(new_n8854), .Y(new_n9269));
  nand_4 g08893(.A(new_n8867), .B(new_n8857), .Y(new_n9270));
  nand_4 g08894(.A(new_n9270), .B(new_n9269), .Y(new_n9271));
  xor_3  g08895(.A(new_n9271), .B(new_n9268), .Y(new_n9272));
  nand_4 g08896(.A(new_n8983), .B(new_n8980), .Y(new_n9273));
  not_3  g08897(.A(new_n8998), .Y(new_n9274));
  nand_4 g08898(.A(new_n9274), .B(new_n8985), .Y(new_n9275));
  nand_4 g08899(.A(new_n9275), .B(new_n9273), .Y(new_n9276));
  nand_4 g08900(.A(n10545), .B(n6254), .Y(new_n9277));
  nand_4 g08901(.A(new_n8988), .B(new_n8986), .Y(new_n9278));
  nand_4 g08902(.A(new_n8997), .B(new_n8989), .Y(new_n9279));
  nand_4 g08903(.A(new_n9279), .B(new_n9278), .Y(new_n9280));
  nand_4 g08904(.A(n8759), .B(n1198), .Y(new_n9281));
  not_3  g08905(.A(new_n9281), .Y(new_n9282));
  xnor_3 g08906(.A(new_n9282), .B(new_n9280), .Y(new_n9283));
  xnor_3 g08907(.A(new_n9283), .B(new_n9277), .Y(new_n9284));
  xnor_3 g08908(.A(new_n9284), .B(new_n9276), .Y(new_n9285));
  nand_4 g08909(.A(n12705), .B(n4370), .Y(new_n9286));
  not_3  g08910(.A(new_n9286), .Y(new_n9287));
  nand_4 g08911(.A(n9725), .B(n5964), .Y(new_n9288));
  nand_4 g08912(.A(n12000), .B(n1097), .Y(new_n9289));
  xor_3  g08913(.A(new_n9289), .B(new_n9288), .Y(new_n9290));
  nand_4 g08914(.A(n5320), .B(n4312), .Y(new_n9291));
  nand_4 g08915(.A(n12025), .B(n11877), .Y(new_n9292));
  xor_3  g08916(.A(new_n9292), .B(new_n9291), .Y(new_n9293));
  xnor_3 g08917(.A(new_n9293), .B(new_n9290), .Y(new_n9294));
  xnor_3 g08918(.A(new_n9294), .B(new_n9287), .Y(new_n9295));
  not_3  g08919(.A(new_n8628), .Y(new_n9296));
  nor_4  g08920(.A(new_n8630), .B(new_n9296), .Y(new_n9297));
  not_3  g08921(.A(new_n8627), .Y(new_n9298));
  nor_4  g08922(.A(new_n8631), .B(new_n9298), .Y(new_n9299));
  nor_4  g08923(.A(new_n9299), .B(new_n9297), .Y(new_n9300));
  not_3  g08924(.A(new_n8639), .Y(new_n9301));
  nor_4  g08925(.A(new_n8641), .B(new_n9301), .Y(new_n9302));
  not_3  g08926(.A(new_n8638), .Y(new_n9303));
  nor_4  g08927(.A(new_n8642), .B(new_n9303), .Y(new_n9304));
  nor_4  g08928(.A(new_n9304), .B(new_n9302), .Y(new_n9305));
  xnor_3 g08929(.A(new_n9305), .B(new_n9300), .Y(new_n9306));
  xnor_3 g08930(.A(new_n9306), .B(new_n9295), .Y(new_n9307));
  not_3  g08931(.A(new_n8976), .Y(new_n9308));
  nor_4  g08932(.A(new_n8978), .B(new_n9308), .Y(new_n9309));
  not_3  g08933(.A(new_n8975), .Y(new_n9310));
  nor_4  g08934(.A(new_n8979), .B(new_n9310), .Y(new_n9311));
  nor_4  g08935(.A(new_n9311), .B(new_n9309), .Y(new_n9312));
  nand_4 g08936(.A(n11407), .B(n10547), .Y(new_n9313));
  nand_4 g08937(.A(n6604), .B(n5305), .Y(new_n9314));
  not_3  g08938(.A(new_n9314), .Y(new_n9315));
  xor_3  g08939(.A(new_n9315), .B(new_n9313), .Y(new_n9316));
  xnor_3 g08940(.A(new_n9316), .B(new_n9312), .Y(new_n9317));
  not_3  g08941(.A(new_n8636), .Y(new_n9318));
  or_4   g08942(.A(new_n9318), .B(new_n8635), .Y(new_n9319));
  not_3  g08943(.A(new_n8637), .Y(new_n9320));
  nand_4 g08944(.A(new_n8643), .B(new_n9320), .Y(new_n9321));
  nand_4 g08945(.A(new_n9321), .B(new_n9319), .Y(new_n9322));
  xnor_3 g08946(.A(new_n9322), .B(new_n9317), .Y(new_n9323));
  xnor_3 g08947(.A(new_n9323), .B(new_n9307), .Y(new_n9324));
  xnor_3 g08948(.A(new_n9324), .B(new_n9285), .Y(new_n9325));
  xnor_3 g08949(.A(new_n9325), .B(new_n9272), .Y(new_n9326));
  xnor_3 g08950(.A(new_n9326), .B(new_n9266), .Y(new_n9327));
  xnor_3 g08951(.A(new_n9327), .B(new_n9263), .Y(new_n9328));
  nand_4 g08952(.A(new_n8652), .B(new_n8621), .Y(new_n9329));
  nand_4 g08953(.A(new_n8670), .B(new_n8653), .Y(new_n9330));
  nand_4 g08954(.A(new_n9330), .B(new_n9329), .Y(new_n9331));
  nand_4 g08955(.A(new_n9002), .B(new_n9001), .Y(new_n9332));
  not_3  g08956(.A(new_n8999), .Y(new_n9333));
  nand_4 g08957(.A(new_n9004), .B(new_n9333), .Y(new_n9334));
  nand_4 g08958(.A(new_n9334), .B(new_n9332), .Y(new_n9335));
  not_3  g08959(.A(new_n8871), .Y(new_n9336));
  nor_4  g08960(.A(new_n8876), .B(new_n9336), .Y(new_n9337));
  nor_4  g08961(.A(new_n8879), .B(new_n9337), .Y(new_n9338));
  xnor_3 g08962(.A(new_n9338), .B(new_n9335), .Y(new_n9339));
  xnor_3 g08963(.A(new_n9339), .B(new_n9331), .Y(new_n9340));
  xnor_3 g08964(.A(new_n9340), .B(new_n9328), .Y(new_n9341));
  xnor_3 g08965(.A(new_n9341), .B(new_n9218), .Y(new_n9342));
  xnor_3 g08966(.A(new_n9342), .B(new_n9212), .Y(new_n9343));
  xnor_3 g08967(.A(new_n9343), .B(new_n9145), .Y(n3287));
  xnor_3 g08968(.A(new_n9141), .B(new_n9117), .Y(n3339));
  not_3  g08969(.A(new_n4119), .Y(new_n9346));
  xor_3  g08970(.A(new_n9346), .B(new_n4117), .Y(n3456));
  nand_4 g08971(.A(n6687), .B(n4005), .Y(new_n9348));
  not_3  g08972(.A(new_n9348), .Y(new_n9349));
  nand_4 g08973(.A(n12720), .B(n6770), .Y(new_n9350));
  not_3  g08974(.A(new_n9350), .Y(new_n9351));
  nand_4 g08975(.A(n9920), .B(n2509), .Y(new_n9352));
  nand_4 g08976(.A(n6038), .B(n3627), .Y(new_n9353));
  xor_3  g08977(.A(new_n9353), .B(new_n9352), .Y(new_n9354));
  xnor_3 g08978(.A(new_n9354), .B(new_n9351), .Y(new_n9355));
  nand_4 g08979(.A(n9920), .B(n6038), .Y(new_n9356));
  not_3  g08980(.A(new_n9356), .Y(new_n9357));
  nand_4 g08981(.A(n12720), .B(n4189), .Y(new_n9358));
  not_3  g08982(.A(new_n9358), .Y(new_n9359));
  nor_4  g08983(.A(new_n9359), .B(new_n9357), .Y(new_n9360));
  nand_4 g08984(.A(n6770), .B(n2509), .Y(new_n9361));
  not_3  g08985(.A(new_n9361), .Y(new_n9362));
  xnor_3 g08986(.A(new_n9358), .B(new_n9356), .Y(new_n9363));
  nor_4  g08987(.A(new_n9363), .B(new_n9362), .Y(new_n9364));
  nor_4  g08988(.A(new_n9364), .B(new_n9360), .Y(new_n9365));
  not_3  g08989(.A(new_n9365), .Y(new_n9366));
  xnor_3 g08990(.A(new_n9366), .B(new_n9355), .Y(new_n9367));
  nand_4 g08991(.A(n2564), .B(n2508), .Y(new_n9368));
  not_3  g08992(.A(new_n9368), .Y(new_n9369));
  nand_4 g08993(.A(n6770), .B(n6038), .Y(new_n9370));
  not_3  g08994(.A(new_n9370), .Y(new_n9371));
  nand_4 g08995(.A(n4189), .B(n2509), .Y(new_n9372));
  not_3  g08996(.A(new_n9372), .Y(new_n9373));
  nor_4  g08997(.A(new_n9373), .B(new_n9371), .Y(new_n9374));
  nand_4 g08998(.A(n12720), .B(n2564), .Y(new_n9375));
  not_3  g08999(.A(new_n9375), .Y(new_n9376));
  xnor_3 g09000(.A(new_n9372), .B(new_n9370), .Y(new_n9377));
  nor_4  g09001(.A(new_n9377), .B(new_n9376), .Y(new_n9378));
  nor_4  g09002(.A(new_n9378), .B(new_n9374), .Y(new_n9379));
  nand_4 g09003(.A(new_n9379), .B(new_n9369), .Y(new_n9380));
  xnor_3 g09004(.A(new_n9363), .B(new_n9362), .Y(new_n9381));
  xnor_3 g09005(.A(new_n9379), .B(new_n9368), .Y(new_n9382));
  nand_4 g09006(.A(new_n9382), .B(new_n9381), .Y(new_n9383));
  nand_4 g09007(.A(new_n9383), .B(new_n9380), .Y(new_n9384));
  nand_4 g09008(.A(n2585), .B(n2564), .Y(new_n9385));
  nand_4 g09009(.A(n4189), .B(n2508), .Y(new_n9386));
  xor_3  g09010(.A(new_n9386), .B(new_n9385), .Y(new_n9387_1));
  xnor_3 g09011(.A(new_n9387_1), .B(new_n9384), .Y(new_n9388));
  xnor_3 g09012(.A(new_n9388), .B(new_n9367), .Y(new_n9389));
  nand_4 g09013(.A(n6687), .B(n2585), .Y(new_n9390));
  not_3  g09014(.A(new_n9390), .Y(new_n9391));
  nand_4 g09015(.A(n6687), .B(n2508), .Y(new_n9392));
  nand_4 g09016(.A(new_n9359), .B(new_n378), .Y(new_n9393));
  nand_4 g09017(.A(n6038), .B(n4189), .Y(new_n9394));
  nand_4 g09018(.A(n12720), .B(n6687), .Y(new_n9395));
  nand_4 g09019(.A(new_n9395), .B(new_n9394), .Y(new_n9396));
  nand_4 g09020(.A(n2564), .B(n2509), .Y(new_n9397));
  not_3  g09021(.A(new_n9397), .Y(new_n9398));
  nand_4 g09022(.A(new_n9398), .B(new_n9396), .Y(new_n9399));
  nand_4 g09023(.A(new_n9399), .B(new_n9393), .Y(new_n9400_1));
  not_3  g09024(.A(new_n9400_1), .Y(new_n9401));
  nor_4  g09025(.A(new_n9401), .B(new_n9392), .Y(new_n9402));
  not_3  g09026(.A(new_n9402), .Y(new_n9403));
  not_3  g09027(.A(new_n9392), .Y(new_n9404));
  xor_3  g09028(.A(new_n9400_1), .B(new_n9404), .Y(new_n9405));
  xor_3  g09029(.A(new_n9377), .B(new_n9375), .Y(new_n9406));
  nand_4 g09030(.A(new_n9406), .B(new_n9405), .Y(new_n9407));
  nand_4 g09031(.A(new_n9407), .B(new_n9403), .Y(new_n9408));
  nor_4  g09032(.A(new_n9408), .B(new_n9391), .Y(new_n9409));
  not_3  g09033(.A(new_n9409), .Y(new_n9410));
  xor_3  g09034(.A(new_n9382), .B(new_n9381), .Y(new_n9411));
  not_3  g09035(.A(new_n9408), .Y(new_n9412));
  xor_3  g09036(.A(new_n9412), .B(new_n9391), .Y(new_n9413));
  nor_4  g09037(.A(new_n9413), .B(new_n9411), .Y(new_n9414));
  not_3  g09038(.A(new_n9414), .Y(new_n9415));
  nand_4 g09039(.A(new_n9415), .B(new_n9410), .Y(new_n9416));
  nor_4  g09040(.A(new_n9416), .B(new_n9389), .Y(new_n9417));
  not_3  g09041(.A(new_n9389), .Y(new_n9418));
  nor_4  g09042(.A(new_n9414), .B(new_n9409), .Y(new_n9419));
  nor_4  g09043(.A(new_n9419), .B(new_n9418), .Y(new_n9420));
  nor_4  g09044(.A(new_n9420), .B(new_n9417), .Y(new_n9421));
  nand_4 g09045(.A(new_n9421), .B(new_n9349), .Y(new_n9422));
  not_3  g09046(.A(new_n9393), .Y(new_n9423));
  not_3  g09047(.A(new_n9396), .Y(new_n9424));
  nor_4  g09048(.A(new_n9424), .B(new_n9423), .Y(new_n9425));
  nand_4 g09049(.A(n6038), .B(n2564), .Y(new_n9426));
  nand_4 g09050(.A(n6687), .B(n2509), .Y(new_n9427));
  nor_4  g09051(.A(new_n9427), .B(new_n9426), .Y(new_n9428));
  not_3  g09052(.A(new_n9428), .Y(new_n9429));
  nor_4  g09053(.A(new_n9429), .B(new_n9425), .Y(new_n9430));
  xor_3  g09054(.A(new_n9406), .B(new_n9405), .Y(new_n9431));
  nand_4 g09055(.A(new_n9431), .B(new_n9430), .Y(new_n9432));
  not_3  g09056(.A(new_n9411), .Y(new_n9433));
  not_3  g09057(.A(new_n9413), .Y(new_n9434));
  nor_4  g09058(.A(new_n9434), .B(new_n9433), .Y(new_n9435));
  nor_4  g09059(.A(new_n9435), .B(new_n9414), .Y(new_n9436));
  nor_4  g09060(.A(new_n9436), .B(new_n9432), .Y(new_n9437));
  xnor_3 g09061(.A(new_n9421), .B(new_n9348), .Y(new_n9438));
  nand_4 g09062(.A(new_n9438), .B(new_n9437), .Y(new_n9439));
  nand_4 g09063(.A(new_n9439), .B(new_n9422), .Y(new_n9440));
  nor_4  g09064(.A(new_n9354), .B(new_n9351), .Y(new_n9441));
  not_3  g09065(.A(new_n9441), .Y(new_n9442));
  nor_4  g09066(.A(new_n9365), .B(new_n9355), .Y(new_n9443));
  not_3  g09067(.A(new_n9443), .Y(new_n9444));
  nand_4 g09068(.A(new_n9444), .B(new_n9442), .Y(new_n9445));
  nand_4 g09069(.A(n4005), .B(n2564), .Y(new_n9446));
  nand_4 g09070(.A(n4189), .B(n2585), .Y(new_n9447));
  nand_4 g09071(.A(n12706), .B(n6687), .Y(new_n9448));
  not_3  g09072(.A(new_n9448), .Y(new_n9449));
  xor_3  g09073(.A(new_n9449), .B(new_n9447), .Y(new_n9450));
  xnor_3 g09074(.A(new_n9450), .B(new_n9446), .Y(new_n9451));
  not_3  g09075(.A(new_n9451), .Y(new_n9452));
  xnor_3 g09076(.A(new_n9452), .B(new_n9445), .Y(new_n9453));
  nor_4  g09077(.A(new_n9353), .B(new_n9352), .Y(new_n9454));
  nand_4 g09078(.A(n6770), .B(n2508), .Y(new_n9455));
  not_3  g09079(.A(new_n9455), .Y(new_n9456));
  xor_3  g09080(.A(new_n9456), .B(new_n9454), .Y(new_n9457_1));
  not_3  g09081(.A(new_n9457_1), .Y(new_n9458));
  nand_4 g09082(.A(n3627), .B(n2509), .Y(new_n9459));
  not_3  g09083(.A(new_n9459), .Y(new_n9460));
  nand_4 g09084(.A(n12720), .B(n9920), .Y(new_n9461));
  nand_4 g09085(.A(n6038), .B(n4516), .Y(new_n9462));
  nand_4 g09086(.A(new_n9462), .B(new_n9461), .Y(new_n9463));
  not_3  g09087(.A(new_n9461), .Y(new_n9464));
  not_3  g09088(.A(new_n9462), .Y(new_n9465));
  nand_4 g09089(.A(new_n9465), .B(new_n9464), .Y(new_n9466));
  nand_4 g09090(.A(new_n9466), .B(new_n9463), .Y(new_n9467));
  xor_3  g09091(.A(new_n9467), .B(new_n9460), .Y(new_n9468));
  xnor_3 g09092(.A(new_n9468), .B(new_n9458), .Y(new_n9469));
  xnor_3 g09093(.A(new_n9469), .B(new_n9453), .Y(new_n9470));
  nand_4 g09094(.A(new_n9387_1), .B(new_n9384), .Y(new_n9471));
  nor_4  g09095(.A(new_n9386), .B(new_n9385), .Y(new_n9472));
  nor_4  g09096(.A(new_n9388), .B(new_n9367), .Y(new_n9473));
  xnor_3 g09097(.A(new_n9473), .B(new_n9472), .Y(new_n9474));
  nand_4 g09098(.A(new_n9474), .B(new_n9471), .Y(new_n9475));
  xnor_3 g09099(.A(new_n9475), .B(new_n9470), .Y(new_n9476));
  xnor_3 g09100(.A(new_n9476), .B(new_n9417), .Y(new_n9477));
  xnor_3 g09101(.A(new_n9477), .B(new_n9440), .Y(new_n9478));
  not_3  g09102(.A(new_n9478), .Y(new_n9479));
  nand_4 g09103(.A(n8336), .B(n1209), .Y(new_n9480));
  nand_4 g09104(.A(n7354), .B(n6986), .Y(new_n9481));
  nand_4 g09105(.A(new_n9481), .B(new_n9480), .Y(new_n9482));
  not_3  g09106(.A(new_n9482), .Y(new_n9483));
  not_3  g09107(.A(new_n9480), .Y(new_n9484));
  not_3  g09108(.A(new_n9481), .Y(new_n9485));
  nand_4 g09109(.A(new_n9485), .B(new_n9484), .Y(new_n9486));
  not_3  g09110(.A(new_n9486), .Y(new_n9487));
  nor_4  g09111(.A(new_n9487), .B(new_n9483), .Y(new_n9488));
  nand_4 g09112(.A(n10928), .B(n7354), .Y(new_n9489));
  nand_4 g09113(.A(n8336), .B(n7500), .Y(new_n9490));
  nor_4  g09114(.A(new_n9490), .B(new_n9489), .Y(new_n9491));
  not_3  g09115(.A(new_n9491), .Y(new_n9492));
  nor_4  g09116(.A(new_n9492), .B(new_n9488), .Y(new_n9493));
  not_3  g09117(.A(new_n9493), .Y(new_n9494));
  nand_4 g09118(.A(n8336), .B(n5105), .Y(new_n9495));
  not_3  g09119(.A(new_n9495), .Y(new_n9496));
  nand_4 g09120(.A(n10928), .B(n7500), .Y(new_n9497));
  not_3  g09121(.A(new_n9497), .Y(new_n9498));
  nand_4 g09122(.A(new_n9498), .B(new_n9482), .Y(new_n9499));
  nand_4 g09123(.A(new_n9499), .B(new_n9486), .Y(new_n9500));
  xor_3  g09124(.A(new_n9500), .B(new_n9496), .Y(new_n9501));
  nand_4 g09125(.A(n7500), .B(n6986), .Y(new_n9502));
  not_3  g09126(.A(new_n9502), .Y(new_n9503));
  nand_4 g09127(.A(n7354), .B(n2226), .Y(new_n9504));
  not_3  g09128(.A(new_n9504), .Y(new_n9505));
  nand_4 g09129(.A(n10928), .B(n1209), .Y(new_n9506));
  not_3  g09130(.A(new_n9506), .Y(new_n9507));
  nor_4  g09131(.A(new_n9507), .B(new_n9505), .Y(new_n9508));
  nor_4  g09132(.A(new_n9506), .B(new_n9504), .Y(new_n9509));
  nor_4  g09133(.A(new_n9509), .B(new_n9508), .Y(new_n9510));
  xor_3  g09134(.A(new_n9510), .B(new_n9503), .Y(new_n9511));
  xnor_3 g09135(.A(new_n9511), .B(new_n9501), .Y(new_n9512));
  nor_4  g09136(.A(new_n9512), .B(new_n9494), .Y(new_n9513));
  nand_4 g09137(.A(n8336), .B(n4141), .Y(new_n9514));
  not_3  g09138(.A(new_n9514), .Y(new_n9515));
  not_3  g09139(.A(new_n9500), .Y(new_n9516));
  nor_4  g09140(.A(new_n9516), .B(new_n9495), .Y(new_n9517));
  not_3  g09141(.A(new_n9517), .Y(new_n9518));
  nand_4 g09142(.A(new_n9511), .B(new_n9501), .Y(new_n9519));
  nand_4 g09143(.A(new_n9519), .B(new_n9518), .Y(new_n9520));
  not_3  g09144(.A(new_n9520), .Y(new_n9521));
  xor_3  g09145(.A(new_n9521), .B(new_n9515), .Y(new_n9522));
  nand_4 g09146(.A(n10928), .B(n5105), .Y(new_n9523));
  not_3  g09147(.A(new_n9523), .Y(new_n9524));
  nor_4  g09148(.A(new_n9509), .B(new_n9503), .Y(new_n9525));
  nor_4  g09149(.A(new_n9525), .B(new_n9508), .Y(new_n9526));
  xor_3  g09150(.A(new_n9526), .B(new_n9524), .Y(new_n9527));
  nand_4 g09151(.A(n6986), .B(n1209), .Y(new_n9528));
  not_3  g09152(.A(new_n9528), .Y(new_n9529));
  nand_4 g09153(.A(n7500), .B(n2226), .Y(new_n9530));
  nand_4 g09154(.A(n7354), .B(n1094), .Y(new_n9531));
  xnor_3 g09155(.A(new_n9531), .B(new_n9530), .Y(new_n9532));
  xor_3  g09156(.A(new_n9532), .B(new_n9529), .Y(new_n9533));
  xnor_3 g09157(.A(new_n9533), .B(new_n9527), .Y(new_n9534));
  xnor_3 g09158(.A(new_n9534), .B(new_n9522), .Y(new_n9535));
  nand_4 g09159(.A(new_n9535), .B(new_n9513), .Y(new_n9536));
  not_3  g09160(.A(new_n9536), .Y(new_n9537));
  nand_4 g09161(.A(n8336), .B(n4928), .Y(new_n9538));
  not_3  g09162(.A(new_n9538), .Y(new_n9539));
  nand_4 g09163(.A(n2226), .B(n1209), .Y(new_n9540));
  not_3  g09164(.A(new_n9540), .Y(new_n9541));
  not_3  g09165(.A(new_n9530), .Y(new_n9542));
  not_3  g09166(.A(new_n9531), .Y(new_n9543));
  nor_4  g09167(.A(new_n9543), .B(new_n9542), .Y(new_n9544));
  nor_4  g09168(.A(new_n9532), .B(new_n9529), .Y(new_n9545));
  nor_4  g09169(.A(new_n9545), .B(new_n9544), .Y(new_n9546));
  xnor_3 g09170(.A(new_n9546), .B(new_n9541), .Y(new_n9547));
  nand_4 g09171(.A(n7500), .B(n1094), .Y(new_n9548));
  nand_4 g09172(.A(n10678), .B(n7354), .Y(new_n9549));
  not_3  g09173(.A(new_n9549), .Y(new_n9550));
  xor_3  g09174(.A(new_n9550), .B(new_n9548), .Y(new_n9551));
  xnor_3 g09175(.A(new_n9551), .B(new_n9547), .Y(new_n9552));
  not_3  g09176(.A(new_n9552), .Y(new_n9553));
  nand_4 g09177(.A(n10928), .B(n4141), .Y(new_n9554));
  nand_4 g09178(.A(n6986), .B(n5105), .Y(new_n9555));
  xor_3  g09179(.A(new_n9555), .B(new_n9554), .Y(new_n9556));
  not_3  g09180(.A(new_n9556), .Y(new_n9557));
  xor_3  g09181(.A(new_n9557), .B(new_n9553), .Y(new_n9558));
  and_4  g09182(.A(new_n9526), .B(new_n9524), .Y(new_n9559));
  not_3  g09183(.A(new_n9527), .Y(new_n9560));
  nor_4  g09184(.A(new_n9533), .B(new_n9560), .Y(new_n9561));
  nor_4  g09185(.A(new_n9561), .B(new_n9559), .Y(new_n9562));
  xnor_3 g09186(.A(new_n9562), .B(new_n9558), .Y(new_n9563));
  not_3  g09187(.A(new_n9563), .Y(new_n9564));
  nor_4  g09188(.A(new_n9520), .B(new_n9515), .Y(new_n9565));
  nor_4  g09189(.A(new_n9534), .B(new_n9522), .Y(new_n9566));
  nor_4  g09190(.A(new_n9566), .B(new_n9565), .Y(new_n9567));
  xnor_3 g09191(.A(new_n9567), .B(new_n9564), .Y(new_n9568));
  xnor_3 g09192(.A(new_n9568), .B(new_n9539), .Y(new_n9569));
  xnor_3 g09193(.A(new_n9569), .B(new_n9537), .Y(new_n9570));
  nand_4 g09194(.A(n8028), .B(n5314), .Y(new_n9571_1));
  not_3  g09195(.A(new_n9571_1), .Y(new_n9572));
  nand_4 g09196(.A(n11222), .B(n1980), .Y(new_n9573));
  not_3  g09197(.A(new_n9573), .Y(new_n9574));
  nand_4 g09198(.A(new_n9574), .B(new_n9572), .Y(new_n9575));
  nand_4 g09199(.A(new_n9573), .B(new_n9571_1), .Y(new_n9576));
  nand_4 g09200(.A(new_n9576), .B(new_n9575), .Y(new_n9577));
  nand_4 g09201(.A(n11153), .B(n8028), .Y(new_n9578_1));
  nand_4 g09202(.A(n11222), .B(n10848), .Y(new_n9579));
  nor_4  g09203(.A(new_n9579), .B(new_n9578_1), .Y(new_n9580));
  and_4  g09204(.A(new_n9580), .B(new_n9577), .Y(new_n9581));
  not_3  g09205(.A(new_n9581), .Y(new_n9582));
  nand_4 g09206(.A(n11222), .B(n7294), .Y(new_n9583_1));
  nand_4 g09207(.A(n11153), .B(n10848), .Y(new_n9584));
  not_3  g09208(.A(new_n9584), .Y(new_n9585));
  nand_4 g09209(.A(new_n9585), .B(new_n9576), .Y(new_n9586));
  nand_4 g09210(.A(new_n9586), .B(new_n9575), .Y(new_n9587));
  not_3  g09211(.A(new_n9587), .Y(new_n9588));
  xnor_3 g09212(.A(new_n9588), .B(new_n9583_1), .Y(new_n9589));
  nand_4 g09213(.A(n10848), .B(n5314), .Y(new_n9590));
  not_3  g09214(.A(new_n9590), .Y(new_n9591));
  nand_4 g09215(.A(n8028), .B(n996), .Y(new_n9592));
  not_3  g09216(.A(new_n9592), .Y(new_n9593));
  nand_4 g09217(.A(n11153), .B(n1980), .Y(new_n9594));
  not_3  g09218(.A(new_n9594), .Y(new_n9595));
  nor_4  g09219(.A(new_n9595), .B(new_n9593), .Y(new_n9596));
  nor_4  g09220(.A(new_n9594), .B(new_n9592), .Y(new_n9597));
  nor_4  g09221(.A(new_n9597), .B(new_n9596), .Y(new_n9598));
  xnor_3 g09222(.A(new_n9598), .B(new_n9591), .Y(new_n9599));
  xnor_3 g09223(.A(new_n9599), .B(new_n9589), .Y(new_n9600));
  nor_4  g09224(.A(new_n9600), .B(new_n9582), .Y(new_n9601));
  not_3  g09225(.A(new_n9601), .Y(new_n9602));
  nor_4  g09226(.A(new_n9588), .B(new_n9583_1), .Y(new_n9603));
  nor_4  g09227(.A(new_n9599), .B(new_n9589), .Y(new_n9604));
  nor_4  g09228(.A(new_n9604), .B(new_n9603), .Y(new_n9605));
  nand_4 g09229(.A(n12704), .B(n11222), .Y(new_n9606));
  not_3  g09230(.A(new_n9606), .Y(new_n9607));
  nand_4 g09231(.A(n11153), .B(n7294), .Y(new_n9608));
  not_3  g09232(.A(new_n9608), .Y(new_n9609));
  nor_4  g09233(.A(new_n9597), .B(new_n9591), .Y(new_n9610));
  nor_4  g09234(.A(new_n9610), .B(new_n9596), .Y(new_n9611));
  xnor_3 g09235(.A(new_n9611), .B(new_n9609), .Y(new_n9612));
  nand_4 g09236(.A(n10848), .B(n996), .Y(new_n9613));
  not_3  g09237(.A(new_n9613), .Y(new_n9614));
  nand_4 g09238(.A(n5314), .B(n1980), .Y(new_n9615));
  not_3  g09239(.A(new_n9615), .Y(new_n9616));
  nand_4 g09240(.A(n8028), .B(n5767), .Y(new_n9617));
  not_3  g09241(.A(new_n9617), .Y(new_n9618));
  nor_4  g09242(.A(new_n9618), .B(new_n9616), .Y(new_n9619));
  not_3  g09243(.A(new_n9619), .Y(new_n9620));
  nor_4  g09244(.A(new_n9617), .B(new_n9615), .Y(new_n9621));
  not_3  g09245(.A(new_n9621), .Y(new_n9622));
  nand_4 g09246(.A(new_n9622), .B(new_n9620), .Y(new_n9623));
  xnor_3 g09247(.A(new_n9623), .B(new_n9614), .Y(new_n9624));
  xnor_3 g09248(.A(new_n9624), .B(new_n9612), .Y(new_n9625));
  nor_4  g09249(.A(new_n9625), .B(new_n9607), .Y(new_n9626));
  not_3  g09250(.A(new_n9625), .Y(new_n9627));
  nor_4  g09251(.A(new_n9627), .B(new_n9606), .Y(new_n9628));
  nor_4  g09252(.A(new_n9628), .B(new_n9626), .Y(new_n9629));
  xnor_3 g09253(.A(new_n9629), .B(new_n9605), .Y(new_n9630));
  not_3  g09254(.A(new_n9630), .Y(new_n9631));
  nor_4  g09255(.A(new_n9631), .B(new_n9602), .Y(new_n9632));
  nor_4  g09256(.A(new_n9630), .B(new_n9601), .Y(new_n9633));
  nor_4  g09257(.A(new_n9633), .B(new_n9632), .Y(new_n9634));
  nand_4 g09258(.A(n7891), .B(n1564), .Y(new_n9635));
  nand_4 g09259(.A(n12069), .B(n533), .Y(new_n9636));
  nand_4 g09260(.A(new_n9636), .B(new_n9635), .Y(new_n9637_1));
  nor_4  g09261(.A(new_n9636), .B(new_n9635), .Y(new_n9638));
  not_3  g09262(.A(new_n9638), .Y(new_n9639));
  nand_4 g09263(.A(new_n9639), .B(new_n9637_1), .Y(new_n9640_1));
  not_3  g09264(.A(new_n9640_1), .Y(new_n9641));
  nand_4 g09265(.A(n12391), .B(n1564), .Y(new_n9642));
  nand_4 g09266(.A(n12069), .B(n1512), .Y(new_n9643));
  nor_4  g09267(.A(new_n9643), .B(new_n9642), .Y(new_n9644));
  not_3  g09268(.A(new_n9644), .Y(new_n9645));
  nor_4  g09269(.A(new_n9645), .B(new_n9641), .Y(new_n9646));
  not_3  g09270(.A(new_n9646), .Y(new_n9647));
  nand_4 g09271(.A(n12069), .B(n2802), .Y(new_n9648));
  nand_4 g09272(.A(n12391), .B(n1512), .Y(new_n9649));
  not_3  g09273(.A(new_n9649), .Y(new_n9650));
  nand_4 g09274(.A(new_n9650), .B(new_n9637_1), .Y(new_n9651));
  nand_4 g09275(.A(new_n9651), .B(new_n9639), .Y(new_n9652));
  not_3  g09276(.A(new_n9652), .Y(new_n9653));
  nor_4  g09277(.A(new_n9653), .B(new_n9648), .Y(new_n9654));
  not_3  g09278(.A(new_n9648), .Y(new_n9655));
  nor_4  g09279(.A(new_n9652), .B(new_n9655), .Y(new_n9656));
  nor_4  g09280(.A(new_n9656), .B(new_n9654), .Y(new_n9657));
  nand_4 g09281(.A(n7891), .B(n1512), .Y(new_n9658));
  nand_4 g09282(.A(n7160), .B(n1564), .Y(new_n9659));
  nand_4 g09283(.A(n12391), .B(n533), .Y(new_n9660));
  xnor_3 g09284(.A(new_n9660), .B(new_n9659), .Y(new_n9661));
  xnor_3 g09285(.A(new_n9661), .B(new_n9658), .Y(new_n9662));
  not_3  g09286(.A(new_n9662), .Y(new_n9663));
  xnor_3 g09287(.A(new_n9663), .B(new_n9657), .Y(new_n9664));
  nor_4  g09288(.A(new_n9664), .B(new_n9647), .Y(new_n9665));
  not_3  g09289(.A(new_n9664), .Y(new_n9666));
  nor_4  g09290(.A(new_n9666), .B(new_n9646), .Y(new_n9667));
  nor_4  g09291(.A(new_n9667), .B(new_n9665), .Y(new_n9668));
  not_3  g09292(.A(new_n9600), .Y(new_n9669));
  nor_4  g09293(.A(new_n9669), .B(new_n9581), .Y(new_n9670));
  nor_4  g09294(.A(new_n9670), .B(new_n9601), .Y(new_n9671));
  nor_4  g09295(.A(new_n9671), .B(new_n9668), .Y(new_n9672));
  nand_4 g09296(.A(new_n9650), .B(new_n382), .Y(new_n9673));
  nand_4 g09297(.A(new_n9673), .B(new_n9640_1), .Y(new_n9674));
  not_3  g09298(.A(new_n9651), .Y(new_n9675));
  nand_4 g09299(.A(new_n9675), .B(new_n382), .Y(new_n9676));
  nand_4 g09300(.A(new_n9676), .B(new_n9674), .Y(new_n9677));
  not_3  g09301(.A(new_n381_1), .Y(new_n9678));
  nor_4  g09302(.A(new_n9584), .B(new_n9678), .Y(new_n9679));
  not_3  g09303(.A(new_n9679), .Y(new_n9680));
  nand_4 g09304(.A(new_n9680), .B(new_n9577), .Y(new_n9681));
  nand_4 g09305(.A(new_n9679), .B(new_n9576), .Y(new_n9682));
  nand_4 g09306(.A(new_n9682), .B(new_n9681), .Y(new_n9683));
  and_4  g09307(.A(new_n9683), .B(new_n9677), .Y(new_n9684));
  nor_4  g09308(.A(new_n382), .B(new_n381_1), .Y(new_n9685));
  xnor_3 g09309(.A(new_n9579), .B(new_n9578_1), .Y(new_n9686));
  not_3  g09310(.A(new_n9686), .Y(new_n9687));
  nor_4  g09311(.A(new_n9687), .B(new_n9685), .Y(new_n9688));
  xor_3  g09312(.A(new_n9686), .B(new_n9685), .Y(new_n9689));
  xor_3  g09313(.A(new_n9643), .B(new_n9642), .Y(new_n9690));
  nor_4  g09314(.A(new_n9690), .B(new_n9689), .Y(new_n9691));
  nor_4  g09315(.A(new_n9691), .B(new_n9688), .Y(new_n9692));
  xnor_3 g09316(.A(new_n9683), .B(new_n9677), .Y(new_n9693));
  nor_4  g09317(.A(new_n9693), .B(new_n9692), .Y(new_n9694));
  nor_4  g09318(.A(new_n9694), .B(new_n9684), .Y(new_n9695));
  xnor_3 g09319(.A(new_n9671), .B(new_n9668), .Y(new_n9696));
  nor_4  g09320(.A(new_n9696), .B(new_n9695), .Y(new_n9697));
  nor_4  g09321(.A(new_n9697), .B(new_n9672), .Y(new_n9698));
  nor_4  g09322(.A(new_n9698), .B(new_n9634), .Y(new_n9699));
  nand_4 g09323(.A(n12069), .B(n6806), .Y(new_n9700));
  nand_4 g09324(.A(n12391), .B(n2802), .Y(new_n9701));
  not_3  g09325(.A(new_n9701), .Y(new_n9702));
  not_3  g09326(.A(new_n9659), .Y(new_n9703));
  not_3  g09327(.A(new_n9660), .Y(new_n9704));
  nor_4  g09328(.A(new_n9704), .B(new_n9703), .Y(new_n9705));
  not_3  g09329(.A(new_n9658), .Y(new_n9706_1));
  nor_4  g09330(.A(new_n9661), .B(new_n9706_1), .Y(new_n9707));
  nor_4  g09331(.A(new_n9707), .B(new_n9705), .Y(new_n9708));
  xnor_3 g09332(.A(new_n9708), .B(new_n9702), .Y(new_n9709));
  nand_4 g09333(.A(n7891), .B(n533), .Y(new_n9710));
  nand_4 g09334(.A(n4828), .B(n1564), .Y(new_n9711));
  nand_4 g09335(.A(n7160), .B(n1512), .Y(new_n9712));
  xnor_3 g09336(.A(new_n9712), .B(new_n9711), .Y(new_n9713));
  xnor_3 g09337(.A(new_n9713), .B(new_n9710), .Y(new_n9714));
  xnor_3 g09338(.A(new_n9714), .B(new_n9709), .Y(new_n9715));
  nand_4 g09339(.A(new_n9715), .B(new_n9700), .Y(new_n9716));
  not_3  g09340(.A(new_n9716), .Y(new_n9717));
  nor_4  g09341(.A(new_n9715), .B(new_n9700), .Y(new_n9718));
  nor_4  g09342(.A(new_n9718), .B(new_n9717), .Y(new_n9719));
  not_3  g09343(.A(new_n9654), .Y(new_n9720));
  nand_4 g09344(.A(new_n9663), .B(new_n9657), .Y(new_n9721));
  nand_4 g09345(.A(new_n9721), .B(new_n9720), .Y(new_n9722));
  not_3  g09346(.A(new_n9722), .Y(new_n9723));
  xnor_3 g09347(.A(new_n9723), .B(new_n9719), .Y(new_n9724));
  nand_4 g09348(.A(new_n9724), .B(new_n9665), .Y(new_n9725_1));
  not_3  g09349(.A(new_n9725_1), .Y(new_n9726));
  nor_4  g09350(.A(new_n9724), .B(new_n9665), .Y(new_n9727));
  nor_4  g09351(.A(new_n9727), .B(new_n9726), .Y(new_n9728));
  xnor_3 g09352(.A(new_n9698), .B(new_n9634), .Y(new_n9729));
  nor_4  g09353(.A(new_n9729), .B(new_n9728), .Y(new_n9730));
  nor_4  g09354(.A(new_n9730), .B(new_n9699), .Y(new_n9731));
  not_3  g09355(.A(new_n9731), .Y(new_n9732));
  nand_4 g09356(.A(n11222), .B(n5814), .Y(new_n9733));
  nand_4 g09357(.A(n1980), .B(n996), .Y(new_n9734));
  nand_4 g09358(.A(n8028), .B(n5319), .Y(new_n9735));
  nand_4 g09359(.A(n10848), .B(n5767), .Y(new_n9736));
  xnor_3 g09360(.A(new_n9736), .B(new_n9735), .Y(new_n9737));
  nor_4  g09361(.A(new_n9737), .B(new_n9734), .Y(new_n9738));
  not_3  g09362(.A(new_n9734), .Y(new_n9739));
  not_3  g09363(.A(new_n9737), .Y(new_n9740));
  nor_4  g09364(.A(new_n9740), .B(new_n9739), .Y(new_n9741));
  nor_4  g09365(.A(new_n9741), .B(new_n9738), .Y(new_n9742));
  nor_4  g09366(.A(new_n9621), .B(new_n9614), .Y(new_n9743));
  nor_4  g09367(.A(new_n9743), .B(new_n9619), .Y(new_n9744));
  xnor_3 g09368(.A(new_n9744), .B(new_n9742), .Y(new_n9745));
  nand_4 g09369(.A(n12704), .B(n11153), .Y(new_n9746));
  nand_4 g09370(.A(n7294), .B(n5314), .Y(new_n9747));
  xor_3  g09371(.A(new_n9747), .B(new_n9746), .Y(new_n9748));
  xnor_3 g09372(.A(new_n9748), .B(new_n9745), .Y(new_n9749));
  and_4  g09373(.A(new_n9611), .B(new_n9609), .Y(new_n9750));
  not_3  g09374(.A(new_n9624), .Y(new_n9751));
  nor_4  g09375(.A(new_n9751), .B(new_n9612), .Y(new_n9752));
  nor_4  g09376(.A(new_n9752), .B(new_n9750), .Y(new_n9753));
  xnor_3 g09377(.A(new_n9753), .B(new_n9749), .Y(new_n9754));
  not_3  g09378(.A(new_n9628), .Y(new_n9755));
  nor_4  g09379(.A(new_n9626), .B(new_n9605), .Y(new_n9756_1));
  not_3  g09380(.A(new_n9756_1), .Y(new_n9757));
  nand_4 g09381(.A(new_n9757), .B(new_n9755), .Y(new_n9758));
  xnor_3 g09382(.A(new_n9758), .B(new_n9754), .Y(new_n9759));
  xnor_3 g09383(.A(new_n9759), .B(new_n9733), .Y(new_n9760));
  xnor_3 g09384(.A(new_n9760), .B(new_n9632), .Y(new_n9761));
  nand_4 g09385(.A(n12069), .B(n5069), .Y(new_n9762));
  nand_4 g09386(.A(n7160), .B(n533), .Y(new_n9763_1));
  nand_4 g09387(.A(n2515), .B(n1564), .Y(new_n9764));
  nand_4 g09388(.A(n4828), .B(n1512), .Y(new_n9765));
  xnor_3 g09389(.A(new_n9765), .B(new_n9764), .Y(new_n9766));
  nor_4  g09390(.A(new_n9766), .B(new_n9763_1), .Y(new_n9767_1));
  not_3  g09391(.A(new_n9763_1), .Y(new_n9768));
  not_3  g09392(.A(new_n9766), .Y(new_n9769));
  nor_4  g09393(.A(new_n9769), .B(new_n9768), .Y(new_n9770));
  nor_4  g09394(.A(new_n9770), .B(new_n9767_1), .Y(new_n9771));
  and_4  g09395(.A(new_n9712), .B(new_n9711), .Y(new_n9772));
  not_3  g09396(.A(new_n9710), .Y(new_n9773));
  nor_4  g09397(.A(new_n9713), .B(new_n9773), .Y(new_n9774));
  nor_4  g09398(.A(new_n9774), .B(new_n9772), .Y(new_n9775));
  xnor_3 g09399(.A(new_n9775), .B(new_n9771), .Y(new_n9776));
  nand_4 g09400(.A(n7891), .B(n2802), .Y(new_n9777));
  nand_4 g09401(.A(n12391), .B(n6806), .Y(new_n9778));
  xor_3  g09402(.A(new_n9778), .B(new_n9777), .Y(new_n9779));
  not_3  g09403(.A(new_n9779), .Y(new_n9780));
  nor_4  g09404(.A(new_n9780), .B(new_n9776), .Y(new_n9781));
  not_3  g09405(.A(new_n9776), .Y(new_n9782));
  nor_4  g09406(.A(new_n9779), .B(new_n9782), .Y(new_n9783));
  nor_4  g09407(.A(new_n9783), .B(new_n9781), .Y(new_n9784));
  nand_4 g09408(.A(new_n9708), .B(new_n9702), .Y(new_n9785));
  not_3  g09409(.A(new_n9785), .Y(new_n9786));
  nor_4  g09410(.A(new_n9714), .B(new_n9709), .Y(new_n9787));
  nor_4  g09411(.A(new_n9787), .B(new_n9786), .Y(new_n9788));
  not_3  g09412(.A(new_n9788), .Y(new_n9789));
  xnor_3 g09413(.A(new_n9789), .B(new_n9784), .Y(new_n9790));
  nand_4 g09414(.A(new_n9723), .B(new_n9719), .Y(new_n9791));
  nand_4 g09415(.A(new_n9791), .B(new_n9716), .Y(new_n9792));
  xnor_3 g09416(.A(new_n9792), .B(new_n9790), .Y(new_n9793));
  nand_4 g09417(.A(new_n9793), .B(new_n9762), .Y(new_n9794));
  not_3  g09418(.A(new_n9762), .Y(new_n9795));
  not_3  g09419(.A(new_n9792), .Y(new_n9796));
  xnor_3 g09420(.A(new_n9796), .B(new_n9790), .Y(new_n9797));
  nand_4 g09421(.A(new_n9797), .B(new_n9795), .Y(new_n9798));
  nand_4 g09422(.A(new_n9798), .B(new_n9794), .Y(new_n9799));
  xnor_3 g09423(.A(new_n9799), .B(new_n9725_1), .Y(new_n9800));
  not_3  g09424(.A(new_n9800), .Y(new_n9801));
  nand_4 g09425(.A(new_n9801), .B(new_n9761), .Y(new_n9802));
  not_3  g09426(.A(new_n9761), .Y(new_n9803));
  nand_4 g09427(.A(new_n9800), .B(new_n9803), .Y(new_n9804));
  nand_4 g09428(.A(new_n9804), .B(new_n9802), .Y(new_n9805));
  xnor_3 g09429(.A(new_n9805), .B(new_n9732), .Y(new_n9806));
  nor_4  g09430(.A(new_n9806), .B(new_n9570), .Y(new_n9807));
  xnor_3 g09431(.A(new_n9806), .B(new_n9570), .Y(new_n9808));
  nor_4  g09432(.A(new_n9535), .B(new_n9513), .Y(new_n9809));
  nor_4  g09433(.A(new_n9809), .B(new_n9537), .Y(new_n9810));
  xnor_3 g09434(.A(new_n9729), .B(new_n9728), .Y(new_n9811));
  nand_4 g09435(.A(new_n9811), .B(new_n9810), .Y(new_n9812));
  not_3  g09436(.A(new_n9812), .Y(new_n9813));
  not_3  g09437(.A(new_n9810), .Y(new_n9814));
  not_3  g09438(.A(new_n9728), .Y(new_n9815));
  xnor_3 g09439(.A(new_n9729), .B(new_n9815), .Y(new_n9816));
  nand_4 g09440(.A(new_n9816), .B(new_n9814), .Y(new_n9817));
  nand_4 g09441(.A(new_n9817), .B(new_n9812), .Y(new_n9818));
  not_3  g09442(.A(new_n9512), .Y(new_n9819));
  xor_3  g09443(.A(new_n9819), .B(new_n9494), .Y(new_n9820_1));
  not_3  g09444(.A(new_n9696), .Y(new_n9821));
  xnor_3 g09445(.A(new_n9821), .B(new_n9695), .Y(new_n9822));
  nor_4  g09446(.A(new_n9822), .B(new_n9820_1), .Y(new_n9823));
  xnor_3 g09447(.A(new_n9822), .B(new_n9820_1), .Y(new_n9824));
  xnor_3 g09448(.A(new_n9693), .B(new_n9692), .Y(new_n9825));
  nor_4  g09449(.A(new_n9497), .B(new_n380), .Y(new_n9826));
  not_3  g09450(.A(new_n9826), .Y(new_n9827));
  nor_4  g09451(.A(new_n9827), .B(new_n9482), .Y(new_n9828));
  not_3  g09452(.A(new_n9488), .Y(new_n9829));
  nor_4  g09453(.A(new_n9826), .B(new_n9829), .Y(new_n9830));
  nor_4  g09454(.A(new_n9830), .B(new_n9828), .Y(new_n9831));
  not_3  g09455(.A(new_n9831), .Y(new_n9832));
  nor_4  g09456(.A(new_n9832), .B(new_n9825), .Y(new_n9833));
  not_3  g09457(.A(new_n9833), .Y(new_n9834));
  not_3  g09458(.A(new_n9825), .Y(new_n9835));
  xor_3  g09459(.A(new_n9831), .B(new_n9835), .Y(new_n9836));
  xnor_3 g09460(.A(new_n9690), .B(new_n9689), .Y(new_n9837));
  xor_3  g09461(.A(new_n9490), .B(new_n9489), .Y(new_n9838));
  nand_4 g09462(.A(new_n9838), .B(new_n9837), .Y(new_n9839));
  not_3  g09463(.A(new_n9839), .Y(new_n9840));
  nor_4  g09464(.A(new_n384), .B(new_n379), .Y(new_n9841));
  not_3  g09465(.A(new_n9841), .Y(new_n9842));
  xnor_3 g09466(.A(new_n9838), .B(new_n9837), .Y(new_n9843));
  nor_4  g09467(.A(new_n9843), .B(new_n9842), .Y(new_n9844));
  nor_4  g09468(.A(new_n9844), .B(new_n9840), .Y(new_n9845));
  nand_4 g09469(.A(new_n9845), .B(new_n9836), .Y(new_n9846));
  nand_4 g09470(.A(new_n9846), .B(new_n9834), .Y(new_n9847));
  nor_4  g09471(.A(new_n9847), .B(new_n9824), .Y(new_n9848));
  nor_4  g09472(.A(new_n9848), .B(new_n9823), .Y(new_n9849));
  nor_4  g09473(.A(new_n9849), .B(new_n9818), .Y(new_n9850));
  nor_4  g09474(.A(new_n9850), .B(new_n9813), .Y(new_n9851));
  nor_4  g09475(.A(new_n9851), .B(new_n9808), .Y(new_n9852));
  nor_4  g09476(.A(new_n9852), .B(new_n9807), .Y(new_n9853));
  nand_4 g09477(.A(new_n9567), .B(new_n9564), .Y(new_n9854));
  and_4  g09478(.A(new_n9546), .B(new_n9541), .Y(new_n9855));
  nor_4  g09479(.A(new_n9551), .B(new_n9547), .Y(new_n9856));
  nor_4  g09480(.A(new_n9856), .B(new_n9855), .Y(new_n9857));
  nand_4 g09481(.A(n10928), .B(n4928), .Y(new_n9858));
  nand_4 g09482(.A(n6986), .B(n4141), .Y(new_n9859));
  nand_4 g09483(.A(n8336), .B(n8236), .Y(new_n9860));
  xor_3  g09484(.A(new_n9860), .B(new_n9859), .Y(new_n9861));
  not_3  g09485(.A(new_n9861), .Y(new_n9862));
  xor_3  g09486(.A(new_n9862), .B(new_n9858), .Y(new_n9863));
  not_3  g09487(.A(new_n9863), .Y(new_n9864));
  xnor_3 g09488(.A(new_n9864), .B(new_n9857), .Y(new_n9865));
  nor_4  g09489(.A(new_n9549), .B(new_n9548), .Y(new_n9866));
  not_3  g09490(.A(new_n9866), .Y(new_n9867));
  nand_4 g09491(.A(n5105), .B(n2226), .Y(new_n9868));
  xor_3  g09492(.A(new_n9868), .B(new_n9867), .Y(new_n9869));
  nand_4 g09493(.A(n10678), .B(n7500), .Y(new_n9870));
  nand_4 g09494(.A(n7354), .B(n7320), .Y(new_n9871));
  nand_4 g09495(.A(n1209), .B(n1094), .Y(new_n9872));
  not_3  g09496(.A(new_n9872), .Y(new_n9873));
  xor_3  g09497(.A(new_n9873), .B(new_n9871), .Y(new_n9874));
  xnor_3 g09498(.A(new_n9874), .B(new_n9870), .Y(new_n9875));
  xnor_3 g09499(.A(new_n9875), .B(new_n9869), .Y(new_n9876));
  xnor_3 g09500(.A(new_n9876), .B(new_n9865), .Y(new_n9877));
  nand_4 g09501(.A(new_n9556), .B(new_n9553), .Y(new_n9878));
  nor_4  g09502(.A(new_n9555), .B(new_n9554), .Y(new_n9879));
  nor_4  g09503(.A(new_n9562), .B(new_n9558), .Y(new_n9880));
  xnor_3 g09504(.A(new_n9880), .B(new_n9879), .Y(new_n9881));
  nand_4 g09505(.A(new_n9881), .B(new_n9878), .Y(new_n9882));
  xnor_3 g09506(.A(new_n9882), .B(new_n9877), .Y(new_n9883));
  xnor_3 g09507(.A(new_n9883), .B(new_n9854), .Y(new_n9884));
  nand_4 g09508(.A(new_n9568), .B(new_n9538), .Y(new_n9885));
  nand_4 g09509(.A(new_n9569), .B(new_n9536), .Y(new_n9886));
  nand_4 g09510(.A(new_n9886), .B(new_n9885), .Y(new_n9887));
  xnor_3 g09511(.A(new_n9887), .B(new_n9884), .Y(new_n9888));
  not_3  g09512(.A(new_n9888), .Y(new_n9889));
  not_3  g09513(.A(new_n9754), .Y(new_n9890));
  not_3  g09514(.A(new_n9758), .Y(new_n9891));
  nor_4  g09515(.A(new_n9891), .B(new_n9890), .Y(new_n9892));
  not_3  g09516(.A(new_n9892), .Y(new_n9893));
  nand_4 g09517(.A(new_n9744), .B(new_n9742), .Y(new_n9894));
  not_3  g09518(.A(new_n9894), .Y(new_n9895));
  nor_4  g09519(.A(new_n9895), .B(new_n9738), .Y(new_n9896));
  not_3  g09520(.A(new_n9896), .Y(new_n9897));
  nand_4 g09521(.A(n11153), .B(n5814), .Y(new_n9898));
  nand_4 g09522(.A(n12704), .B(n5314), .Y(new_n9899));
  nand_4 g09523(.A(n11222), .B(n4903), .Y(new_n9900));
  not_3  g09524(.A(new_n9900), .Y(new_n9901));
  xor_3  g09525(.A(new_n9901), .B(new_n9899), .Y(new_n9902));
  xnor_3 g09526(.A(new_n9902), .B(new_n9898), .Y(new_n9903));
  xnor_3 g09527(.A(new_n9903), .B(new_n9897), .Y(new_n9904));
  nor_4  g09528(.A(new_n9736), .B(new_n9735), .Y(new_n9905));
  nand_4 g09529(.A(n7294), .B(n996), .Y(new_n9906));
  not_3  g09530(.A(new_n9906), .Y(new_n9907));
  xor_3  g09531(.A(new_n9907), .B(new_n9905), .Y(new_n9908));
  nand_4 g09532(.A(n10848), .B(n5319), .Y(new_n9909));
  not_3  g09533(.A(new_n9909), .Y(new_n9910));
  nand_4 g09534(.A(n5767), .B(n1980), .Y(new_n9911));
  nand_4 g09535(.A(n9457), .B(n8028), .Y(new_n9912));
  not_3  g09536(.A(new_n9912), .Y(new_n9913));
  xor_3  g09537(.A(new_n9913), .B(new_n9911), .Y(new_n9914));
  xnor_3 g09538(.A(new_n9914), .B(new_n9910), .Y(new_n9915));
  xnor_3 g09539(.A(new_n9915), .B(new_n9908), .Y(new_n9916));
  xnor_3 g09540(.A(new_n9916), .B(new_n9904), .Y(new_n9917));
  not_3  g09541(.A(new_n9917), .Y(new_n9918));
  not_3  g09542(.A(new_n9745), .Y(new_n9919));
  nand_4 g09543(.A(new_n9748), .B(new_n9919), .Y(new_n9920_1));
  nor_4  g09544(.A(new_n9747), .B(new_n9746), .Y(new_n9921));
  not_3  g09545(.A(new_n9749), .Y(new_n9922));
  nor_4  g09546(.A(new_n9753), .B(new_n9922), .Y(new_n9923));
  xnor_3 g09547(.A(new_n9923), .B(new_n9921), .Y(new_n9924));
  nand_4 g09548(.A(new_n9924), .B(new_n9920_1), .Y(new_n9925));
  xnor_3 g09549(.A(new_n9925), .B(new_n9918), .Y(new_n9926));
  xnor_3 g09550(.A(new_n9926), .B(new_n9893), .Y(new_n9927));
  not_3  g09551(.A(new_n9733), .Y(new_n9928));
  not_3  g09552(.A(new_n9759), .Y(new_n9929));
  nor_4  g09553(.A(new_n9929), .B(new_n9928), .Y(new_n9930));
  nor_4  g09554(.A(new_n9759), .B(new_n9733), .Y(new_n9931));
  nor_4  g09555(.A(new_n9931), .B(new_n9632), .Y(new_n9932));
  nor_4  g09556(.A(new_n9932), .B(new_n9930), .Y(new_n9933));
  xnor_3 g09557(.A(new_n9933), .B(new_n9927), .Y(new_n9934));
  nor_4  g09558(.A(new_n9792), .B(new_n9790), .Y(new_n9935));
  not_3  g09559(.A(new_n9935), .Y(new_n9936));
  not_3  g09560(.A(new_n9781), .Y(new_n9937));
  nor_4  g09561(.A(new_n9778), .B(new_n9777), .Y(new_n9938_1));
  nand_4 g09562(.A(new_n9789), .B(new_n9784), .Y(new_n9939));
  not_3  g09563(.A(new_n9939), .Y(new_n9940));
  xnor_3 g09564(.A(new_n9940), .B(new_n9938_1), .Y(new_n9941));
  nand_4 g09565(.A(new_n9941), .B(new_n9937), .Y(new_n9942));
  nor_4  g09566(.A(new_n9765), .B(new_n9764), .Y(new_n9943));
  nand_4 g09567(.A(n7160), .B(n2802), .Y(new_n9944));
  not_3  g09568(.A(new_n9944), .Y(new_n9945));
  xor_3  g09569(.A(new_n9945), .B(new_n9943), .Y(new_n9946));
  nand_4 g09570(.A(n2515), .B(n1512), .Y(new_n9947));
  not_3  g09571(.A(new_n9947), .Y(new_n9948));
  nand_4 g09572(.A(n1564), .B(n1199), .Y(new_n9949));
  nand_4 g09573(.A(n4828), .B(n533), .Y(new_n9950));
  nand_4 g09574(.A(new_n9950), .B(new_n9949), .Y(new_n9951));
  not_3  g09575(.A(new_n9949), .Y(new_n9952));
  not_3  g09576(.A(new_n9950), .Y(new_n9953));
  nand_4 g09577(.A(new_n9953), .B(new_n9952), .Y(new_n9954));
  nand_4 g09578(.A(new_n9954), .B(new_n9951), .Y(new_n9955));
  xor_3  g09579(.A(new_n9955), .B(new_n9948), .Y(new_n9956_1));
  not_3  g09580(.A(new_n9956_1), .Y(new_n9957));
  nor_4  g09581(.A(new_n9957), .B(new_n9946), .Y(new_n9958));
  not_3  g09582(.A(new_n9946), .Y(new_n9959));
  nor_4  g09583(.A(new_n9956_1), .B(new_n9959), .Y(new_n9960));
  nor_4  g09584(.A(new_n9960), .B(new_n9958), .Y(new_n9961));
  not_3  g09585(.A(new_n9767_1), .Y(new_n9962));
  nand_4 g09586(.A(new_n9775), .B(new_n9771), .Y(new_n9963));
  nand_4 g09587(.A(new_n9963), .B(new_n9962), .Y(new_n9964));
  nand_4 g09588(.A(n12391), .B(n5069), .Y(new_n9965));
  nand_4 g09589(.A(n7891), .B(n6806), .Y(new_n9966));
  nand_4 g09590(.A(n12069), .B(n12044), .Y(new_n9967));
  not_3  g09591(.A(new_n9967), .Y(new_n9968));
  xor_3  g09592(.A(new_n9968), .B(new_n9966), .Y(new_n9969));
  xnor_3 g09593(.A(new_n9969), .B(new_n9965), .Y(new_n9970));
  xnor_3 g09594(.A(new_n9970), .B(new_n9964), .Y(new_n9971));
  xnor_3 g09595(.A(new_n9971), .B(new_n9961), .Y(new_n9972));
  xnor_3 g09596(.A(new_n9972), .B(new_n9942), .Y(new_n9973));
  xnor_3 g09597(.A(new_n9973), .B(new_n9936), .Y(new_n9974));
  nand_4 g09598(.A(new_n9794), .B(new_n9726), .Y(new_n9975));
  nand_4 g09599(.A(new_n9975), .B(new_n9798), .Y(new_n9976));
  xnor_3 g09600(.A(new_n9976), .B(new_n9974), .Y(new_n9977));
  nand_4 g09601(.A(new_n9804), .B(new_n9731), .Y(new_n9978));
  nand_4 g09602(.A(new_n9978), .B(new_n9802), .Y(new_n9979));
  xnor_3 g09603(.A(new_n9979), .B(new_n9977), .Y(new_n9980));
  xnor_3 g09604(.A(new_n9980), .B(new_n9934), .Y(new_n9981));
  nand_4 g09605(.A(new_n9981), .B(new_n9889), .Y(new_n9982));
  not_3  g09606(.A(new_n9934), .Y(new_n9983));
  xnor_3 g09607(.A(new_n9980), .B(new_n9983), .Y(new_n9984));
  nand_4 g09608(.A(new_n9984), .B(new_n9888), .Y(new_n9985));
  nand_4 g09609(.A(new_n9985), .B(new_n9982), .Y(new_n9986));
  xnor_3 g09610(.A(new_n9986), .B(new_n9853), .Y(new_n9987));
  not_3  g09611(.A(new_n9987), .Y(new_n9988));
  nand_4 g09612(.A(new_n9988), .B(new_n9479), .Y(new_n9989));
  nand_4 g09613(.A(new_n9987), .B(new_n9478), .Y(new_n9990));
  not_3  g09614(.A(new_n9439), .Y(new_n9991));
  nor_4  g09615(.A(new_n9438), .B(new_n9437), .Y(new_n9992));
  nor_4  g09616(.A(new_n9992), .B(new_n9991), .Y(new_n9993));
  xnor_3 g09617(.A(new_n9436), .B(new_n9432), .Y(new_n9994));
  not_3  g09618(.A(new_n9994), .Y(new_n9995));
  xnor_3 g09619(.A(new_n9849), .B(new_n9818), .Y(new_n9996));
  not_3  g09620(.A(new_n9996), .Y(new_n9997));
  nand_4 g09621(.A(new_n9997), .B(new_n9995), .Y(new_n9998));
  nand_4 g09622(.A(new_n9996), .B(new_n9994), .Y(new_n9999));
  not_3  g09623(.A(new_n9430), .Y(new_n10000));
  xnor_3 g09624(.A(new_n9431), .B(new_n10000), .Y(new_n10001));
  not_3  g09625(.A(new_n9824), .Y(new_n10002));
  xnor_3 g09626(.A(new_n9847), .B(new_n10002), .Y(new_n10003));
  nor_4  g09627(.A(new_n10003), .B(new_n10001), .Y(new_n10004));
  xnor_3 g09628(.A(new_n10003), .B(new_n10001), .Y(new_n10005));
  xnor_3 g09629(.A(new_n9845), .B(new_n9836), .Y(new_n10006));
  nor_4  g09630(.A(new_n9397), .B(new_n378), .Y(new_n10007));
  nor_4  g09631(.A(new_n10007), .B(new_n9425), .Y(new_n10008));
  not_3  g09632(.A(new_n10007), .Y(new_n10009));
  nor_4  g09633(.A(new_n10009), .B(new_n9424), .Y(new_n10010));
  nor_4  g09634(.A(new_n10010), .B(new_n10008), .Y(new_n10011));
  nor_4  g09635(.A(new_n10011), .B(new_n10006), .Y(new_n10012));
  xnor_3 g09636(.A(new_n10011), .B(new_n10006), .Y(new_n10013));
  not_3  g09637(.A(new_n386), .Y(new_n10014));
  nor_4  g09638(.A(new_n10014), .B(new_n377), .Y(new_n10015));
  xor_3  g09639(.A(new_n9427), .B(new_n9426), .Y(new_n10016));
  nor_4  g09640(.A(new_n10016), .B(new_n10015), .Y(new_n10017));
  xnor_3 g09641(.A(new_n9843), .B(new_n9841), .Y(new_n10018));
  xnor_3 g09642(.A(new_n10016), .B(new_n10015), .Y(new_n10019));
  nor_4  g09643(.A(new_n10019), .B(new_n10018), .Y(new_n10020));
  nor_4  g09644(.A(new_n10020), .B(new_n10017), .Y(new_n10021));
  nor_4  g09645(.A(new_n10021), .B(new_n10013), .Y(new_n10022_1));
  nor_4  g09646(.A(new_n10022_1), .B(new_n10012), .Y(new_n10023));
  nor_4  g09647(.A(new_n10023), .B(new_n10005), .Y(new_n10024));
  nor_4  g09648(.A(new_n10024), .B(new_n10004), .Y(new_n10025));
  nand_4 g09649(.A(new_n10025), .B(new_n9999), .Y(new_n10026));
  nand_4 g09650(.A(new_n10026), .B(new_n9998), .Y(new_n10027));
  nor_4  g09651(.A(new_n10027), .B(new_n9993), .Y(new_n10028));
  not_3  g09652(.A(new_n9851), .Y(new_n10029));
  xnor_3 g09653(.A(new_n10029), .B(new_n9808), .Y(new_n10030));
  xnor_3 g09654(.A(new_n10027), .B(new_n9993), .Y(new_n10031));
  nor_4  g09655(.A(new_n10031), .B(new_n10030), .Y(new_n10032));
  nor_4  g09656(.A(new_n10032), .B(new_n10028), .Y(new_n10033));
  nand_4 g09657(.A(new_n10033), .B(new_n9990), .Y(new_n10034));
  nand_4 g09658(.A(new_n10034), .B(new_n9989), .Y(new_n10035));
  nor_4  g09659(.A(new_n9883), .B(new_n9854), .Y(new_n10036));
  nor_4  g09660(.A(new_n9887), .B(new_n9884), .Y(new_n10037));
  nor_4  g09661(.A(new_n10037), .B(new_n10036), .Y(new_n10038));
  nand_4 g09662(.A(new_n9973), .B(new_n9935), .Y(new_n10039));
  nand_4 g09663(.A(new_n9976), .B(new_n9974), .Y(new_n10040));
  nand_4 g09664(.A(new_n10040), .B(new_n10039), .Y(new_n10041));
  nand_4 g09665(.A(new_n9907), .B(new_n9905), .Y(new_n10042));
  nand_4 g09666(.A(new_n9915), .B(new_n9908), .Y(new_n10043));
  nand_4 g09667(.A(new_n10043), .B(new_n10042), .Y(new_n10044));
  nand_4 g09668(.A(n10848), .B(n9457), .Y(new_n10045));
  nand_4 g09669(.A(n11222), .B(n1906), .Y(new_n10046));
  not_3  g09670(.A(new_n10046), .Y(new_n10047));
  xor_3  g09671(.A(new_n10047), .B(new_n10045), .Y(new_n10048));
  xor_3  g09672(.A(new_n10048), .B(new_n10044), .Y(new_n10049));
  not_3  g09673(.A(new_n9911), .Y(new_n10050));
  nor_4  g09674(.A(new_n9913), .B(new_n10050), .Y(new_n10051));
  nor_4  g09675(.A(new_n9914), .B(new_n9910), .Y(new_n10052));
  nor_4  g09676(.A(new_n10052), .B(new_n10051), .Y(new_n10053));
  nand_4 g09677(.A(n8028), .B(n4817), .Y(new_n10054));
  not_3  g09678(.A(new_n10054), .Y(new_n10055));
  nand_4 g09679(.A(n6578), .B(n1564), .Y(new_n10056));
  nand_4 g09680(.A(n5814), .B(n5314), .Y(new_n10057));
  xor_3  g09681(.A(new_n10057), .B(new_n10056), .Y(new_n10058));
  xor_3  g09682(.A(new_n10058), .B(new_n10055), .Y(new_n10059));
  xnor_3 g09683(.A(new_n10059), .B(new_n10053), .Y(new_n10060));
  not_3  g09684(.A(new_n9899), .Y(new_n10061));
  nor_4  g09685(.A(new_n9901), .B(new_n10061), .Y(new_n10062));
  not_3  g09686(.A(new_n9898), .Y(new_n10063));
  nor_4  g09687(.A(new_n9902), .B(new_n10063), .Y(new_n10064));
  nor_4  g09688(.A(new_n10064), .B(new_n10062), .Y(new_n10065));
  nand_4 g09689(.A(n7294), .B(n5767), .Y(new_n10066));
  nand_4 g09690(.A(n12069), .B(n5694), .Y(new_n10067));
  nand_4 g09691(.A(n11153), .B(n4903), .Y(new_n10068));
  xor_3  g09692(.A(new_n10068), .B(new_n10067), .Y(new_n10069));
  xor_3  g09693(.A(new_n10069), .B(new_n10066), .Y(new_n10070));
  xnor_3 g09694(.A(new_n10070), .B(new_n10065), .Y(new_n10071));
  xnor_3 g09695(.A(new_n10071), .B(new_n10060), .Y(new_n10072));
  xnor_3 g09696(.A(new_n10072), .B(new_n10049), .Y(new_n10073));
  xnor_3 g09697(.A(new_n10073), .B(new_n10041), .Y(new_n10074));
  xnor_3 g09698(.A(new_n10074), .B(new_n10038), .Y(new_n10075));
  not_3  g09699(.A(new_n9476), .Y(new_n10076));
  nand_4 g09700(.A(new_n10076), .B(new_n9417), .Y(new_n10077));
  nand_4 g09701(.A(new_n9477), .B(new_n9440), .Y(new_n10078));
  nand_4 g09702(.A(new_n10078), .B(new_n10077), .Y(new_n10079));
  nand_4 g09703(.A(new_n9923), .B(new_n9921), .Y(new_n10080));
  nand_4 g09704(.A(new_n9925), .B(new_n9917), .Y(new_n10081));
  nand_4 g09705(.A(new_n10081), .B(new_n10080), .Y(new_n10082));
  nand_4 g09706(.A(n5319), .B(n1980), .Y(new_n10083));
  xnor_3 g09707(.A(new_n10083), .B(new_n10082), .Y(new_n10084));
  nand_4 g09708(.A(n12720), .B(n3627), .Y(new_n10085));
  nand_4 g09709(.A(n4516), .B(n2509), .Y(new_n10086));
  xor_3  g09710(.A(new_n10086), .B(new_n10085), .Y(new_n10087));
  nand_4 g09711(.A(new_n9463), .B(new_n9460), .Y(new_n10088));
  and_4  g09712(.A(new_n10088), .B(new_n9466), .Y(new_n10089));
  xnor_3 g09713(.A(new_n10089), .B(new_n10087), .Y(new_n10090));
  nand_4 g09714(.A(n12706), .B(n2564), .Y(new_n10091));
  not_3  g09715(.A(new_n10091), .Y(new_n10092));
  nand_4 g09716(.A(n9920), .B(n2508), .Y(new_n10093));
  nand_4 g09717(.A(n4189), .B(n4005), .Y(new_n10094));
  xor_3  g09718(.A(new_n10094), .B(new_n10093), .Y(new_n10095));
  xnor_3 g09719(.A(new_n10095), .B(new_n10092), .Y(new_n10096));
  xnor_3 g09720(.A(new_n10096), .B(new_n10090), .Y(new_n10097));
  not_3  g09721(.A(new_n9447), .Y(new_n10098));
  nor_4  g09722(.A(new_n9449), .B(new_n10098), .Y(new_n10099));
  not_3  g09723(.A(new_n9446), .Y(new_n10100));
  nor_4  g09724(.A(new_n9450), .B(new_n10100), .Y(new_n10101));
  nor_4  g09725(.A(new_n10101), .B(new_n10099), .Y(new_n10102));
  or_4   g09726(.A(new_n9456), .B(new_n9454), .Y(new_n10103));
  nand_4 g09727(.A(new_n9468), .B(new_n9457_1), .Y(new_n10104));
  nand_4 g09728(.A(new_n10104), .B(new_n10103), .Y(new_n10105));
  xnor_3 g09729(.A(new_n10105), .B(new_n10102), .Y(new_n10106));
  xnor_3 g09730(.A(new_n10106), .B(new_n10097), .Y(new_n10107));
  xnor_3 g09731(.A(new_n10107), .B(new_n10084), .Y(new_n10108));
  nand_4 g09732(.A(new_n9473), .B(new_n9472), .Y(new_n10109));
  nand_4 g09733(.A(new_n9475), .B(new_n9470), .Y(new_n10110));
  nand_4 g09734(.A(new_n10110), .B(new_n10109), .Y(new_n10111));
  nand_4 g09735(.A(new_n9451), .B(new_n9445), .Y(new_n10112));
  nand_4 g09736(.A(new_n9469), .B(new_n9453), .Y(new_n10113));
  nand_4 g09737(.A(new_n10113), .B(new_n10112), .Y(new_n10114));
  nand_4 g09738(.A(n6770), .B(n2585), .Y(new_n10115));
  nand_4 g09739(.A(new_n9951), .B(new_n9948), .Y(new_n10116));
  and_4  g09740(.A(new_n10116), .B(new_n9954), .Y(new_n10117));
  nand_4 g09741(.A(n6687), .B(n615), .Y(new_n10118));
  nand_4 g09742(.A(n6038), .B(n2087), .Y(new_n10119));
  xor_3  g09743(.A(new_n10119), .B(new_n10118), .Y(new_n10120));
  xnor_3 g09744(.A(new_n10120), .B(new_n10117), .Y(new_n10121));
  xnor_3 g09745(.A(new_n10121), .B(new_n10115), .Y(new_n10122));
  xnor_3 g09746(.A(new_n10122), .B(new_n10114), .Y(new_n10123));
  xnor_3 g09747(.A(new_n10123), .B(new_n10111), .Y(new_n10124));
  xnor_3 g09748(.A(new_n10124), .B(new_n10108), .Y(new_n10125));
  nand_4 g09749(.A(new_n9940), .B(new_n9938_1), .Y(new_n10126));
  not_3  g09750(.A(new_n9972), .Y(new_n10127));
  nand_4 g09751(.A(new_n10127), .B(new_n9942), .Y(new_n10128));
  nand_4 g09752(.A(new_n10128), .B(new_n10126), .Y(new_n10129));
  not_3  g09753(.A(new_n9964), .Y(new_n10130));
  nand_4 g09754(.A(new_n9970), .B(new_n10130), .Y(new_n10131));
  not_3  g09755(.A(new_n9961), .Y(new_n10132));
  nand_4 g09756(.A(new_n9971), .B(new_n10132), .Y(new_n10133));
  nand_4 g09757(.A(new_n10133), .B(new_n10131), .Y(new_n10134));
  nand_4 g09758(.A(new_n9945), .B(new_n9943), .Y(new_n10135));
  not_3  g09759(.A(new_n9960), .Y(new_n10136));
  nand_4 g09760(.A(new_n10136), .B(new_n10135), .Y(new_n10137));
  nand_4 g09761(.A(n12391), .B(n12044), .Y(new_n10138));
  nand_4 g09762(.A(n1512), .B(n1199), .Y(new_n10139));
  nand_4 g09763(.A(n7160), .B(n6806), .Y(new_n10140));
  xor_3  g09764(.A(new_n10140), .B(new_n10139), .Y(new_n10141));
  nand_4 g09765(.A(n2515), .B(n533), .Y(new_n10142));
  nand_4 g09766(.A(n4828), .B(n2802), .Y(new_n10143));
  xor_3  g09767(.A(new_n10143), .B(new_n10142), .Y(new_n10144));
  xnor_3 g09768(.A(new_n10144), .B(new_n10141), .Y(new_n10145));
  xnor_3 g09769(.A(new_n10145), .B(new_n10138), .Y(new_n10146));
  nand_4 g09770(.A(n7891), .B(n5069), .Y(new_n10147));
  not_3  g09771(.A(new_n10147), .Y(new_n10148));
  not_3  g09772(.A(new_n9966), .Y(new_n10149));
  nor_4  g09773(.A(new_n9968), .B(new_n10149), .Y(new_n10150));
  not_3  g09774(.A(new_n9965), .Y(new_n10151));
  nor_4  g09775(.A(new_n9969), .B(new_n10151), .Y(new_n10152));
  nor_4  g09776(.A(new_n10152), .B(new_n10150), .Y(new_n10153));
  xnor_3 g09777(.A(new_n10153), .B(new_n10148), .Y(new_n10154));
  xnor_3 g09778(.A(new_n10154), .B(new_n10146), .Y(new_n10155));
  xnor_3 g09779(.A(new_n10155), .B(new_n10137), .Y(new_n10156));
  xnor_3 g09780(.A(new_n10156), .B(new_n10134), .Y(new_n10157));
  xnor_3 g09781(.A(new_n10157), .B(new_n10129), .Y(new_n10158));
  xnor_3 g09782(.A(new_n10158), .B(new_n10125), .Y(new_n10159));
  xnor_3 g09783(.A(new_n10159), .B(new_n10079), .Y(new_n10160));
  xnor_3 g09784(.A(new_n10160), .B(new_n10075), .Y(new_n10161));
  not_3  g09785(.A(new_n9979), .Y(new_n10162));
  nand_4 g09786(.A(new_n10162), .B(new_n9977), .Y(new_n10163));
  nand_4 g09787(.A(new_n9980), .B(new_n9934), .Y(new_n10164));
  nand_4 g09788(.A(new_n10164), .B(new_n10163), .Y(new_n10165));
  nand_4 g09789(.A(new_n9926), .B(new_n9892), .Y(new_n10166));
  nand_4 g09790(.A(new_n9933), .B(new_n9927), .Y(new_n10167));
  nand_4 g09791(.A(new_n10167), .B(new_n10166), .Y(new_n10168));
  nand_4 g09792(.A(new_n9864), .B(new_n9857), .Y(new_n10169));
  not_3  g09793(.A(new_n9865), .Y(new_n10170));
  not_3  g09794(.A(new_n9876), .Y(new_n10171));
  nand_4 g09795(.A(new_n10171), .B(new_n10170), .Y(new_n10172));
  nand_4 g09796(.A(new_n10172), .B(new_n10169), .Y(new_n10173));
  xnor_3 g09797(.A(new_n10173), .B(new_n10168), .Y(new_n10174_1));
  nand_4 g09798(.A(new_n9880), .B(new_n9879), .Y(new_n10175));
  nand_4 g09799(.A(new_n9882), .B(new_n9877), .Y(new_n10176));
  nand_4 g09800(.A(new_n10176), .B(new_n10175), .Y(new_n10177));
  nand_4 g09801(.A(n7500), .B(n7320), .Y(new_n10178));
  nand_4 g09802(.A(n7523), .B(n7354), .Y(new_n10179));
  xor_3  g09803(.A(new_n10179), .B(new_n10178), .Y(new_n10180));
  nand_4 g09804(.A(n4141), .B(n2226), .Y(new_n10181));
  nand_4 g09805(.A(n8336), .B(n783), .Y(new_n10182));
  not_3  g09806(.A(new_n10182), .Y(new_n10183));
  xor_3  g09807(.A(new_n10183), .B(new_n10181), .Y(new_n10184));
  xor_3  g09808(.A(new_n10184), .B(new_n10180), .Y(new_n10185));
  nor_4  g09809(.A(new_n9868), .B(new_n9867), .Y(new_n10186));
  not_3  g09810(.A(new_n9869), .Y(new_n10187));
  nor_4  g09811(.A(new_n9875), .B(new_n10187), .Y(new_n10188));
  nor_4  g09812(.A(new_n10188), .B(new_n10186), .Y(new_n10189));
  nand_4 g09813(.A(n12704), .B(n996), .Y(new_n10190));
  not_3  g09814(.A(new_n10190), .Y(new_n10191));
  not_3  g09815(.A(new_n9871), .Y(new_n10192));
  nor_4  g09816(.A(new_n9873), .B(new_n10192), .Y(new_n10193));
  not_3  g09817(.A(new_n9870), .Y(new_n10194));
  nor_4  g09818(.A(new_n9874), .B(new_n10194), .Y(new_n10195));
  nor_4  g09819(.A(new_n10195), .B(new_n10193), .Y(new_n10196));
  nand_4 g09820(.A(n6986), .B(n4928), .Y(new_n10197));
  nand_4 g09821(.A(n10678), .B(n1209), .Y(new_n10198));
  xor_3  g09822(.A(new_n10198), .B(new_n10197), .Y(new_n10199));
  nand_4 g09823(.A(n10928), .B(n8236), .Y(new_n10200));
  nand_4 g09824(.A(n5105), .B(n1094), .Y(new_n10201));
  xor_3  g09825(.A(new_n10201), .B(new_n10200), .Y(new_n10202));
  xnor_3 g09826(.A(new_n10202), .B(new_n10199), .Y(new_n10203));
  xnor_3 g09827(.A(new_n10203), .B(new_n10196), .Y(new_n10204));
  xnor_3 g09828(.A(new_n10204), .B(new_n10191), .Y(new_n10205));
  xnor_3 g09829(.A(new_n10205), .B(new_n10189), .Y(new_n10206));
  xnor_3 g09830(.A(new_n10206), .B(new_n10185), .Y(new_n10207));
  nand_4 g09831(.A(new_n9903), .B(new_n9896), .Y(new_n10208));
  nand_4 g09832(.A(new_n9916), .B(new_n9904), .Y(new_n10209));
  nand_4 g09833(.A(new_n10209), .B(new_n10208), .Y(new_n10210));
  and_4  g09834(.A(new_n9860), .B(new_n9859), .Y(new_n10211));
  not_3  g09835(.A(new_n9858), .Y(new_n10212));
  nor_4  g09836(.A(new_n9862), .B(new_n10212), .Y(new_n10213));
  or_4   g09837(.A(new_n10213), .B(new_n10211), .Y(new_n10214));
  xnor_3 g09838(.A(new_n10214), .B(new_n10210), .Y(new_n10215));
  xnor_3 g09839(.A(new_n10215), .B(new_n10207), .Y(new_n10216));
  xnor_3 g09840(.A(new_n10216), .B(new_n10177), .Y(new_n10217_1));
  xnor_3 g09841(.A(new_n10217_1), .B(new_n10174_1), .Y(new_n10218));
  xnor_3 g09842(.A(new_n10218), .B(new_n10165), .Y(new_n10219));
  xnor_3 g09843(.A(new_n10219), .B(new_n10161), .Y(new_n10220));
  nand_4 g09844(.A(new_n9982), .B(new_n9853), .Y(new_n10221));
  nand_4 g09845(.A(new_n10221), .B(new_n9985), .Y(new_n10222));
  xnor_3 g09846(.A(new_n10222), .B(new_n10220), .Y(new_n10223_1));
  xnor_3 g09847(.A(new_n10223_1), .B(new_n10035), .Y(n3654));
  xnor_3 g09848(.A(new_n10031), .B(new_n10030), .Y(n3661));
  nor_4  g09849(.A(new_n6538), .B(new_n6537), .Y(new_n10226));
  not_3  g09850(.A(new_n10226), .Y(new_n10227));
  nand_4 g09851(.A(n1798), .B(n1097), .Y(new_n10228));
  nand_4 g09852(.A(n12591), .B(n5305), .Y(new_n10229));
  nand_4 g09853(.A(new_n10229), .B(new_n10228), .Y(new_n10230));
  not_3  g09854(.A(new_n10230), .Y(new_n10231));
  not_3  g09855(.A(new_n10228), .Y(new_n10232));
  not_3  g09856(.A(new_n10229), .Y(new_n10233));
  nand_4 g09857(.A(new_n10233), .B(new_n10232), .Y(new_n10234));
  not_3  g09858(.A(new_n10234), .Y(new_n10235));
  nor_4  g09859(.A(new_n10235), .B(new_n10231), .Y(new_n10236));
  nor_4  g09860(.A(new_n10236), .B(new_n10227), .Y(new_n10237));
  nand_4 g09861(.A(n7456), .B(n5305), .Y(new_n10238));
  nand_4 g09862(.A(n5964), .B(n3932), .Y(new_n10239));
  not_3  g09863(.A(new_n10239), .Y(new_n10240));
  nand_4 g09864(.A(new_n10240), .B(new_n10230), .Y(new_n10241));
  nand_4 g09865(.A(new_n10241), .B(new_n10234), .Y(new_n10242));
  xor_3  g09866(.A(new_n10242), .B(new_n10238), .Y(new_n10243));
  nand_4 g09867(.A(n3932), .B(n1097), .Y(new_n10244));
  not_3  g09868(.A(new_n10244), .Y(new_n10245));
  nand_4 g09869(.A(n4312), .B(n1798), .Y(new_n10246));
  nand_4 g09870(.A(n12591), .B(n5964), .Y(new_n10247));
  xnor_3 g09871(.A(new_n10247), .B(new_n10246), .Y(new_n10248));
  xor_3  g09872(.A(new_n10248), .B(new_n10245), .Y(new_n10249));
  nor_4  g09873(.A(new_n10249), .B(new_n10243), .Y(new_n10250));
  not_3  g09874(.A(new_n10238), .Y(new_n10251));
  xor_3  g09875(.A(new_n10242), .B(new_n10251), .Y(new_n10252));
  xor_3  g09876(.A(new_n10248), .B(new_n10244), .Y(new_n10253));
  nor_4  g09877(.A(new_n10253), .B(new_n10252), .Y(new_n10254));
  nor_4  g09878(.A(new_n10254), .B(new_n10250), .Y(new_n10255));
  nand_4 g09879(.A(new_n10255), .B(new_n10237), .Y(new_n10256));
  nand_4 g09880(.A(n11662), .B(n5305), .Y(new_n10257));
  nand_4 g09881(.A(n7456), .B(n5964), .Y(new_n10258));
  nand_4 g09882(.A(n4312), .B(n3932), .Y(new_n10259));
  nand_4 g09883(.A(n12591), .B(n1097), .Y(new_n10260));
  nand_4 g09884(.A(n12705), .B(n1798), .Y(new_n10261));
  xnor_3 g09885(.A(new_n10261), .B(new_n10260), .Y(new_n10262));
  not_3  g09886(.A(new_n10262), .Y(new_n10263));
  nor_4  g09887(.A(new_n10263), .B(new_n10259), .Y(new_n10264));
  not_3  g09888(.A(new_n10259), .Y(new_n10265));
  nor_4  g09889(.A(new_n10262), .B(new_n10265), .Y(new_n10266));
  nor_4  g09890(.A(new_n10266), .B(new_n10264), .Y(new_n10267));
  xnor_3 g09891(.A(new_n10267), .B(new_n10258), .Y(new_n10268));
  and_4  g09892(.A(new_n10247), .B(new_n10246), .Y(new_n10269));
  nor_4  g09893(.A(new_n10248), .B(new_n10245), .Y(new_n10270));
  nor_4  g09894(.A(new_n10270), .B(new_n10269), .Y(new_n10271));
  xnor_3 g09895(.A(new_n10271), .B(new_n10268), .Y(new_n10272));
  not_3  g09896(.A(new_n10272), .Y(new_n10273));
  nor_4  g09897(.A(new_n10273), .B(new_n10257), .Y(new_n10274));
  not_3  g09898(.A(new_n10257), .Y(new_n10275));
  nor_4  g09899(.A(new_n10272), .B(new_n10275), .Y(new_n10276));
  nor_4  g09900(.A(new_n10276), .B(new_n10274), .Y(new_n10277));
  not_3  g09901(.A(new_n10242), .Y(new_n10278_1));
  nor_4  g09902(.A(new_n10278_1), .B(new_n10238), .Y(new_n10279));
  not_3  g09903(.A(new_n10279), .Y(new_n10280));
  nand_4 g09904(.A(new_n10253), .B(new_n10252), .Y(new_n10281));
  nand_4 g09905(.A(new_n10281), .B(new_n10280), .Y(new_n10282));
  xnor_3 g09906(.A(new_n10282), .B(new_n10277), .Y(new_n10283));
  xor_3  g09907(.A(new_n10283), .B(new_n10256), .Y(new_n10284));
  not_3  g09908(.A(new_n10255), .Y(new_n10285));
  xor_3  g09909(.A(new_n10285), .B(new_n10237), .Y(new_n10286));
  not_3  g09910(.A(new_n10286), .Y(new_n10287));
  nand_4 g09911(.A(n11023), .B(n8759), .Y(new_n10288));
  not_3  g09912(.A(new_n10288), .Y(new_n10289));
  nand_4 g09913(.A(n8759), .B(n3022), .Y(new_n10290));
  nand_4 g09914(.A(n12299), .B(n6703), .Y(new_n10291));
  nand_4 g09915(.A(new_n10291), .B(new_n10290), .Y(new_n10292));
  nand_4 g09916(.A(n9640), .B(n6776), .Y(new_n10293));
  not_3  g09917(.A(new_n10293), .Y(new_n10294));
  nand_4 g09918(.A(new_n10294), .B(new_n10292), .Y(new_n10295));
  not_3  g09919(.A(new_n10290), .Y(new_n10296));
  not_3  g09920(.A(new_n10291), .Y(new_n10297));
  nand_4 g09921(.A(new_n10297), .B(new_n10296), .Y(new_n10298));
  nand_4 g09922(.A(new_n10298), .B(new_n10295), .Y(new_n10299));
  xor_3  g09923(.A(new_n10299), .B(new_n10289), .Y(new_n10300));
  nand_4 g09924(.A(n12299), .B(n9640), .Y(new_n10301));
  not_3  g09925(.A(new_n10301), .Y(new_n10302));
  nand_4 g09926(.A(n6776), .B(n3022), .Y(new_n10303));
  not_3  g09927(.A(new_n10303), .Y(new_n10304));
  nand_4 g09928(.A(n7436), .B(n6703), .Y(new_n10305));
  not_3  g09929(.A(new_n10305), .Y(new_n10306));
  nor_4  g09930(.A(new_n10306), .B(new_n10304), .Y(new_n10307));
  nor_4  g09931(.A(new_n10305), .B(new_n10303), .Y(new_n10308));
  nor_4  g09932(.A(new_n10308), .B(new_n10307), .Y(new_n10309));
  xor_3  g09933(.A(new_n10309), .B(new_n10302), .Y(new_n10310));
  xnor_3 g09934(.A(new_n10310), .B(new_n10300), .Y(new_n10311));
  nor_4  g09935(.A(new_n10293), .B(new_n6530), .Y(new_n10312));
  and_4  g09936(.A(new_n10298), .B(new_n10292), .Y(new_n10313));
  nor_4  g09937(.A(new_n10313), .B(new_n10312), .Y(new_n10314));
  not_3  g09938(.A(new_n10314), .Y(new_n10315));
  nor_4  g09939(.A(new_n10315), .B(new_n10293), .Y(new_n10316));
  not_3  g09940(.A(new_n10316), .Y(new_n10317));
  xnor_3 g09941(.A(new_n10317), .B(new_n10311), .Y(new_n10318));
  nor_4  g09942(.A(new_n6556), .B(new_n6555), .Y(new_n10319));
  not_3  g09943(.A(new_n10319), .Y(new_n10320));
  nand_4 g09944(.A(n5645), .B(n2530), .Y(new_n10321));
  not_3  g09945(.A(new_n10321), .Y(new_n10322));
  nand_4 g09946(.A(n8665), .B(n5331), .Y(new_n10323));
  not_3  g09947(.A(new_n10323), .Y(new_n10324));
  nor_4  g09948(.A(new_n10324), .B(new_n10322), .Y(new_n10325));
  nor_4  g09949(.A(new_n10323), .B(new_n10321), .Y(new_n10326));
  nor_4  g09950(.A(new_n10326), .B(new_n10325), .Y(new_n10327_1));
  nor_4  g09951(.A(new_n10327_1), .B(new_n10320), .Y(new_n10328));
  not_3  g09952(.A(new_n10328), .Y(new_n10329));
  nand_4 g09953(.A(n11922), .B(n5331), .Y(new_n10330));
  nand_4 g09954(.A(n2530), .B(n1067), .Y(new_n10331));
  nand_4 g09955(.A(n8665), .B(n8476), .Y(new_n10332));
  not_3  g09956(.A(new_n10332), .Y(new_n10333));
  nand_4 g09957(.A(n12648), .B(n5645), .Y(new_n10334));
  not_3  g09958(.A(new_n10334), .Y(new_n10335));
  nor_4  g09959(.A(new_n10335), .B(new_n10333), .Y(new_n10336));
  nor_4  g09960(.A(new_n10334), .B(new_n10332), .Y(new_n10337));
  nor_4  g09961(.A(new_n10337), .B(new_n10336), .Y(new_n10338));
  xnor_3 g09962(.A(new_n10338), .B(new_n10331), .Y(new_n10339));
  not_3  g09963(.A(new_n10339), .Y(new_n10340));
  xnor_3 g09964(.A(new_n10340), .B(new_n10330), .Y(new_n10341));
  not_3  g09965(.A(new_n10325), .Y(new_n10342));
  nand_4 g09966(.A(n8476), .B(n1067), .Y(new_n10343));
  not_3  g09967(.A(new_n10343), .Y(new_n10344));
  nand_4 g09968(.A(new_n10344), .B(new_n10342), .Y(new_n10345));
  not_3  g09969(.A(new_n10345), .Y(new_n10346));
  nor_4  g09970(.A(new_n10346), .B(new_n10326), .Y(new_n10347));
  xnor_3 g09971(.A(new_n10347), .B(new_n10341), .Y(new_n10348));
  xnor_3 g09972(.A(new_n10348), .B(new_n10329), .Y(new_n10349));
  not_3  g09973(.A(new_n10349), .Y(new_n10350));
  nand_4 g09974(.A(n7965), .B(n2749), .Y(new_n10351));
  nand_4 g09975(.A(n7965), .B(n3754), .Y(new_n10352));
  nand_4 g09976(.A(n11892), .B(n11876), .Y(new_n10353));
  nor_4  g09977(.A(new_n10353), .B(new_n10352), .Y(new_n10354));
  not_3  g09978(.A(new_n10354), .Y(new_n10355));
  nand_4 g09979(.A(new_n10353), .B(new_n10352), .Y(new_n10356));
  nand_4 g09980(.A(n10898), .B(n7388), .Y(new_n10357));
  not_3  g09981(.A(new_n10357), .Y(new_n10358));
  nand_4 g09982(.A(new_n10358), .B(new_n10356), .Y(new_n10359));
  nand_4 g09983(.A(new_n10359), .B(new_n10355), .Y(new_n10360));
  not_3  g09984(.A(new_n10360), .Y(new_n10361));
  nor_4  g09985(.A(new_n10361), .B(new_n10351), .Y(new_n10362));
  not_3  g09986(.A(new_n10351), .Y(new_n10363));
  nor_4  g09987(.A(new_n10360), .B(new_n10363), .Y(new_n10364));
  nor_4  g09988(.A(new_n10364), .B(new_n10362), .Y(new_n10365));
  nand_4 g09989(.A(n11892), .B(n10898), .Y(new_n10366));
  nand_4 g09990(.A(n7388), .B(n3754), .Y(new_n10367));
  nand_4 g09991(.A(n11876), .B(n2393), .Y(new_n10368));
  xnor_3 g09992(.A(new_n10368), .B(new_n10367), .Y(new_n10369));
  xnor_3 g09993(.A(new_n10369), .B(new_n10366), .Y(new_n10370));
  not_3  g09994(.A(new_n10370), .Y(new_n10371));
  xnor_3 g09995(.A(new_n10371), .B(new_n10365), .Y(new_n10372));
  not_3  g09996(.A(new_n6532), .Y(new_n10373));
  nor_4  g09997(.A(new_n10357), .B(new_n10373), .Y(new_n10374));
  nand_4 g09998(.A(new_n10356), .B(new_n10355), .Y(new_n10375));
  not_3  g09999(.A(new_n10375), .Y(new_n10376));
  nor_4  g10000(.A(new_n10376), .B(new_n10374), .Y(new_n10377));
  not_3  g10001(.A(new_n10377), .Y(new_n10378));
  nor_4  g10002(.A(new_n10378), .B(new_n10357), .Y(new_n10379));
  not_3  g10003(.A(new_n10379), .Y(new_n10380));
  xnor_3 g10004(.A(new_n10380), .B(new_n10372), .Y(new_n10381));
  not_3  g10005(.A(new_n10381), .Y(new_n10382));
  nor_4  g10006(.A(new_n10382), .B(new_n10350), .Y(new_n10383));
  nor_4  g10007(.A(new_n10381), .B(new_n10349), .Y(new_n10384));
  nor_4  g10008(.A(new_n10384), .B(new_n10383), .Y(new_n10385));
  not_3  g10009(.A(new_n10385), .Y(new_n10386));
  not_3  g10010(.A(new_n6551), .Y(new_n10387));
  nand_4 g10011(.A(new_n6557), .B(new_n6554), .Y(new_n10388));
  nand_4 g10012(.A(new_n10388), .B(new_n10387), .Y(new_n10389));
  nand_4 g10013(.A(new_n10374), .B(new_n10356), .Y(new_n10390));
  nand_4 g10014(.A(new_n10390), .B(new_n10378), .Y(new_n10391_1));
  not_3  g10015(.A(new_n10391_1), .Y(new_n10392));
  nor_4  g10016(.A(new_n10392), .B(new_n10389), .Y(new_n10393));
  xnor_3 g10017(.A(new_n10392), .B(new_n10389), .Y(new_n10394));
  not_3  g10018(.A(new_n6531), .Y(new_n10395));
  nor_4  g10019(.A(new_n10343), .B(new_n10395), .Y(new_n10396));
  not_3  g10020(.A(new_n10396), .Y(new_n10397));
  nor_4  g10021(.A(new_n10397), .B(new_n10342), .Y(new_n10398));
  not_3  g10022(.A(new_n10327_1), .Y(new_n10399));
  nor_4  g10023(.A(new_n10396), .B(new_n10399), .Y(new_n10400));
  nor_4  g10024(.A(new_n10400), .B(new_n10398), .Y(new_n10401));
  not_3  g10025(.A(new_n10401), .Y(new_n10402));
  nor_4  g10026(.A(new_n10402), .B(new_n10394), .Y(new_n10403));
  nor_4  g10027(.A(new_n10403), .B(new_n10393), .Y(new_n10404));
  xnor_3 g10028(.A(new_n10404), .B(new_n10386), .Y(new_n10405));
  not_3  g10029(.A(new_n10405), .Y(new_n10406));
  nor_4  g10030(.A(new_n10406), .B(new_n10318), .Y(new_n10407));
  not_3  g10031(.A(new_n10318), .Y(new_n10408));
  nor_4  g10032(.A(new_n10405), .B(new_n10408), .Y(new_n10409));
  nor_4  g10033(.A(new_n10409), .B(new_n10407), .Y(new_n10410));
  nand_4 g10034(.A(new_n6544), .B(new_n6541), .Y(new_n10411));
  not_3  g10035(.A(new_n10411), .Y(new_n10412));
  nor_4  g10036(.A(new_n6559), .B(new_n10412), .Y(new_n10413));
  not_3  g10037(.A(new_n10413), .Y(new_n10414));
  nor_4  g10038(.A(new_n10295), .B(new_n6530), .Y(new_n10415));
  nor_4  g10039(.A(new_n10415), .B(new_n10314), .Y(new_n10416));
  nor_4  g10040(.A(new_n10416), .B(new_n10414), .Y(new_n10417));
  not_3  g10041(.A(new_n10417), .Y(new_n10418));
  not_3  g10042(.A(new_n10394), .Y(new_n10419));
  xor_3  g10043(.A(new_n10401), .B(new_n10419), .Y(new_n10420));
  not_3  g10044(.A(new_n10416), .Y(new_n10421));
  nor_4  g10045(.A(new_n10421), .B(new_n10413), .Y(new_n10422));
  nor_4  g10046(.A(new_n10422), .B(new_n10417), .Y(new_n10423));
  nand_4 g10047(.A(new_n10423), .B(new_n10420), .Y(new_n10424));
  nand_4 g10048(.A(new_n10424), .B(new_n10418), .Y(new_n10425));
  xnor_3 g10049(.A(new_n10425), .B(new_n10410), .Y(new_n10426));
  nand_4 g10050(.A(new_n10426), .B(new_n10287), .Y(new_n10427));
  not_3  g10051(.A(new_n10427), .Y(new_n10428));
  nor_4  g10052(.A(new_n10426), .B(new_n10287), .Y(new_n10429));
  nor_4  g10053(.A(new_n10429), .B(new_n10428), .Y(new_n10430));
  xor_3  g10054(.A(new_n10402), .B(new_n10419), .Y(new_n10431));
  not_3  g10055(.A(new_n10423), .Y(new_n10432));
  xnor_3 g10056(.A(new_n10432), .B(new_n10431), .Y(new_n10433));
  not_3  g10057(.A(new_n6528), .Y(new_n10434));
  nor_4  g10058(.A(new_n10239), .B(new_n10434), .Y(new_n10435));
  not_3  g10059(.A(new_n10435), .Y(new_n10436));
  nor_4  g10060(.A(new_n10436), .B(new_n10230), .Y(new_n10437));
  not_3  g10061(.A(new_n10236), .Y(new_n10438));
  nor_4  g10062(.A(new_n10435), .B(new_n10438), .Y(new_n10439_1));
  nor_4  g10063(.A(new_n10439_1), .B(new_n10437), .Y(new_n10440));
  not_3  g10064(.A(new_n10440), .Y(new_n10441));
  nor_4  g10065(.A(new_n10441), .B(new_n10433), .Y(new_n10442));
  nand_4 g10066(.A(new_n6539), .B(new_n6536), .Y(new_n10443));
  nand_4 g10067(.A(new_n6561), .B(new_n6540), .Y(new_n10444));
  nand_4 g10068(.A(new_n10444), .B(new_n10443), .Y(new_n10445));
  xnor_3 g10069(.A(new_n10441), .B(new_n10433), .Y(new_n10446));
  nor_4  g10070(.A(new_n10446), .B(new_n10445), .Y(new_n10447));
  nor_4  g10071(.A(new_n10447), .B(new_n10442), .Y(new_n10448));
  nand_4 g10072(.A(new_n10448), .B(new_n10430), .Y(new_n10449));
  nand_4 g10073(.A(new_n10449), .B(new_n10427), .Y(new_n10450));
  xnor_3 g10074(.A(new_n10450), .B(new_n10284), .Y(new_n10451_1));
  nor_4  g10075(.A(new_n10317), .B(new_n10311), .Y(new_n10452));
  nand_4 g10076(.A(n10451), .B(n8759), .Y(new_n10453));
  nand_4 g10077(.A(n11023), .B(n6776), .Y(new_n10454));
  not_3  g10078(.A(new_n10454), .Y(new_n10455));
  nor_4  g10079(.A(new_n10308), .B(new_n10302), .Y(new_n10456));
  nor_4  g10080(.A(new_n10456), .B(new_n10307), .Y(new_n10457));
  xnor_3 g10081(.A(new_n10457), .B(new_n10455), .Y(new_n10458));
  nand_4 g10082(.A(n9640), .B(n7436), .Y(new_n10459));
  nand_4 g10083(.A(n12299), .B(n3022), .Y(new_n10460));
  not_3  g10084(.A(new_n10460), .Y(new_n10461));
  nand_4 g10085(.A(n8276), .B(n6703), .Y(new_n10462));
  not_3  g10086(.A(new_n10462), .Y(new_n10463));
  nor_4  g10087(.A(new_n10463), .B(new_n10461), .Y(new_n10464));
  not_3  g10088(.A(new_n10464), .Y(new_n10465));
  nor_4  g10089(.A(new_n10462), .B(new_n10460), .Y(new_n10466));
  not_3  g10090(.A(new_n10466), .Y(new_n10467));
  nand_4 g10091(.A(new_n10467), .B(new_n10465), .Y(new_n10468));
  xnor_3 g10092(.A(new_n10468), .B(new_n10459), .Y(new_n10469));
  xnor_3 g10093(.A(new_n10469), .B(new_n10458), .Y(new_n10470));
  nor_4  g10094(.A(new_n10470), .B(new_n10453), .Y(new_n10471));
  not_3  g10095(.A(new_n10453), .Y(new_n10472));
  not_3  g10096(.A(new_n10470), .Y(new_n10473));
  nor_4  g10097(.A(new_n10473), .B(new_n10472), .Y(new_n10474));
  nor_4  g10098(.A(new_n10474), .B(new_n10471), .Y(new_n10475));
  not_3  g10099(.A(new_n10475), .Y(new_n10476_1));
  not_3  g10100(.A(new_n10299), .Y(new_n10477));
  nor_4  g10101(.A(new_n10477), .B(new_n10288), .Y(new_n10478));
  not_3  g10102(.A(new_n10478), .Y(new_n10479));
  nand_4 g10103(.A(new_n10310), .B(new_n10300), .Y(new_n10480));
  nand_4 g10104(.A(new_n10480), .B(new_n10479), .Y(new_n10481));
  xnor_3 g10105(.A(new_n10481), .B(new_n10476_1), .Y(new_n10482));
  xnor_3 g10106(.A(new_n10482), .B(new_n10452), .Y(new_n10483));
  not_3  g10107(.A(new_n10483), .Y(new_n10484));
  nor_4  g10108(.A(new_n10380), .B(new_n10372), .Y(new_n10485));
  nand_4 g10109(.A(n7965), .B(n159), .Y(new_n10486));
  not_3  g10110(.A(new_n10362), .Y(new_n10487));
  nand_4 g10111(.A(new_n10371), .B(new_n10365), .Y(new_n10488));
  nand_4 g10112(.A(new_n10488), .B(new_n10487), .Y(new_n10489));
  not_3  g10113(.A(new_n10489), .Y(new_n10490));
  xnor_3 g10114(.A(new_n10490), .B(new_n10486), .Y(new_n10491));
  nand_4 g10115(.A(n7388), .B(n2749), .Y(new_n10492));
  not_3  g10116(.A(new_n10492), .Y(new_n10493));
  not_3  g10117(.A(new_n10367), .Y(new_n10494));
  not_3  g10118(.A(new_n10368), .Y(new_n10495));
  nor_4  g10119(.A(new_n10495), .B(new_n10494), .Y(new_n10496));
  not_3  g10120(.A(new_n10366), .Y(new_n10497));
  nor_4  g10121(.A(new_n10369), .B(new_n10497), .Y(new_n10498));
  nor_4  g10122(.A(new_n10498), .B(new_n10496), .Y(new_n10499));
  nand_4 g10123(.A(new_n10499), .B(new_n10493), .Y(new_n10500));
  not_3  g10124(.A(new_n10500), .Y(new_n10501));
  nor_4  g10125(.A(new_n10499), .B(new_n10493), .Y(new_n10502));
  nor_4  g10126(.A(new_n10502), .B(new_n10501), .Y(new_n10503));
  nand_4 g10127(.A(n11892), .B(n3754), .Y(new_n10504));
  not_3  g10128(.A(new_n10504), .Y(new_n10505));
  nand_4 g10129(.A(n11876), .B(n5860), .Y(new_n10506));
  nand_4 g10130(.A(n10898), .B(n2393), .Y(new_n10507));
  xnor_3 g10131(.A(new_n10507), .B(new_n10506), .Y(new_n10508));
  xnor_3 g10132(.A(new_n10508), .B(new_n10505), .Y(new_n10509));
  xnor_3 g10133(.A(new_n10509), .B(new_n10503), .Y(new_n10510_1));
  xnor_3 g10134(.A(new_n10510_1), .B(new_n10491), .Y(new_n10511));
  xnor_3 g10135(.A(new_n10511), .B(new_n10485), .Y(new_n10512));
  nor_4  g10136(.A(new_n10348), .B(new_n10329), .Y(new_n10513));
  nand_4 g10137(.A(n5331), .B(n2551), .Y(new_n10514));
  nand_4 g10138(.A(n11922), .B(n8476), .Y(new_n10515));
  not_3  g10139(.A(new_n10515), .Y(new_n10516));
  not_3  g10140(.A(new_n10331), .Y(new_n10517));
  nor_4  g10141(.A(new_n10337), .B(new_n10517), .Y(new_n10518));
  nor_4  g10142(.A(new_n10518), .B(new_n10336), .Y(new_n10519));
  xnor_3 g10143(.A(new_n10519), .B(new_n10516), .Y(new_n10520));
  nand_4 g10144(.A(n12648), .B(n1067), .Y(new_n10521));
  not_3  g10145(.A(new_n10521), .Y(new_n10522));
  nand_4 g10146(.A(n8665), .B(n2530), .Y(new_n10523));
  not_3  g10147(.A(new_n10523), .Y(new_n10524));
  nand_4 g10148(.A(n10545), .B(n5645), .Y(new_n10525));
  not_3  g10149(.A(new_n10525), .Y(new_n10526));
  nor_4  g10150(.A(new_n10526), .B(new_n10524), .Y(new_n10527));
  not_3  g10151(.A(new_n10527), .Y(new_n10528));
  nor_4  g10152(.A(new_n10525), .B(new_n10523), .Y(new_n10529));
  not_3  g10153(.A(new_n10529), .Y(new_n10530));
  nand_4 g10154(.A(new_n10530), .B(new_n10528), .Y(new_n10531));
  xnor_3 g10155(.A(new_n10531), .B(new_n10522), .Y(new_n10532));
  xnor_3 g10156(.A(new_n10532), .B(new_n10520), .Y(new_n10533));
  not_3  g10157(.A(new_n10533), .Y(new_n10534));
  nor_4  g10158(.A(new_n10534), .B(new_n10514), .Y(new_n10535));
  not_3  g10159(.A(new_n10514), .Y(new_n10536));
  nor_4  g10160(.A(new_n10533), .B(new_n10536), .Y(new_n10537));
  nor_4  g10161(.A(new_n10537), .B(new_n10535), .Y(new_n10538));
  nor_4  g10162(.A(new_n10340), .B(new_n10330), .Y(new_n10539));
  nor_4  g10163(.A(new_n10347), .B(new_n10341), .Y(new_n10540));
  nor_4  g10164(.A(new_n10540), .B(new_n10539), .Y(new_n10541));
  not_3  g10165(.A(new_n10541), .Y(new_n10542));
  xnor_3 g10166(.A(new_n10542), .B(new_n10538), .Y(new_n10543));
  not_3  g10167(.A(new_n10543), .Y(new_n10544));
  nor_4  g10168(.A(new_n10544), .B(new_n10513), .Y(new_n10545_1));
  not_3  g10169(.A(new_n10513), .Y(new_n10546));
  nor_4  g10170(.A(new_n10543), .B(new_n10546), .Y(new_n10547_1));
  nor_4  g10171(.A(new_n10547_1), .B(new_n10545_1), .Y(new_n10548));
  xnor_3 g10172(.A(new_n10548), .B(new_n10512), .Y(new_n10549));
  not_3  g10173(.A(new_n10549), .Y(new_n10550));
  not_3  g10174(.A(new_n10383), .Y(new_n10551));
  not_3  g10175(.A(new_n10404), .Y(new_n10552));
  nand_4 g10176(.A(new_n10552), .B(new_n10385), .Y(new_n10553));
  nand_4 g10177(.A(new_n10553), .B(new_n10551), .Y(new_n10554));
  xnor_3 g10178(.A(new_n10554), .B(new_n10550), .Y(new_n10555));
  xnor_3 g10179(.A(new_n10555), .B(new_n10484), .Y(new_n10556));
  not_3  g10180(.A(new_n10409), .Y(new_n10557));
  nand_4 g10181(.A(new_n10425), .B(new_n10410), .Y(new_n10558));
  nand_4 g10182(.A(new_n10558), .B(new_n10557), .Y(new_n10559));
  xnor_3 g10183(.A(new_n10559), .B(new_n10556), .Y(new_n10560));
  xor_3  g10184(.A(new_n10560), .B(new_n10451_1), .Y(n3677));
  not_3  g10185(.A(new_n9136), .Y(new_n10562));
  xor_3  g10186(.A(new_n9137_1), .B(new_n10562), .Y(n3849));
  xor_3  g10187(.A(new_n6524), .B(new_n6523), .Y(n4088));
  xor_3  g10188(.A(new_n1197), .B(new_n1095), .Y(n4155));
  not_3  g10189(.A(new_n3091), .Y(new_n10566));
  nand_4 g10190(.A(new_n3049), .B(new_n3048), .Y(new_n10567));
  xnor_3 g10191(.A(new_n10567), .B(new_n10566), .Y(n4159));
  xor_3  g10192(.A(new_n6511), .B(new_n6313), .Y(n4226));
  nand_4 g10193(.A(n12591), .B(n4312), .Y(new_n10570));
  not_3  g10194(.A(new_n10570), .Y(new_n10571));
  nand_4 g10195(.A(new_n10261), .B(new_n10260), .Y(new_n10572));
  not_3  g10196(.A(new_n10572), .Y(new_n10573));
  nor_4  g10197(.A(new_n10266), .B(new_n10573), .Y(new_n10574));
  xnor_3 g10198(.A(new_n10574), .B(new_n10571), .Y(new_n10575));
  not_3  g10199(.A(new_n10575), .Y(new_n10576));
  nand_4 g10200(.A(n12705), .B(n3932), .Y(new_n10577));
  nand_4 g10201(.A(n12025), .B(n1798), .Y(new_n10578));
  not_3  g10202(.A(new_n10578), .Y(new_n10579));
  xor_3  g10203(.A(new_n10579), .B(new_n10577), .Y(new_n10580));
  xnor_3 g10204(.A(new_n10580), .B(new_n10576), .Y(new_n10581));
  nand_4 g10205(.A(n11662), .B(n5964), .Y(new_n10582));
  nand_4 g10206(.A(n7456), .B(n1097), .Y(new_n10583));
  xor_3  g10207(.A(new_n10583), .B(new_n10582), .Y(new_n10584));
  xnor_3 g10208(.A(new_n10584), .B(new_n10581), .Y(new_n10585));
  nor_4  g10209(.A(new_n10267), .B(new_n10258), .Y(new_n10586));
  not_3  g10210(.A(new_n10271), .Y(new_n10587));
  nor_4  g10211(.A(new_n10587), .B(new_n10268), .Y(new_n10588));
  nor_4  g10212(.A(new_n10588), .B(new_n10586), .Y(new_n10589_1));
  xnor_3 g10213(.A(new_n10589_1), .B(new_n10585), .Y(new_n10590));
  not_3  g10214(.A(new_n10590), .Y(new_n10591));
  not_3  g10215(.A(new_n10274), .Y(new_n10592));
  nand_4 g10216(.A(new_n10282), .B(new_n10277), .Y(new_n10593));
  nand_4 g10217(.A(new_n10593), .B(new_n10592), .Y(new_n10594));
  nand_4 g10218(.A(new_n10594), .B(new_n10591), .Y(new_n10595));
  nor_4  g10219(.A(new_n10574), .B(new_n10571), .Y(new_n10596));
  not_3  g10220(.A(new_n10596), .Y(new_n10597));
  nand_4 g10221(.A(new_n10580), .B(new_n10576), .Y(new_n10598));
  nand_4 g10222(.A(new_n10598), .B(new_n10597), .Y(new_n10599));
  nand_4 g10223(.A(n10327), .B(n5964), .Y(new_n10600));
  nand_4 g10224(.A(n11662), .B(n1097), .Y(new_n10601));
  nand_4 g10225(.A(n9583), .B(n5305), .Y(new_n10602));
  not_3  g10226(.A(new_n10602), .Y(new_n10603));
  xor_3  g10227(.A(new_n10603), .B(new_n10601), .Y(new_n10604));
  xnor_3 g10228(.A(new_n10604), .B(new_n10600), .Y(new_n10605));
  xnor_3 g10229(.A(new_n10605), .B(new_n10599), .Y(new_n10606));
  nor_4  g10230(.A(new_n10578), .B(new_n10577), .Y(new_n10607));
  nand_4 g10231(.A(n7456), .B(n4312), .Y(new_n10608));
  not_3  g10232(.A(new_n10608), .Y(new_n10609));
  xor_3  g10233(.A(new_n10609), .B(new_n10607), .Y(new_n10610));
  not_3  g10234(.A(new_n10610), .Y(new_n10611));
  nand_4 g10235(.A(n12025), .B(n3932), .Y(new_n10612));
  nand_4 g10236(.A(n12705), .B(n12591), .Y(new_n10613));
  nand_4 g10237(.A(n11257), .B(n1798), .Y(new_n10614));
  not_3  g10238(.A(new_n10614), .Y(new_n10615));
  xor_3  g10239(.A(new_n10615), .B(new_n10613), .Y(new_n10616));
  xnor_3 g10240(.A(new_n10616), .B(new_n10612), .Y(new_n10617));
  not_3  g10241(.A(new_n10617), .Y(new_n10618));
  nor_4  g10242(.A(new_n10618), .B(new_n10611), .Y(new_n10619));
  nor_4  g10243(.A(new_n10617), .B(new_n10610), .Y(new_n10620));
  nor_4  g10244(.A(new_n10620), .B(new_n10619), .Y(new_n10621));
  xnor_3 g10245(.A(new_n10621), .B(new_n10606), .Y(new_n10622));
  nand_4 g10246(.A(new_n10584), .B(new_n10581), .Y(new_n10623));
  nor_4  g10247(.A(new_n10583), .B(new_n10582), .Y(new_n10624));
  nor_4  g10248(.A(new_n10589_1), .B(new_n10585), .Y(new_n10625));
  xnor_3 g10249(.A(new_n10625), .B(new_n10624), .Y(new_n10626));
  nand_4 g10250(.A(new_n10626), .B(new_n10623), .Y(new_n10627));
  xnor_3 g10251(.A(new_n10627), .B(new_n10622), .Y(new_n10628));
  xnor_3 g10252(.A(new_n10628), .B(new_n10595), .Y(new_n10629));
  nand_4 g10253(.A(n10327), .B(n5305), .Y(new_n10630));
  not_3  g10254(.A(new_n10630), .Y(new_n10631));
  xnor_3 g10255(.A(new_n10594), .B(new_n10590), .Y(new_n10632));
  nor_4  g10256(.A(new_n10632), .B(new_n10631), .Y(new_n10633));
  nor_4  g10257(.A(new_n10283), .B(new_n10256), .Y(new_n10634));
  xnor_3 g10258(.A(new_n10632), .B(new_n10631), .Y(new_n10635));
  nor_4  g10259(.A(new_n10635), .B(new_n10634), .Y(new_n10636));
  nor_4  g10260(.A(new_n10636), .B(new_n10633), .Y(new_n10637));
  xnor_3 g10261(.A(new_n10637), .B(new_n10629), .Y(new_n10638));
  nand_4 g10262(.A(new_n10457), .B(new_n10455), .Y(new_n10639));
  not_3  g10263(.A(new_n10458), .Y(new_n10640));
  not_3  g10264(.A(new_n10469), .Y(new_n10641));
  nand_4 g10265(.A(new_n10641), .B(new_n10640), .Y(new_n10642));
  nand_4 g10266(.A(new_n10642), .B(new_n10639), .Y(new_n10643));
  nand_4 g10267(.A(n10451), .B(n6776), .Y(new_n10644_1));
  nand_4 g10268(.A(n12299), .B(n11023), .Y(new_n10645));
  xor_3  g10269(.A(new_n10645), .B(new_n10644_1), .Y(new_n10646));
  xnor_3 g10270(.A(new_n10646), .B(new_n10643), .Y(new_n10647));
  not_3  g10271(.A(new_n10647), .Y(new_n10648));
  nand_4 g10272(.A(n7436), .B(n3022), .Y(new_n10649));
  not_3  g10273(.A(new_n10649), .Y(new_n10650));
  nand_4 g10274(.A(n9640), .B(n8276), .Y(new_n10651));
  nand_4 g10275(.A(n9241), .B(n6703), .Y(new_n10652));
  not_3  g10276(.A(new_n10652), .Y(new_n10653));
  xor_3  g10277(.A(new_n10653), .B(new_n10651), .Y(new_n10654));
  xnor_3 g10278(.A(new_n10654), .B(new_n10650), .Y(new_n10655));
  not_3  g10279(.A(new_n10459), .Y(new_n10656));
  nor_4  g10280(.A(new_n10466), .B(new_n10656), .Y(new_n10657));
  nor_4  g10281(.A(new_n10657), .B(new_n10464), .Y(new_n10658));
  xnor_3 g10282(.A(new_n10658), .B(new_n10655), .Y(new_n10659));
  xnor_3 g10283(.A(new_n10659), .B(new_n10648), .Y(new_n10660));
  not_3  g10284(.A(new_n10471), .Y(new_n10661));
  nand_4 g10285(.A(new_n10481), .B(new_n10475), .Y(new_n10662));
  nand_4 g10286(.A(new_n10662), .B(new_n10661), .Y(new_n10663));
  nand_4 g10287(.A(new_n10663), .B(new_n10660), .Y(new_n10664));
  nand_4 g10288(.A(new_n10654), .B(new_n10649), .Y(new_n10665));
  not_3  g10289(.A(new_n10658), .Y(new_n10666));
  nand_4 g10290(.A(new_n10666), .B(new_n10655), .Y(new_n10667));
  nand_4 g10291(.A(new_n10667), .B(new_n10665), .Y(new_n10668));
  nand_4 g10292(.A(n10278), .B(n6776), .Y(new_n10669));
  nand_4 g10293(.A(n12299), .B(n10451), .Y(new_n10670));
  nand_4 g10294(.A(n11423), .B(n8759), .Y(new_n10671));
  not_3  g10295(.A(new_n10671), .Y(new_n10672));
  xor_3  g10296(.A(new_n10672), .B(new_n10670), .Y(new_n10673));
  xnor_3 g10297(.A(new_n10673), .B(new_n10669), .Y(new_n10674));
  not_3  g10298(.A(new_n10674), .Y(new_n10675));
  xnor_3 g10299(.A(new_n10675), .B(new_n10668), .Y(new_n10676));
  nor_4  g10300(.A(new_n10652), .B(new_n10651), .Y(new_n10677));
  nand_4 g10301(.A(n11023), .B(n7436), .Y(new_n10678_1));
  not_3  g10302(.A(new_n10678_1), .Y(new_n10679));
  xor_3  g10303(.A(new_n10679), .B(new_n10677), .Y(new_n10680));
  nand_4 g10304(.A(n9640), .B(n9241), .Y(new_n10681));
  nand_4 g10305(.A(n8276), .B(n3022), .Y(new_n10682));
  nand_4 g10306(.A(n10510), .B(n6703), .Y(new_n10683));
  not_3  g10307(.A(new_n10683), .Y(new_n10684));
  xor_3  g10308(.A(new_n10684), .B(new_n10682), .Y(new_n10685_1));
  xnor_3 g10309(.A(new_n10685_1), .B(new_n10681), .Y(new_n10686));
  not_3  g10310(.A(new_n10686), .Y(new_n10687));
  nor_4  g10311(.A(new_n10687), .B(new_n10680), .Y(new_n10688));
  not_3  g10312(.A(new_n10680), .Y(new_n10689));
  nor_4  g10313(.A(new_n10686), .B(new_n10689), .Y(new_n10690));
  nor_4  g10314(.A(new_n10690), .B(new_n10688), .Y(new_n10691));
  not_3  g10315(.A(new_n10691), .Y(new_n10692));
  xnor_3 g10316(.A(new_n10692), .B(new_n10676), .Y(new_n10693));
  nand_4 g10317(.A(new_n10646), .B(new_n10643), .Y(new_n10694));
  nor_4  g10318(.A(new_n10645), .B(new_n10644_1), .Y(new_n10695_1));
  nor_4  g10319(.A(new_n10659), .B(new_n10647), .Y(new_n10696));
  xnor_3 g10320(.A(new_n10696), .B(new_n10695_1), .Y(new_n10697));
  nand_4 g10321(.A(new_n10697), .B(new_n10694), .Y(new_n10698));
  xnor_3 g10322(.A(new_n10698), .B(new_n10693), .Y(new_n10699));
  xnor_3 g10323(.A(new_n10699), .B(new_n10664), .Y(new_n10700));
  nand_4 g10324(.A(n10278), .B(n8759), .Y(new_n10701));
  xnor_3 g10325(.A(new_n10663), .B(new_n10660), .Y(new_n10702));
  nor_4  g10326(.A(new_n10702), .B(new_n10701), .Y(new_n10703));
  nand_4 g10327(.A(new_n10482), .B(new_n10452), .Y(new_n10704));
  xnor_3 g10328(.A(new_n10702), .B(new_n10701), .Y(new_n10705));
  nor_4  g10329(.A(new_n10705), .B(new_n10704), .Y(new_n10706));
  nor_4  g10330(.A(new_n10706), .B(new_n10703), .Y(new_n10707));
  xnor_3 g10331(.A(new_n10707), .B(new_n10700), .Y(new_n10708));
  nand_4 g10332(.A(n12648), .B(n8665), .Y(new_n10709));
  nand_4 g10333(.A(n10545), .B(n1067), .Y(new_n10710));
  nand_4 g10334(.A(n7690), .B(n5645), .Y(new_n10711));
  xnor_3 g10335(.A(new_n10711), .B(new_n10710), .Y(new_n10712));
  nor_4  g10336(.A(new_n10712), .B(new_n10709), .Y(new_n10713));
  not_3  g10337(.A(new_n10709), .Y(new_n10714));
  not_3  g10338(.A(new_n10712), .Y(new_n10715));
  nor_4  g10339(.A(new_n10715), .B(new_n10714), .Y(new_n10716));
  nor_4  g10340(.A(new_n10716), .B(new_n10713), .Y(new_n10717));
  nor_4  g10341(.A(new_n10529), .B(new_n10522), .Y(new_n10718));
  nor_4  g10342(.A(new_n10718), .B(new_n10527), .Y(new_n10719));
  xnor_3 g10343(.A(new_n10719), .B(new_n10717), .Y(new_n10720));
  not_3  g10344(.A(new_n10720), .Y(new_n10721));
  nand_4 g10345(.A(n8476), .B(n2551), .Y(new_n10722));
  nand_4 g10346(.A(n11922), .B(n2530), .Y(new_n10723));
  xor_3  g10347(.A(new_n10723), .B(new_n10722), .Y(new_n10724));
  xnor_3 g10348(.A(new_n10724), .B(new_n10721), .Y(new_n10725));
  and_4  g10349(.A(new_n10519), .B(new_n10516), .Y(new_n10726));
  not_3  g10350(.A(new_n10532), .Y(new_n10727));
  nor_4  g10351(.A(new_n10727), .B(new_n10520), .Y(new_n10728));
  nor_4  g10352(.A(new_n10728), .B(new_n10726), .Y(new_n10729));
  xnor_3 g10353(.A(new_n10729), .B(new_n10725), .Y(new_n10730));
  not_3  g10354(.A(new_n10535), .Y(new_n10731));
  not_3  g10355(.A(new_n10537), .Y(new_n10732));
  nand_4 g10356(.A(new_n10542), .B(new_n10732), .Y(new_n10733));
  nand_4 g10357(.A(new_n10733), .B(new_n10731), .Y(new_n10734));
  not_3  g10358(.A(new_n10734), .Y(new_n10735));
  nor_4  g10359(.A(new_n10735), .B(new_n10730), .Y(new_n10736));
  nor_4  g10360(.A(new_n10711), .B(new_n10710), .Y(new_n10737));
  nand_4 g10361(.A(n12648), .B(n11922), .Y(new_n10738));
  not_3  g10362(.A(new_n10738), .Y(new_n10739));
  xor_3  g10363(.A(new_n10739), .B(new_n10737), .Y(new_n10740));
  nand_4 g10364(.A(n7690), .B(n1067), .Y(new_n10741));
  not_3  g10365(.A(new_n10741), .Y(new_n10742));
  nand_4 g10366(.A(n10545), .B(n8665), .Y(new_n10743));
  nand_4 g10367(.A(n5645), .B(n3616), .Y(new_n10744));
  xnor_3 g10368(.A(new_n10744), .B(new_n10743), .Y(new_n10745));
  xnor_3 g10369(.A(new_n10745), .B(new_n10742), .Y(new_n10746));
  xnor_3 g10370(.A(new_n10746), .B(new_n10740), .Y(new_n10747));
  not_3  g10371(.A(new_n10747), .Y(new_n10748));
  nand_4 g10372(.A(new_n10719), .B(new_n10717), .Y(new_n10749));
  not_3  g10373(.A(new_n10749), .Y(new_n10750));
  nor_4  g10374(.A(new_n10750), .B(new_n10713), .Y(new_n10751));
  not_3  g10375(.A(new_n10751), .Y(new_n10752));
  nand_4 g10376(.A(n12826), .B(n8476), .Y(new_n10753));
  not_3  g10377(.A(new_n10753), .Y(new_n10754));
  nand_4 g10378(.A(n2551), .B(n2530), .Y(new_n10755));
  nand_4 g10379(.A(n5331), .B(n4094), .Y(new_n10756));
  xnor_3 g10380(.A(new_n10756), .B(new_n10755), .Y(new_n10757));
  xor_3  g10381(.A(new_n10757), .B(new_n10754), .Y(new_n10758));
  xnor_3 g10382(.A(new_n10758), .B(new_n10752), .Y(new_n10759));
  xnor_3 g10383(.A(new_n10759), .B(new_n10748), .Y(new_n10760));
  nand_4 g10384(.A(new_n10724), .B(new_n10721), .Y(new_n10761));
  nor_4  g10385(.A(new_n10723), .B(new_n10722), .Y(new_n10762));
  nor_4  g10386(.A(new_n10729), .B(new_n10725), .Y(new_n10763));
  xnor_3 g10387(.A(new_n10763), .B(new_n10762), .Y(new_n10764));
  nand_4 g10388(.A(new_n10764), .B(new_n10761), .Y(new_n10765));
  xnor_3 g10389(.A(new_n10765), .B(new_n10760), .Y(new_n10766));
  xnor_3 g10390(.A(new_n10766), .B(new_n10736), .Y(new_n10767));
  nand_4 g10391(.A(n12826), .B(n5331), .Y(new_n10768));
  not_3  g10392(.A(new_n10768), .Y(new_n10769));
  xnor_3 g10393(.A(new_n10734), .B(new_n10730), .Y(new_n10770));
  nand_4 g10394(.A(new_n10770), .B(new_n10769), .Y(new_n10771));
  not_3  g10395(.A(new_n10770), .Y(new_n10772));
  nand_4 g10396(.A(new_n10772), .B(new_n10768), .Y(new_n10773));
  nand_4 g10397(.A(new_n10773), .B(new_n10547_1), .Y(new_n10774));
  nand_4 g10398(.A(new_n10774), .B(new_n10771), .Y(new_n10775));
  xnor_3 g10399(.A(new_n10775), .B(new_n10767), .Y(new_n10776));
  not_3  g10400(.A(new_n10776), .Y(new_n10777));
  nand_4 g10401(.A(n7965), .B(n1510), .Y(new_n10778));
  not_3  g10402(.A(new_n10778), .Y(new_n10779));
  nand_4 g10403(.A(new_n10509), .B(new_n10503), .Y(new_n10780));
  nand_4 g10404(.A(new_n10780), .B(new_n10500), .Y(new_n10781));
  nand_4 g10405(.A(n7388), .B(n159), .Y(new_n10782));
  nand_4 g10406(.A(n11892), .B(n2749), .Y(new_n10783));
  xor_3  g10407(.A(new_n10783), .B(new_n10782), .Y(new_n10784));
  xnor_3 g10408(.A(new_n10784), .B(new_n10781), .Y(new_n10785));
  nand_4 g10409(.A(n3754), .B(n2393), .Y(new_n10786));
  nand_4 g10410(.A(n10898), .B(n5860), .Y(new_n10787));
  nand_4 g10411(.A(n11876), .B(n3986), .Y(new_n10788));
  xnor_3 g10412(.A(new_n10788), .B(new_n10787), .Y(new_n10789_1));
  nor_4  g10413(.A(new_n10789_1), .B(new_n10786), .Y(new_n10790));
  not_3  g10414(.A(new_n10786), .Y(new_n10791));
  not_3  g10415(.A(new_n10789_1), .Y(new_n10792));
  nor_4  g10416(.A(new_n10792), .B(new_n10791), .Y(new_n10793));
  nor_4  g10417(.A(new_n10793), .B(new_n10790), .Y(new_n10794));
  and_4  g10418(.A(new_n10507), .B(new_n10506), .Y(new_n10795));
  nor_4  g10419(.A(new_n10508), .B(new_n10505), .Y(new_n10796));
  nor_4  g10420(.A(new_n10796), .B(new_n10795), .Y(new_n10797));
  nand_4 g10421(.A(new_n10797), .B(new_n10794), .Y(new_n10798));
  not_3  g10422(.A(new_n10798), .Y(new_n10799));
  nor_4  g10423(.A(new_n10797), .B(new_n10794), .Y(new_n10800));
  nor_4  g10424(.A(new_n10800), .B(new_n10799), .Y(new_n10801));
  xnor_3 g10425(.A(new_n10801), .B(new_n10785), .Y(new_n10802));
  nor_4  g10426(.A(new_n10490), .B(new_n10486), .Y(new_n10803));
  nor_4  g10427(.A(new_n10510_1), .B(new_n10491), .Y(new_n10804));
  nor_4  g10428(.A(new_n10804), .B(new_n10803), .Y(new_n10805));
  xnor_3 g10429(.A(new_n10805), .B(new_n10802), .Y(new_n10806));
  nand_4 g10430(.A(new_n10806), .B(new_n10779), .Y(new_n10807));
  not_3  g10431(.A(new_n10485), .Y(new_n10808));
  nor_4  g10432(.A(new_n10511), .B(new_n10808), .Y(new_n10809));
  xnor_3 g10433(.A(new_n10806), .B(new_n10778), .Y(new_n10810));
  nand_4 g10434(.A(new_n10810), .B(new_n10809), .Y(new_n10811));
  nand_4 g10435(.A(new_n10811), .B(new_n10807), .Y(new_n10812));
  not_3  g10436(.A(new_n10802), .Y(new_n10813));
  nor_4  g10437(.A(new_n10805), .B(new_n10813), .Y(new_n10814));
  nor_4  g10438(.A(new_n10783), .B(new_n10782), .Y(new_n10815));
  nor_4  g10439(.A(new_n10784), .B(new_n10781), .Y(new_n10816));
  nor_4  g10440(.A(new_n10801), .B(new_n10785), .Y(new_n10817));
  nor_4  g10441(.A(new_n10817), .B(new_n10816), .Y(new_n10818));
  xnor_3 g10442(.A(new_n10818), .B(new_n10815), .Y(new_n10819));
  not_3  g10443(.A(new_n10790), .Y(new_n10820));
  nand_4 g10444(.A(new_n10798), .B(new_n10820), .Y(new_n10821));
  nand_4 g10445(.A(n7388), .B(n1510), .Y(new_n10822));
  not_3  g10446(.A(new_n10822), .Y(new_n10823));
  nand_4 g10447(.A(n11892), .B(n159), .Y(new_n10824));
  not_3  g10448(.A(new_n10824), .Y(new_n10825));
  nand_4 g10449(.A(n12247), .B(n7965), .Y(new_n10826));
  not_3  g10450(.A(new_n10826), .Y(new_n10827));
  nand_4 g10451(.A(new_n10827), .B(new_n10825), .Y(new_n10828));
  nand_4 g10452(.A(new_n10826), .B(new_n10824), .Y(new_n10829));
  nand_4 g10453(.A(new_n10829), .B(new_n10828), .Y(new_n10830));
  xor_3  g10454(.A(new_n10830), .B(new_n10823), .Y(new_n10831));
  xnor_3 g10455(.A(new_n10831), .B(new_n10821), .Y(new_n10832));
  nor_4  g10456(.A(new_n10788), .B(new_n10787), .Y(new_n10833));
  nand_4 g10457(.A(n2749), .B(n2393), .Y(new_n10834));
  not_3  g10458(.A(new_n10834), .Y(new_n10835));
  xor_3  g10459(.A(new_n10835), .B(new_n10833), .Y(new_n10836));
  not_3  g10460(.A(new_n10836), .Y(new_n10837));
  nand_4 g10461(.A(n10898), .B(n3986), .Y(new_n10838));
  not_3  g10462(.A(new_n10838), .Y(new_n10839));
  nand_4 g10463(.A(n11876), .B(n5857), .Y(new_n10840));
  nand_4 g10464(.A(n5860), .B(n3754), .Y(new_n10841));
  not_3  g10465(.A(new_n10841), .Y(new_n10842));
  xor_3  g10466(.A(new_n10842), .B(new_n10840), .Y(new_n10843));
  xnor_3 g10467(.A(new_n10843), .B(new_n10839), .Y(new_n10844));
  xnor_3 g10468(.A(new_n10844), .B(new_n10837), .Y(new_n10845));
  xnor_3 g10469(.A(new_n10845), .B(new_n10832), .Y(new_n10846));
  xnor_3 g10470(.A(new_n10846), .B(new_n10819), .Y(new_n10847));
  xnor_3 g10471(.A(new_n10847), .B(new_n10814), .Y(new_n10848_1));
  xnor_3 g10472(.A(new_n10848_1), .B(new_n10812), .Y(new_n10849));
  xnor_3 g10473(.A(new_n10849), .B(new_n10777), .Y(new_n10850));
  xnor_3 g10474(.A(new_n10810), .B(new_n10809), .Y(new_n10851_1));
  nand_4 g10475(.A(new_n10773), .B(new_n10771), .Y(new_n10852));
  xnor_3 g10476(.A(new_n10852), .B(new_n10547_1), .Y(new_n10853));
  not_3  g10477(.A(new_n10853), .Y(new_n10854));
  nand_4 g10478(.A(new_n10854), .B(new_n10851_1), .Y(new_n10855));
  nor_4  g10479(.A(new_n10548), .B(new_n10512), .Y(new_n10856));
  not_3  g10480(.A(new_n10856), .Y(new_n10857));
  nand_4 g10481(.A(new_n10554), .B(new_n10550), .Y(new_n10858));
  nand_4 g10482(.A(new_n10858), .B(new_n10857), .Y(new_n10859));
  xnor_3 g10483(.A(new_n10853), .B(new_n10851_1), .Y(new_n10860));
  nand_4 g10484(.A(new_n10860), .B(new_n10859), .Y(new_n10861));
  nand_4 g10485(.A(new_n10861), .B(new_n10855), .Y(new_n10862));
  xnor_3 g10486(.A(new_n10862), .B(new_n10850), .Y(new_n10863));
  xnor_3 g10487(.A(new_n10863), .B(new_n10708), .Y(new_n10864));
  not_3  g10488(.A(new_n10704), .Y(new_n10865));
  not_3  g10489(.A(new_n10705), .Y(new_n10866));
  nor_4  g10490(.A(new_n10866), .B(new_n10865), .Y(new_n10867));
  nor_4  g10491(.A(new_n10867), .B(new_n10706), .Y(new_n10868));
  not_3  g10492(.A(new_n10868), .Y(new_n10869));
  not_3  g10493(.A(new_n10860), .Y(new_n10870));
  xnor_3 g10494(.A(new_n10870), .B(new_n10859), .Y(new_n10871));
  nand_4 g10495(.A(new_n10871), .B(new_n10869), .Y(new_n10872));
  nand_4 g10496(.A(new_n10555), .B(new_n10484), .Y(new_n10873));
  not_3  g10497(.A(new_n10873), .Y(new_n10874));
  nor_4  g10498(.A(new_n10559), .B(new_n10556), .Y(new_n10875));
  nor_4  g10499(.A(new_n10875), .B(new_n10874), .Y(new_n10876));
  xnor_3 g10500(.A(new_n10871), .B(new_n10868), .Y(new_n10877));
  nand_4 g10501(.A(new_n10877), .B(new_n10876), .Y(new_n10878));
  nand_4 g10502(.A(new_n10878), .B(new_n10872), .Y(new_n10879));
  xnor_3 g10503(.A(new_n10879), .B(new_n10864), .Y(new_n10880));
  nand_4 g10504(.A(new_n10880), .B(new_n10638), .Y(new_n10881));
  not_3  g10505(.A(new_n10638), .Y(new_n10882));
  xnor_3 g10506(.A(new_n10880), .B(new_n10882), .Y(new_n10883));
  not_3  g10507(.A(new_n10635), .Y(new_n10884));
  xor_3  g10508(.A(new_n10884), .B(new_n10634), .Y(new_n10885));
  not_3  g10509(.A(new_n10885), .Y(new_n10886));
  not_3  g10510(.A(new_n10877), .Y(new_n10887));
  xnor_3 g10511(.A(new_n10887), .B(new_n10876), .Y(new_n10888));
  nand_4 g10512(.A(new_n10888), .B(new_n10886), .Y(new_n10889));
  not_3  g10513(.A(new_n10889), .Y(new_n10890));
  nor_4  g10514(.A(new_n10888), .B(new_n10886), .Y(new_n10891));
  nor_4  g10515(.A(new_n10891), .B(new_n10890), .Y(new_n10892));
  not_3  g10516(.A(new_n10284), .Y(new_n10893));
  not_3  g10517(.A(new_n10450), .Y(new_n10894));
  nor_4  g10518(.A(new_n10894), .B(new_n10893), .Y(new_n10895));
  nor_4  g10519(.A(new_n10560), .B(new_n10451_1), .Y(new_n10896));
  nor_4  g10520(.A(new_n10896), .B(new_n10895), .Y(new_n10897));
  nand_4 g10521(.A(new_n10897), .B(new_n10892), .Y(new_n10898_1));
  nand_4 g10522(.A(new_n10898_1), .B(new_n10889), .Y(new_n10899));
  nand_4 g10523(.A(new_n10899), .B(new_n10883), .Y(new_n10900));
  nand_4 g10524(.A(new_n10900), .B(new_n10881), .Y(new_n10901));
  nand_4 g10525(.A(new_n10863), .B(new_n10708), .Y(new_n10902));
  not_3  g10526(.A(new_n10708), .Y(new_n10903));
  xnor_3 g10527(.A(new_n10863), .B(new_n10903), .Y(new_n10904));
  nand_4 g10528(.A(new_n10879), .B(new_n10904), .Y(new_n10905));
  nand_4 g10529(.A(new_n10905), .B(new_n10902), .Y(new_n10906));
  nand_4 g10530(.A(new_n10696), .B(new_n10695_1), .Y(new_n10907));
  nand_4 g10531(.A(new_n10698), .B(new_n10693), .Y(new_n10908));
  nand_4 g10532(.A(new_n10908), .B(new_n10907), .Y(new_n10909));
  and_4  g10533(.A(new_n10679), .B(new_n10677), .Y(new_n10910));
  or_4   g10534(.A(new_n10690), .B(new_n10910), .Y(new_n10911));
  not_3  g10535(.A(new_n10670), .Y(new_n10912));
  nor_4  g10536(.A(new_n10672), .B(new_n10912), .Y(new_n10913_1));
  not_3  g10537(.A(new_n10669), .Y(new_n10914));
  nor_4  g10538(.A(new_n10673), .B(new_n10914), .Y(new_n10915));
  nor_4  g10539(.A(new_n10915), .B(new_n10913_1), .Y(new_n10916));
  nand_4 g10540(.A(n12511), .B(n7965), .Y(new_n10917));
  xor_3  g10541(.A(new_n10917), .B(new_n10916), .Y(new_n10918));
  nand_4 g10542(.A(n8759), .B(n2278), .Y(new_n10919));
  nand_4 g10543(.A(n10510), .B(n9640), .Y(new_n10920));
  xor_3  g10544(.A(new_n10920), .B(new_n10919), .Y(new_n10921));
  xnor_3 g10545(.A(new_n10921), .B(new_n10918), .Y(new_n10922));
  xnor_3 g10546(.A(new_n10922), .B(new_n10911), .Y(new_n10923));
  xnor_3 g10547(.A(new_n10923), .B(new_n10909), .Y(new_n10924));
  xnor_3 g10548(.A(new_n10924), .B(new_n10906), .Y(new_n10925));
  nand_4 g10549(.A(new_n10849), .B(new_n10777), .Y(new_n10926));
  not_3  g10550(.A(new_n10850), .Y(new_n10927));
  nand_4 g10551(.A(new_n10862), .B(new_n10927), .Y(new_n10928_1));
  nand_4 g10552(.A(new_n10928_1), .B(new_n10926), .Y(new_n10929));
  not_3  g10553(.A(new_n10847), .Y(new_n10930));
  nand_4 g10554(.A(new_n10930), .B(new_n10814), .Y(new_n10931));
  nand_4 g10555(.A(new_n10848_1), .B(new_n10812), .Y(new_n10932));
  nand_4 g10556(.A(new_n10932), .B(new_n10931), .Y(new_n10933));
  nor_4  g10557(.A(new_n10699), .B(new_n10664), .Y(new_n10934));
  nor_4  g10558(.A(new_n10707), .B(new_n10700), .Y(new_n10935));
  nor_4  g10559(.A(new_n10935), .B(new_n10934), .Y(new_n10936));
  nand_4 g10560(.A(new_n10766), .B(new_n10736), .Y(new_n10937));
  not_3  g10561(.A(new_n10767), .Y(new_n10938));
  nand_4 g10562(.A(new_n10775), .B(new_n10938), .Y(new_n10939));
  nand_4 g10563(.A(new_n10939), .B(new_n10937), .Y(new_n10940));
  not_3  g10564(.A(new_n10821), .Y(new_n10941));
  nand_4 g10565(.A(new_n10831), .B(new_n10941), .Y(new_n10942));
  not_3  g10566(.A(new_n10845), .Y(new_n10943));
  nand_4 g10567(.A(new_n10943), .B(new_n10832), .Y(new_n10944));
  nand_4 g10568(.A(new_n10944), .B(new_n10942), .Y(new_n10945));
  nand_4 g10569(.A(new_n10829), .B(new_n10823), .Y(new_n10946));
  and_4  g10570(.A(new_n10946), .B(new_n10828), .Y(new_n10947));
  nand_4 g10571(.A(n11892), .B(n1510), .Y(new_n10948));
  nand_4 g10572(.A(n2393), .B(n159), .Y(new_n10949_1));
  xor_3  g10573(.A(new_n10949_1), .B(new_n10948), .Y(new_n10950));
  xnor_3 g10574(.A(new_n10950), .B(new_n10947), .Y(new_n10951));
  not_3  g10575(.A(new_n10840), .Y(new_n10952));
  nor_4  g10576(.A(new_n10842), .B(new_n10952), .Y(new_n10953));
  nor_4  g10577(.A(new_n10843), .B(new_n10839), .Y(new_n10954));
  nor_4  g10578(.A(new_n10954), .B(new_n10953), .Y(new_n10955));
  nand_4 g10579(.A(n5860), .B(n2749), .Y(new_n10956));
  nand_4 g10580(.A(n10685), .B(n5331), .Y(new_n10957));
  nand_4 g10581(.A(n5645), .B(n4499), .Y(new_n10958));
  xor_3  g10582(.A(new_n10958), .B(new_n10957), .Y(new_n10959));
  xnor_3 g10583(.A(new_n10959), .B(new_n10956), .Y(new_n10960));
  xnor_3 g10584(.A(new_n10960), .B(new_n10955), .Y(new_n10961));
  xnor_3 g10585(.A(new_n10961), .B(new_n10951), .Y(new_n10962));
  nand_4 g10586(.A(new_n10835), .B(new_n10833), .Y(new_n10963));
  nand_4 g10587(.A(new_n10844), .B(new_n10836), .Y(new_n10964));
  nand_4 g10588(.A(new_n10964), .B(new_n10963), .Y(new_n10965_1));
  nand_4 g10589(.A(n12247), .B(n7388), .Y(new_n10966));
  not_3  g10590(.A(new_n10966), .Y(new_n10967));
  xnor_3 g10591(.A(new_n10967), .B(new_n10965_1), .Y(new_n10968));
  xnor_3 g10592(.A(new_n10968), .B(new_n10962), .Y(new_n10969));
  xnor_3 g10593(.A(new_n10969), .B(new_n10945), .Y(new_n10970));
  xnor_3 g10594(.A(new_n10970), .B(new_n10940), .Y(new_n10971));
  xnor_3 g10595(.A(new_n10971), .B(new_n10936), .Y(new_n10972));
  xnor_3 g10596(.A(new_n10972), .B(new_n10933), .Y(new_n10973));
  xnor_3 g10597(.A(new_n10973), .B(new_n10929), .Y(new_n10974));
  nand_4 g10598(.A(new_n10758), .B(new_n10751), .Y(new_n10975));
  nand_4 g10599(.A(new_n10759), .B(new_n10747), .Y(new_n10976));
  nand_4 g10600(.A(new_n10976), .B(new_n10975), .Y(new_n10977));
  nand_4 g10601(.A(n12648), .B(n2551), .Y(new_n10978));
  not_3  g10602(.A(new_n10978), .Y(new_n10979));
  and_4  g10603(.A(new_n10756), .B(new_n10755), .Y(new_n10980));
  nor_4  g10604(.A(new_n10757), .B(new_n10754), .Y(new_n10981));
  nor_4  g10605(.A(new_n10981), .B(new_n10980), .Y(new_n10982));
  xnor_3 g10606(.A(new_n10982), .B(new_n10979), .Y(new_n10983));
  and_4  g10607(.A(new_n10744), .B(new_n10743), .Y(new_n10984));
  nor_4  g10608(.A(new_n10745), .B(new_n10742), .Y(new_n10985));
  nor_4  g10609(.A(new_n10985), .B(new_n10984), .Y(new_n10986));
  nand_4 g10610(.A(n11922), .B(n10545), .Y(new_n10987));
  nand_4 g10611(.A(n8665), .B(n7690), .Y(new_n10988));
  xnor_3 g10612(.A(new_n10988), .B(new_n10987), .Y(new_n10989));
  nand_4 g10613(.A(n8476), .B(n4094), .Y(new_n10990_1));
  nand_4 g10614(.A(n12826), .B(n2530), .Y(new_n10991));
  xnor_3 g10615(.A(new_n10991), .B(new_n10990_1), .Y(new_n10992));
  xnor_3 g10616(.A(new_n10992), .B(new_n10989), .Y(new_n10993));
  xnor_3 g10617(.A(new_n10993), .B(new_n10986), .Y(new_n10994));
  xnor_3 g10618(.A(new_n10994), .B(new_n10983), .Y(new_n10995));
  nand_4 g10619(.A(new_n10739), .B(new_n10737), .Y(new_n10996));
  nand_4 g10620(.A(new_n10746), .B(new_n10740), .Y(new_n10997));
  nand_4 g10621(.A(new_n10997), .B(new_n10996), .Y(new_n10998));
  nand_4 g10622(.A(n10547), .B(n1798), .Y(new_n10999));
  not_3  g10623(.A(new_n10999), .Y(new_n11000));
  xnor_3 g10624(.A(new_n11000), .B(new_n10998), .Y(new_n11001));
  xnor_3 g10625(.A(new_n11001), .B(new_n10995), .Y(new_n11002));
  xnor_3 g10626(.A(new_n11002), .B(new_n10977), .Y(new_n11003));
  nand_4 g10627(.A(n3616), .B(n1067), .Y(new_n11004));
  nand_4 g10628(.A(n5305), .B(n753), .Y(new_n11005));
  xor_3  g10629(.A(new_n11005), .B(new_n11004), .Y(new_n11006));
  xnor_3 g10630(.A(new_n11006), .B(new_n11003), .Y(new_n11007));
  nand_4 g10631(.A(new_n10763), .B(new_n10762), .Y(new_n11008));
  not_3  g10632(.A(new_n10760), .Y(new_n11009));
  nand_4 g10633(.A(new_n10765), .B(new_n11009), .Y(new_n11010));
  nand_4 g10634(.A(new_n11010), .B(new_n11008), .Y(new_n11011));
  xnor_3 g10635(.A(new_n11011), .B(new_n11007), .Y(new_n11012));
  not_3  g10636(.A(new_n10682), .Y(new_n11013));
  nor_4  g10637(.A(new_n10684), .B(new_n11013), .Y(new_n11014));
  not_3  g10638(.A(new_n10681), .Y(new_n11015));
  nor_4  g10639(.A(new_n10685_1), .B(new_n11015), .Y(new_n11016));
  nor_4  g10640(.A(new_n11016), .B(new_n11014), .Y(new_n11017));
  nand_4 g10641(.A(n10451), .B(n7436), .Y(new_n11018));
  nand_4 g10642(.A(n9241), .B(n3022), .Y(new_n11019));
  xor_3  g10643(.A(new_n11019), .B(new_n11018), .Y(new_n11020));
  nand_4 g10644(.A(n11423), .B(n6776), .Y(new_n11021));
  nand_4 g10645(.A(n11023), .B(n8276), .Y(new_n11022));
  not_3  g10646(.A(new_n11022), .Y(new_n11023_1));
  xor_3  g10647(.A(new_n11023_1), .B(new_n11021), .Y(new_n11024));
  xor_3  g10648(.A(new_n11024), .B(new_n11020), .Y(new_n11025));
  xnor_3 g10649(.A(new_n11025), .B(new_n11017), .Y(new_n11026));
  nand_4 g10650(.A(n12299), .B(n10278), .Y(new_n11027));
  nand_4 g10651(.A(n10644), .B(n6703), .Y(new_n11028));
  not_3  g10652(.A(new_n11028), .Y(new_n11029));
  xor_3  g10653(.A(new_n11029), .B(new_n11027), .Y(new_n11030));
  xnor_3 g10654(.A(new_n11030), .B(new_n11026), .Y(new_n11031));
  xnor_3 g10655(.A(new_n11031), .B(new_n11012), .Y(new_n11032));
  nand_4 g10656(.A(new_n10625), .B(new_n10624), .Y(new_n11033));
  not_3  g10657(.A(new_n10622), .Y(new_n11034));
  nand_4 g10658(.A(new_n10627), .B(new_n11034), .Y(new_n11035));
  nand_4 g10659(.A(new_n11035), .B(new_n11033), .Y(new_n11036));
  nand_4 g10660(.A(new_n10674), .B(new_n10668), .Y(new_n11037));
  nand_4 g10661(.A(new_n10692), .B(new_n10676), .Y(new_n11038));
  nand_4 g10662(.A(new_n11038), .B(new_n11037), .Y(new_n11039));
  xnor_3 g10663(.A(new_n11039), .B(new_n11036), .Y(new_n11040));
  xnor_3 g10664(.A(new_n11040), .B(new_n11032), .Y(new_n11041));
  and_4  g10665(.A(new_n10605), .B(new_n10599), .Y(new_n11042));
  not_3  g10666(.A(new_n10621), .Y(new_n11043));
  nor_4  g10667(.A(new_n11043), .B(new_n10606), .Y(new_n11044));
  nor_4  g10668(.A(new_n11044), .B(new_n11042), .Y(new_n11045));
  not_3  g10669(.A(new_n10595), .Y(new_n11046));
  nand_4 g10670(.A(new_n10628), .B(new_n11046), .Y(new_n11047));
  nand_4 g10671(.A(new_n10637), .B(new_n10629), .Y(new_n11048));
  nand_4 g10672(.A(new_n11048), .B(new_n11047), .Y(new_n11049));
  xnor_3 g10673(.A(new_n11049), .B(new_n11045), .Y(new_n11050));
  xnor_3 g10674(.A(new_n11050), .B(new_n11041), .Y(new_n11051));
  nand_4 g10675(.A(new_n10818), .B(new_n10815), .Y(new_n11052));
  not_3  g10676(.A(new_n10819), .Y(new_n11053));
  not_3  g10677(.A(new_n10846), .Y(new_n11054));
  nand_4 g10678(.A(new_n11054), .B(new_n11053), .Y(new_n11055));
  nand_4 g10679(.A(new_n11055), .B(new_n11052), .Y(new_n11056));
  nor_4  g10680(.A(new_n10609), .B(new_n10607), .Y(new_n11057));
  nor_4  g10681(.A(new_n10619), .B(new_n11057), .Y(new_n11058));
  nand_4 g10682(.A(n10898), .B(n5857), .Y(new_n11059));
  nand_4 g10683(.A(n11257), .B(n3932), .Y(new_n11060));
  not_3  g10684(.A(new_n11060), .Y(new_n11061));
  xor_3  g10685(.A(new_n11061), .B(new_n11059), .Y(new_n11062));
  xor_3  g10686(.A(new_n11062), .B(new_n11058), .Y(new_n11063));
  nand_4 g10687(.A(n11876), .B(n45), .Y(new_n11064));
  nand_4 g10688(.A(n3986), .B(n3754), .Y(new_n11065));
  not_3  g10689(.A(new_n11065), .Y(new_n11066));
  xor_3  g10690(.A(new_n11066), .B(new_n11064), .Y(new_n11067));
  nand_4 g10691(.A(n10327), .B(n1097), .Y(new_n11068));
  nand_4 g10692(.A(n12705), .B(n7456), .Y(new_n11069));
  xor_3  g10693(.A(new_n11069), .B(new_n11068), .Y(new_n11070));
  nand_4 g10694(.A(n12591), .B(n12025), .Y(new_n11071));
  nand_4 g10695(.A(n9583), .B(n5964), .Y(new_n11072));
  nand_4 g10696(.A(n11662), .B(n4312), .Y(new_n11073));
  xor_3  g10697(.A(new_n11073), .B(new_n11072), .Y(new_n11074));
  xor_3  g10698(.A(new_n11074), .B(new_n11071), .Y(new_n11075));
  xnor_3 g10699(.A(new_n11075), .B(new_n11070), .Y(new_n11076));
  not_3  g10700(.A(new_n10601), .Y(new_n11077));
  nor_4  g10701(.A(new_n10603), .B(new_n11077), .Y(new_n11078));
  not_3  g10702(.A(new_n10600), .Y(new_n11079));
  nor_4  g10703(.A(new_n10604), .B(new_n11079), .Y(new_n11080));
  nor_4  g10704(.A(new_n11080), .B(new_n11078), .Y(new_n11081));
  not_3  g10705(.A(new_n10613), .Y(new_n11082));
  nor_4  g10706(.A(new_n10615), .B(new_n11082), .Y(new_n11083));
  not_3  g10707(.A(new_n10612), .Y(new_n11084));
  nor_4  g10708(.A(new_n10616), .B(new_n11084), .Y(new_n11085));
  nor_4  g10709(.A(new_n11085), .B(new_n11083), .Y(new_n11086));
  xnor_3 g10710(.A(new_n11086), .B(new_n11081), .Y(new_n11087));
  xnor_3 g10711(.A(new_n11087), .B(new_n11076), .Y(new_n11088));
  xnor_3 g10712(.A(new_n11088), .B(new_n11067), .Y(new_n11089));
  xnor_3 g10713(.A(new_n11089), .B(new_n11063), .Y(new_n11090));
  xnor_3 g10714(.A(new_n11090), .B(new_n11056), .Y(new_n11091));
  xnor_3 g10715(.A(new_n11091), .B(new_n11051), .Y(new_n11092));
  xnor_3 g10716(.A(new_n11092), .B(new_n10974), .Y(new_n11093));
  xnor_3 g10717(.A(new_n11093), .B(new_n10925), .Y(new_n11094));
  xnor_3 g10718(.A(new_n11094), .B(new_n10901), .Y(n4230));
  not_3  g10719(.A(new_n6285), .Y(new_n11096));
  xor_3  g10720(.A(new_n11096), .B(new_n6284), .Y(n4300));
  not_3  g10721(.A(new_n3830), .Y(new_n11098));
  xor_3  g10722(.A(new_n11098), .B(new_n3829), .Y(n4326));
  not_3  g10723(.A(new_n1324), .Y(new_n11100));
  nor_4  g10724(.A(new_n11100), .B(new_n1317), .Y(new_n11101));
  not_3  g10725(.A(new_n11101), .Y(new_n11102));
  nand_4 g10726(.A(n6687), .B(n5320), .Y(new_n11103));
  not_3  g10727(.A(new_n1300), .Y(new_n11104));
  nand_4 g10728(.A(new_n1309), .B(new_n11104), .Y(new_n11105));
  not_3  g10729(.A(new_n11105), .Y(new_n11106));
  nor_4  g10730(.A(new_n1316), .B(new_n1310), .Y(new_n11107));
  nor_4  g10731(.A(new_n11107), .B(new_n11106), .Y(new_n11108));
  xnor_3 g10732(.A(new_n11108), .B(new_n11103), .Y(new_n11109));
  nand_4 g10733(.A(n4370), .B(n2564), .Y(new_n11110));
  not_3  g10734(.A(new_n11110), .Y(new_n11111));
  and_4  g10735(.A(new_n1314), .B(new_n1313), .Y(new_n11112));
  nor_4  g10736(.A(new_n1315), .B(new_n1312), .Y(new_n11113));
  nor_4  g10737(.A(new_n11113), .B(new_n11112), .Y(new_n11114));
  nand_4 g10738(.A(new_n11114), .B(new_n11111), .Y(new_n11115));
  not_3  g10739(.A(new_n11115), .Y(new_n11116));
  nor_4  g10740(.A(new_n11114), .B(new_n11111), .Y(new_n11117));
  nor_4  g10741(.A(new_n11117), .B(new_n11116), .Y(new_n11118));
  nand_4 g10742(.A(n6770), .B(n5212), .Y(new_n11119));
  nand_4 g10743(.A(n11877), .B(n4189), .Y(new_n11120));
  nand_4 g10744(.A(n11407), .B(n9920), .Y(new_n11121));
  xnor_3 g10745(.A(new_n11121), .B(new_n11120), .Y(new_n11122));
  xor_3  g10746(.A(new_n11122), .B(new_n11119), .Y(new_n11123));
  nand_4 g10747(.A(new_n11123), .B(new_n11118), .Y(new_n11124));
  not_3  g10748(.A(new_n11124), .Y(new_n11125));
  nor_4  g10749(.A(new_n11123), .B(new_n11118), .Y(new_n11126));
  nor_4  g10750(.A(new_n11126), .B(new_n11125), .Y(new_n11127));
  not_3  g10751(.A(new_n11127), .Y(new_n11128));
  xnor_3 g10752(.A(new_n11128), .B(new_n11109), .Y(new_n11129));
  not_3  g10753(.A(new_n11129), .Y(new_n11130));
  xor_3  g10754(.A(new_n11130), .B(new_n11102), .Y(new_n11131));
  not_3  g10755(.A(new_n1444), .Y(new_n11132));
  nor_4  g10756(.A(new_n11132), .B(new_n1443), .Y(new_n11133));
  nand_4 g10757(.A(n8336), .B(n2433), .Y(new_n11134));
  nand_4 g10758(.A(n10928), .B(n8819), .Y(new_n11135));
  not_3  g10759(.A(new_n11135), .Y(new_n11136));
  not_3  g10760(.A(new_n1434), .Y(new_n11137));
  not_3  g10761(.A(new_n1435), .Y(new_n11138));
  nor_4  g10762(.A(new_n11138), .B(new_n11137), .Y(new_n11139));
  nor_4  g10763(.A(new_n1435), .B(new_n1434), .Y(new_n11140));
  nor_4  g10764(.A(new_n11140), .B(new_n1433), .Y(new_n11141));
  nor_4  g10765(.A(new_n11141), .B(new_n11139), .Y(new_n11142));
  xnor_3 g10766(.A(new_n11142), .B(new_n11136), .Y(new_n11143));
  nand_4 g10767(.A(n11728), .B(n2226), .Y(new_n11144));
  not_3  g10768(.A(new_n11144), .Y(new_n11145));
  nand_4 g10769(.A(n6986), .B(n6429), .Y(new_n11146));
  not_3  g10770(.A(new_n11146), .Y(new_n11147));
  nand_4 g10771(.A(n12709), .B(n1094), .Y(new_n11148));
  not_3  g10772(.A(new_n11148), .Y(new_n11149));
  nor_4  g10773(.A(new_n11149), .B(new_n11147), .Y(new_n11150));
  nor_4  g10774(.A(new_n11148), .B(new_n11146), .Y(new_n11151));
  nor_4  g10775(.A(new_n11151), .B(new_n11150), .Y(new_n11152));
  xnor_3 g10776(.A(new_n11152), .B(new_n11145), .Y(new_n11153_1));
  xnor_3 g10777(.A(new_n11153_1), .B(new_n11143), .Y(new_n11154));
  nor_4  g10778(.A(new_n11154), .B(new_n11134), .Y(new_n11155));
  not_3  g10779(.A(new_n11134), .Y(new_n11156));
  not_3  g10780(.A(new_n11154), .Y(new_n11157));
  nor_4  g10781(.A(new_n11157), .B(new_n11156), .Y(new_n11158));
  nor_4  g10782(.A(new_n11158), .B(new_n11155), .Y(new_n11159));
  nor_4  g10783(.A(new_n1438), .B(new_n1431), .Y(new_n11160));
  not_3  g10784(.A(new_n11160), .Y(new_n11161));
  nand_4 g10785(.A(new_n1442), .B(new_n1439), .Y(new_n11162));
  nand_4 g10786(.A(new_n11162), .B(new_n11161), .Y(new_n11163));
  xnor_3 g10787(.A(new_n11163), .B(new_n11159), .Y(new_n11164));
  xnor_3 g10788(.A(new_n11164), .B(new_n11133), .Y(new_n11165));
  nand_4 g10789(.A(new_n1491), .B(new_n1445), .Y(new_n11166));
  nand_4 g10790(.A(new_n1496), .B(new_n1499), .Y(new_n11167));
  nand_4 g10791(.A(new_n11167), .B(new_n11166), .Y(new_n11168));
  nand_4 g10792(.A(new_n11168), .B(new_n11165), .Y(new_n11169));
  not_3  g10793(.A(new_n11165), .Y(new_n11170));
  not_3  g10794(.A(new_n11166), .Y(new_n11171));
  nor_4  g10795(.A(new_n1498), .B(new_n11171), .Y(new_n11172));
  nand_4 g10796(.A(new_n11172), .B(new_n11170), .Y(new_n11173));
  nand_4 g10797(.A(new_n11173), .B(new_n11169), .Y(new_n11174));
  nand_4 g10798(.A(n12069), .B(n11967), .Y(new_n11175));
  nand_4 g10799(.A(n12391), .B(n6254), .Y(new_n11176));
  not_3  g10800(.A(new_n11176), .Y(new_n11177));
  not_3  g10801(.A(new_n1453), .Y(new_n11178));
  nor_4  g10802(.A(new_n1459), .B(new_n11178), .Y(new_n11179));
  nor_4  g10803(.A(new_n11179), .B(new_n1458), .Y(new_n11180));
  xnor_3 g10804(.A(new_n11180), .B(new_n11177), .Y(new_n11181));
  nand_4 g10805(.A(n7160), .B(n7159), .Y(new_n11182));
  not_3  g10806(.A(new_n11182), .Y(new_n11183));
  nand_4 g10807(.A(n12777), .B(n7891), .Y(new_n11184));
  not_3  g10808(.A(new_n11184), .Y(new_n11185));
  nand_4 g10809(.A(n12489), .B(n4828), .Y(new_n11186));
  not_3  g10810(.A(new_n11186), .Y(new_n11187));
  nor_4  g10811(.A(new_n11187), .B(new_n11185), .Y(new_n11188));
  nor_4  g10812(.A(new_n11186), .B(new_n11184), .Y(new_n11189));
  nor_4  g10813(.A(new_n11189), .B(new_n11188), .Y(new_n11190));
  xnor_3 g10814(.A(new_n11190), .B(new_n11183), .Y(new_n11191));
  xnor_3 g10815(.A(new_n11191), .B(new_n11181), .Y(new_n11192));
  nor_4  g10816(.A(new_n11192), .B(new_n11175), .Y(new_n11193));
  not_3  g10817(.A(new_n11175), .Y(new_n11194));
  not_3  g10818(.A(new_n11192), .Y(new_n11195));
  nor_4  g10819(.A(new_n11195), .B(new_n11194), .Y(new_n11196));
  nor_4  g10820(.A(new_n11196), .B(new_n11193), .Y(new_n11197));
  nand_4 g10821(.A(new_n1451), .B(new_n1447), .Y(new_n11198));
  nor_4  g10822(.A(new_n1462), .B(new_n1452), .Y(new_n11199));
  not_3  g10823(.A(new_n11199), .Y(new_n11200));
  nand_4 g10824(.A(new_n11200), .B(new_n11198), .Y(new_n11201));
  xnor_3 g10825(.A(new_n11201), .B(new_n11197), .Y(new_n11202));
  not_3  g10826(.A(new_n11202), .Y(new_n11203));
  nor_4  g10827(.A(new_n11203), .B(new_n1466), .Y(new_n11204));
  not_3  g10828(.A(new_n1466), .Y(new_n11205));
  nor_4  g10829(.A(new_n11202), .B(new_n11205), .Y(new_n11206));
  nor_4  g10830(.A(new_n11206), .B(new_n11204), .Y(new_n11207));
  not_3  g10831(.A(new_n11207), .Y(new_n11208));
  nand_4 g10832(.A(n12947), .B(n11222), .Y(new_n11209));
  nand_4 g10833(.A(n11791), .B(n11153), .Y(new_n11210));
  not_3  g10834(.A(new_n1475), .Y(new_n11211));
  not_3  g10835(.A(new_n1476), .Y(new_n11212));
  nor_4  g10836(.A(new_n11212), .B(new_n11211), .Y(new_n11213));
  not_3  g10837(.A(new_n1474), .Y(new_n11214));
  nor_4  g10838(.A(new_n1477), .B(new_n11214), .Y(new_n11215));
  nor_4  g10839(.A(new_n11215), .B(new_n11213), .Y(new_n11216_1));
  xnor_3 g10840(.A(new_n11216_1), .B(new_n11210), .Y(new_n11217));
  nand_4 g10841(.A(n5760), .B(n996), .Y(new_n11218));
  nand_4 g10842(.A(n5314), .B(n1478), .Y(new_n11219));
  nand_4 g10843(.A(n10990), .B(n5767), .Y(new_n11220));
  nand_4 g10844(.A(new_n11220), .B(new_n11219), .Y(new_n11221));
  not_3  g10845(.A(new_n11221), .Y(new_n11222_1));
  not_3  g10846(.A(new_n11219), .Y(new_n11223));
  not_3  g10847(.A(new_n11220), .Y(new_n11224));
  nand_4 g10848(.A(new_n11224), .B(new_n11223), .Y(new_n11225));
  not_3  g10849(.A(new_n11225), .Y(new_n11226));
  nor_4  g10850(.A(new_n11226), .B(new_n11222_1), .Y(new_n11227));
  xnor_3 g10851(.A(new_n11227), .B(new_n11218), .Y(new_n11228));
  xnor_3 g10852(.A(new_n11228), .B(new_n11217), .Y(new_n11229));
  xnor_3 g10853(.A(new_n11229), .B(new_n11209), .Y(new_n11230));
  nor_4  g10854(.A(new_n1472), .B(new_n1470), .Y(new_n11231));
  nor_4  g10855(.A(new_n1478_1), .B(new_n1473), .Y(new_n11232));
  nor_4  g10856(.A(new_n11232), .B(new_n11231), .Y(new_n11233));
  xnor_3 g10857(.A(new_n11233), .B(new_n11230), .Y(new_n11234));
  not_3  g10858(.A(new_n11234), .Y(new_n11235));
  xor_3  g10859(.A(new_n11235), .B(new_n1482), .Y(new_n11236));
  nor_4  g10860(.A(new_n1485), .B(new_n1469), .Y(new_n11237));
  nor_4  g10861(.A(new_n1490), .B(new_n1486), .Y(new_n11238));
  nor_4  g10862(.A(new_n11238), .B(new_n11237), .Y(new_n11239));
  nand_4 g10863(.A(new_n11239), .B(new_n11236), .Y(new_n11240));
  not_3  g10864(.A(new_n1482), .Y(new_n11241));
  xor_3  g10865(.A(new_n11235), .B(new_n11241), .Y(new_n11242));
  not_3  g10866(.A(new_n11239), .Y(new_n11243));
  nand_4 g10867(.A(new_n11243), .B(new_n11242), .Y(new_n11244));
  nand_4 g10868(.A(new_n11244), .B(new_n11240), .Y(new_n11245));
  xnor_3 g10869(.A(new_n11245), .B(new_n11208), .Y(new_n11246));
  xnor_3 g10870(.A(new_n11246), .B(new_n11174), .Y(new_n11247));
  nor_4  g10871(.A(new_n11247), .B(new_n11131), .Y(new_n11248));
  nand_4 g10872(.A(new_n11247), .B(new_n11131), .Y(new_n11249));
  not_3  g10873(.A(new_n11249), .Y(new_n11250));
  nor_4  g10874(.A(new_n11250), .B(new_n11248), .Y(new_n11251));
  not_3  g10875(.A(new_n1427), .Y(new_n11252));
  nand_4 g10876(.A(new_n1501), .B(new_n1430), .Y(new_n11253));
  nand_4 g10877(.A(new_n11253), .B(new_n11252), .Y(new_n11254));
  xor_3  g10878(.A(new_n11254), .B(new_n11251), .Y(n4333));
  nand_4 g10879(.A(n11877), .B(n11757), .Y(new_n11256));
  not_3  g10880(.A(new_n11256), .Y(new_n11257_1));
  nand_4 g10881(.A(n5240), .B(n5212), .Y(new_n11258));
  nand_4 g10882(.A(n11821), .B(n11407), .Y(new_n11259));
  xnor_3 g10883(.A(new_n11259), .B(new_n11258), .Y(new_n11260));
  not_3  g10884(.A(new_n11260), .Y(new_n11261));
  nor_4  g10885(.A(new_n11261), .B(new_n11257_1), .Y(new_n11262));
  nor_4  g10886(.A(new_n11260), .B(new_n11256), .Y(new_n11263));
  nor_4  g10887(.A(new_n11263), .B(new_n11262), .Y(new_n11264));
  not_3  g10888(.A(new_n11264), .Y(new_n11265));
  nand_4 g10889(.A(n11407), .B(n5240), .Y(new_n11266));
  nand_4 g10890(.A(n11877), .B(n3172), .Y(new_n11267));
  nand_4 g10891(.A(new_n11267), .B(new_n11266), .Y(new_n11268));
  not_3  g10892(.A(new_n11268), .Y(new_n11269));
  nand_4 g10893(.A(n11757), .B(n5212), .Y(new_n11270));
  not_3  g10894(.A(new_n11270), .Y(new_n11271));
  xnor_3 g10895(.A(new_n11267), .B(new_n11266), .Y(new_n11272));
  nor_4  g10896(.A(new_n11272), .B(new_n11271), .Y(new_n11273));
  nor_4  g10897(.A(new_n11273), .B(new_n11269), .Y(new_n11274));
  nor_4  g10898(.A(new_n11274), .B(new_n11265), .Y(new_n11275));
  not_3  g10899(.A(new_n11274), .Y(new_n11276));
  nor_4  g10900(.A(new_n11276), .B(new_n11264), .Y(new_n11277));
  nor_4  g10901(.A(new_n11277), .B(new_n11275), .Y(new_n11278));
  nand_4 g10902(.A(n5320), .B(n1333), .Y(new_n11279));
  nand_4 g10903(.A(n4370), .B(n3172), .Y(new_n11280));
  xor_3  g10904(.A(new_n11280), .B(new_n11279), .Y(new_n11281));
  xnor_3 g10905(.A(new_n11281), .B(new_n11278), .Y(new_n11282));
  nand_4 g10906(.A(n4370), .B(n1333), .Y(new_n11283));
  not_3  g10907(.A(new_n11283), .Y(new_n11284));
  nand_4 g10908(.A(n11877), .B(n1333), .Y(new_n11285));
  not_3  g10909(.A(new_n11285), .Y(new_n11286));
  nand_4 g10910(.A(n11757), .B(n11407), .Y(new_n11287));
  not_3  g10911(.A(new_n11287), .Y(new_n11288));
  nor_4  g10912(.A(new_n11288), .B(new_n11286), .Y(new_n11289));
  nand_4 g10913(.A(n5212), .B(n3172), .Y(new_n11290));
  not_3  g10914(.A(new_n11290), .Y(new_n11291));
  xnor_3 g10915(.A(new_n11287), .B(new_n11285), .Y(new_n11292));
  nor_4  g10916(.A(new_n11292), .B(new_n11291), .Y(new_n11293));
  nor_4  g10917(.A(new_n11293), .B(new_n11289), .Y(new_n11294));
  nand_4 g10918(.A(new_n11294), .B(new_n11284), .Y(new_n11295));
  not_3  g10919(.A(new_n11295), .Y(new_n11296_1));
  nor_4  g10920(.A(new_n11294), .B(new_n11284), .Y(new_n11297));
  nor_4  g10921(.A(new_n11297), .B(new_n11296_1), .Y(new_n11298));
  xor_3  g10922(.A(new_n11272), .B(new_n11270), .Y(new_n11299));
  nand_4 g10923(.A(new_n11299), .B(new_n11298), .Y(new_n11300));
  nand_4 g10924(.A(new_n11300), .B(new_n11295), .Y(new_n11301));
  nand_4 g10925(.A(new_n11301), .B(new_n11282), .Y(new_n11302));
  not_3  g10926(.A(new_n11302), .Y(new_n11303));
  nor_4  g10927(.A(new_n11301), .B(new_n11282), .Y(new_n11304));
  nor_4  g10928(.A(new_n11304), .B(new_n11303), .Y(new_n11305));
  not_3  g10929(.A(new_n11305), .Y(new_n11306));
  nand_4 g10930(.A(n7862), .B(n5320), .Y(new_n11307));
  xnor_3 g10931(.A(new_n11299), .B(new_n11298), .Y(new_n11308));
  nand_4 g10932(.A(new_n11308), .B(new_n11307), .Y(new_n11309));
  xnor_3 g10933(.A(new_n11308), .B(new_n11307), .Y(new_n11310));
  not_3  g10934(.A(new_n11310), .Y(new_n11311_1));
  nand_4 g10935(.A(n7862), .B(n4370), .Y(new_n11312));
  not_3  g10936(.A(new_n11312), .Y(new_n11313));
  nand_4 g10937(.A(n11407), .B(n3172), .Y(new_n11314));
  not_3  g10938(.A(new_n11314), .Y(new_n11315));
  nand_4 g10939(.A(n11877), .B(n7862), .Y(new_n11316));
  not_3  g10940(.A(new_n11316), .Y(new_n11317));
  nor_4  g10941(.A(new_n11317), .B(new_n11315), .Y(new_n11318));
  nand_4 g10942(.A(n11407), .B(n7862), .Y(new_n11319));
  nor_4  g10943(.A(new_n11319), .B(new_n11267), .Y(new_n11320));
  nand_4 g10944(.A(n5212), .B(n1333), .Y(new_n11321));
  not_3  g10945(.A(new_n11321), .Y(new_n11322));
  nor_4  g10946(.A(new_n11322), .B(new_n11320), .Y(new_n11323));
  nor_4  g10947(.A(new_n11323), .B(new_n11318), .Y(new_n11324));
  and_4  g10948(.A(new_n11324), .B(new_n11313), .Y(new_n11325));
  not_3  g10949(.A(new_n11325), .Y(new_n11326_1));
  xor_3  g10950(.A(new_n11324), .B(new_n11312), .Y(new_n11327));
  xor_3  g10951(.A(new_n11292), .B(new_n11291), .Y(new_n11328));
  nor_4  g10952(.A(new_n11328), .B(new_n11327), .Y(new_n11329));
  not_3  g10953(.A(new_n11329), .Y(new_n11330));
  nand_4 g10954(.A(new_n11330), .B(new_n11326_1), .Y(new_n11331));
  not_3  g10955(.A(new_n11331), .Y(new_n11332));
  nand_4 g10956(.A(new_n11332), .B(new_n11311_1), .Y(new_n11333));
  nand_4 g10957(.A(new_n11333), .B(new_n11309), .Y(new_n11334));
  nor_4  g10958(.A(new_n11334), .B(new_n11306), .Y(new_n11335));
  not_3  g10959(.A(new_n11335), .Y(new_n11336));
  not_3  g10960(.A(new_n11278), .Y(new_n11337));
  nand_4 g10961(.A(new_n11281), .B(new_n11337), .Y(new_n11338));
  nor_4  g10962(.A(new_n11280), .B(new_n11279), .Y(new_n11339));
  xnor_3 g10963(.A(new_n11303), .B(new_n11339), .Y(new_n11340));
  nand_4 g10964(.A(new_n11340), .B(new_n11338), .Y(new_n11341));
  nor_4  g10965(.A(new_n11259), .B(new_n11258), .Y(new_n11342));
  nand_4 g10966(.A(n11757), .B(n4370), .Y(new_n11343));
  not_3  g10967(.A(new_n11343), .Y(new_n11344));
  xor_3  g10968(.A(new_n11344), .B(new_n11342), .Y(new_n11345));
  nand_4 g10969(.A(n11821), .B(n5212), .Y(new_n11346));
  not_3  g10970(.A(new_n11346), .Y(new_n11347));
  nand_4 g10971(.A(n11877), .B(n5240), .Y(new_n11348));
  nand_4 g10972(.A(n11407), .B(n9080), .Y(new_n11349));
  not_3  g10973(.A(new_n11349), .Y(new_n11350));
  xor_3  g10974(.A(new_n11350), .B(new_n11348), .Y(new_n11351));
  xnor_3 g10975(.A(new_n11351), .B(new_n11347), .Y(new_n11352));
  xnor_3 g10976(.A(new_n11352), .B(new_n11345), .Y(new_n11353));
  nor_4  g10977(.A(new_n11275), .B(new_n11262), .Y(new_n11354));
  nand_4 g10978(.A(n12000), .B(n1333), .Y(new_n11355));
  nand_4 g10979(.A(n5320), .B(n3172), .Y(new_n11356));
  nand_4 g10980(.A(n9725), .B(n7862), .Y(new_n11357));
  not_3  g10981(.A(new_n11357), .Y(new_n11358));
  xor_3  g10982(.A(new_n11358), .B(new_n11356), .Y(new_n11359));
  xnor_3 g10983(.A(new_n11359), .B(new_n11355), .Y(new_n11360));
  xnor_3 g10984(.A(new_n11360), .B(new_n11354), .Y(new_n11361));
  xnor_3 g10985(.A(new_n11361), .B(new_n11353), .Y(new_n11362));
  xor_3  g10986(.A(new_n11362), .B(new_n11341), .Y(new_n11363));
  xnor_3 g10987(.A(new_n11363), .B(new_n11336), .Y(new_n11364));
  nand_4 g10988(.A(n12000), .B(n7862), .Y(new_n11365));
  not_3  g10989(.A(new_n11365), .Y(new_n11366));
  not_3  g10990(.A(new_n11334), .Y(new_n11367));
  nor_4  g10991(.A(new_n11367), .B(new_n11305), .Y(new_n11368));
  nor_4  g10992(.A(new_n11368), .B(new_n11335), .Y(new_n11369));
  nor_4  g10993(.A(new_n11369), .B(new_n11366), .Y(new_n11370));
  nor_4  g10994(.A(new_n11320), .B(new_n11318), .Y(new_n11371));
  nand_4 g10995(.A(n11407), .B(n1333), .Y(new_n11372));
  nand_4 g10996(.A(n7862), .B(n5212), .Y(new_n11373));
  nor_4  g10997(.A(new_n11373), .B(new_n11372), .Y(new_n11374));
  not_3  g10998(.A(new_n11374), .Y(new_n11375));
  nor_4  g10999(.A(new_n11375), .B(new_n11371), .Y(new_n11376));
  not_3  g11000(.A(new_n11376), .Y(new_n11377));
  xnor_3 g11001(.A(new_n11328), .B(new_n11327), .Y(new_n11378));
  nor_4  g11002(.A(new_n11378), .B(new_n11377), .Y(new_n11379));
  xor_3  g11003(.A(new_n11331), .B(new_n11311_1), .Y(new_n11380));
  nand_4 g11004(.A(new_n11380), .B(new_n11379), .Y(new_n11381));
  not_3  g11005(.A(new_n11381), .Y(new_n11382));
  xnor_3 g11006(.A(new_n11369), .B(new_n11366), .Y(new_n11383));
  nor_4  g11007(.A(new_n11383), .B(new_n11382), .Y(new_n11384));
  nor_4  g11008(.A(new_n11384), .B(new_n11370), .Y(new_n11385));
  xnor_3 g11009(.A(new_n11385), .B(new_n11364), .Y(new_n11386));
  nand_4 g11010(.A(n11311), .B(n6429), .Y(new_n11387));
  nand_4 g11011(.A(n12709), .B(n4203), .Y(new_n11388));
  nand_4 g11012(.A(n11728), .B(n4187), .Y(new_n11389));
  xnor_3 g11013(.A(new_n11389), .B(new_n11388), .Y(new_n11390));
  nor_4  g11014(.A(new_n11390), .B(new_n11387), .Y(new_n11391));
  not_3  g11015(.A(new_n11387), .Y(new_n11392));
  not_3  g11016(.A(new_n11390), .Y(new_n11393));
  nor_4  g11017(.A(new_n11393), .B(new_n11392), .Y(new_n11394));
  nor_4  g11018(.A(new_n11394), .B(new_n11391), .Y(new_n11395));
  nand_4 g11019(.A(n12709), .B(n4187), .Y(new_n11396));
  nand_4 g11020(.A(n6429), .B(n2464), .Y(new_n11397));
  and_4  g11021(.A(new_n11397), .B(new_n11396), .Y(new_n11398));
  nand_4 g11022(.A(n11728), .B(n11311), .Y(new_n11399));
  not_3  g11023(.A(new_n11399), .Y(new_n11400));
  xnor_3 g11024(.A(new_n11397), .B(new_n11396), .Y(new_n11401));
  nor_4  g11025(.A(new_n11401), .B(new_n11400), .Y(new_n11402));
  nor_4  g11026(.A(new_n11402), .B(new_n11398), .Y(new_n11403));
  xnor_3 g11027(.A(new_n11403), .B(new_n11395), .Y(new_n11404));
  nand_4 g11028(.A(n9400), .B(n2433), .Y(new_n11405));
  nand_4 g11029(.A(n8819), .B(n2464), .Y(new_n11406));
  xor_3  g11030(.A(new_n11406), .B(new_n11405), .Y(new_n11407_1));
  not_3  g11031(.A(new_n11407_1), .Y(new_n11408));
  nor_4  g11032(.A(new_n11408), .B(new_n11404), .Y(new_n11409));
  not_3  g11033(.A(new_n11404), .Y(new_n11410));
  nor_4  g11034(.A(new_n11407_1), .B(new_n11410), .Y(new_n11411));
  nor_4  g11035(.A(new_n11411), .B(new_n11409), .Y(new_n11412));
  nand_4 g11036(.A(n9400), .B(n8819), .Y(new_n11413));
  not_3  g11037(.A(new_n11413), .Y(new_n11414));
  nand_4 g11038(.A(n12709), .B(n11311), .Y(new_n11415));
  not_3  g11039(.A(new_n11415), .Y(new_n11416));
  nand_4 g11040(.A(n9400), .B(n6429), .Y(new_n11417));
  not_3  g11041(.A(new_n11417), .Y(new_n11418));
  nor_4  g11042(.A(new_n11418), .B(new_n11416), .Y(new_n11419));
  nand_4 g11043(.A(n11728), .B(n2464), .Y(new_n11420));
  not_3  g11044(.A(new_n11420), .Y(new_n11421));
  xnor_3 g11045(.A(new_n11417), .B(new_n11415), .Y(new_n11422));
  nor_4  g11046(.A(new_n11422), .B(new_n11421), .Y(new_n11423_1));
  nor_4  g11047(.A(new_n11423_1), .B(new_n11419), .Y(new_n11424));
  nand_4 g11048(.A(new_n11424), .B(new_n11414), .Y(new_n11425));
  not_3  g11049(.A(new_n11425), .Y(new_n11426));
  xnor_3 g11050(.A(new_n11424), .B(new_n11414), .Y(new_n11427));
  xnor_3 g11051(.A(new_n11401), .B(new_n11399), .Y(new_n11428));
  nor_4  g11052(.A(new_n11428), .B(new_n11427), .Y(new_n11429));
  nor_4  g11053(.A(new_n11429), .B(new_n11426), .Y(new_n11430));
  not_3  g11054(.A(new_n11430), .Y(new_n11431));
  xnor_3 g11055(.A(new_n11431), .B(new_n11412), .Y(new_n11432));
  nand_4 g11056(.A(n6877), .B(n2433), .Y(new_n11433));
  xnor_3 g11057(.A(new_n11428), .B(new_n11427), .Y(new_n11434));
  nor_4  g11058(.A(new_n11434), .B(new_n11433), .Y(new_n11435));
  not_3  g11059(.A(new_n11435), .Y(new_n11436));
  not_3  g11060(.A(new_n11433), .Y(new_n11437));
  not_3  g11061(.A(new_n11434), .Y(new_n11438));
  nor_4  g11062(.A(new_n11438), .B(new_n11437), .Y(new_n11439));
  nor_4  g11063(.A(new_n11439), .B(new_n11435), .Y(new_n11440));
  nand_4 g11064(.A(n8819), .B(n6877), .Y(new_n11441));
  not_3  g11065(.A(new_n11441), .Y(new_n11442));
  nand_4 g11066(.A(n12709), .B(n2464), .Y(new_n11443));
  not_3  g11067(.A(new_n11443), .Y(new_n11444));
  nand_4 g11068(.A(n6877), .B(n6429), .Y(new_n11445));
  not_3  g11069(.A(new_n11445), .Y(new_n11446));
  nor_4  g11070(.A(new_n11446), .B(new_n11444), .Y(new_n11447));
  nor_4  g11071(.A(new_n11445), .B(new_n11443), .Y(new_n11448));
  nand_4 g11072(.A(n11728), .B(n9400), .Y(new_n11449));
  not_3  g11073(.A(new_n11449), .Y(new_n11450));
  nor_4  g11074(.A(new_n11450), .B(new_n11448), .Y(new_n11451));
  nor_4  g11075(.A(new_n11451), .B(new_n11447), .Y(new_n11452));
  nand_4 g11076(.A(new_n11452), .B(new_n11442), .Y(new_n11453));
  not_3  g11077(.A(new_n11453), .Y(new_n11454));
  xnor_3 g11078(.A(new_n11452), .B(new_n11442), .Y(new_n11455));
  and_4  g11079(.A(new_n11422), .B(new_n11421), .Y(new_n11456));
  nor_4  g11080(.A(new_n11456), .B(new_n11423_1), .Y(new_n11457));
  nor_4  g11081(.A(new_n11457), .B(new_n11455), .Y(new_n11458));
  nor_4  g11082(.A(new_n11458), .B(new_n11454), .Y(new_n11459));
  not_3  g11083(.A(new_n11459), .Y(new_n11460));
  nand_4 g11084(.A(new_n11460), .B(new_n11440), .Y(new_n11461));
  nand_4 g11085(.A(new_n11461), .B(new_n11436), .Y(new_n11462));
  not_3  g11086(.A(new_n11462), .Y(new_n11463));
  nor_4  g11087(.A(new_n11463), .B(new_n11432), .Y(new_n11464));
  not_3  g11088(.A(new_n11409), .Y(new_n11465));
  nor_4  g11089(.A(new_n11406), .B(new_n11405), .Y(new_n11466));
  nand_4 g11090(.A(new_n11431), .B(new_n11412), .Y(new_n11467));
  not_3  g11091(.A(new_n11467), .Y(new_n11468));
  xnor_3 g11092(.A(new_n11468), .B(new_n11466), .Y(new_n11469));
  nand_4 g11093(.A(new_n11469), .B(new_n11465), .Y(new_n11470));
  not_3  g11094(.A(new_n11391), .Y(new_n11471));
  nand_4 g11095(.A(new_n11403), .B(new_n11395), .Y(new_n11472));
  nand_4 g11096(.A(new_n11472), .B(new_n11471), .Y(new_n11473));
  nand_4 g11097(.A(n9400), .B(n8717), .Y(new_n11474));
  not_3  g11098(.A(new_n11474), .Y(new_n11475));
  nand_4 g11099(.A(n2464), .B(n2433), .Y(new_n11476));
  nand_4 g11100(.A(n7730), .B(n6877), .Y(new_n11477));
  not_3  g11101(.A(new_n11477), .Y(new_n11478_1));
  xor_3  g11102(.A(new_n11478_1), .B(new_n11476), .Y(new_n11479));
  xnor_3 g11103(.A(new_n11479), .B(new_n11475), .Y(new_n11480));
  xnor_3 g11104(.A(new_n11480), .B(new_n11473), .Y(new_n11481));
  nor_4  g11105(.A(new_n11389), .B(new_n11388), .Y(new_n11482));
  not_3  g11106(.A(new_n11482), .Y(new_n11483));
  nand_4 g11107(.A(n11311), .B(n8819), .Y(new_n11484));
  xor_3  g11108(.A(new_n11484), .B(new_n11483), .Y(new_n11485));
  nand_4 g11109(.A(n11728), .B(n4203), .Y(new_n11486));
  nand_4 g11110(.A(n6429), .B(n4187), .Y(new_n11487));
  nand_4 g11111(.A(n12753), .B(n12709), .Y(new_n11488));
  not_3  g11112(.A(new_n11488), .Y(new_n11489));
  xor_3  g11113(.A(new_n11489), .B(new_n11487), .Y(new_n11490));
  xnor_3 g11114(.A(new_n11490), .B(new_n11486), .Y(new_n11491));
  xnor_3 g11115(.A(new_n11491), .B(new_n11485), .Y(new_n11492));
  xnor_3 g11116(.A(new_n11492), .B(new_n11481), .Y(new_n11493));
  xnor_3 g11117(.A(new_n11493), .B(new_n11470), .Y(new_n11494));
  xnor_3 g11118(.A(new_n11494), .B(new_n11464), .Y(new_n11495));
  not_3  g11119(.A(new_n11495), .Y(new_n11496));
  nand_4 g11120(.A(n8717), .B(n6877), .Y(new_n11497));
  not_3  g11121(.A(new_n11497), .Y(new_n11498));
  not_3  g11122(.A(new_n11432), .Y(new_n11499));
  nor_4  g11123(.A(new_n11462), .B(new_n11499), .Y(new_n11500));
  nor_4  g11124(.A(new_n11500), .B(new_n11464), .Y(new_n11501));
  nand_4 g11125(.A(new_n11501), .B(new_n11498), .Y(new_n11502));
  nor_4  g11126(.A(new_n11448), .B(new_n11447), .Y(new_n11503));
  nand_4 g11127(.A(n12709), .B(n9400), .Y(new_n11504));
  nand_4 g11128(.A(n11728), .B(n6877), .Y(new_n11505));
  nor_4  g11129(.A(new_n11505), .B(new_n11504), .Y(new_n11506));
  not_3  g11130(.A(new_n11506), .Y(new_n11507));
  nor_4  g11131(.A(new_n11507), .B(new_n11503), .Y(new_n11508));
  not_3  g11132(.A(new_n11508), .Y(new_n11509));
  xnor_3 g11133(.A(new_n11457), .B(new_n11455), .Y(new_n11510));
  nor_4  g11134(.A(new_n11510), .B(new_n11509), .Y(new_n11511));
  not_3  g11135(.A(new_n11511), .Y(new_n11512));
  xnor_3 g11136(.A(new_n11460), .B(new_n11440), .Y(new_n11513));
  nor_4  g11137(.A(new_n11513), .B(new_n11512), .Y(new_n11514));
  xnor_3 g11138(.A(new_n11501), .B(new_n11497), .Y(new_n11515));
  nand_4 g11139(.A(new_n11515), .B(new_n11514), .Y(new_n11516));
  nand_4 g11140(.A(new_n11516), .B(new_n11502), .Y(new_n11517));
  xnor_3 g11141(.A(new_n11517), .B(new_n11496), .Y(new_n11518));
  nand_4 g11142(.A(n11478), .B(n6254), .Y(new_n11519));
  not_3  g11143(.A(new_n11519), .Y(new_n11520));
  nand_4 g11144(.A(n12489), .B(n137), .Y(new_n11521));
  not_3  g11145(.A(new_n11521), .Y(new_n11522));
  nand_4 g11146(.A(n12777), .B(n11478), .Y(new_n11523));
  not_3  g11147(.A(new_n11523), .Y(new_n11524));
  nor_4  g11148(.A(new_n11524), .B(new_n11522), .Y(new_n11525));
  nand_4 g11149(.A(n7159), .B(n5283), .Y(new_n11526));
  not_3  g11150(.A(new_n11526), .Y(new_n11527));
  xnor_3 g11151(.A(new_n11523), .B(new_n11521), .Y(new_n11528));
  nor_4  g11152(.A(new_n11528), .B(new_n11527), .Y(new_n11529));
  nor_4  g11153(.A(new_n11529), .B(new_n11525), .Y(new_n11530));
  nand_4 g11154(.A(new_n11530), .B(new_n11520), .Y(new_n11531));
  nand_4 g11155(.A(n7159), .B(n137), .Y(new_n11532));
  not_3  g11156(.A(new_n11532), .Y(new_n11533));
  nand_4 g11157(.A(n12489), .B(n6294), .Y(new_n11534));
  nand_4 g11158(.A(n12777), .B(n5283), .Y(new_n11535));
  xnor_3 g11159(.A(new_n11535), .B(new_n11534), .Y(new_n11536_1));
  xnor_3 g11160(.A(new_n11536_1), .B(new_n11533), .Y(new_n11537));
  xnor_3 g11161(.A(new_n11530), .B(new_n11519), .Y(new_n11538));
  nand_4 g11162(.A(new_n11538), .B(new_n11537), .Y(new_n11539));
  nand_4 g11163(.A(new_n11539), .B(new_n11531), .Y(new_n11540));
  nand_4 g11164(.A(n11967), .B(n11478), .Y(new_n11541));
  nand_4 g11165(.A(n6254), .B(n5283), .Y(new_n11542));
  nor_4  g11166(.A(new_n11542), .B(new_n11541), .Y(new_n11543));
  and_4  g11167(.A(new_n11542), .B(new_n11541), .Y(new_n11544));
  nor_4  g11168(.A(new_n11544), .B(new_n11543), .Y(new_n11545));
  not_3  g11169(.A(new_n11545), .Y(new_n11546));
  xnor_3 g11170(.A(new_n11546), .B(new_n11540), .Y(new_n11547));
  nand_4 g11171(.A(n12777), .B(n137), .Y(new_n11548));
  nand_4 g11172(.A(n7159), .B(n6294), .Y(new_n11549));
  nand_4 g11173(.A(n12489), .B(n6797), .Y(new_n11550));
  xnor_3 g11174(.A(new_n11550), .B(new_n11549), .Y(new_n11551));
  nor_4  g11175(.A(new_n11551), .B(new_n11548), .Y(new_n11552));
  not_3  g11176(.A(new_n11548), .Y(new_n11553));
  not_3  g11177(.A(new_n11551), .Y(new_n11554));
  nor_4  g11178(.A(new_n11554), .B(new_n11553), .Y(new_n11555));
  nor_4  g11179(.A(new_n11555), .B(new_n11552), .Y(new_n11556));
  and_4  g11180(.A(new_n11535), .B(new_n11534), .Y(new_n11557));
  nor_4  g11181(.A(new_n11536_1), .B(new_n11533), .Y(new_n11558));
  nor_4  g11182(.A(new_n11558), .B(new_n11557), .Y(new_n11559));
  nand_4 g11183(.A(new_n11559), .B(new_n11556), .Y(new_n11560));
  not_3  g11184(.A(new_n11560), .Y(new_n11561));
  nor_4  g11185(.A(new_n11559), .B(new_n11556), .Y(new_n11562));
  nor_4  g11186(.A(new_n11562), .B(new_n11561), .Y(new_n11563));
  nand_4 g11187(.A(new_n11563), .B(new_n11547), .Y(new_n11564));
  xnor_3 g11188(.A(new_n11545), .B(new_n11540), .Y(new_n11565));
  xnor_3 g11189(.A(new_n11559), .B(new_n11556), .Y(new_n11566));
  nand_4 g11190(.A(new_n11566), .B(new_n11565), .Y(new_n11567));
  nand_4 g11191(.A(new_n11567), .B(new_n11564), .Y(new_n11568));
  nand_4 g11192(.A(n11967), .B(n4805), .Y(new_n11569));
  not_3  g11193(.A(new_n11569), .Y(new_n11570));
  nand_4 g11194(.A(n6254), .B(n4805), .Y(new_n11571));
  not_3  g11195(.A(new_n11571), .Y(new_n11572));
  nand_4 g11196(.A(n12489), .B(n5283), .Y(new_n11573));
  not_3  g11197(.A(new_n11573), .Y(new_n11574));
  nand_4 g11198(.A(n12777), .B(n4805), .Y(new_n11575));
  not_3  g11199(.A(new_n11575), .Y(new_n11576));
  nor_4  g11200(.A(new_n11576), .B(new_n11574), .Y(new_n11577));
  nor_4  g11201(.A(new_n11575), .B(new_n11573), .Y(new_n11578));
  nand_4 g11202(.A(n11478), .B(n7159), .Y(new_n11579));
  not_3  g11203(.A(new_n11579), .Y(new_n11580));
  nor_4  g11204(.A(new_n11580), .B(new_n11578), .Y(new_n11581));
  nor_4  g11205(.A(new_n11581), .B(new_n11577), .Y(new_n11582));
  nand_4 g11206(.A(new_n11582), .B(new_n11572), .Y(new_n11583));
  not_3  g11207(.A(new_n11583), .Y(new_n11584));
  nor_4  g11208(.A(new_n11582), .B(new_n11572), .Y(new_n11585));
  nor_4  g11209(.A(new_n11585), .B(new_n11584), .Y(new_n11586));
  xnor_3 g11210(.A(new_n11528), .B(new_n11526), .Y(new_n11587));
  not_3  g11211(.A(new_n11587), .Y(new_n11588));
  nand_4 g11212(.A(new_n11588), .B(new_n11586), .Y(new_n11589));
  nand_4 g11213(.A(new_n11589), .B(new_n11583), .Y(new_n11590));
  nor_4  g11214(.A(new_n11590), .B(new_n11570), .Y(new_n11591));
  not_3  g11215(.A(new_n11591), .Y(new_n11592));
  not_3  g11216(.A(new_n11539), .Y(new_n11593));
  nor_4  g11217(.A(new_n11538), .B(new_n11537), .Y(new_n11594));
  nor_4  g11218(.A(new_n11594), .B(new_n11593), .Y(new_n11595));
  not_3  g11219(.A(new_n11595), .Y(new_n11596));
  xnor_3 g11220(.A(new_n11590), .B(new_n11569), .Y(new_n11597));
  nand_4 g11221(.A(new_n11597), .B(new_n11596), .Y(new_n11598));
  nand_4 g11222(.A(new_n11598), .B(new_n11592), .Y(new_n11599));
  nor_4  g11223(.A(new_n11599), .B(new_n11568), .Y(new_n11600));
  not_3  g11224(.A(new_n11552), .Y(new_n11601));
  nand_4 g11225(.A(new_n11560), .B(new_n11601), .Y(new_n11602));
  nand_4 g11226(.A(n11478), .B(n447), .Y(new_n11603));
  nand_4 g11227(.A(n11967), .B(n5283), .Y(new_n11604));
  nand_4 g11228(.A(n4805), .B(n1353), .Y(new_n11605));
  nand_4 g11229(.A(new_n11605), .B(new_n11604), .Y(new_n11606));
  not_3  g11230(.A(new_n11604), .Y(new_n11607));
  not_3  g11231(.A(new_n11605), .Y(new_n11608));
  nand_4 g11232(.A(new_n11608), .B(new_n11607), .Y(new_n11609));
  nand_4 g11233(.A(new_n11609), .B(new_n11606), .Y(new_n11610));
  xnor_3 g11234(.A(new_n11610), .B(new_n11603), .Y(new_n11611));
  xnor_3 g11235(.A(new_n11611), .B(new_n11602), .Y(new_n11612));
  nor_4  g11236(.A(new_n11550), .B(new_n11549), .Y(new_n11613));
  not_3  g11237(.A(new_n11613), .Y(new_n11614));
  nand_4 g11238(.A(n6254), .B(n137), .Y(new_n11615));
  xor_3  g11239(.A(new_n11615), .B(new_n11614), .Y(new_n11616));
  nand_4 g11240(.A(n7159), .B(n6797), .Y(new_n11617));
  nand_4 g11241(.A(n12777), .B(n6294), .Y(new_n11618));
  nand_4 g11242(.A(n12489), .B(n3146), .Y(new_n11619));
  xnor_3 g11243(.A(new_n11619), .B(new_n11618), .Y(new_n11620));
  xnor_3 g11244(.A(new_n11620), .B(new_n11617), .Y(new_n11621));
  xnor_3 g11245(.A(new_n11621), .B(new_n11616), .Y(new_n11622));
  xnor_3 g11246(.A(new_n11622), .B(new_n11612), .Y(new_n11623));
  not_3  g11247(.A(new_n11540), .Y(new_n11624));
  nor_4  g11248(.A(new_n11546), .B(new_n11624), .Y(new_n11625));
  not_3  g11249(.A(new_n11625), .Y(new_n11626));
  not_3  g11250(.A(new_n11543), .Y(new_n11627));
  xnor_3 g11251(.A(new_n11564), .B(new_n11627), .Y(new_n11628));
  nand_4 g11252(.A(new_n11628), .B(new_n11626), .Y(new_n11629));
  xnor_3 g11253(.A(new_n11629), .B(new_n11623), .Y(new_n11630));
  xnor_3 g11254(.A(new_n11630), .B(new_n11600), .Y(new_n11631));
  nand_4 g11255(.A(n4805), .B(n447), .Y(new_n11632));
  not_3  g11256(.A(new_n11632), .Y(new_n11633));
  xnor_3 g11257(.A(new_n11590), .B(new_n11570), .Y(new_n11634));
  nor_4  g11258(.A(new_n11634), .B(new_n11595), .Y(new_n11635));
  nor_4  g11259(.A(new_n11635), .B(new_n11591), .Y(new_n11636));
  xnor_3 g11260(.A(new_n11636), .B(new_n11568), .Y(new_n11637));
  nand_4 g11261(.A(new_n11637), .B(new_n11633), .Y(new_n11638));
  nor_4  g11262(.A(new_n11578), .B(new_n11577), .Y(new_n11639));
  nand_4 g11263(.A(n12489), .B(n11478), .Y(new_n11640));
  nand_4 g11264(.A(n7159), .B(n4805), .Y(new_n11641));
  nor_4  g11265(.A(new_n11641), .B(new_n11640), .Y(new_n11642));
  not_3  g11266(.A(new_n11642), .Y(new_n11643));
  nor_4  g11267(.A(new_n11643), .B(new_n11639), .Y(new_n11644));
  not_3  g11268(.A(new_n11644), .Y(new_n11645));
  xnor_3 g11269(.A(new_n11588), .B(new_n11586), .Y(new_n11646));
  nor_4  g11270(.A(new_n11646), .B(new_n11645), .Y(new_n11647));
  xnor_3 g11271(.A(new_n11634), .B(new_n11595), .Y(new_n11648));
  nand_4 g11272(.A(new_n11648), .B(new_n11647), .Y(new_n11649));
  not_3  g11273(.A(new_n11649), .Y(new_n11650));
  xnor_3 g11274(.A(new_n11637), .B(new_n11632), .Y(new_n11651));
  nand_4 g11275(.A(new_n11651), .B(new_n11650), .Y(new_n11652));
  nand_4 g11276(.A(new_n11652), .B(new_n11638), .Y(new_n11653));
  xnor_3 g11277(.A(new_n11653), .B(new_n11631), .Y(new_n11654));
  nand_4 g11278(.A(n11791), .B(n3992), .Y(new_n11655));
  not_3  g11279(.A(new_n11655), .Y(new_n11656));
  nand_4 g11280(.A(n10990), .B(n6358), .Y(new_n11657));
  not_3  g11281(.A(new_n11657), .Y(new_n11658));
  nand_4 g11282(.A(n3992), .B(n1478), .Y(new_n11659));
  not_3  g11283(.A(new_n11659), .Y(new_n11660));
  nor_4  g11284(.A(new_n11660), .B(new_n11658), .Y(new_n11661));
  nand_4 g11285(.A(n8384), .B(n5760), .Y(new_n11662_1));
  not_3  g11286(.A(new_n11662_1), .Y(new_n11663));
  xnor_3 g11287(.A(new_n11659), .B(new_n11657), .Y(new_n11664));
  nor_4  g11288(.A(new_n11664), .B(new_n11663), .Y(new_n11665));
  nor_4  g11289(.A(new_n11665), .B(new_n11661), .Y(new_n11666));
  nand_4 g11290(.A(new_n11666), .B(new_n11656), .Y(new_n11667));
  nand_4 g11291(.A(n6358), .B(n5760), .Y(new_n11668));
  not_3  g11292(.A(new_n11668), .Y(new_n11669));
  nand_4 g11293(.A(n10990), .B(n5198), .Y(new_n11670));
  nand_4 g11294(.A(n8384), .B(n1478), .Y(new_n11671));
  xnor_3 g11295(.A(new_n11671), .B(new_n11670), .Y(new_n11672));
  xnor_3 g11296(.A(new_n11672), .B(new_n11669), .Y(new_n11673));
  xnor_3 g11297(.A(new_n11666), .B(new_n11655), .Y(new_n11674));
  nand_4 g11298(.A(new_n11674), .B(new_n11673), .Y(new_n11675));
  nand_4 g11299(.A(new_n11675), .B(new_n11667), .Y(new_n11676));
  nand_4 g11300(.A(n12947), .B(n3992), .Y(new_n11677));
  not_3  g11301(.A(new_n11677), .Y(new_n11678));
  nand_4 g11302(.A(n11791), .B(n8384), .Y(new_n11679));
  not_3  g11303(.A(new_n11679), .Y(new_n11680));
  nor_4  g11304(.A(new_n11680), .B(new_n11678), .Y(new_n11681));
  nor_4  g11305(.A(new_n11679), .B(new_n11677), .Y(new_n11682));
  nor_4  g11306(.A(new_n11682), .B(new_n11681), .Y(new_n11683));
  not_3  g11307(.A(new_n11683), .Y(new_n11684));
  xnor_3 g11308(.A(new_n11684), .B(new_n11676), .Y(new_n11685));
  nand_4 g11309(.A(n6358), .B(n1478), .Y(new_n11686));
  nand_4 g11310(.A(n5760), .B(n5198), .Y(new_n11687));
  nand_4 g11311(.A(n10990), .B(n1471), .Y(new_n11688));
  xnor_3 g11312(.A(new_n11688), .B(new_n11687), .Y(new_n11689));
  nor_4  g11313(.A(new_n11689), .B(new_n11686), .Y(new_n11690));
  not_3  g11314(.A(new_n11686), .Y(new_n11691));
  not_3  g11315(.A(new_n11689), .Y(new_n11692));
  nor_4  g11316(.A(new_n11692), .B(new_n11691), .Y(new_n11693));
  nor_4  g11317(.A(new_n11693), .B(new_n11690), .Y(new_n11694));
  not_3  g11318(.A(new_n11694), .Y(new_n11695));
  and_4  g11319(.A(new_n11671), .B(new_n11670), .Y(new_n11696));
  nor_4  g11320(.A(new_n11672), .B(new_n11669), .Y(new_n11697));
  nor_4  g11321(.A(new_n11697), .B(new_n11696), .Y(new_n11698));
  xnor_3 g11322(.A(new_n11698), .B(new_n11695), .Y(new_n11699));
  nand_4 g11323(.A(new_n11699), .B(new_n11685), .Y(new_n11700));
  xnor_3 g11324(.A(new_n11683), .B(new_n11676), .Y(new_n11701));
  xnor_3 g11325(.A(new_n11698), .B(new_n11694), .Y(new_n11702));
  nand_4 g11326(.A(new_n11702), .B(new_n11701), .Y(new_n11703));
  nand_4 g11327(.A(new_n11703), .B(new_n11700), .Y(new_n11704));
  nand_4 g11328(.A(n12947), .B(n7236), .Y(new_n11705));
  not_3  g11329(.A(new_n11705), .Y(new_n11706));
  nand_4 g11330(.A(n11791), .B(n7236), .Y(new_n11707_1));
  not_3  g11331(.A(new_n11707_1), .Y(new_n11708));
  nand_4 g11332(.A(n10990), .B(n8384), .Y(new_n11709));
  nand_4 g11333(.A(n7236), .B(n1478), .Y(new_n11710));
  nand_4 g11334(.A(new_n11710), .B(new_n11709), .Y(new_n11711));
  not_3  g11335(.A(new_n11711), .Y(new_n11712));
  nor_4  g11336(.A(new_n11710), .B(new_n11709), .Y(new_n11713));
  nand_4 g11337(.A(n5760), .B(n3992), .Y(new_n11714));
  not_3  g11338(.A(new_n11714), .Y(new_n11715));
  nor_4  g11339(.A(new_n11715), .B(new_n11713), .Y(new_n11716));
  nor_4  g11340(.A(new_n11716), .B(new_n11712), .Y(new_n11717));
  nand_4 g11341(.A(new_n11717), .B(new_n11708), .Y(new_n11718));
  not_3  g11342(.A(new_n11718), .Y(new_n11719));
  nor_4  g11343(.A(new_n11717), .B(new_n11708), .Y(new_n11720));
  nor_4  g11344(.A(new_n11720), .B(new_n11719), .Y(new_n11721));
  xnor_3 g11345(.A(new_n11664), .B(new_n11662_1), .Y(new_n11722));
  not_3  g11346(.A(new_n11722), .Y(new_n11723));
  nand_4 g11347(.A(new_n11723), .B(new_n11721), .Y(new_n11724));
  nand_4 g11348(.A(new_n11724), .B(new_n11718), .Y(new_n11725));
  nor_4  g11349(.A(new_n11725), .B(new_n11706), .Y(new_n11726));
  not_3  g11350(.A(new_n11726), .Y(new_n11727));
  not_3  g11351(.A(new_n11675), .Y(new_n11728_1));
  nor_4  g11352(.A(new_n11674), .B(new_n11673), .Y(new_n11729));
  nor_4  g11353(.A(new_n11729), .B(new_n11728_1), .Y(new_n11730));
  not_3  g11354(.A(new_n11730), .Y(new_n11731));
  xnor_3 g11355(.A(new_n11725), .B(new_n11705), .Y(new_n11732));
  nand_4 g11356(.A(new_n11732), .B(new_n11731), .Y(new_n11733));
  nand_4 g11357(.A(new_n11733), .B(new_n11727), .Y(new_n11734));
  nor_4  g11358(.A(new_n11734), .B(new_n11704), .Y(new_n11735));
  not_3  g11359(.A(new_n11690), .Y(new_n11736));
  nand_4 g11360(.A(new_n11698), .B(new_n11694), .Y(new_n11737));
  nand_4 g11361(.A(new_n11737), .B(new_n11736), .Y(new_n11738));
  nand_4 g11362(.A(n6441), .B(n3992), .Y(new_n11739));
  not_3  g11363(.A(new_n11739), .Y(new_n11740));
  nand_4 g11364(.A(n12947), .B(n8384), .Y(new_n11741));
  nand_4 g11365(.A(n11999), .B(n7236), .Y(new_n11742));
  xnor_3 g11366(.A(new_n11742), .B(new_n11741), .Y(new_n11743));
  and_4  g11367(.A(new_n11743), .B(new_n11740), .Y(new_n11744));
  nor_4  g11368(.A(new_n11743), .B(new_n11740), .Y(new_n11745));
  nor_4  g11369(.A(new_n11745), .B(new_n11744), .Y(new_n11746));
  xnor_3 g11370(.A(new_n11746), .B(new_n11738), .Y(new_n11747));
  nor_4  g11371(.A(new_n11688), .B(new_n11687), .Y(new_n11748));
  nand_4 g11372(.A(n11791), .B(n6358), .Y(new_n11749));
  not_3  g11373(.A(new_n11749), .Y(new_n11750));
  xor_3  g11374(.A(new_n11750), .B(new_n11748), .Y(new_n11751));
  nand_4 g11375(.A(n5760), .B(n1471), .Y(new_n11752));
  not_3  g11376(.A(new_n11752), .Y(new_n11753));
  nand_4 g11377(.A(n5198), .B(n1478), .Y(new_n11754));
  nand_4 g11378(.A(n10990), .B(n7646), .Y(new_n11755_1));
  xnor_3 g11379(.A(new_n11755_1), .B(new_n11754), .Y(new_n11756));
  and_4  g11380(.A(new_n11756), .B(new_n11753), .Y(new_n11757_1));
  nor_4  g11381(.A(new_n11756), .B(new_n11753), .Y(new_n11758));
  nor_4  g11382(.A(new_n11758), .B(new_n11757_1), .Y(new_n11759));
  xnor_3 g11383(.A(new_n11759), .B(new_n11751), .Y(new_n11760));
  xnor_3 g11384(.A(new_n11760), .B(new_n11747), .Y(new_n11761));
  not_3  g11385(.A(new_n11676), .Y(new_n11762));
  nor_4  g11386(.A(new_n11684), .B(new_n11762), .Y(new_n11763));
  not_3  g11387(.A(new_n11763), .Y(new_n11764));
  not_3  g11388(.A(new_n11682), .Y(new_n11765));
  xnor_3 g11389(.A(new_n11700), .B(new_n11765), .Y(new_n11766));
  nand_4 g11390(.A(new_n11766), .B(new_n11764), .Y(new_n11767));
  xnor_3 g11391(.A(new_n11767), .B(new_n11761), .Y(new_n11768));
  xnor_3 g11392(.A(new_n11768), .B(new_n11735), .Y(new_n11769));
  nand_4 g11393(.A(n7236), .B(n6441), .Y(new_n11770));
  not_3  g11394(.A(new_n11770), .Y(new_n11771));
  xnor_3 g11395(.A(new_n11725), .B(new_n11706), .Y(new_n11772));
  nor_4  g11396(.A(new_n11772), .B(new_n11730), .Y(new_n11773));
  nor_4  g11397(.A(new_n11773), .B(new_n11726), .Y(new_n11774));
  xnor_3 g11398(.A(new_n11774), .B(new_n11704), .Y(new_n11775));
  nand_4 g11399(.A(new_n11775), .B(new_n11771), .Y(new_n11776));
  xnor_3 g11400(.A(new_n11723), .B(new_n11721), .Y(new_n11777));
  nand_4 g11401(.A(n10990), .B(n7236), .Y(new_n11778));
  not_3  g11402(.A(new_n11778), .Y(new_n11779));
  nor_4  g11403(.A(new_n11779), .B(new_n11714), .Y(new_n11780_1));
  nor_4  g11404(.A(new_n11780_1), .B(new_n11711), .Y(new_n11781));
  nor_4  g11405(.A(new_n11781), .B(new_n11713), .Y(new_n11782));
  nor_4  g11406(.A(new_n11782), .B(new_n11714), .Y(new_n11783));
  not_3  g11407(.A(new_n11783), .Y(new_n11784));
  nor_4  g11408(.A(new_n11784), .B(new_n11777), .Y(new_n11785));
  xnor_3 g11409(.A(new_n11772), .B(new_n11730), .Y(new_n11786));
  nand_4 g11410(.A(new_n11786), .B(new_n11785), .Y(new_n11787));
  not_3  g11411(.A(new_n11787), .Y(new_n11788));
  xnor_3 g11412(.A(new_n11775), .B(new_n11770), .Y(new_n11789));
  nand_4 g11413(.A(new_n11789), .B(new_n11788), .Y(new_n11790));
  nand_4 g11414(.A(new_n11790), .B(new_n11776), .Y(new_n11791_1));
  xnor_3 g11415(.A(new_n11791_1), .B(new_n11769), .Y(new_n11792));
  nand_4 g11416(.A(new_n11792), .B(new_n11654), .Y(new_n11793));
  not_3  g11417(.A(new_n11600), .Y(new_n11794));
  xnor_3 g11418(.A(new_n11630), .B(new_n11794), .Y(new_n11795));
  xnor_3 g11419(.A(new_n11653), .B(new_n11795), .Y(new_n11796));
  not_3  g11420(.A(new_n11735), .Y(new_n11797));
  xnor_3 g11421(.A(new_n11768), .B(new_n11797), .Y(new_n11798));
  xnor_3 g11422(.A(new_n11791_1), .B(new_n11798), .Y(new_n11799));
  nand_4 g11423(.A(new_n11799), .B(new_n11796), .Y(new_n11800));
  nand_4 g11424(.A(new_n11800), .B(new_n11793), .Y(new_n11801));
  xnor_3 g11425(.A(new_n11599), .B(new_n11568), .Y(new_n11802));
  nand_4 g11426(.A(new_n11802), .B(new_n11632), .Y(new_n11803));
  nand_4 g11427(.A(new_n11803), .B(new_n11638), .Y(new_n11804));
  xnor_3 g11428(.A(new_n11804), .B(new_n11650), .Y(new_n11805));
  not_3  g11429(.A(new_n11805), .Y(new_n11806));
  xnor_3 g11430(.A(new_n11648), .B(new_n11647), .Y(new_n11807));
  xnor_3 g11431(.A(new_n11786), .B(new_n11785), .Y(new_n11808));
  nor_4  g11432(.A(new_n11808), .B(new_n11807), .Y(new_n11809));
  xnor_3 g11433(.A(new_n11808), .B(new_n11807), .Y(new_n11810));
  xnor_3 g11434(.A(new_n11646), .B(new_n11644), .Y(new_n11811));
  xnor_3 g11435(.A(new_n11783), .B(new_n11777), .Y(new_n11812));
  nor_4  g11436(.A(new_n11812), .B(new_n11811), .Y(new_n11813));
  not_3  g11437(.A(new_n11813), .Y(new_n11814));
  nand_4 g11438(.A(n12489), .B(n4805), .Y(new_n11815));
  not_3  g11439(.A(new_n11815), .Y(new_n11816));
  nand_4 g11440(.A(new_n11816), .B(new_n11779), .Y(new_n11817));
  xnor_3 g11441(.A(new_n11641), .B(new_n11640), .Y(new_n11818));
  nand_4 g11442(.A(new_n11818), .B(new_n11817), .Y(new_n11819));
  not_3  g11443(.A(new_n11819), .Y(new_n11820));
  xnor_3 g11444(.A(new_n11818), .B(new_n11817), .Y(new_n11821_1));
  nand_4 g11445(.A(n10990), .B(n3992), .Y(new_n11822));
  nand_4 g11446(.A(n7236), .B(n5760), .Y(new_n11823));
  not_3  g11447(.A(new_n11823), .Y(new_n11824));
  xnor_3 g11448(.A(new_n11824), .B(new_n11822), .Y(new_n11825));
  nor_4  g11449(.A(new_n11825), .B(new_n11821_1), .Y(new_n11826));
  nor_4  g11450(.A(new_n11826), .B(new_n11820), .Y(new_n11827));
  nand_4 g11451(.A(new_n11780_1), .B(new_n11711), .Y(new_n11828));
  nand_4 g11452(.A(new_n11828), .B(new_n11782), .Y(new_n11829));
  not_3  g11453(.A(new_n11829), .Y(new_n11830));
  nor_4  g11454(.A(new_n11830), .B(new_n11827), .Y(new_n11831));
  not_3  g11455(.A(new_n11831), .Y(new_n11832));
  xnor_3 g11456(.A(new_n11829), .B(new_n11827), .Y(new_n11833));
  nor_4  g11457(.A(new_n11816), .B(new_n11579), .Y(new_n11834));
  and_4  g11458(.A(new_n11834), .B(new_n11577), .Y(new_n11835));
  not_3  g11459(.A(new_n11639), .Y(new_n11836));
  nor_4  g11460(.A(new_n11834), .B(new_n11836), .Y(new_n11837));
  nor_4  g11461(.A(new_n11837), .B(new_n11835), .Y(new_n11838));
  nand_4 g11462(.A(new_n11838), .B(new_n11833), .Y(new_n11839));
  nand_4 g11463(.A(new_n11839), .B(new_n11832), .Y(new_n11840));
  not_3  g11464(.A(new_n11812), .Y(new_n11841));
  xnor_3 g11465(.A(new_n11841), .B(new_n11811), .Y(new_n11842));
  nand_4 g11466(.A(new_n11842), .B(new_n11840), .Y(new_n11843));
  nand_4 g11467(.A(new_n11843), .B(new_n11814), .Y(new_n11844));
  nor_4  g11468(.A(new_n11844), .B(new_n11810), .Y(new_n11845));
  nor_4  g11469(.A(new_n11845), .B(new_n11809), .Y(new_n11846));
  nand_4 g11470(.A(new_n11846), .B(new_n11806), .Y(new_n11847));
  xnor_3 g11471(.A(new_n11789), .B(new_n11788), .Y(new_n11848));
  xnor_3 g11472(.A(new_n11846), .B(new_n11805), .Y(new_n11849));
  nand_4 g11473(.A(new_n11849), .B(new_n11848), .Y(new_n11850));
  nand_4 g11474(.A(new_n11850), .B(new_n11847), .Y(new_n11851));
  xnor_3 g11475(.A(new_n11851), .B(new_n11801), .Y(new_n11852));
  xnor_3 g11476(.A(new_n11852), .B(new_n11518), .Y(new_n11853));
  xnor_3 g11477(.A(new_n11501), .B(new_n11498), .Y(new_n11854));
  xnor_3 g11478(.A(new_n11854), .B(new_n11514), .Y(new_n11855));
  xnor_3 g11479(.A(new_n11513), .B(new_n11512), .Y(new_n11856));
  xnor_3 g11480(.A(new_n11510), .B(new_n11509), .Y(new_n11857));
  not_3  g11481(.A(new_n11857), .Y(new_n11858));
  xnor_3 g11482(.A(new_n11842), .B(new_n11840), .Y(new_n11859));
  nand_4 g11483(.A(new_n11859), .B(new_n11858), .Y(new_n11860));
  not_3  g11484(.A(new_n11860), .Y(new_n11861));
  xnor_3 g11485(.A(new_n11859), .B(new_n11858), .Y(new_n11862));
  xnor_3 g11486(.A(new_n11838), .B(new_n11833), .Y(new_n11863));
  nand_4 g11487(.A(n12709), .B(n6877), .Y(new_n11864));
  not_3  g11488(.A(new_n11864), .Y(new_n11865));
  nor_4  g11489(.A(new_n11865), .B(new_n11449), .Y(new_n11866));
  and_4  g11490(.A(new_n11866), .B(new_n11447), .Y(new_n11867));
  not_3  g11491(.A(new_n11503), .Y(new_n11868));
  nor_4  g11492(.A(new_n11866), .B(new_n11868), .Y(new_n11869));
  nor_4  g11493(.A(new_n11869), .B(new_n11867), .Y(new_n11870));
  not_3  g11494(.A(new_n11870), .Y(new_n11871));
  nand_4 g11495(.A(new_n11871), .B(new_n11863), .Y(new_n11872));
  not_3  g11496(.A(new_n11872), .Y(new_n11873));
  xnor_3 g11497(.A(new_n11871), .B(new_n11863), .Y(new_n11874));
  xnor_3 g11498(.A(new_n11825), .B(new_n11821_1), .Y(new_n11875));
  xor_3  g11499(.A(new_n11505), .B(new_n11504), .Y(new_n11876_1));
  nand_4 g11500(.A(new_n11876_1), .B(new_n11875), .Y(new_n11877_1));
  not_3  g11501(.A(new_n11877_1), .Y(new_n11878));
  xor_3  g11502(.A(new_n11816), .B(new_n11778), .Y(new_n11879));
  nor_4  g11503(.A(new_n11879), .B(new_n11864), .Y(new_n11880));
  not_3  g11504(.A(new_n11880), .Y(new_n11881));
  xnor_3 g11505(.A(new_n11876_1), .B(new_n11875), .Y(new_n11882));
  nor_4  g11506(.A(new_n11882), .B(new_n11881), .Y(new_n11883));
  nor_4  g11507(.A(new_n11883), .B(new_n11878), .Y(new_n11884));
  nor_4  g11508(.A(new_n11884), .B(new_n11874), .Y(new_n11885));
  nor_4  g11509(.A(new_n11885), .B(new_n11873), .Y(new_n11886));
  nor_4  g11510(.A(new_n11886), .B(new_n11862), .Y(new_n11887));
  nor_4  g11511(.A(new_n11887), .B(new_n11861), .Y(new_n11888));
  nand_4 g11512(.A(new_n11888), .B(new_n11856), .Y(new_n11889));
  not_3  g11513(.A(new_n11856), .Y(new_n11890));
  xnor_3 g11514(.A(new_n11888), .B(new_n11890), .Y(new_n11891));
  xnor_3 g11515(.A(new_n11844), .B(new_n11810), .Y(new_n11892_1));
  nand_4 g11516(.A(new_n11892_1), .B(new_n11891), .Y(new_n11893));
  nand_4 g11517(.A(new_n11893), .B(new_n11889), .Y(new_n11894));
  not_3  g11518(.A(new_n11894), .Y(new_n11895));
  nor_4  g11519(.A(new_n11895), .B(new_n11855), .Y(new_n11896));
  not_3  g11520(.A(new_n11896), .Y(new_n11897));
  not_3  g11521(.A(new_n11850), .Y(new_n11898));
  nor_4  g11522(.A(new_n11849), .B(new_n11848), .Y(new_n11899));
  nor_4  g11523(.A(new_n11899), .B(new_n11898), .Y(new_n11900));
  xnor_3 g11524(.A(new_n11894), .B(new_n11855), .Y(new_n11901));
  nand_4 g11525(.A(new_n11901), .B(new_n11900), .Y(new_n11902));
  nand_4 g11526(.A(new_n11902), .B(new_n11897), .Y(new_n11903));
  nand_4 g11527(.A(new_n11903), .B(new_n11853), .Y(new_n11904));
  xnor_3 g11528(.A(new_n11517), .B(new_n11495), .Y(new_n11905));
  xnor_3 g11529(.A(new_n11852), .B(new_n11905), .Y(new_n11906));
  not_3  g11530(.A(new_n11900), .Y(new_n11907));
  xnor_3 g11531(.A(new_n11515), .B(new_n11514), .Y(new_n11908));
  xnor_3 g11532(.A(new_n11894), .B(new_n11908), .Y(new_n11909));
  nor_4  g11533(.A(new_n11909), .B(new_n11907), .Y(new_n11910));
  nor_4  g11534(.A(new_n11910), .B(new_n11896), .Y(new_n11911));
  nand_4 g11535(.A(new_n11911), .B(new_n11906), .Y(new_n11912));
  nand_4 g11536(.A(new_n11912), .B(new_n11904), .Y(new_n11913));
  not_3  g11537(.A(new_n11913), .Y(new_n11914));
  nand_4 g11538(.A(new_n11914), .B(new_n11386), .Y(new_n11915));
  xnor_3 g11539(.A(new_n11913), .B(new_n11386), .Y(new_n11916));
  xnor_3 g11540(.A(new_n11383), .B(new_n11382), .Y(new_n11917_1));
  not_3  g11541(.A(new_n11917_1), .Y(new_n11918));
  xnor_3 g11542(.A(new_n11380), .B(new_n11379), .Y(new_n11919_1));
  not_3  g11543(.A(new_n11892_1), .Y(new_n11920));
  xnor_3 g11544(.A(new_n11920), .B(new_n11891), .Y(new_n11921));
  nand_4 g11545(.A(new_n11921), .B(new_n11919_1), .Y(new_n11922_1));
  not_3  g11546(.A(new_n11919_1), .Y(new_n11923));
  xnor_3 g11547(.A(new_n11921), .B(new_n11923), .Y(new_n11924));
  not_3  g11548(.A(new_n11378), .Y(new_n11925));
  xor_3  g11549(.A(new_n11925), .B(new_n11376), .Y(new_n11926));
  xnor_3 g11550(.A(new_n11886), .B(new_n11862), .Y(new_n11927));
  not_3  g11551(.A(new_n11927), .Y(new_n11928));
  nor_4  g11552(.A(new_n11928), .B(new_n11926), .Y(new_n11929));
  not_3  g11553(.A(new_n11929), .Y(new_n11930));
  xnor_3 g11554(.A(new_n11884), .B(new_n11874), .Y(new_n11931));
  not_3  g11555(.A(new_n11931), .Y(new_n11932));
  not_3  g11556(.A(new_n11319), .Y(new_n11933));
  nor_4  g11557(.A(new_n11321), .B(new_n11933), .Y(new_n11934));
  nor_4  g11558(.A(new_n11934), .B(new_n11371), .Y(new_n11935));
  not_3  g11559(.A(new_n11934), .Y(new_n11936));
  nor_4  g11560(.A(new_n11936), .B(new_n11318), .Y(new_n11937));
  nor_4  g11561(.A(new_n11937), .B(new_n11935), .Y(new_n11938));
  nor_4  g11562(.A(new_n11938), .B(new_n11932), .Y(new_n11939));
  not_3  g11563(.A(new_n11939), .Y(new_n11940));
  not_3  g11564(.A(new_n11938), .Y(new_n11941));
  nor_4  g11565(.A(new_n11941), .B(new_n11931), .Y(new_n11942));
  nor_4  g11566(.A(new_n11942), .B(new_n11939), .Y(new_n11943));
  xor_3  g11567(.A(new_n11815), .B(new_n11778), .Y(new_n11944));
  nor_4  g11568(.A(new_n11944), .B(new_n11865), .Y(new_n11945));
  nor_4  g11569(.A(new_n11945), .B(new_n11880), .Y(new_n11946));
  nand_4 g11570(.A(new_n11946), .B(new_n11933), .Y(new_n11947));
  not_3  g11571(.A(new_n11947), .Y(new_n11948));
  xor_3  g11572(.A(new_n11373), .B(new_n11372), .Y(new_n11949));
  nor_4  g11573(.A(new_n11949), .B(new_n11948), .Y(new_n11950));
  not_3  g11574(.A(new_n11950), .Y(new_n11951));
  not_3  g11575(.A(new_n11882), .Y(new_n11952));
  xor_3  g11576(.A(new_n11952), .B(new_n11881), .Y(new_n11953));
  xor_3  g11577(.A(new_n11949), .B(new_n11948), .Y(new_n11954));
  nand_4 g11578(.A(new_n11954), .B(new_n11953), .Y(new_n11955));
  nand_4 g11579(.A(new_n11955), .B(new_n11951), .Y(new_n11956));
  nand_4 g11580(.A(new_n11956), .B(new_n11943), .Y(new_n11957));
  nand_4 g11581(.A(new_n11957), .B(new_n11940), .Y(new_n11958));
  not_3  g11582(.A(new_n11926), .Y(new_n11959));
  nor_4  g11583(.A(new_n11927), .B(new_n11959), .Y(new_n11960));
  nor_4  g11584(.A(new_n11960), .B(new_n11929), .Y(new_n11961));
  nand_4 g11585(.A(new_n11961), .B(new_n11958), .Y(new_n11962));
  nand_4 g11586(.A(new_n11962), .B(new_n11930), .Y(new_n11963));
  nand_4 g11587(.A(new_n11963), .B(new_n11924), .Y(new_n11964));
  nand_4 g11588(.A(new_n11964), .B(new_n11922_1), .Y(new_n11965));
  nand_4 g11589(.A(new_n11965), .B(new_n11918), .Y(new_n11966));
  nor_4  g11590(.A(new_n11901), .B(new_n11900), .Y(new_n11967_1));
  nor_4  g11591(.A(new_n11967_1), .B(new_n11910), .Y(new_n11968));
  xnor_3 g11592(.A(new_n11965), .B(new_n11917_1), .Y(new_n11969));
  nand_4 g11593(.A(new_n11969), .B(new_n11968), .Y(new_n11970));
  nand_4 g11594(.A(new_n11970), .B(new_n11966), .Y(new_n11971));
  nand_4 g11595(.A(new_n11971), .B(new_n11916), .Y(new_n11972));
  nand_4 g11596(.A(new_n11972), .B(new_n11915), .Y(new_n11973));
  not_3  g11597(.A(new_n11852), .Y(new_n11974));
  nor_4  g11598(.A(new_n11974), .B(new_n11518), .Y(new_n11975));
  not_3  g11599(.A(new_n11904), .Y(new_n11976));
  nor_4  g11600(.A(new_n11976), .B(new_n11975), .Y(new_n11977));
  xnor_3 g11601(.A(new_n11977), .B(new_n11973), .Y(new_n11978));
  nand_4 g11602(.A(new_n11768), .B(new_n11735), .Y(new_n11979));
  nand_4 g11603(.A(new_n11791_1), .B(new_n11798), .Y(new_n11980));
  nand_4 g11604(.A(new_n11980), .B(new_n11979), .Y(new_n11981));
  not_3  g11605(.A(new_n11494), .Y(new_n11982));
  nand_4 g11606(.A(new_n11982), .B(new_n11464), .Y(new_n11983));
  nand_4 g11607(.A(new_n11517), .B(new_n11495), .Y(new_n11984));
  nand_4 g11608(.A(new_n11984), .B(new_n11983), .Y(new_n11985));
  xnor_3 g11609(.A(new_n11985), .B(new_n11981), .Y(new_n11986));
  nand_4 g11610(.A(new_n11363), .B(new_n11335), .Y(new_n11987));
  nand_4 g11611(.A(new_n11385), .B(new_n11364), .Y(new_n11988));
  nand_4 g11612(.A(new_n11988), .B(new_n11987), .Y(new_n11989));
  not_3  g11613(.A(new_n11354), .Y(new_n11990));
  nand_4 g11614(.A(new_n11360), .B(new_n11990), .Y(new_n11991));
  nand_4 g11615(.A(new_n11361), .B(new_n11353), .Y(new_n11992));
  nand_4 g11616(.A(new_n11992), .B(new_n11991), .Y(new_n11993));
  nand_4 g11617(.A(n6877), .B(n1198), .Y(new_n11994));
  nand_4 g11618(.A(n12753), .B(n11728), .Y(new_n11995));
  xor_3  g11619(.A(new_n11995), .B(new_n11994), .Y(new_n11996));
  nand_4 g11620(.A(n10990), .B(n4722), .Y(new_n11997));
  nand_4 g11621(.A(n1478), .B(n1471), .Y(new_n11998));
  xor_3  g11622(.A(new_n11998), .B(new_n11997), .Y(new_n11999_1));
  xor_3  g11623(.A(new_n11999_1), .B(new_n11996), .Y(new_n12000_1));
  xnor_3 g11624(.A(new_n12000_1), .B(new_n11993), .Y(new_n12001));
  nand_4 g11625(.A(n6429), .B(n4203), .Y(new_n12002));
  not_3  g11626(.A(new_n12002), .Y(new_n12003));
  nand_4 g11627(.A(new_n11480), .B(new_n11473), .Y(new_n12004));
  not_3  g11628(.A(new_n11481), .Y(new_n12005_1));
  nand_4 g11629(.A(new_n11492), .B(new_n12005_1), .Y(new_n12006));
  nand_4 g11630(.A(new_n12006), .B(new_n12004), .Y(new_n12007));
  xnor_3 g11631(.A(new_n12007), .B(new_n12003), .Y(new_n12008));
  xnor_3 g11632(.A(new_n12008), .B(new_n12001), .Y(new_n12009));
  nand_4 g11633(.A(n8819), .B(n4187), .Y(new_n12010));
  not_3  g11634(.A(new_n11476), .Y(new_n12011));
  nor_4  g11635(.A(new_n11478_1), .B(new_n12011), .Y(new_n12012));
  nor_4  g11636(.A(new_n11479), .B(new_n11475), .Y(new_n12013));
  nor_4  g11637(.A(new_n12013), .B(new_n12012), .Y(new_n12014_1));
  xor_3  g11638(.A(new_n12014_1), .B(new_n12010), .Y(new_n12015));
  xnor_3 g11639(.A(new_n12015), .B(new_n12009), .Y(new_n12016));
  nand_4 g11640(.A(new_n11468), .B(new_n11466), .Y(new_n12017));
  nand_4 g11641(.A(new_n11493), .B(new_n11470), .Y(new_n12018));
  nand_4 g11642(.A(new_n12018), .B(new_n12017), .Y(new_n12019));
  nor_4  g11643(.A(new_n11344), .B(new_n11342), .Y(new_n12020_1));
  not_3  g11644(.A(new_n11345), .Y(new_n12021));
  nor_4  g11645(.A(new_n11352), .B(new_n12021), .Y(new_n12022));
  nor_4  g11646(.A(new_n12022), .B(new_n12020_1), .Y(new_n12023));
  nand_4 g11647(.A(n9080), .B(n5212), .Y(new_n12024));
  xor_3  g11648(.A(new_n12024), .B(new_n12023), .Y(new_n12025_1));
  not_3  g11649(.A(new_n11356), .Y(new_n12026));
  nor_4  g11650(.A(new_n11358), .B(new_n12026), .Y(new_n12027));
  not_3  g11651(.A(new_n11355), .Y(new_n12028));
  nor_4  g11652(.A(new_n11359), .B(new_n12028), .Y(new_n12029));
  nor_4  g11653(.A(new_n12029), .B(new_n12027), .Y(new_n12030));
  nand_4 g11654(.A(n12709), .B(n10174), .Y(new_n12031));
  not_3  g11655(.A(new_n12031), .Y(new_n12032));
  nand_4 g11656(.A(n12000), .B(n3172), .Y(new_n12033));
  nand_4 g11657(.A(n5240), .B(n4370), .Y(new_n12034));
  xor_3  g11658(.A(new_n12034), .B(new_n12033), .Y(new_n12035));
  xnor_3 g11659(.A(new_n12035), .B(new_n12032), .Y(new_n12036));
  xnor_3 g11660(.A(new_n12036), .B(new_n12030), .Y(new_n12037));
  nand_4 g11661(.A(n9725), .B(n1333), .Y(new_n12038));
  not_3  g11662(.A(new_n12038), .Y(new_n12039));
  nand_4 g11663(.A(n11757), .B(n5320), .Y(new_n12040));
  nand_4 g11664(.A(n11877), .B(n11821), .Y(new_n12041));
  xor_3  g11665(.A(new_n12041), .B(new_n12040), .Y(new_n12042));
  xnor_3 g11666(.A(new_n12042), .B(new_n12039), .Y(new_n12043));
  not_3  g11667(.A(new_n11348), .Y(new_n12044_1));
  nor_4  g11668(.A(new_n11350), .B(new_n12044_1), .Y(new_n12045));
  nor_4  g11669(.A(new_n11351), .B(new_n11347), .Y(new_n12046));
  nor_4  g11670(.A(new_n12046), .B(new_n12045), .Y(new_n12047));
  xnor_3 g11671(.A(new_n12047), .B(new_n12043), .Y(new_n12048));
  xnor_3 g11672(.A(new_n12048), .B(new_n12037), .Y(new_n12049));
  nand_4 g11673(.A(n7646), .B(n5760), .Y(new_n12050));
  nand_4 g11674(.A(n10022), .B(n7236), .Y(new_n12051));
  not_3  g11675(.A(new_n12051), .Y(new_n12052));
  xor_3  g11676(.A(new_n12052), .B(new_n12050), .Y(new_n12053));
  xnor_3 g11677(.A(new_n12053), .B(new_n12049), .Y(new_n12054));
  xnor_3 g11678(.A(new_n12054), .B(new_n12025_1), .Y(new_n12055));
  xnor_3 g11679(.A(new_n12055), .B(new_n12019), .Y(new_n12056));
  xnor_3 g11680(.A(new_n12056), .B(new_n12016), .Y(new_n12057));
  xnor_3 g11681(.A(new_n12057), .B(new_n11989), .Y(new_n12058));
  xnor_3 g11682(.A(new_n12058), .B(new_n11986), .Y(new_n12059));
  not_3  g11683(.A(new_n11801), .Y(new_n12060));
  not_3  g11684(.A(new_n11851), .Y(new_n12061));
  nand_4 g11685(.A(new_n12061), .B(new_n12060), .Y(new_n12062));
  nand_4 g11686(.A(new_n12062), .B(new_n11793), .Y(new_n12063));
  nor_4  g11687(.A(new_n11615), .B(new_n11614), .Y(new_n12064));
  xor_3  g11688(.A(new_n11615), .B(new_n11613), .Y(new_n12065));
  nor_4  g11689(.A(new_n11621), .B(new_n12065), .Y(new_n12066));
  nor_4  g11690(.A(new_n12066), .B(new_n12064), .Y(new_n12067));
  and_4  g11691(.A(new_n11742), .B(new_n11741), .Y(new_n12068));
  nor_4  g11692(.A(new_n11745), .B(new_n12068), .Y(new_n12069_1));
  nand_4 g11693(.A(n4805), .B(n4436), .Y(new_n12070));
  not_3  g11694(.A(new_n12070), .Y(new_n12071));
  not_3  g11695(.A(new_n11603), .Y(new_n12072));
  nand_4 g11696(.A(new_n11606), .B(new_n12072), .Y(new_n12073));
  nand_4 g11697(.A(new_n12073), .B(new_n11609), .Y(new_n12074));
  xor_3  g11698(.A(new_n12074), .B(new_n12071), .Y(new_n12075));
  xor_3  g11699(.A(new_n12075), .B(new_n12069_1), .Y(new_n12076_1));
  xnor_3 g11700(.A(new_n12076_1), .B(new_n12067), .Y(new_n12077));
  nand_4 g11701(.A(new_n11750), .B(new_n11748), .Y(new_n12078));
  not_3  g11702(.A(new_n11759), .Y(new_n12079));
  nand_4 g11703(.A(new_n12079), .B(new_n11751), .Y(new_n12080));
  nand_4 g11704(.A(new_n12080), .B(new_n12078), .Y(new_n12081));
  nand_4 g11705(.A(n7159), .B(n3146), .Y(new_n12082));
  not_3  g11706(.A(new_n12082), .Y(new_n12083));
  nand_4 g11707(.A(n11967), .B(n137), .Y(new_n12084));
  nand_4 g11708(.A(n8384), .B(n6441), .Y(new_n12085));
  xor_3  g11709(.A(new_n12085), .B(new_n12084), .Y(new_n12086));
  xor_3  g11710(.A(new_n12086), .B(new_n12083), .Y(new_n12087));
  nand_4 g11711(.A(n12777), .B(n6797), .Y(new_n12088));
  nand_4 g11712(.A(n6294), .B(n6254), .Y(new_n12089));
  xor_3  g11713(.A(new_n12089), .B(new_n12088), .Y(new_n12090));
  nand_4 g11714(.A(n12947), .B(n6358), .Y(new_n12091));
  nand_4 g11715(.A(n11999), .B(n3992), .Y(new_n12092));
  not_3  g11716(.A(new_n12092), .Y(new_n12093));
  xor_3  g11717(.A(new_n12093), .B(new_n12091), .Y(new_n12094));
  xor_3  g11718(.A(new_n12094), .B(new_n12090), .Y(new_n12095));
  xnor_3 g11719(.A(new_n12095), .B(new_n12087), .Y(new_n12096));
  xnor_3 g11720(.A(new_n12096), .B(new_n12081), .Y(new_n12097));
  nand_4 g11721(.A(n11478), .B(n1353), .Y(new_n12098));
  nand_4 g11722(.A(n7862), .B(n6604), .Y(new_n12099));
  nand_4 g11723(.A(n11407), .B(n6826), .Y(new_n12100));
  xor_3  g11724(.A(new_n12100), .B(new_n12099), .Y(new_n12101));
  xor_3  g11725(.A(new_n12101), .B(new_n12098), .Y(new_n12102));
  nor_4  g11726(.A(new_n11619), .B(new_n11618), .Y(new_n12103));
  not_3  g11727(.A(new_n11617), .Y(new_n12104));
  nand_4 g11728(.A(new_n11619), .B(new_n11618), .Y(new_n12105));
  nand_4 g11729(.A(new_n12105), .B(new_n12104), .Y(new_n12106));
  not_3  g11730(.A(new_n12106), .Y(new_n12107));
  nor_4  g11731(.A(new_n12107), .B(new_n12103), .Y(new_n12108));
  xnor_3 g11732(.A(new_n12108), .B(new_n12102), .Y(new_n12109));
  xnor_3 g11733(.A(new_n12109), .B(new_n12097), .Y(new_n12110));
  xnor_3 g11734(.A(new_n12110), .B(new_n12077), .Y(new_n12111_1));
  not_3  g11735(.A(new_n11602), .Y(new_n12112));
  nand_4 g11736(.A(new_n11611), .B(new_n12112), .Y(new_n12113));
  xnor_3 g11737(.A(new_n11621), .B(new_n12065), .Y(new_n12114));
  nand_4 g11738(.A(new_n12114), .B(new_n11612), .Y(new_n12115));
  nand_4 g11739(.A(new_n12115), .B(new_n12113), .Y(new_n12116));
  not_3  g11740(.A(new_n11746), .Y(new_n12117));
  nor_4  g11741(.A(new_n12117), .B(new_n11738), .Y(new_n12118));
  not_3  g11742(.A(new_n11747), .Y(new_n12119));
  nor_4  g11743(.A(new_n11760), .B(new_n12119), .Y(new_n12120));
  nor_4  g11744(.A(new_n12120), .B(new_n12118), .Y(new_n12121));
  xor_3  g11745(.A(new_n12121), .B(new_n12116), .Y(new_n12122));
  xnor_3 g11746(.A(new_n12122), .B(new_n12111_1), .Y(new_n12123));
  nand_4 g11747(.A(new_n11630), .B(new_n11600), .Y(new_n12124));
  nand_4 g11748(.A(new_n11653), .B(new_n11795), .Y(new_n12125));
  nand_4 g11749(.A(new_n12125), .B(new_n12124), .Y(new_n12126));
  nor_4  g11750(.A(new_n11700), .B(new_n11765), .Y(new_n12127));
  not_3  g11751(.A(new_n11767), .Y(new_n12128));
  nor_4  g11752(.A(new_n12128), .B(new_n11761), .Y(new_n12129));
  nor_4  g11753(.A(new_n12129), .B(new_n12127), .Y(new_n12130));
  xnor_3 g11754(.A(new_n12130), .B(new_n12126), .Y(new_n12131));
  nor_4  g11755(.A(new_n11564), .B(new_n11627), .Y(new_n12132));
  not_3  g11756(.A(new_n11629), .Y(new_n12133));
  nor_4  g11757(.A(new_n12133), .B(new_n11623), .Y(new_n12134));
  nor_4  g11758(.A(new_n12134), .B(new_n12132), .Y(new_n12135));
  nand_4 g11759(.A(new_n11303), .B(new_n11339), .Y(new_n12136));
  nand_4 g11760(.A(new_n11362), .B(new_n11341), .Y(new_n12137));
  nand_4 g11761(.A(new_n12137), .B(new_n12136), .Y(new_n12138));
  and_4  g11762(.A(new_n11755_1), .B(new_n11754), .Y(new_n12139));
  nor_4  g11763(.A(new_n11758), .B(new_n12139), .Y(new_n12140));
  nand_4 g11764(.A(n5283), .B(n447), .Y(new_n12141));
  nand_4 g11765(.A(n12489), .B(n4938), .Y(new_n12142));
  nand_4 g11766(.A(n11791), .B(n5198), .Y(new_n12143));
  xor_3  g11767(.A(new_n12143), .B(new_n12142), .Y(new_n12144));
  xor_3  g11768(.A(new_n12144), .B(new_n12141), .Y(new_n12145_1));
  xnor_3 g11769(.A(new_n12145_1), .B(new_n12140), .Y(new_n12146));
  xnor_3 g11770(.A(new_n12146), .B(new_n12138), .Y(new_n12147));
  nand_4 g11771(.A(n8717), .B(n2464), .Y(new_n12148));
  not_3  g11772(.A(new_n12148), .Y(new_n12149));
  nor_4  g11773(.A(new_n11484), .B(new_n11483), .Y(new_n12150));
  not_3  g11774(.A(new_n11485), .Y(new_n12151));
  nor_4  g11775(.A(new_n11491), .B(new_n12151), .Y(new_n12152));
  nor_4  g11776(.A(new_n12152), .B(new_n12150), .Y(new_n12153));
  not_3  g11777(.A(new_n11487), .Y(new_n12154));
  nor_4  g11778(.A(new_n11489), .B(new_n12154), .Y(new_n12155));
  not_3  g11779(.A(new_n11486), .Y(new_n12156));
  nor_4  g11780(.A(new_n11490), .B(new_n12156), .Y(new_n12157));
  nor_4  g11781(.A(new_n12157), .B(new_n12155), .Y(new_n12158));
  nand_4 g11782(.A(n11311), .B(n2433), .Y(new_n12159));
  nand_4 g11783(.A(n9400), .B(n7730), .Y(new_n12160));
  not_3  g11784(.A(new_n12160), .Y(new_n12161));
  xor_3  g11785(.A(new_n12161), .B(new_n12159), .Y(new_n12162));
  xnor_3 g11786(.A(new_n12162), .B(new_n12158), .Y(new_n12163));
  xnor_3 g11787(.A(new_n12163), .B(new_n12153), .Y(new_n12164));
  xnor_3 g11788(.A(new_n12164), .B(new_n12149), .Y(new_n12165));
  xnor_3 g11789(.A(new_n12165), .B(new_n12147), .Y(new_n12166));
  xnor_3 g11790(.A(new_n12166), .B(new_n12135), .Y(new_n12167));
  xnor_3 g11791(.A(new_n12167), .B(new_n12131), .Y(new_n12168));
  xnor_3 g11792(.A(new_n12168), .B(new_n12123), .Y(new_n12169));
  xnor_3 g11793(.A(new_n12169), .B(new_n12063), .Y(new_n12170));
  xnor_3 g11794(.A(new_n12170), .B(new_n12059), .Y(new_n12171));
  xnor_3 g11795(.A(new_n12171), .B(new_n11978), .Y(n4378));
  xor_3  g11796(.A(new_n4109), .B(new_n4021), .Y(n4397));
  xor_3  g11797(.A(new_n4453), .B(new_n4442), .Y(n4553));
  xor_3  g11798(.A(new_n1043), .B(new_n1033), .Y(n4686));
  xnor_3 g11799(.A(new_n10023), .B(new_n10005), .Y(n4689));
  not_3  g11800(.A(new_n5277), .Y(new_n12177));
  nand_4 g11801(.A(new_n5232), .B(new_n5231), .Y(new_n12178));
  xnor_3 g11802(.A(new_n12178), .B(new_n12177), .Y(n4733));
  xnor_3 g11803(.A(new_n2184), .B(new_n2176), .Y(n4757));
  not_3  g11804(.A(new_n5273), .Y(new_n12181));
  xor_3  g11805(.A(new_n12181), .B(new_n5271), .Y(n4971));
  xnor_3 g11806(.A(new_n7035), .B(new_n7034), .Y(n5030));
  not_3  g11807(.A(new_n3089), .Y(new_n12184));
  xor_3  g11808(.A(new_n12184), .B(new_n3056), .Y(n5034));
  not_3  g11809(.A(new_n3073), .Y(new_n12186));
  xor_3  g11810(.A(new_n3082), .B(new_n12186), .Y(n5094));
  nand_4 g11811(.A(new_n11124), .B(new_n11115), .Y(new_n12188));
  nand_4 g11812(.A(n5320), .B(n2564), .Y(new_n12189));
  nand_4 g11813(.A(n4370), .B(n4189), .Y(new_n12190));
  xor_3  g11814(.A(new_n12190), .B(new_n12189), .Y(new_n12191));
  xnor_3 g11815(.A(new_n12191), .B(new_n12188), .Y(new_n12192));
  nand_4 g11816(.A(n11877), .B(n6770), .Y(new_n12193));
  not_3  g11817(.A(new_n12193), .Y(new_n12194));
  and_4  g11818(.A(new_n11121), .B(new_n11120), .Y(new_n12195));
  not_3  g11819(.A(new_n11119), .Y(new_n12196));
  nor_4  g11820(.A(new_n11122), .B(new_n12196), .Y(new_n12197));
  nor_4  g11821(.A(new_n12197), .B(new_n12195), .Y(new_n12198));
  nand_4 g11822(.A(new_n12198), .B(new_n12194), .Y(new_n12199));
  not_3  g11823(.A(new_n12199), .Y(new_n12200));
  nor_4  g11824(.A(new_n12198), .B(new_n12194), .Y(new_n12201));
  nor_4  g11825(.A(new_n12201), .B(new_n12200), .Y(new_n12202));
  nand_4 g11826(.A(n9920), .B(n5212), .Y(new_n12203));
  nand_4 g11827(.A(n11407), .B(n3627), .Y(new_n12204));
  xor_3  g11828(.A(new_n12204), .B(new_n12203), .Y(new_n12205));
  xnor_3 g11829(.A(new_n12205), .B(new_n12202), .Y(new_n12206));
  xnor_3 g11830(.A(new_n12206), .B(new_n12192), .Y(new_n12207));
  not_3  g11831(.A(new_n12207), .Y(new_n12208));
  nor_4  g11832(.A(new_n11108), .B(new_n11103), .Y(new_n12209));
  not_3  g11833(.A(new_n12209), .Y(new_n12210));
  not_3  g11834(.A(new_n11103), .Y(new_n12211));
  xnor_3 g11835(.A(new_n11108), .B(new_n12211), .Y(new_n12212));
  nand_4 g11836(.A(new_n11127), .B(new_n12212), .Y(new_n12213));
  nand_4 g11837(.A(new_n12213), .B(new_n12210), .Y(new_n12214));
  nand_4 g11838(.A(new_n12214), .B(new_n12208), .Y(new_n12215));
  nand_4 g11839(.A(new_n12205), .B(new_n12202), .Y(new_n12216));
  nand_4 g11840(.A(new_n12216), .B(new_n12199), .Y(new_n12217));
  nand_4 g11841(.A(n12000), .B(n2564), .Y(new_n12218));
  not_3  g11842(.A(new_n12218), .Y(new_n12219));
  nand_4 g11843(.A(n5320), .B(n4189), .Y(new_n12220));
  nand_4 g11844(.A(n9725), .B(n6687), .Y(new_n12221_1));
  xor_3  g11845(.A(new_n12221_1), .B(new_n12220), .Y(new_n12222));
  xnor_3 g11846(.A(new_n12222), .B(new_n12219), .Y(new_n12223));
  xnor_3 g11847(.A(new_n12223), .B(new_n12217), .Y(new_n12224));
  nor_4  g11848(.A(new_n12204), .B(new_n12203), .Y(new_n12225));
  nand_4 g11849(.A(n6770), .B(n4370), .Y(new_n12226));
  not_3  g11850(.A(new_n12226), .Y(new_n12227));
  xor_3  g11851(.A(new_n12227), .B(new_n12225), .Y(new_n12228));
  nand_4 g11852(.A(n5212), .B(n3627), .Y(new_n12229));
  nand_4 g11853(.A(n11877), .B(n9920), .Y(new_n12230));
  nand_4 g11854(.A(n11407), .B(n4516), .Y(new_n12231));
  nand_4 g11855(.A(new_n12231), .B(new_n12230), .Y(new_n12232));
  not_3  g11856(.A(new_n12230), .Y(new_n12233));
  not_3  g11857(.A(new_n12231), .Y(new_n12234));
  nand_4 g11858(.A(new_n12234), .B(new_n12233), .Y(new_n12235));
  nand_4 g11859(.A(new_n12235), .B(new_n12232), .Y(new_n12236));
  xor_3  g11860(.A(new_n12236), .B(new_n12229), .Y(new_n12237));
  xnor_3 g11861(.A(new_n12237), .B(new_n12228), .Y(new_n12238));
  not_3  g11862(.A(new_n12238), .Y(new_n12239));
  xnor_3 g11863(.A(new_n12239), .B(new_n12224), .Y(new_n12240));
  not_3  g11864(.A(new_n12240), .Y(new_n12241));
  not_3  g11865(.A(new_n12188), .Y(new_n12242));
  not_3  g11866(.A(new_n12191), .Y(new_n12243));
  nor_4  g11867(.A(new_n12243), .B(new_n12242), .Y(new_n12244));
  not_3  g11868(.A(new_n12244), .Y(new_n12245));
  nor_4  g11869(.A(new_n12190), .B(new_n12189), .Y(new_n12246));
  nor_4  g11870(.A(new_n12206), .B(new_n12192), .Y(new_n12247_1));
  xnor_3 g11871(.A(new_n12247_1), .B(new_n12246), .Y(new_n12248));
  nand_4 g11872(.A(new_n12248), .B(new_n12245), .Y(new_n12249));
  nor_4  g11873(.A(new_n12249), .B(new_n12241), .Y(new_n12250));
  nand_4 g11874(.A(new_n12249), .B(new_n12241), .Y(new_n12251));
  not_3  g11875(.A(new_n12251), .Y(new_n12252));
  nor_4  g11876(.A(new_n12252), .B(new_n12250), .Y(new_n12253));
  xnor_3 g11877(.A(new_n12253), .B(new_n12215), .Y(new_n12254));
  nand_4 g11878(.A(n12000), .B(n6687), .Y(new_n12255));
  not_3  g11879(.A(new_n12255), .Y(new_n12256));
  xnor_3 g11880(.A(new_n12214), .B(new_n12208), .Y(new_n12257));
  not_3  g11881(.A(new_n12257), .Y(new_n12258));
  nand_4 g11882(.A(new_n12258), .B(new_n12256), .Y(new_n12259));
  nor_4  g11883(.A(new_n11129), .B(new_n11102), .Y(new_n12260));
  xnor_3 g11884(.A(new_n12257), .B(new_n12256), .Y(new_n12261));
  nand_4 g11885(.A(new_n12261), .B(new_n12260), .Y(new_n12262));
  nand_4 g11886(.A(new_n12262), .B(new_n12259), .Y(new_n12263));
  xnor_3 g11887(.A(new_n12263), .B(new_n12254), .Y(new_n12264));
  not_3  g11888(.A(new_n12264), .Y(new_n12265));
  nand_4 g11889(.A(n8717), .B(n8336), .Y(new_n12266));
  nand_4 g11890(.A(n6429), .B(n2226), .Y(new_n12267));
  nand_4 g11891(.A(n11728), .B(n1094), .Y(new_n12268));
  nand_4 g11892(.A(n12709), .B(n10678), .Y(new_n12269));
  xnor_3 g11893(.A(new_n12269), .B(new_n12268), .Y(new_n12270));
  nor_4  g11894(.A(new_n12270), .B(new_n12267), .Y(new_n12271));
  not_3  g11895(.A(new_n12267), .Y(new_n12272));
  not_3  g11896(.A(new_n12270), .Y(new_n12273));
  nor_4  g11897(.A(new_n12273), .B(new_n12272), .Y(new_n12274));
  nor_4  g11898(.A(new_n12274), .B(new_n12271), .Y(new_n12275));
  nor_4  g11899(.A(new_n11151), .B(new_n11145), .Y(new_n12276));
  nor_4  g11900(.A(new_n12276), .B(new_n11150), .Y(new_n12277));
  xnor_3 g11901(.A(new_n12277), .B(new_n12275), .Y(new_n12278));
  nand_4 g11902(.A(n10928), .B(n2433), .Y(new_n12279));
  nand_4 g11903(.A(n8819), .B(n6986), .Y(new_n12280));
  xor_3  g11904(.A(new_n12280), .B(new_n12279), .Y(new_n12281));
  xnor_3 g11905(.A(new_n12281), .B(new_n12278), .Y(new_n12282));
  nand_4 g11906(.A(new_n11142), .B(new_n11136), .Y(new_n12283));
  not_3  g11907(.A(new_n12283), .Y(new_n12284));
  nor_4  g11908(.A(new_n11153_1), .B(new_n11143), .Y(new_n12285));
  nor_4  g11909(.A(new_n12285), .B(new_n12284), .Y(new_n12286));
  not_3  g11910(.A(new_n12286), .Y(new_n12287));
  nand_4 g11911(.A(new_n12287), .B(new_n12282), .Y(new_n12288));
  not_3  g11912(.A(new_n12288), .Y(new_n12289));
  nor_4  g11913(.A(new_n12287), .B(new_n12282), .Y(new_n12290));
  nor_4  g11914(.A(new_n12290), .B(new_n12289), .Y(new_n12291));
  not_3  g11915(.A(new_n11155), .Y(new_n12292));
  nand_4 g11916(.A(new_n11163), .B(new_n11159), .Y(new_n12293));
  nand_4 g11917(.A(new_n12293), .B(new_n12292), .Y(new_n12294));
  xnor_3 g11918(.A(new_n12294), .B(new_n12291), .Y(new_n12295));
  nor_4  g11919(.A(new_n12295), .B(new_n12266), .Y(new_n12296));
  not_3  g11920(.A(new_n12296), .Y(new_n12297));
  not_3  g11921(.A(new_n11133), .Y(new_n12298));
  nor_4  g11922(.A(new_n11164), .B(new_n12298), .Y(new_n12299_1));
  not_3  g11923(.A(new_n12266), .Y(new_n12300));
  xnor_3 g11924(.A(new_n12295), .B(new_n12300), .Y(new_n12301));
  nand_4 g11925(.A(new_n12301), .B(new_n12299_1), .Y(new_n12302));
  nand_4 g11926(.A(new_n12302), .B(new_n12297), .Y(new_n12303));
  nand_4 g11927(.A(new_n12294), .B(new_n12291), .Y(new_n12304));
  not_3  g11928(.A(new_n12271), .Y(new_n12305));
  nand_4 g11929(.A(new_n12277), .B(new_n12275), .Y(new_n12306));
  and_4  g11930(.A(new_n12306), .B(new_n12305), .Y(new_n12307));
  nand_4 g11931(.A(n10928), .B(n8717), .Y(new_n12308));
  not_3  g11932(.A(new_n12308), .Y(new_n12309));
  nand_4 g11933(.A(n6986), .B(n2433), .Y(new_n12310));
  nand_4 g11934(.A(n8336), .B(n7730), .Y(new_n12311));
  not_3  g11935(.A(new_n12311), .Y(new_n12312));
  xor_3  g11936(.A(new_n12312), .B(new_n12310), .Y(new_n12313));
  xnor_3 g11937(.A(new_n12313), .B(new_n12309), .Y(new_n12314));
  xnor_3 g11938(.A(new_n12314), .B(new_n12307), .Y(new_n12315));
  nor_4  g11939(.A(new_n12269), .B(new_n12268), .Y(new_n12316));
  not_3  g11940(.A(new_n12316), .Y(new_n12317));
  nand_4 g11941(.A(n8819), .B(n2226), .Y(new_n12318));
  xor_3  g11942(.A(new_n12318), .B(new_n12317), .Y(new_n12319));
  nand_4 g11943(.A(n11728), .B(n10678), .Y(new_n12320));
  nand_4 g11944(.A(n6429), .B(n1094), .Y(new_n12321));
  nand_4 g11945(.A(n12709), .B(n7320), .Y(new_n12322));
  not_3  g11946(.A(new_n12322), .Y(new_n12323));
  xor_3  g11947(.A(new_n12323), .B(new_n12321), .Y(new_n12324));
  xnor_3 g11948(.A(new_n12324), .B(new_n12320), .Y(new_n12325));
  xnor_3 g11949(.A(new_n12325), .B(new_n12319), .Y(new_n12326));
  xnor_3 g11950(.A(new_n12326), .B(new_n12315), .Y(new_n12327));
  not_3  g11951(.A(new_n12278), .Y(new_n12328));
  nand_4 g11952(.A(new_n12281), .B(new_n12328), .Y(new_n12329));
  nor_4  g11953(.A(new_n12280), .B(new_n12279), .Y(new_n12330));
  xnor_3 g11954(.A(new_n12289), .B(new_n12330), .Y(new_n12331));
  nand_4 g11955(.A(new_n12331), .B(new_n12329), .Y(new_n12332));
  xnor_3 g11956(.A(new_n12332), .B(new_n12327), .Y(new_n12333));
  xnor_3 g11957(.A(new_n12333), .B(new_n12304), .Y(new_n12334));
  xnor_3 g11958(.A(new_n12334), .B(new_n12303), .Y(new_n12335));
  xnor_3 g11959(.A(new_n12301), .B(new_n12299_1), .Y(new_n12336));
  not_3  g11960(.A(new_n11169), .Y(new_n12337));
  not_3  g11961(.A(new_n11173), .Y(new_n12338));
  nor_4  g11962(.A(new_n11246), .B(new_n12338), .Y(new_n12339));
  nor_4  g11963(.A(new_n12339), .B(new_n12337), .Y(new_n12340));
  nor_4  g11964(.A(new_n12340), .B(new_n12336), .Y(new_n12341));
  not_3  g11965(.A(new_n12341), .Y(new_n12342));
  nand_4 g11966(.A(new_n12340), .B(new_n12336), .Y(new_n12343));
  nor_4  g11967(.A(new_n11234), .B(new_n11241), .Y(new_n12344));
  not_3  g11968(.A(new_n12344), .Y(new_n12345));
  nand_4 g11969(.A(n11222), .B(n6441), .Y(new_n12346));
  not_3  g11970(.A(new_n11210), .Y(new_n12347));
  nand_4 g11971(.A(new_n11216_1), .B(new_n12347), .Y(new_n12348));
  nand_4 g11972(.A(new_n11228), .B(new_n11217), .Y(new_n12349));
  nand_4 g11973(.A(new_n12349), .B(new_n12348), .Y(new_n12350));
  nand_4 g11974(.A(n12947), .B(n11153), .Y(new_n12351));
  nand_4 g11975(.A(n11791), .B(n5314), .Y(new_n12352));
  xor_3  g11976(.A(new_n12352), .B(new_n12351), .Y(new_n12353));
  xnor_3 g11977(.A(new_n12353), .B(new_n12350), .Y(new_n12354));
  nand_4 g11978(.A(n1478), .B(n996), .Y(new_n12355));
  nand_4 g11979(.A(n10990), .B(n5319), .Y(new_n12356));
  nand_4 g11980(.A(n5767), .B(n5760), .Y(new_n12357));
  xnor_3 g11981(.A(new_n12357), .B(new_n12356), .Y(new_n12358));
  nor_4  g11982(.A(new_n12358), .B(new_n12355), .Y(new_n12359));
  not_3  g11983(.A(new_n12355), .Y(new_n12360));
  not_3  g11984(.A(new_n12358), .Y(new_n12361));
  nor_4  g11985(.A(new_n12361), .B(new_n12360), .Y(new_n12362));
  nor_4  g11986(.A(new_n12362), .B(new_n12359), .Y(new_n12363));
  nand_4 g11987(.A(new_n11225), .B(new_n11218), .Y(new_n12364));
  nand_4 g11988(.A(new_n12364), .B(new_n11221), .Y(new_n12365));
  xor_3  g11989(.A(new_n12365), .B(new_n12363), .Y(new_n12366));
  xnor_3 g11990(.A(new_n12366), .B(new_n12354), .Y(new_n12367));
  nor_4  g11991(.A(new_n11229), .B(new_n11209), .Y(new_n12368));
  nor_4  g11992(.A(new_n11233), .B(new_n11230), .Y(new_n12369));
  nor_4  g11993(.A(new_n12369), .B(new_n12368), .Y(new_n12370));
  nor_4  g11994(.A(new_n12370), .B(new_n12367), .Y(new_n12371));
  not_3  g11995(.A(new_n12367), .Y(new_n12372));
  not_3  g11996(.A(new_n12370), .Y(new_n12373));
  nor_4  g11997(.A(new_n12373), .B(new_n12372), .Y(new_n12374));
  nor_4  g11998(.A(new_n12374), .B(new_n12371), .Y(new_n12375));
  xnor_3 g11999(.A(new_n12375), .B(new_n12346), .Y(new_n12376));
  xnor_3 g12000(.A(new_n12376), .B(new_n12345), .Y(new_n12377));
  not_3  g12001(.A(new_n11206), .Y(new_n12378));
  nand_4 g12002(.A(n12069), .B(n447), .Y(new_n12379));
  nand_4 g12003(.A(n12777), .B(n7160), .Y(new_n12380));
  nand_4 g12004(.A(n7159), .B(n4828), .Y(new_n12381));
  nand_4 g12005(.A(n12489), .B(n2515), .Y(new_n12382));
  xnor_3 g12006(.A(new_n12382), .B(new_n12381), .Y(new_n12383));
  nor_4  g12007(.A(new_n12383), .B(new_n12380), .Y(new_n12384));
  not_3  g12008(.A(new_n12380), .Y(new_n12385));
  not_3  g12009(.A(new_n12383), .Y(new_n12386));
  nor_4  g12010(.A(new_n12386), .B(new_n12385), .Y(new_n12387));
  nor_4  g12011(.A(new_n12387), .B(new_n12384), .Y(new_n12388));
  nor_4  g12012(.A(new_n11189), .B(new_n11183), .Y(new_n12389));
  nor_4  g12013(.A(new_n12389), .B(new_n11188), .Y(new_n12390));
  xnor_3 g12014(.A(new_n12390), .B(new_n12388), .Y(new_n12391_1));
  nand_4 g12015(.A(n12391), .B(n11967), .Y(new_n12392));
  nand_4 g12016(.A(n7891), .B(n6254), .Y(new_n12393));
  not_3  g12017(.A(new_n12393), .Y(new_n12394));
  xor_3  g12018(.A(new_n12394), .B(new_n12392), .Y(new_n12395));
  xnor_3 g12019(.A(new_n12395), .B(new_n12391_1), .Y(new_n12396));
  and_4  g12020(.A(new_n11180), .B(new_n11177), .Y(new_n12397));
  nor_4  g12021(.A(new_n11191), .B(new_n11181), .Y(new_n12398));
  nor_4  g12022(.A(new_n12398), .B(new_n12397), .Y(new_n12399));
  not_3  g12023(.A(new_n12399), .Y(new_n12400));
  xnor_3 g12024(.A(new_n12400), .B(new_n12396), .Y(new_n12401));
  not_3  g12025(.A(new_n11193), .Y(new_n12402));
  nand_4 g12026(.A(new_n11201), .B(new_n11197), .Y(new_n12403));
  nand_4 g12027(.A(new_n12403), .B(new_n12402), .Y(new_n12404));
  xnor_3 g12028(.A(new_n12404), .B(new_n12401), .Y(new_n12405));
  xnor_3 g12029(.A(new_n12405), .B(new_n12379), .Y(new_n12406));
  not_3  g12030(.A(new_n12406), .Y(new_n12407));
  nor_4  g12031(.A(new_n12407), .B(new_n12378), .Y(new_n12408));
  nor_4  g12032(.A(new_n12406), .B(new_n11206), .Y(new_n12409));
  nor_4  g12033(.A(new_n12409), .B(new_n12408), .Y(new_n12410));
  not_3  g12034(.A(new_n12410), .Y(new_n12411));
  nand_4 g12035(.A(new_n11244), .B(new_n11207), .Y(new_n12412));
  nand_4 g12036(.A(new_n12412), .B(new_n11240), .Y(new_n12413));
  xnor_3 g12037(.A(new_n12413), .B(new_n12411), .Y(new_n12414));
  xnor_3 g12038(.A(new_n12414), .B(new_n12377), .Y(new_n12415));
  nand_4 g12039(.A(new_n12415), .B(new_n12343), .Y(new_n12416));
  nand_4 g12040(.A(new_n12416), .B(new_n12342), .Y(new_n12417));
  xnor_3 g12041(.A(new_n12417), .B(new_n12335), .Y(new_n12418));
  not_3  g12042(.A(new_n12363), .Y(new_n12419));
  nor_4  g12043(.A(new_n12365), .B(new_n12419), .Y(new_n12420));
  nor_4  g12044(.A(new_n12420), .B(new_n12359), .Y(new_n12421));
  not_3  g12045(.A(new_n12421), .Y(new_n12422));
  nand_4 g12046(.A(n11153), .B(n6441), .Y(new_n12423));
  nand_4 g12047(.A(n12947), .B(n5314), .Y(new_n12424));
  nand_4 g12048(.A(n11999), .B(n11222), .Y(new_n12425));
  not_3  g12049(.A(new_n12425), .Y(new_n12426));
  xor_3  g12050(.A(new_n12426), .B(new_n12424), .Y(new_n12427));
  xnor_3 g12051(.A(new_n12427), .B(new_n12423), .Y(new_n12428));
  xnor_3 g12052(.A(new_n12428), .B(new_n12422), .Y(new_n12429));
  nor_4  g12053(.A(new_n12357), .B(new_n12356), .Y(new_n12430));
  nand_4 g12054(.A(n11791), .B(n996), .Y(new_n12431));
  xor_3  g12055(.A(new_n12431), .B(new_n12430), .Y(new_n12432));
  nand_4 g12056(.A(n5760), .B(n5319), .Y(new_n12433));
  nand_4 g12057(.A(n5767), .B(n1478), .Y(new_n12434));
  nand_4 g12058(.A(n10990), .B(n9457), .Y(new_n12435));
  not_3  g12059(.A(new_n12435), .Y(new_n12436));
  xor_3  g12060(.A(new_n12436), .B(new_n12434), .Y(new_n12437));
  xnor_3 g12061(.A(new_n12437), .B(new_n12433), .Y(new_n12438));
  xnor_3 g12062(.A(new_n12438), .B(new_n12432), .Y(new_n12439));
  not_3  g12063(.A(new_n12439), .Y(new_n12440));
  xnor_3 g12064(.A(new_n12440), .B(new_n12429), .Y(new_n12441));
  nand_4 g12065(.A(new_n12353), .B(new_n12350), .Y(new_n12442));
  nor_4  g12066(.A(new_n12352), .B(new_n12351), .Y(new_n12443));
  nor_4  g12067(.A(new_n12366), .B(new_n12354), .Y(new_n12444_1));
  xnor_3 g12068(.A(new_n12444_1), .B(new_n12443), .Y(new_n12445));
  nand_4 g12069(.A(new_n12445), .B(new_n12442), .Y(new_n12446));
  xnor_3 g12070(.A(new_n12446), .B(new_n12441), .Y(new_n12447));
  xnor_3 g12071(.A(new_n12447), .B(new_n12371), .Y(new_n12448));
  not_3  g12072(.A(new_n12346), .Y(new_n12449));
  nand_4 g12073(.A(new_n12375), .B(new_n12449), .Y(new_n12450));
  nand_4 g12074(.A(new_n12376), .B(new_n12344), .Y(new_n12451));
  nand_4 g12075(.A(new_n12451), .B(new_n12450), .Y(new_n12452));
  xnor_3 g12076(.A(new_n12452), .B(new_n12448), .Y(new_n12453));
  not_3  g12077(.A(new_n12401), .Y(new_n12454));
  not_3  g12078(.A(new_n12404), .Y(new_n12455));
  nor_4  g12079(.A(new_n12455), .B(new_n12454), .Y(new_n12456));
  not_3  g12080(.A(new_n12456), .Y(new_n12457));
  nand_4 g12081(.A(new_n12390), .B(new_n12388), .Y(new_n12458));
  not_3  g12082(.A(new_n12458), .Y(new_n12459));
  nor_4  g12083(.A(new_n12459), .B(new_n12384), .Y(new_n12460));
  not_3  g12084(.A(new_n12460), .Y(new_n12461));
  nand_4 g12085(.A(n12391), .B(n447), .Y(new_n12462));
  not_3  g12086(.A(new_n12462), .Y(new_n12463));
  nand_4 g12087(.A(n11967), .B(n7891), .Y(new_n12464));
  nand_4 g12088(.A(n12069), .B(n1353), .Y(new_n12465));
  nand_4 g12089(.A(new_n12465), .B(new_n12464), .Y(new_n12466));
  not_3  g12090(.A(new_n12464), .Y(new_n12467));
  not_3  g12091(.A(new_n12465), .Y(new_n12468));
  nand_4 g12092(.A(new_n12468), .B(new_n12467), .Y(new_n12469));
  nand_4 g12093(.A(new_n12469), .B(new_n12466), .Y(new_n12470));
  xor_3  g12094(.A(new_n12470), .B(new_n12463), .Y(new_n12471));
  xnor_3 g12095(.A(new_n12471), .B(new_n12461), .Y(new_n12472));
  nor_4  g12096(.A(new_n12382), .B(new_n12381), .Y(new_n12473));
  nand_4 g12097(.A(n7160), .B(n6254), .Y(new_n12474));
  xor_3  g12098(.A(new_n12474), .B(new_n12473), .Y(new_n12475));
  nand_4 g12099(.A(n7159), .B(n2515), .Y(new_n12476));
  not_3  g12100(.A(new_n12476), .Y(new_n12477));
  nand_4 g12101(.A(n12777), .B(n4828), .Y(new_n12478));
  nand_4 g12102(.A(n12489), .B(n1199), .Y(new_n12479));
  nand_4 g12103(.A(new_n12479), .B(new_n12478), .Y(new_n12480));
  not_3  g12104(.A(new_n12478), .Y(new_n12481));
  not_3  g12105(.A(new_n12479), .Y(new_n12482));
  nand_4 g12106(.A(new_n12482), .B(new_n12481), .Y(new_n12483));
  nand_4 g12107(.A(new_n12483), .B(new_n12480), .Y(new_n12484));
  xor_3  g12108(.A(new_n12484), .B(new_n12477), .Y(new_n12485));
  xnor_3 g12109(.A(new_n12485), .B(new_n12475), .Y(new_n12486));
  not_3  g12110(.A(new_n12486), .Y(new_n12487));
  xnor_3 g12111(.A(new_n12487), .B(new_n12472), .Y(new_n12488));
  nor_4  g12112(.A(new_n12395), .B(new_n12391_1), .Y(new_n12489_1));
  not_3  g12113(.A(new_n12489_1), .Y(new_n12490));
  nor_4  g12114(.A(new_n12393), .B(new_n12392), .Y(new_n12491));
  nor_4  g12115(.A(new_n12399), .B(new_n12396), .Y(new_n12492));
  xnor_3 g12116(.A(new_n12492), .B(new_n12491), .Y(new_n12493));
  nand_4 g12117(.A(new_n12493), .B(new_n12490), .Y(new_n12494));
  xnor_3 g12118(.A(new_n12494), .B(new_n12488), .Y(new_n12495));
  xnor_3 g12119(.A(new_n12495), .B(new_n12457), .Y(new_n12496));
  not_3  g12120(.A(new_n12379), .Y(new_n12497));
  not_3  g12121(.A(new_n12405), .Y(new_n12498));
  nor_4  g12122(.A(new_n12498), .B(new_n12497), .Y(new_n12499));
  nor_4  g12123(.A(new_n12409), .B(new_n12499), .Y(new_n12500));
  xnor_3 g12124(.A(new_n12500), .B(new_n12496), .Y(new_n12501));
  xnor_3 g12125(.A(new_n12501), .B(new_n12453), .Y(new_n12502));
  nand_4 g12126(.A(new_n12413), .B(new_n12411), .Y(new_n12503));
  xnor_3 g12127(.A(new_n12413), .B(new_n12410), .Y(new_n12504));
  nand_4 g12128(.A(new_n12504), .B(new_n12377), .Y(new_n12505));
  nand_4 g12129(.A(new_n12505), .B(new_n12503), .Y(new_n12506));
  xnor_3 g12130(.A(new_n12506), .B(new_n12502), .Y(new_n12507));
  not_3  g12131(.A(new_n12507), .Y(new_n12508));
  xnor_3 g12132(.A(new_n12508), .B(new_n12418), .Y(new_n12509));
  not_3  g12133(.A(new_n12509), .Y(new_n12510));
  nand_4 g12134(.A(new_n12510), .B(new_n12265), .Y(new_n12511_1));
  nand_4 g12135(.A(new_n12509), .B(new_n12264), .Y(new_n12512));
  nand_4 g12136(.A(new_n12512), .B(new_n12511_1), .Y(new_n12513));
  not_3  g12137(.A(new_n12262), .Y(new_n12514));
  nor_4  g12138(.A(new_n12261), .B(new_n12260), .Y(new_n12515));
  nor_4  g12139(.A(new_n12515), .B(new_n12514), .Y(new_n12516));
  nor_4  g12140(.A(new_n11254), .B(new_n11248), .Y(new_n12517));
  nor_4  g12141(.A(new_n12517), .B(new_n11250), .Y(new_n12518));
  nor_4  g12142(.A(new_n12518), .B(new_n12516), .Y(new_n12519));
  xnor_3 g12143(.A(new_n12518), .B(new_n12516), .Y(new_n12520));
  xnor_3 g12144(.A(new_n12504), .B(new_n12377), .Y(new_n12521));
  not_3  g12145(.A(new_n12336), .Y(new_n12522));
  xnor_3 g12146(.A(new_n11245), .B(new_n11207), .Y(new_n12523));
  nand_4 g12147(.A(new_n12523), .B(new_n11173), .Y(new_n12524));
  nand_4 g12148(.A(new_n12524), .B(new_n11169), .Y(new_n12525));
  nor_4  g12149(.A(new_n12525), .B(new_n12522), .Y(new_n12526));
  nor_4  g12150(.A(new_n12526), .B(new_n12341), .Y(new_n12527));
  xnor_3 g12151(.A(new_n12527), .B(new_n12521), .Y(new_n12528));
  nor_4  g12152(.A(new_n12528), .B(new_n12520), .Y(new_n12529));
  nor_4  g12153(.A(new_n12529), .B(new_n12519), .Y(new_n12530));
  xnor_3 g12154(.A(new_n12530), .B(new_n12513), .Y(n5132));
  xor_3  g12155(.A(new_n11946), .B(new_n11933), .Y(n5191));
  nor_4  g12156(.A(new_n3991), .B(new_n3845), .Y(new_n12533));
  nor_4  g12157(.A(new_n12533), .B(new_n3848), .Y(new_n12534));
  nor_4  g12158(.A(new_n3977), .B(new_n3940), .Y(new_n12535));
  nor_4  g12159(.A(new_n3982), .B(new_n3978), .Y(new_n12536));
  nor_4  g12160(.A(new_n12536), .B(new_n12535), .Y(new_n12537));
  not_3  g12161(.A(new_n12537), .Y(new_n12538));
  not_3  g12162(.A(new_n3352), .Y(new_n12539));
  nand_4 g12163(.A(new_n3384), .B(new_n12539), .Y(new_n12540));
  nand_4 g12164(.A(new_n3407), .B(new_n3385), .Y(new_n12541));
  nand_4 g12165(.A(new_n12541), .B(new_n12540), .Y(new_n12542));
  nor_4  g12166(.A(new_n3906), .B(new_n3903), .Y(new_n12543));
  nor_4  g12167(.A(new_n3921), .B(new_n3907), .Y(new_n12544));
  nor_4  g12168(.A(new_n12544), .B(new_n12543), .Y(new_n12545));
  xnor_3 g12169(.A(new_n12545), .B(new_n12542), .Y(new_n12546));
  nand_4 g12170(.A(n1835), .B(n1333), .Y(new_n12547));
  nand_4 g12171(.A(n9637), .B(n3172), .Y(new_n12548));
  xor_3  g12172(.A(new_n12548), .B(new_n12547), .Y(new_n12549));
  nand_4 g12173(.A(n9080), .B(n4921), .Y(new_n12550));
  nand_4 g12174(.A(n11917), .B(n11821), .Y(new_n12551));
  xor_3  g12175(.A(new_n12551), .B(new_n12550), .Y(new_n12552));
  xor_3  g12176(.A(new_n12552), .B(new_n12549), .Y(new_n12553));
  xnor_3 g12177(.A(new_n12553), .B(new_n12546), .Y(new_n12554));
  xnor_3 g12178(.A(new_n12554), .B(new_n12538), .Y(new_n12555));
  nor_4  g12179(.A(new_n3887), .B(new_n3851), .Y(new_n12556));
  nor_4  g12180(.A(new_n3501), .B(new_n3466), .Y(new_n12557));
  nor_4  g12181(.A(new_n3890), .B(new_n12557), .Y(new_n12558));
  nand_4 g12182(.A(new_n12558), .B(new_n3465), .Y(new_n12559));
  nand_4 g12183(.A(new_n12559), .B(new_n3889), .Y(new_n12560));
  nor_4  g12184(.A(new_n12560), .B(new_n3888), .Y(new_n12561));
  nor_4  g12185(.A(new_n12561), .B(new_n12556), .Y(new_n12562));
  nand_4 g12186(.A(new_n3970), .B(new_n3969), .Y(new_n12563));
  not_3  g12187(.A(new_n3967), .Y(new_n12564));
  nand_4 g12188(.A(new_n3972), .B(new_n12564), .Y(new_n12565));
  nand_4 g12189(.A(new_n12565), .B(new_n12563), .Y(new_n12566));
  nand_4 g12190(.A(n10174), .B(n3719), .Y(new_n12567));
  nand_4 g12191(.A(n6877), .B(n4190), .Y(new_n12568));
  nand_4 g12192(.A(n12753), .B(n3602), .Y(new_n12569));
  xor_3  g12193(.A(new_n12569), .B(new_n12568), .Y(new_n12570));
  nand_4 g12194(.A(n4086), .B(n1471), .Y(new_n12571));
  nand_4 g12195(.A(n8065), .B(n2464), .Y(new_n12572));
  nand_4 g12196(.A(n11311), .B(n10439), .Y(new_n12573));
  xor_3  g12197(.A(new_n12573), .B(new_n12572), .Y(new_n12574));
  xnor_3 g12198(.A(new_n12574), .B(new_n12571), .Y(new_n12575));
  nand_4 g12199(.A(n7236), .B(n1357), .Y(new_n12576));
  nand_4 g12200(.A(n7646), .B(n405), .Y(new_n12577));
  xnor_3 g12201(.A(new_n12577), .B(new_n12576), .Y(new_n12578));
  nand_4 g12202(.A(n6126), .B(n4203), .Y(new_n12579));
  nand_4 g12203(.A(n10391), .B(n9400), .Y(new_n12580));
  xnor_3 g12204(.A(new_n12580), .B(new_n12579), .Y(new_n12581));
  xnor_3 g12205(.A(new_n12581), .B(new_n12578), .Y(new_n12582));
  nor_4  g12206(.A(new_n3858), .B(new_n3857), .Y(new_n12583));
  nand_4 g12207(.A(new_n3858), .B(new_n3857), .Y(new_n12584));
  nand_4 g12208(.A(new_n12584), .B(new_n3856), .Y(new_n12585));
  not_3  g12209(.A(new_n12585), .Y(new_n12586));
  nor_4  g12210(.A(new_n12586), .B(new_n12583), .Y(new_n12587));
  xnor_3 g12211(.A(new_n12587), .B(new_n12582), .Y(new_n12588));
  xnor_3 g12212(.A(new_n12588), .B(new_n12575), .Y(new_n12589));
  xnor_3 g12213(.A(new_n12589), .B(new_n12570), .Y(new_n12590));
  nand_4 g12214(.A(n5240), .B(n3842), .Y(new_n12591_1));
  not_3  g12215(.A(new_n12591_1), .Y(new_n12592));
  nand_4 g12216(.A(n8595), .B(n4187), .Y(new_n12593));
  nand_4 g12217(.A(n8433), .B(n4722), .Y(new_n12594));
  xor_3  g12218(.A(new_n12594), .B(new_n12593), .Y(new_n12595));
  xnor_3 g12219(.A(new_n12595), .B(new_n12592), .Y(new_n12596));
  nand_4 g12220(.A(new_n3865_1), .B(new_n3863), .Y(new_n12597));
  nand_4 g12221(.A(new_n3872), .B(new_n3866), .Y(new_n12598));
  nand_4 g12222(.A(new_n12598), .B(new_n12597), .Y(new_n12599));
  and_4  g12223(.A(new_n3870), .B(new_n3869), .Y(new_n12600));
  nor_4  g12224(.A(new_n3871), .B(new_n3868), .Y(new_n12601));
  nor_4  g12225(.A(new_n12601), .B(new_n12600), .Y(new_n12602));
  xnor_3 g12226(.A(new_n12602), .B(new_n12599), .Y(new_n12603));
  xnor_3 g12227(.A(new_n12603), .B(new_n12596), .Y(new_n12604));
  xnor_3 g12228(.A(new_n12604), .B(new_n12590), .Y(new_n12605));
  not_3  g12229(.A(new_n3854), .Y(new_n12606));
  nand_4 g12230(.A(new_n3860), .B(new_n12606), .Y(new_n12607));
  nand_4 g12231(.A(new_n3873), .B(new_n3861), .Y(new_n12608));
  nand_4 g12232(.A(new_n12608), .B(new_n12607), .Y(new_n12609));
  nor_4  g12233(.A(new_n3359), .B(new_n3358), .Y(new_n12610));
  nand_4 g12234(.A(new_n3359), .B(new_n3358), .Y(new_n12611));
  nand_4 g12235(.A(new_n12611), .B(new_n3357), .Y(new_n12612));
  not_3  g12236(.A(new_n12612), .Y(new_n12613));
  nor_4  g12237(.A(new_n12613), .B(new_n12610), .Y(new_n12614));
  xnor_3 g12238(.A(new_n12614), .B(new_n12609), .Y(new_n12615));
  xnor_3 g12239(.A(new_n12615), .B(new_n12605), .Y(new_n12616));
  xnor_3 g12240(.A(new_n12616), .B(new_n12567), .Y(new_n12617));
  xnor_3 g12241(.A(new_n12617), .B(new_n12566), .Y(new_n12618));
  nor_4  g12242(.A(new_n3886), .B(new_n3875), .Y(new_n12619));
  nor_4  g12243(.A(new_n12619), .B(new_n3882), .Y(new_n12620));
  not_3  g12244(.A(new_n3355), .Y(new_n12621));
  nand_4 g12245(.A(new_n3361), .B(new_n12621), .Y(new_n12622));
  not_3  g12246(.A(new_n3377), .Y(new_n12623));
  nand_4 g12247(.A(new_n12623), .B(new_n3362), .Y(new_n12624));
  nand_4 g12248(.A(new_n12624), .B(new_n12622), .Y(new_n12625));
  nor_4  g12249(.A(new_n3365), .B(new_n3364), .Y(new_n12626));
  nor_4  g12250(.A(new_n3376), .B(new_n12626), .Y(new_n12627));
  not_3  g12251(.A(new_n3368), .Y(new_n12628));
  nor_4  g12252(.A(new_n3370), .B(new_n12628), .Y(new_n12629));
  not_3  g12253(.A(new_n3367), .Y(new_n12630));
  nor_4  g12254(.A(new_n3371), .B(new_n12630), .Y(new_n12631));
  nor_4  g12255(.A(new_n12631), .B(new_n12629), .Y(new_n12632));
  nand_4 g12256(.A(n11757), .B(n2577), .Y(new_n12633));
  not_3  g12257(.A(new_n12633), .Y(new_n12634));
  xnor_3 g12258(.A(new_n12634), .B(new_n12632), .Y(new_n12635));
  xnor_3 g12259(.A(new_n12635), .B(new_n12627), .Y(new_n12636));
  xnor_3 g12260(.A(new_n12636), .B(new_n12625), .Y(new_n12637));
  xnor_3 g12261(.A(new_n12637), .B(new_n12620), .Y(new_n12638));
  xnor_3 g12262(.A(new_n12638), .B(new_n12618), .Y(new_n12639));
  xnor_3 g12263(.A(new_n12639), .B(new_n12562), .Y(new_n12640));
  nand_4 g12264(.A(new_n3973), .B(new_n3943), .Y(new_n12641));
  not_3  g12265(.A(new_n3974), .Y(new_n12642));
  not_3  g12266(.A(new_n3976), .Y(new_n12643));
  nand_4 g12267(.A(new_n12643), .B(new_n12642), .Y(new_n12644));
  nand_4 g12268(.A(new_n12644), .B(new_n12641), .Y(new_n12645));
  or_4   g12269(.A(new_n3917), .B(new_n3912), .Y(new_n12646));
  not_3  g12270(.A(new_n12646), .Y(new_n12647));
  nor_4  g12271(.A(new_n12647), .B(new_n3918), .Y(new_n12648_1));
  xnor_3 g12272(.A(new_n12648_1), .B(new_n12645), .Y(new_n12649));
  xnor_3 g12273(.A(new_n12649), .B(new_n12640), .Y(new_n12650));
  xnor_3 g12274(.A(new_n12650), .B(new_n12555), .Y(new_n12651));
  not_3  g12275(.A(new_n3893), .Y(new_n12652));
  nand_4 g12276(.A(new_n3983), .B(new_n12652), .Y(new_n12653));
  nand_4 g12277(.A(new_n3990), .B(new_n3984), .Y(new_n12654));
  nand_4 g12278(.A(new_n12654), .B(new_n12653), .Y(new_n12655));
  nor_4  g12279(.A(new_n3930), .B(new_n3896), .Y(new_n12656));
  nor_4  g12280(.A(new_n3939), .B(new_n3931), .Y(new_n12657));
  nor_4  g12281(.A(new_n12657), .B(new_n12656), .Y(new_n12658));
  not_3  g12282(.A(new_n3949), .Y(new_n12659));
  nor_4  g12283(.A(new_n3954), .B(new_n12659), .Y(new_n12660));
  not_3  g12284(.A(new_n3955), .Y(new_n12661));
  nor_4  g12285(.A(new_n3966), .B(new_n12661), .Y(new_n12662));
  nor_4  g12286(.A(new_n12662), .B(new_n12660), .Y(new_n12663));
  nand_4 g12287(.A(new_n3381), .B(new_n3380), .Y(new_n12664));
  not_3  g12288(.A(new_n3378), .Y(new_n12665));
  nand_4 g12289(.A(new_n3383), .B(new_n12665), .Y(new_n12666));
  nand_4 g12290(.A(new_n12666), .B(new_n12664), .Y(new_n12667));
  nand_4 g12291(.A(new_n3927), .B(new_n3925), .Y(new_n12668));
  nand_4 g12292(.A(new_n3929), .B(new_n3922), .Y(new_n12669));
  nand_4 g12293(.A(new_n12669), .B(new_n12668), .Y(new_n12670));
  nand_4 g12294(.A(new_n3910), .B(new_n3908), .Y(new_n12671));
  not_3  g12295(.A(new_n3920), .Y(new_n12672));
  nand_4 g12296(.A(new_n12672), .B(new_n3911), .Y(new_n12673));
  nand_4 g12297(.A(new_n12673), .B(new_n12671), .Y(new_n12674));
  nand_4 g12298(.A(n5283), .B(n503), .Y(new_n12675));
  not_3  g12299(.A(new_n12675), .Y(new_n12676));
  not_3  g12300(.A(new_n3899), .Y(new_n12677));
  nor_4  g12301(.A(new_n3901), .B(new_n12677), .Y(new_n12678));
  nor_4  g12302(.A(new_n3902), .B(new_n3898), .Y(new_n12679));
  nor_4  g12303(.A(new_n12679), .B(new_n12678), .Y(new_n12680));
  xnor_3 g12304(.A(new_n12680), .B(new_n12676), .Y(new_n12681));
  xnor_3 g12305(.A(new_n12681), .B(new_n12674), .Y(new_n12682));
  nor_4  g12306(.A(new_n3958), .B(new_n3957), .Y(new_n12683));
  not_3  g12307(.A(new_n3959), .Y(new_n12684));
  nor_4  g12308(.A(new_n3965), .B(new_n12684), .Y(new_n12685));
  nor_4  g12309(.A(new_n12685), .B(new_n12683), .Y(new_n12686));
  not_3  g12310(.A(new_n3945), .Y(new_n12687));
  nor_4  g12311(.A(new_n3947), .B(new_n12687), .Y(new_n12688));
  not_3  g12312(.A(new_n3944), .Y(new_n12689));
  nor_4  g12313(.A(new_n3948), .B(new_n12689), .Y(new_n12690));
  nor_4  g12314(.A(new_n12690), .B(new_n12688), .Y(new_n12691));
  nand_4 g12315(.A(n5198), .B(n217), .Y(new_n12692));
  not_3  g12316(.A(new_n12692), .Y(new_n12693));
  nand_4 g12317(.A(n11296), .B(n3992), .Y(new_n12694));
  nand_4 g12318(.A(n6611), .B(n6358), .Y(new_n12695));
  xor_3  g12319(.A(new_n12695), .B(new_n12694), .Y(new_n12696));
  xnor_3 g12320(.A(new_n12696), .B(new_n12693), .Y(new_n12697));
  xnor_3 g12321(.A(new_n12697), .B(new_n12691), .Y(new_n12698));
  xnor_3 g12322(.A(new_n12698), .B(new_n12686), .Y(new_n12699));
  nand_4 g12323(.A(n4970), .B(n137), .Y(new_n12700));
  nand_4 g12324(.A(n6797), .B(n4826), .Y(new_n12701));
  nand_4 g12325(.A(n7610), .B(n6294), .Y(new_n12702));
  xor_3  g12326(.A(new_n12702), .B(new_n12701), .Y(new_n12703));
  xnor_3 g12327(.A(new_n12703), .B(new_n12700), .Y(new_n12704_1));
  nor_4  g12328(.A(new_n3963), .B(new_n3962), .Y(new_n12705_1));
  nand_4 g12329(.A(new_n3963), .B(new_n3962), .Y(new_n12706_1));
  nand_4 g12330(.A(new_n12706_1), .B(new_n3961), .Y(new_n12707));
  not_3  g12331(.A(new_n12707), .Y(new_n12708));
  nor_4  g12332(.A(new_n12708), .B(new_n12705_1), .Y(new_n12709_1));
  xnor_3 g12333(.A(new_n12709_1), .B(new_n12704_1), .Y(new_n12710));
  nand_4 g12334(.A(n11478), .B(n10965), .Y(new_n12711));
  not_3  g12335(.A(new_n12711), .Y(new_n12712));
  nand_4 g12336(.A(n11536), .B(n7862), .Y(new_n12713));
  nand_4 g12337(.A(n9956), .B(n6826), .Y(new_n12714));
  xor_3  g12338(.A(new_n12714), .B(new_n12713), .Y(new_n12715));
  xnor_3 g12339(.A(new_n12715), .B(new_n12712), .Y(new_n12716));
  nand_4 g12340(.A(n8384), .B(n6359), .Y(new_n12717));
  nand_4 g12341(.A(n7733), .B(n3146), .Y(new_n12718));
  xor_3  g12342(.A(new_n12718), .B(new_n12717), .Y(new_n12719));
  nand_4 g12343(.A(n12925), .B(n4938), .Y(new_n12720_1));
  nand_4 g12344(.A(n7546), .B(n4805), .Y(new_n12721));
  xor_3  g12345(.A(new_n12721), .B(new_n12720_1), .Y(new_n12722));
  xnor_3 g12346(.A(new_n12722), .B(new_n12719), .Y(new_n12723));
  xnor_3 g12347(.A(new_n12723), .B(new_n12716), .Y(new_n12724));
  xnor_3 g12348(.A(new_n12724), .B(new_n12710), .Y(new_n12725));
  xnor_3 g12349(.A(new_n12725), .B(new_n12699), .Y(new_n12726));
  xnor_3 g12350(.A(new_n12726), .B(new_n12682), .Y(new_n12727));
  xnor_3 g12351(.A(new_n12727), .B(new_n12670), .Y(new_n12728));
  xnor_3 g12352(.A(new_n12728), .B(new_n12667), .Y(new_n12729));
  xnor_3 g12353(.A(new_n12729), .B(new_n12663), .Y(new_n12730));
  xnor_3 g12354(.A(new_n12730), .B(new_n12658), .Y(new_n12731));
  not_3  g12355(.A(new_n12731), .Y(new_n12732));
  xnor_3 g12356(.A(new_n12732), .B(new_n12655), .Y(new_n12733));
  nand_4 g12357(.A(new_n12733), .B(new_n12651), .Y(new_n12734));
  xnor_3 g12358(.A(new_n12554), .B(new_n12537), .Y(new_n12735));
  xnor_3 g12359(.A(new_n12650), .B(new_n12735), .Y(new_n12736));
  xnor_3 g12360(.A(new_n12731), .B(new_n12655), .Y(new_n12737));
  nand_4 g12361(.A(new_n12737), .B(new_n12736), .Y(new_n12738));
  nand_4 g12362(.A(new_n12738), .B(new_n12734), .Y(new_n12739));
  xnor_3 g12363(.A(new_n12739), .B(new_n12534), .Y(n5257));
  not_3  g12364(.A(new_n11956), .Y(new_n12741));
  xor_3  g12365(.A(new_n12741), .B(new_n11943), .Y(n5411));
  xor_3  g12366(.A(new_n3832), .B(new_n3823), .Y(n5435));
  xor_3  g12367(.A(new_n6535), .B(new_n6528), .Y(n5641));
  not_3  g12368(.A(new_n9129), .Y(new_n12745));
  xor_3  g12369(.A(new_n9139), .B(new_n12745), .Y(n5670));
  not_3  g12370(.A(new_n5275), .Y(new_n12747));
  xor_3  g12371(.A(new_n12747), .B(new_n5240_1), .Y(n5693));
  not_3  g12372(.A(new_n1411), .Y(new_n12749));
  xor_3  g12373(.A(new_n1424), .B(new_n12749), .Y(n5934));
  not_3  g12374(.A(new_n11958), .Y(new_n12751));
  xor_3  g12375(.A(new_n11961), .B(new_n12751), .Y(n6089));
  not_3  g12376(.A(new_n8290), .Y(new_n12753_1));
  nand_4 g12377(.A(new_n8292), .B(new_n12753_1), .Y(new_n12754));
  nor_4  g12378(.A(new_n8271), .B(new_n8267), .Y(new_n12755));
  not_3  g12379(.A(new_n12755), .Y(new_n12756));
  nand_4 g12380(.A(new_n8278), .B(new_n8272), .Y(new_n12757));
  nand_4 g12381(.A(new_n12757), .B(new_n12756), .Y(new_n12758));
  nand_4 g12382(.A(n2564), .B(n2253), .Y(new_n12759));
  nand_4 g12383(.A(n9195), .B(n4189), .Y(new_n12760));
  nand_4 g12384(.A(n6687), .B(n3865), .Y(new_n12761));
  nand_4 g12385(.A(new_n12761), .B(new_n12760), .Y(new_n12762));
  not_3  g12386(.A(new_n12760), .Y(new_n12763));
  not_3  g12387(.A(new_n12761), .Y(new_n12764));
  nand_4 g12388(.A(new_n12764), .B(new_n12763), .Y(new_n12765));
  nand_4 g12389(.A(new_n12765), .B(new_n12762), .Y(new_n12766));
  xnor_3 g12390(.A(new_n12766), .B(new_n12759), .Y(new_n12767));
  xnor_3 g12391(.A(new_n12767), .B(new_n12758), .Y(new_n12768));
  not_3  g12392(.A(new_n12768), .Y(new_n12769));
  nor_4  g12393(.A(new_n8270), .B(new_n8269), .Y(new_n12770));
  nand_4 g12394(.A(n6770), .B(n4634), .Y(new_n12771));
  xor_3  g12395(.A(new_n12771), .B(new_n12770), .Y(new_n12772));
  nand_4 g12396(.A(n3627), .B(n2879), .Y(new_n12773));
  not_3  g12397(.A(new_n12773), .Y(new_n12774));
  nand_4 g12398(.A(n10223), .B(n9920), .Y(new_n12775));
  nand_4 g12399(.A(n7265), .B(n4516), .Y(new_n12776));
  xnor_3 g12400(.A(new_n12776), .B(new_n12775), .Y(new_n12777_1));
  xnor_3 g12401(.A(new_n12777_1), .B(new_n12774), .Y(new_n12778));
  not_3  g12402(.A(new_n12778), .Y(new_n12779));
  xnor_3 g12403(.A(new_n12779), .B(new_n12772), .Y(new_n12780));
  not_3  g12404(.A(new_n12780), .Y(new_n12781));
  xor_3  g12405(.A(new_n12781), .B(new_n12769), .Y(new_n12782));
  nand_4 g12406(.A(new_n8283), .B(new_n8280), .Y(new_n12783));
  nor_4  g12407(.A(new_n8282), .B(new_n8281), .Y(new_n12784));
  nor_4  g12408(.A(new_n8289), .B(new_n8285), .Y(new_n12785));
  xnor_3 g12409(.A(new_n12785), .B(new_n12784), .Y(new_n12786));
  nand_4 g12410(.A(new_n12786), .B(new_n12783), .Y(new_n12787));
  xnor_3 g12411(.A(new_n12787), .B(new_n12782), .Y(new_n12788));
  xnor_3 g12412(.A(new_n12788), .B(new_n12754), .Y(new_n12789));
  nor_4  g12413(.A(new_n8293), .B(new_n8266), .Y(new_n12790));
  nor_4  g12414(.A(new_n8294), .B(new_n8264), .Y(new_n12791));
  nor_4  g12415(.A(new_n12791), .B(new_n12790), .Y(new_n12792));
  xnor_3 g12416(.A(new_n12792), .B(new_n12789), .Y(new_n12793));
  nand_4 g12417(.A(new_n8337), .B(new_n8303_1), .Y(new_n12794));
  xnor_3 g12418(.A(new_n8337), .B(new_n8302), .Y(new_n12795));
  nand_4 g12419(.A(new_n12795), .B(new_n8301), .Y(new_n12796));
  nand_4 g12420(.A(new_n12796), .B(new_n12794), .Y(new_n12797));
  not_3  g12421(.A(new_n8308), .Y(new_n12798));
  nand_4 g12422(.A(new_n8317), .B(new_n8312), .Y(new_n12799));
  nand_4 g12423(.A(new_n12799), .B(new_n12798), .Y(new_n12800));
  nand_4 g12424(.A(n12221), .B(n10928), .Y(new_n12801));
  nand_4 g12425(.A(n12145), .B(n6986), .Y(new_n12802));
  nand_4 g12426(.A(n10217), .B(n8336), .Y(new_n12803));
  xnor_3 g12427(.A(new_n12803), .B(new_n12802), .Y(new_n12804));
  xnor_3 g12428(.A(new_n12804), .B(new_n12801), .Y(new_n12805));
  xnor_3 g12429(.A(new_n12805), .B(new_n12800), .Y(new_n12806));
  nor_4  g12430(.A(new_n8306), .B(new_n8305), .Y(new_n12807_1));
  nand_4 g12431(.A(n2522), .B(n2226), .Y(new_n12808));
  xor_3  g12432(.A(new_n12808), .B(new_n12807_1), .Y(new_n12809));
  nand_4 g12433(.A(n10678), .B(n2024), .Y(new_n12810));
  not_3  g12434(.A(new_n12810), .Y(new_n12811));
  nand_4 g12435(.A(n9189), .B(n1094), .Y(new_n12812));
  nand_4 g12436(.A(n7946), .B(n7320), .Y(new_n12813));
  xnor_3 g12437(.A(new_n12813), .B(new_n12812), .Y(new_n12814));
  and_4  g12438(.A(new_n12814), .B(new_n12811), .Y(new_n12815));
  nor_4  g12439(.A(new_n12814), .B(new_n12811), .Y(new_n12816));
  nor_4  g12440(.A(new_n12816), .B(new_n12815), .Y(new_n12817));
  xnor_3 g12441(.A(new_n12817), .B(new_n12809), .Y(new_n12818));
  not_3  g12442(.A(new_n12818), .Y(new_n12819));
  xor_3  g12443(.A(new_n12819), .B(new_n12806), .Y(new_n12820));
  not_3  g12444(.A(new_n12820), .Y(new_n12821));
  nand_4 g12445(.A(new_n8322), .B(new_n8319), .Y(new_n12822));
  nor_4  g12446(.A(new_n8321), .B(new_n8320), .Y(new_n12823));
  nor_4  g12447(.A(new_n8328), .B(new_n8324), .Y(new_n12824));
  xnor_3 g12448(.A(new_n12824), .B(new_n12823), .Y(new_n12825));
  nand_4 g12449(.A(new_n12825), .B(new_n12822), .Y(new_n12826_1));
  xnor_3 g12450(.A(new_n12826_1), .B(new_n12821), .Y(new_n12827));
  xnor_3 g12451(.A(new_n12827), .B(new_n8334), .Y(new_n12828));
  xnor_3 g12452(.A(new_n12828), .B(new_n12797), .Y(new_n12829));
  nor_4  g12453(.A(new_n8372), .B(new_n8369), .Y(new_n12830));
  nor_4  g12454(.A(new_n8358), .B(new_n8357), .Y(new_n12831));
  nand_4 g12455(.A(n7160), .B(n521), .Y(new_n12832));
  not_3  g12456(.A(new_n12832), .Y(new_n12833));
  xor_3  g12457(.A(new_n12833), .B(new_n12831), .Y(new_n12834));
  nand_4 g12458(.A(n2515), .B(n2498), .Y(new_n12835));
  nand_4 g12459(.A(n2558), .B(n1199), .Y(new_n12836));
  nand_4 g12460(.A(n5579), .B(n4828), .Y(new_n12837));
  not_3  g12461(.A(new_n12837), .Y(new_n12838));
  xor_3  g12462(.A(new_n12838), .B(new_n12836), .Y(new_n12839));
  xnor_3 g12463(.A(new_n12839), .B(new_n12835), .Y(new_n12840));
  not_3  g12464(.A(new_n12840), .Y(new_n12841));
  nand_4 g12465(.A(new_n12841), .B(new_n12834), .Y(new_n12842));
  not_3  g12466(.A(new_n12842), .Y(new_n12843));
  nor_4  g12467(.A(new_n12841), .B(new_n12834), .Y(new_n12844));
  nor_4  g12468(.A(new_n12844), .B(new_n12843), .Y(new_n12845));
  not_3  g12469(.A(new_n8355), .Y(new_n12846));
  nand_4 g12470(.A(new_n8359), .B(new_n8356), .Y(new_n12847));
  nand_4 g12471(.A(new_n12847), .B(new_n12846), .Y(new_n12848));
  nand_4 g12472(.A(n12391), .B(n5798), .Y(new_n12849));
  nand_4 g12473(.A(n7891), .B(n6016), .Y(new_n12850));
  nand_4 g12474(.A(n12069), .B(n2347), .Y(new_n12851));
  not_3  g12475(.A(new_n12851), .Y(new_n12852));
  xor_3  g12476(.A(new_n12852), .B(new_n12850), .Y(new_n12853));
  xnor_3 g12477(.A(new_n12853), .B(new_n12849), .Y(new_n12854));
  xnor_3 g12478(.A(new_n12854), .B(new_n12848), .Y(new_n12855));
  xnor_3 g12479(.A(new_n12855), .B(new_n12845), .Y(new_n12856));
  not_3  g12480(.A(new_n8360), .Y(new_n12857));
  not_3  g12481(.A(new_n8364), .Y(new_n12858));
  nand_4 g12482(.A(new_n12858), .B(new_n12857), .Y(new_n12859));
  nor_4  g12483(.A(new_n8362), .B(new_n8361), .Y(new_n12860));
  nor_4  g12484(.A(new_n8368), .B(new_n8365), .Y(new_n12861));
  xnor_3 g12485(.A(new_n12861), .B(new_n12860), .Y(new_n12862));
  nand_4 g12486(.A(new_n12862), .B(new_n12859), .Y(new_n12863));
  xnor_3 g12487(.A(new_n12863), .B(new_n12856), .Y(new_n12864));
  xnor_3 g12488(.A(new_n12864), .B(new_n12830), .Y(new_n12865));
  nor_4  g12489(.A(new_n8373), .B(new_n8349), .Y(new_n12866));
  nor_4  g12490(.A(new_n8374), .B(new_n8348), .Y(new_n12867));
  nor_4  g12491(.A(new_n12867), .B(new_n12866), .Y(new_n12868));
  xnor_3 g12492(.A(new_n12868), .B(new_n12865), .Y(new_n12869));
  nor_4  g12493(.A(new_n8402), .B(new_n8398_1), .Y(new_n12870));
  not_3  g12494(.A(new_n12870), .Y(new_n12871));
  nand_4 g12495(.A(new_n8388), .B(new_n8386), .Y(new_n12872));
  not_3  g12496(.A(new_n12872), .Y(new_n12873));
  nor_4  g12497(.A(new_n12873), .B(new_n8382), .Y(new_n12874));
  not_3  g12498(.A(new_n12874), .Y(new_n12875));
  nand_4 g12499(.A(n11153), .B(n5153), .Y(new_n12876));
  nand_4 g12500(.A(n7270), .B(n5314), .Y(new_n12877));
  nand_4 g12501(.A(n11222), .B(n2507), .Y(new_n12878));
  not_3  g12502(.A(new_n12878), .Y(new_n12879));
  xor_3  g12503(.A(new_n12879), .B(new_n12877), .Y(new_n12880));
  xnor_3 g12504(.A(new_n12880), .B(new_n12876), .Y(new_n12881));
  xnor_3 g12505(.A(new_n12881), .B(new_n12875), .Y(new_n12882));
  nor_4  g12506(.A(new_n8380), .B(new_n8379), .Y(new_n12883));
  not_3  g12507(.A(new_n12883), .Y(new_n12884));
  nand_4 g12508(.A(n996), .B(n806), .Y(new_n12885));
  xor_3  g12509(.A(new_n12885), .B(new_n12884), .Y(new_n12886));
  nand_4 g12510(.A(n9111), .B(n5319), .Y(new_n12887));
  nand_4 g12511(.A(n5767), .B(n3342), .Y(new_n12888));
  nand_4 g12512(.A(n9763), .B(n9457), .Y(new_n12889));
  not_3  g12513(.A(new_n12889), .Y(new_n12890));
  xor_3  g12514(.A(new_n12890), .B(new_n12888), .Y(new_n12891));
  xnor_3 g12515(.A(new_n12891), .B(new_n12887), .Y(new_n12892));
  xnor_3 g12516(.A(new_n12892), .B(new_n12886), .Y(new_n12893));
  xnor_3 g12517(.A(new_n12893), .B(new_n12882), .Y(new_n12894));
  nand_4 g12518(.A(new_n8393), .B(new_n8390), .Y(new_n12895));
  nor_4  g12519(.A(new_n8392), .B(new_n8391), .Y(new_n12896));
  nor_4  g12520(.A(new_n8397), .B(new_n8394), .Y(new_n12897));
  xnor_3 g12521(.A(new_n12897), .B(new_n12896), .Y(new_n12898));
  nand_4 g12522(.A(new_n12898), .B(new_n12895), .Y(new_n12899));
  xnor_3 g12523(.A(new_n12899), .B(new_n12894), .Y(new_n12900));
  xnor_3 g12524(.A(new_n12900), .B(new_n12871), .Y(new_n12901));
  not_3  g12525(.A(new_n8377), .Y(new_n12902));
  not_3  g12526(.A(new_n8403), .Y(new_n12903));
  nor_4  g12527(.A(new_n12903), .B(new_n12902), .Y(new_n12904));
  nor_4  g12528(.A(new_n8407), .B(new_n12904), .Y(new_n12905));
  xnor_3 g12529(.A(new_n12905), .B(new_n12901), .Y(new_n12906));
  xnor_3 g12530(.A(new_n12906), .B(new_n12869), .Y(new_n12907));
  nand_4 g12531(.A(new_n8416), .B(new_n8409), .Y(new_n12908));
  nand_4 g12532(.A(new_n12908), .B(new_n8412), .Y(new_n12909));
  xnor_3 g12533(.A(new_n12909), .B(new_n12907), .Y(new_n12910));
  xnor_3 g12534(.A(new_n12910), .B(new_n12829), .Y(new_n12911));
  nand_4 g12535(.A(new_n8344), .B(new_n8339), .Y(new_n12912));
  nor_4  g12536(.A(new_n8344), .B(new_n8339), .Y(new_n12913));
  not_3  g12537(.A(new_n12912), .Y(new_n12914));
  nor_4  g12538(.A(new_n12914), .B(new_n12913), .Y(new_n12915));
  nand_4 g12539(.A(new_n8417), .B(new_n12915), .Y(new_n12916));
  nand_4 g12540(.A(new_n12916), .B(new_n12912), .Y(new_n12917));
  xnor_3 g12541(.A(new_n12917), .B(new_n12911), .Y(new_n12918));
  not_3  g12542(.A(new_n12918), .Y(new_n12919));
  nand_4 g12543(.A(new_n12919), .B(new_n12793), .Y(new_n12920));
  not_3  g12544(.A(new_n12793), .Y(new_n12921));
  nand_4 g12545(.A(new_n12918), .B(new_n12921), .Y(new_n12922));
  nor_4  g12546(.A(new_n8299), .B(new_n8295), .Y(new_n12923));
  nor_4  g12547(.A(new_n8420), .B(new_n12923), .Y(new_n12924));
  nand_4 g12548(.A(new_n12924), .B(new_n12922), .Y(new_n12925_1));
  nand_4 g12549(.A(new_n12925_1), .B(new_n12920), .Y(new_n12926));
  nor_4  g12550(.A(new_n12910), .B(new_n12829), .Y(new_n12927));
  nor_4  g12551(.A(new_n12917), .B(new_n12911), .Y(new_n12928));
  nor_4  g12552(.A(new_n12928), .B(new_n12927), .Y(new_n12929));
  not_3  g12553(.A(new_n12869), .Y(new_n12930));
  not_3  g12554(.A(new_n12906), .Y(new_n12931));
  nand_4 g12555(.A(new_n12931), .B(new_n12930), .Y(new_n12932));
  nand_4 g12556(.A(new_n12906), .B(new_n12869), .Y(new_n12933));
  nand_4 g12557(.A(new_n12909), .B(new_n12933), .Y(new_n12934));
  nand_4 g12558(.A(new_n12934), .B(new_n12932), .Y(new_n12935));
  nand_4 g12559(.A(new_n12861), .B(new_n12860), .Y(new_n12936));
  not_3  g12560(.A(new_n12856), .Y(new_n12937));
  nand_4 g12561(.A(new_n12863), .B(new_n12937), .Y(new_n12938));
  nand_4 g12562(.A(new_n12938), .B(new_n12936), .Y(new_n12939));
  nand_4 g12563(.A(new_n12785), .B(new_n12784), .Y(new_n12940));
  not_3  g12564(.A(new_n12782), .Y(new_n12941));
  nand_4 g12565(.A(new_n12787), .B(new_n12941), .Y(new_n12942));
  nand_4 g12566(.A(new_n12942), .B(new_n12940), .Y(new_n12943));
  nand_4 g12567(.A(n5579), .B(n2515), .Y(new_n12944));
  nand_4 g12568(.A(n4828), .B(n521), .Y(new_n12945));
  not_3  g12569(.A(new_n12945), .Y(new_n12946));
  xor_3  g12570(.A(new_n12946), .B(new_n12944), .Y(new_n12947_1));
  nor_4  g12571(.A(new_n12837), .B(new_n12836), .Y(new_n12948));
  not_3  g12572(.A(new_n12835), .Y(new_n12949));
  nand_4 g12573(.A(new_n12837), .B(new_n12836), .Y(new_n12950));
  nand_4 g12574(.A(new_n12950), .B(new_n12949), .Y(new_n12951));
  not_3  g12575(.A(new_n12951), .Y(new_n12952));
  nor_4  g12576(.A(new_n12952), .B(new_n12948), .Y(new_n12953));
  nand_4 g12577(.A(n7891), .B(n5798), .Y(new_n12954));
  nand_4 g12578(.A(n12391), .B(n2347), .Y(new_n12955));
  xor_3  g12579(.A(new_n12955), .B(new_n12954), .Y(new_n12956));
  nand_4 g12580(.A(n6687), .B(n2512), .Y(new_n12957));
  nand_4 g12581(.A(n7265), .B(n2087), .Y(new_n12958));
  xor_3  g12582(.A(new_n12958), .B(new_n12957), .Y(new_n12959));
  xnor_3 g12583(.A(new_n12959), .B(new_n12956), .Y(new_n12960));
  xnor_3 g12584(.A(new_n12960), .B(new_n12953), .Y(new_n12961));
  xnor_3 g12585(.A(new_n12961), .B(new_n12947_1), .Y(new_n12962));
  nand_4 g12586(.A(n2498), .B(n1199), .Y(new_n12963));
  nand_4 g12587(.A(new_n12833), .B(new_n12831), .Y(new_n12964));
  nand_4 g12588(.A(new_n12842), .B(new_n12964), .Y(new_n12965));
  xor_3  g12589(.A(new_n12965), .B(new_n12963), .Y(new_n12966));
  xnor_3 g12590(.A(new_n12966), .B(new_n12962), .Y(new_n12967));
  xnor_3 g12591(.A(new_n12967), .B(new_n12943), .Y(new_n12968));
  xnor_3 g12592(.A(new_n12968), .B(new_n12939), .Y(new_n12969));
  xnor_3 g12593(.A(new_n12969), .B(new_n12935), .Y(new_n12970));
  nand_4 g12594(.A(new_n12864), .B(new_n12830), .Y(new_n12971));
  nor_4  g12595(.A(new_n12868), .B(new_n12865), .Y(new_n12972));
  not_3  g12596(.A(new_n12972), .Y(new_n12973));
  nand_4 g12597(.A(new_n12973), .B(new_n12971), .Y(new_n12974));
  nand_4 g12598(.A(new_n12900), .B(new_n12870), .Y(new_n12975));
  nand_4 g12599(.A(new_n12905), .B(new_n12901), .Y(new_n12976));
  nand_4 g12600(.A(new_n12976), .B(new_n12975), .Y(new_n12977));
  nand_4 g12601(.A(new_n12897), .B(new_n12896), .Y(new_n12978));
  not_3  g12602(.A(new_n12894), .Y(new_n12979));
  nand_4 g12603(.A(new_n12899), .B(new_n12979), .Y(new_n12980));
  nand_4 g12604(.A(new_n12980), .B(new_n12978), .Y(new_n12981));
  not_3  g12605(.A(new_n12807_1), .Y(new_n12982));
  nand_4 g12606(.A(new_n12808), .B(new_n12982), .Y(new_n12983));
  not_3  g12607(.A(new_n12809), .Y(new_n12984));
  nand_4 g12608(.A(new_n12817), .B(new_n12984), .Y(new_n12985));
  nand_4 g12609(.A(new_n12985), .B(new_n12983), .Y(new_n12986));
  nand_4 g12610(.A(n9457), .B(n9111), .Y(new_n12987));
  nand_4 g12611(.A(n10678), .B(n9189), .Y(new_n12988));
  nand_4 g12612(.A(n11222), .B(n6431), .Y(new_n12989));
  xor_3  g12613(.A(new_n12989), .B(new_n12988), .Y(new_n12990));
  xnor_3 g12614(.A(new_n12990), .B(new_n12987), .Y(new_n12991));
  xnor_3 g12615(.A(new_n12991), .B(new_n12986), .Y(new_n12992));
  nand_4 g12616(.A(n12145), .B(n2226), .Y(new_n12993));
  nand_4 g12617(.A(n9763), .B(n4817), .Y(new_n12994));
  nand_4 g12618(.A(n5319), .B(n3342), .Y(new_n12995));
  xor_3  g12619(.A(new_n12995), .B(new_n12994), .Y(new_n12996));
  nand_4 g12620(.A(n12221), .B(n6986), .Y(new_n12997));
  nand_4 g12621(.A(n2522), .B(n1094), .Y(new_n12998));
  xor_3  g12622(.A(new_n12998), .B(new_n12997), .Y(new_n12999));
  xnor_3 g12623(.A(new_n12999), .B(new_n12996), .Y(new_n13000));
  xnor_3 g12624(.A(new_n13000), .B(new_n12993), .Y(new_n13001));
  nand_4 g12625(.A(n10928), .B(n10217), .Y(new_n13002));
  not_3  g12626(.A(new_n12812), .Y(new_n13003));
  not_3  g12627(.A(new_n12813), .Y(new_n13004));
  nor_4  g12628(.A(new_n13004), .B(new_n13003), .Y(new_n13005));
  nor_4  g12629(.A(new_n12816), .B(new_n13005), .Y(new_n13006));
  xor_3  g12630(.A(new_n13006), .B(new_n13002), .Y(new_n13007));
  xnor_3 g12631(.A(new_n13007), .B(new_n13001), .Y(new_n13008));
  xnor_3 g12632(.A(new_n13008), .B(new_n12992), .Y(new_n13009));
  xnor_3 g12633(.A(new_n13009), .B(new_n12981), .Y(new_n13010));
  nor_4  g12634(.A(new_n12885), .B(new_n12884), .Y(new_n13011));
  not_3  g12635(.A(new_n12886), .Y(new_n13012));
  nor_4  g12636(.A(new_n12892), .B(new_n13012), .Y(new_n13013));
  nor_4  g12637(.A(new_n13013), .B(new_n13011), .Y(new_n13014));
  not_3  g12638(.A(new_n12888), .Y(new_n13015));
  nor_4  g12639(.A(new_n12890), .B(new_n13015), .Y(new_n13016));
  not_3  g12640(.A(new_n12887), .Y(new_n13017));
  nor_4  g12641(.A(new_n12891), .B(new_n13017), .Y(new_n13018));
  nor_4  g12642(.A(new_n13018), .B(new_n13016), .Y(new_n13019));
  nand_4 g12643(.A(n11153), .B(n2507), .Y(new_n13020));
  nand_4 g12644(.A(n5314), .B(n5153), .Y(new_n13021));
  not_3  g12645(.A(new_n13021), .Y(new_n13022));
  xor_3  g12646(.A(new_n13022), .B(new_n13020), .Y(new_n13023));
  xnor_3 g12647(.A(new_n13023), .B(new_n13019), .Y(new_n13024));
  xnor_3 g12648(.A(new_n13024), .B(new_n13014), .Y(new_n13025));
  nand_4 g12649(.A(n7946), .B(n7523), .Y(new_n13026));
  nand_4 g12650(.A(n9920), .B(n4634), .Y(new_n13027));
  xor_3  g12651(.A(new_n13027), .B(new_n13026), .Y(new_n13028));
  nand_4 g12652(.A(n8336), .B(n7823), .Y(new_n13029));
  nand_4 g12653(.A(n7320), .B(n2024), .Y(new_n13030));
  xor_3  g12654(.A(new_n13030), .B(new_n13029), .Y(new_n13031));
  xnor_3 g12655(.A(new_n13031), .B(new_n13028), .Y(new_n13032));
  not_3  g12656(.A(new_n12759), .Y(new_n13033));
  nand_4 g12657(.A(new_n12762), .B(new_n13033), .Y(new_n13034));
  and_4  g12658(.A(new_n13034), .B(new_n12765), .Y(new_n13035));
  nand_4 g12659(.A(n10223), .B(n3627), .Y(new_n13036));
  nand_4 g12660(.A(n4516), .B(n2879), .Y(new_n13037));
  xor_3  g12661(.A(new_n13037), .B(new_n13036), .Y(new_n13038));
  xnor_3 g12662(.A(new_n13038), .B(new_n13035), .Y(new_n13039));
  xnor_3 g12663(.A(new_n13039), .B(new_n13032), .Y(new_n13040));
  xnor_3 g12664(.A(new_n13040), .B(new_n13025), .Y(new_n13041));
  not_3  g12665(.A(new_n12758), .Y(new_n13042));
  nand_4 g12666(.A(new_n12767), .B(new_n13042), .Y(new_n13043));
  nand_4 g12667(.A(new_n12780), .B(new_n12768), .Y(new_n13044));
  nand_4 g12668(.A(new_n13044), .B(new_n13043), .Y(new_n13045));
  not_3  g12669(.A(new_n12771), .Y(new_n13046));
  nor_4  g12670(.A(new_n13046), .B(new_n12770), .Y(new_n13047));
  nor_4  g12671(.A(new_n12778), .B(new_n12772), .Y(new_n13048));
  nor_4  g12672(.A(new_n13048), .B(new_n13047), .Y(new_n13049));
  nand_4 g12673(.A(n6578), .B(n2558), .Y(new_n13050));
  and_4  g12674(.A(new_n12776), .B(new_n12775), .Y(new_n13051));
  nor_4  g12675(.A(new_n12777_1), .B(new_n12774), .Y(new_n13052));
  nor_4  g12676(.A(new_n13052), .B(new_n13051), .Y(new_n13053));
  nand_4 g12677(.A(n9195), .B(n6770), .Y(new_n13054));
  nand_4 g12678(.A(n4189), .B(n2253), .Y(new_n13055));
  nand_4 g12679(.A(n3865), .B(n2564), .Y(new_n13056));
  xnor_3 g12680(.A(new_n13056), .B(new_n13055), .Y(new_n13057));
  xnor_3 g12681(.A(new_n13057), .B(new_n13054), .Y(new_n13058));
  xnor_3 g12682(.A(new_n13058), .B(new_n13053), .Y(new_n13059));
  xnor_3 g12683(.A(new_n13059), .B(new_n13050), .Y(new_n13060));
  xnor_3 g12684(.A(new_n13060), .B(new_n13049), .Y(new_n13061));
  xnor_3 g12685(.A(new_n13061), .B(new_n13045), .Y(new_n13062));
  not_3  g12686(.A(new_n12800), .Y(new_n13063));
  nand_4 g12687(.A(new_n12805), .B(new_n13063), .Y(new_n13064));
  nand_4 g12688(.A(new_n12818), .B(new_n12806), .Y(new_n13065));
  nand_4 g12689(.A(new_n13065), .B(new_n13064), .Y(new_n13066));
  nor_4  g12690(.A(new_n12803), .B(new_n12802), .Y(new_n13067));
  not_3  g12691(.A(new_n12801), .Y(new_n13068));
  nand_4 g12692(.A(new_n12803), .B(new_n12802), .Y(new_n13069));
  nand_4 g12693(.A(new_n13069), .B(new_n13068), .Y(new_n13070));
  not_3  g12694(.A(new_n13070), .Y(new_n13071));
  nor_4  g12695(.A(new_n13071), .B(new_n13067), .Y(new_n13072));
  xnor_3 g12696(.A(new_n13072), .B(new_n13066), .Y(new_n13073));
  xnor_3 g12697(.A(new_n13073), .B(new_n13062), .Y(new_n13074));
  xnor_3 g12698(.A(new_n13074), .B(new_n13041), .Y(new_n13075));
  xnor_3 g12699(.A(new_n13075), .B(new_n13010), .Y(new_n13076));
  xnor_3 g12700(.A(new_n13076), .B(new_n12977), .Y(new_n13077));
  xnor_3 g12701(.A(new_n13077), .B(new_n12974), .Y(new_n13078));
  not_3  g12702(.A(new_n12754), .Y(new_n13079));
  nand_4 g12703(.A(new_n12788), .B(new_n13079), .Y(new_n13080));
  nand_4 g12704(.A(new_n12792), .B(new_n12789), .Y(new_n13081));
  nand_4 g12705(.A(new_n13081), .B(new_n13080), .Y(new_n13082));
  nand_4 g12706(.A(new_n12824), .B(new_n12823), .Y(new_n13083));
  nand_4 g12707(.A(new_n12826_1), .B(new_n12820), .Y(new_n13084));
  nand_4 g12708(.A(new_n13084), .B(new_n13083), .Y(new_n13085));
  nand_4 g12709(.A(new_n12881), .B(new_n12874), .Y(new_n13086));
  not_3  g12710(.A(new_n12893), .Y(new_n13087));
  nand_4 g12711(.A(new_n13087), .B(new_n12882), .Y(new_n13088));
  nand_4 g12712(.A(new_n13088), .B(new_n13086), .Y(new_n13089));
  not_3  g12713(.A(new_n12877), .Y(new_n13090));
  nor_4  g12714(.A(new_n12879), .B(new_n13090), .Y(new_n13091));
  not_3  g12715(.A(new_n12876), .Y(new_n13092));
  nor_4  g12716(.A(new_n12880), .B(new_n13092), .Y(new_n13093));
  nor_4  g12717(.A(new_n13093), .B(new_n13091), .Y(new_n13094));
  nand_4 g12718(.A(n12069), .B(n1576), .Y(new_n13095));
  nand_4 g12719(.A(n7270), .B(n996), .Y(new_n13096));
  nand_4 g12720(.A(n5767), .B(n806), .Y(new_n13097));
  xor_3  g12721(.A(new_n13097), .B(new_n13096), .Y(new_n13098));
  xor_3  g12722(.A(new_n13098), .B(new_n13095), .Y(new_n13099));
  xnor_3 g12723(.A(new_n13099), .B(new_n13094), .Y(new_n13100));
  xnor_3 g12724(.A(new_n13100), .B(new_n13089), .Y(new_n13101));
  xnor_3 g12725(.A(new_n13101), .B(new_n13085), .Y(new_n13102));
  xnor_3 g12726(.A(new_n13102), .B(new_n13082), .Y(new_n13103));
  xnor_3 g12727(.A(new_n13103), .B(new_n13078), .Y(new_n13104));
  xnor_3 g12728(.A(new_n13104), .B(new_n12970), .Y(new_n13105));
  nand_4 g12729(.A(new_n12827), .B(new_n8334), .Y(new_n13106));
  not_3  g12730(.A(new_n12828), .Y(new_n13107));
  nand_4 g12731(.A(new_n13107), .B(new_n12797), .Y(new_n13108));
  nand_4 g12732(.A(new_n13108), .B(new_n13106), .Y(new_n13109));
  not_3  g12733(.A(new_n12848), .Y(new_n13110));
  nand_4 g12734(.A(new_n12854), .B(new_n13110), .Y(new_n13111));
  not_3  g12735(.A(new_n12845), .Y(new_n13112));
  nand_4 g12736(.A(new_n12855), .B(new_n13112), .Y(new_n13113));
  nand_4 g12737(.A(new_n13113), .B(new_n13111), .Y(new_n13114));
  nand_4 g12738(.A(n7160), .B(n6016), .Y(new_n13115));
  not_3  g12739(.A(new_n12850), .Y(new_n13116));
  nor_4  g12740(.A(new_n12852), .B(new_n13116), .Y(new_n13117));
  not_3  g12741(.A(new_n12849), .Y(new_n13118));
  nor_4  g12742(.A(new_n12853), .B(new_n13118), .Y(new_n13119));
  nor_4  g12743(.A(new_n13119), .B(new_n13117), .Y(new_n13120));
  xor_3  g12744(.A(new_n13120), .B(new_n13115), .Y(new_n13121));
  xor_3  g12745(.A(new_n13121), .B(new_n13114), .Y(new_n13122));
  xnor_3 g12746(.A(new_n13122), .B(new_n13109), .Y(new_n13123));
  xnor_3 g12747(.A(new_n13123), .B(new_n13105), .Y(new_n13124));
  xnor_3 g12748(.A(new_n13124), .B(new_n12929), .Y(new_n13125));
  xnor_3 g12749(.A(new_n13125), .B(new_n12926), .Y(n6192));
  xor_3  g12750(.A(new_n1060), .B(new_n1024), .Y(n6273));
  xnor_3 g12751(.A(new_n8246), .B(new_n8245), .Y(n6445));
  nand_4 g12752(.A(new_n9999), .B(new_n9998), .Y(new_n13129));
  xnor_3 g12753(.A(new_n13129), .B(new_n10025), .Y(n6645));
  not_3  g12754(.A(new_n8472), .Y(new_n13131));
  xor_3  g12755(.A(new_n8475), .B(new_n13131), .Y(n6689));
  xor_3  g12756(.A(new_n1412), .B(new_n1320), .Y(n6742));
  not_3  g12757(.A(new_n2154), .Y(new_n13134));
  xnor_3 g12758(.A(new_n2195), .B(new_n13134), .Y(n6809));
  not_3  g12759(.A(new_n7257), .Y(new_n13136));
  xor_3  g12760(.A(new_n7259), .B(new_n13136), .Y(n6822));
  not_3  g12761(.A(new_n11954), .Y(new_n13138));
  xor_3  g12762(.A(new_n13138), .B(new_n11953), .Y(n6860));
  not_3  g12763(.A(new_n10013), .Y(new_n13140));
  xor_3  g12764(.A(new_n10021), .B(new_n13140), .Y(n7193));
  nand_4 g12765(.A(new_n8237), .B(new_n8236_1), .Y(new_n13142));
  xnor_3 g12766(.A(new_n13142), .B(new_n8248), .Y(n7568));
  not_3  g12767(.A(new_n1422), .Y(new_n13144));
  xor_3  g12768(.A(new_n13144), .B(new_n1421), .Y(n7676));
  nand_4 g12769(.A(new_n471), .B(new_n464), .Y(new_n13146));
  not_3  g12770(.A(new_n483), .Y(new_n13147));
  nand_4 g12771(.A(new_n13147), .B(new_n472), .Y(new_n13148));
  nand_4 g12772(.A(new_n13148), .B(new_n13146), .Y(new_n13149));
  nand_4 g12773(.A(n10644), .B(n7354), .Y(new_n13150));
  xor_3  g12774(.A(new_n13150), .B(new_n13149), .Y(new_n13151));
  nand_4 g12775(.A(new_n969), .B(new_n959), .Y(new_n13152));
  nand_4 g12776(.A(new_n982), .B(new_n970), .Y(new_n13153));
  nand_4 g12777(.A(new_n13153), .B(new_n13152), .Y(new_n13154));
  not_3  g12778(.A(new_n977), .Y(new_n13155));
  nor_4  g12779(.A(new_n979), .B(new_n13155), .Y(new_n13156));
  nor_4  g12780(.A(new_n980), .B(new_n976), .Y(new_n13157));
  nor_4  g12781(.A(new_n13157), .B(new_n13156), .Y(new_n13158));
  xnor_3 g12782(.A(new_n13158), .B(new_n13154), .Y(new_n13159));
  xnor_3 g12783(.A(new_n13159), .B(new_n13151), .Y(new_n13160));
  nor_4  g12784(.A(new_n475), .B(new_n474), .Y(new_n13161));
  not_3  g12785(.A(new_n476), .Y(new_n13162));
  nor_4  g12786(.A(new_n482), .B(new_n13162), .Y(new_n13163));
  nor_4  g12787(.A(new_n13163), .B(new_n13161), .Y(new_n13164));
  nand_4 g12788(.A(n3986), .B(n1980), .Y(new_n13165));
  not_3  g12789(.A(new_n13165), .Y(new_n13166));
  nor_4  g12790(.A(new_n480), .B(new_n479), .Y(new_n13167));
  nand_4 g12791(.A(new_n480), .B(new_n479), .Y(new_n13168));
  nand_4 g12792(.A(new_n13168), .B(new_n478), .Y(new_n13169));
  not_3  g12793(.A(new_n13169), .Y(new_n13170));
  nor_4  g12794(.A(new_n13170), .B(new_n13167), .Y(new_n13171));
  nand_4 g12795(.A(n7436), .B(n4141), .Y(new_n13172));
  nand_4 g12796(.A(n9241), .B(n1209), .Y(new_n13173));
  not_3  g12797(.A(new_n13173), .Y(new_n13174));
  xor_3  g12798(.A(new_n13174), .B(new_n13172), .Y(new_n13175));
  nand_4 g12799(.A(n8276), .B(n5105), .Y(new_n13176));
  nand_4 g12800(.A(n8236), .B(n6776), .Y(new_n13177));
  xor_3  g12801(.A(new_n13177), .B(new_n13176), .Y(new_n13178));
  xor_3  g12802(.A(new_n13178), .B(new_n13175), .Y(new_n13179));
  xnor_3 g12803(.A(new_n13179), .B(new_n13171), .Y(new_n13180));
  xnor_3 g12804(.A(new_n13180), .B(new_n13166), .Y(new_n13181));
  xnor_3 g12805(.A(new_n13181), .B(new_n13164), .Y(new_n13182));
  or_4   g12806(.A(new_n489), .B(new_n488), .Y(new_n13183));
  not_3  g12807(.A(new_n484), .Y(new_n13184));
  nand_4 g12808(.A(new_n491), .B(new_n13184), .Y(new_n13185));
  nand_4 g12809(.A(new_n13185), .B(new_n13183), .Y(new_n13186));
  xnor_3 g12810(.A(new_n13186), .B(new_n13182), .Y(new_n13187));
  xnor_3 g12811(.A(new_n13187), .B(new_n13160), .Y(new_n13188));
  nand_4 g12812(.A(new_n620), .B(new_n586), .Y(new_n13189));
  not_3  g12813(.A(new_n642), .Y(new_n13190));
  nand_4 g12814(.A(new_n13190), .B(new_n621), .Y(new_n13191));
  nand_4 g12815(.A(new_n13191), .B(new_n13189), .Y(new_n13192));
  nand_4 g12816(.A(new_n751), .B(new_n719), .Y(new_n13193));
  not_3  g12817(.A(new_n752), .Y(new_n13194));
  nand_4 g12818(.A(new_n773), .B(new_n13194), .Y(new_n13195));
  nand_4 g12819(.A(new_n13195), .B(new_n13193), .Y(new_n13196));
  nand_4 g12820(.A(n12706), .B(n5964), .Y(new_n13197));
  nand_4 g12821(.A(n4005), .B(n1097), .Y(new_n13198));
  xor_3  g12822(.A(new_n13198), .B(new_n13197), .Y(new_n13199));
  nand_4 g12823(.A(n12720), .B(n12025), .Y(new_n13200));
  nand_4 g12824(.A(n11257), .B(n2509), .Y(new_n13201));
  xor_3  g12825(.A(new_n13201), .B(new_n13200), .Y(new_n13202));
  xor_3  g12826(.A(new_n13202), .B(new_n13199), .Y(new_n13203));
  nand_4 g12827(.A(n12705), .B(n2508), .Y(new_n13204));
  not_3  g12828(.A(new_n961), .Y(new_n13205));
  nand_4 g12829(.A(new_n964), .B(new_n13205), .Y(new_n13206));
  and_4  g12830(.A(new_n13206), .B(new_n967), .Y(new_n13207));
  xor_3  g12831(.A(new_n13207), .B(new_n13204), .Y(new_n13208));
  xnor_3 g12832(.A(new_n13208), .B(new_n13203), .Y(new_n13209));
  xnor_3 g12833(.A(new_n13209), .B(new_n13196), .Y(new_n13210));
  xnor_3 g12834(.A(new_n13210), .B(new_n13192), .Y(new_n13211));
  nand_4 g12835(.A(new_n617), .B(new_n615_1), .Y(new_n13212));
  not_3  g12836(.A(new_n612), .Y(new_n13213));
  nand_4 g12837(.A(new_n619), .B(new_n13213), .Y(new_n13214));
  nand_4 g12838(.A(new_n13214), .B(new_n13212), .Y(new_n13215));
  not_3  g12839(.A(new_n985), .Y(new_n13216));
  nor_4  g12840(.A(new_n986), .B(new_n13216), .Y(new_n13217));
  nor_4  g12841(.A(new_n988), .B(new_n984), .Y(new_n13218));
  nor_4  g12842(.A(new_n13218), .B(new_n13217), .Y(new_n13219));
  xnor_3 g12843(.A(new_n13219), .B(new_n13215), .Y(new_n13220));
  nand_4 g12844(.A(n12704), .B(n2393), .Y(new_n13221));
  not_3  g12845(.A(new_n732), .Y(new_n13222));
  nor_4  g12846(.A(new_n743), .B(new_n13222), .Y(new_n13223));
  nor_4  g12847(.A(new_n13223), .B(new_n731), .Y(new_n13224));
  not_3  g12848(.A(new_n724), .Y(new_n13225));
  nor_4  g12849(.A(new_n726), .B(new_n13225), .Y(new_n13226));
  not_3  g12850(.A(new_n723), .Y(new_n13227));
  nor_4  g12851(.A(new_n727), .B(new_n13227), .Y(new_n13228));
  nor_4  g12852(.A(new_n13228), .B(new_n13226), .Y(new_n13229));
  nand_4 g12853(.A(n4499), .B(n1564), .Y(new_n13230));
  nand_4 g12854(.A(n12648), .B(n6806), .Y(new_n13231));
  xor_3  g12855(.A(new_n13231), .B(new_n13230), .Y(new_n13232));
  nand_4 g12856(.A(n10547), .B(n6038), .Y(new_n13233));
  nand_4 g12857(.A(n5069), .B(n2530), .Y(new_n13234));
  xor_3  g12858(.A(new_n13234), .B(new_n13233), .Y(new_n13235));
  xnor_3 g12859(.A(new_n13235), .B(new_n13232), .Y(new_n13236));
  xnor_3 g12860(.A(new_n13236), .B(new_n13229), .Y(new_n13237));
  nand_4 g12861(.A(n5694), .B(n5331), .Y(new_n13238));
  nand_4 g12862(.A(n7388), .B(n4903), .Y(new_n13239));
  not_3  g12863(.A(new_n13239), .Y(new_n13240));
  xor_3  g12864(.A(new_n13240), .B(new_n13238), .Y(new_n13241));
  xnor_3 g12865(.A(new_n13241), .B(new_n13237), .Y(new_n13242));
  nor_4  g12866(.A(new_n735), .B(new_n734), .Y(new_n13243));
  not_3  g12867(.A(new_n736), .Y(new_n13244));
  nor_4  g12868(.A(new_n742), .B(new_n13244), .Y(new_n13245));
  nor_4  g12869(.A(new_n13245), .B(new_n13243), .Y(new_n13246));
  not_3  g12870(.A(new_n738), .Y(new_n13247));
  nor_4  g12871(.A(new_n740), .B(new_n13247), .Y(new_n13248));
  not_3  g12872(.A(new_n737), .Y(new_n13249));
  nor_4  g12873(.A(new_n741), .B(new_n13249), .Y(new_n13250));
  nor_4  g12874(.A(new_n13250), .B(new_n13248), .Y(new_n13251));
  nand_4 g12875(.A(n7294), .B(n5860), .Y(new_n13252));
  nand_4 g12876(.A(n11892), .B(n5814), .Y(new_n13253));
  xor_3  g12877(.A(new_n13253), .B(new_n13252), .Y(new_n13254));
  xnor_3 g12878(.A(new_n13254), .B(new_n13251), .Y(new_n13255));
  xnor_3 g12879(.A(new_n13255), .B(new_n13246), .Y(new_n13256));
  xnor_3 g12880(.A(new_n13256), .B(new_n13242), .Y(new_n13257));
  xnor_3 g12881(.A(new_n13257), .B(new_n13224), .Y(new_n13258));
  xnor_3 g12882(.A(new_n13258), .B(new_n13221), .Y(new_n13259));
  and_4  g12883(.A(new_n748), .B(new_n747), .Y(new_n13260));
  not_3  g12884(.A(new_n750), .Y(new_n13261));
  nor_4  g12885(.A(new_n13261), .B(new_n744), .Y(new_n13262));
  nor_4  g12886(.A(new_n13262), .B(new_n13260), .Y(new_n13263));
  nand_4 g12887(.A(new_n597), .B(new_n590), .Y(new_n13264));
  not_3  g12888(.A(new_n611), .Y(new_n13265));
  nand_4 g12889(.A(new_n13265), .B(new_n598), .Y(new_n13266));
  nand_4 g12890(.A(new_n13266), .B(new_n13264), .Y(new_n13267));
  not_3  g12891(.A(new_n593), .Y(new_n13268));
  nor_4  g12892(.A(new_n595), .B(new_n13268), .Y(new_n13269));
  not_3  g12893(.A(new_n592), .Y(new_n13270));
  nor_4  g12894(.A(new_n596), .B(new_n13270), .Y(new_n13271));
  nor_4  g12895(.A(new_n13271), .B(new_n13269), .Y(new_n13272));
  not_3  g12896(.A(new_n606), .Y(new_n13273));
  nor_4  g12897(.A(new_n608), .B(new_n13273), .Y(new_n13274));
  nor_4  g12898(.A(new_n609), .B(new_n605), .Y(new_n13275));
  nor_4  g12899(.A(new_n13275), .B(new_n13274), .Y(new_n13276));
  xnor_3 g12900(.A(new_n13276), .B(new_n13272), .Y(new_n13277));
  nand_4 g12901(.A(n10545), .B(n2802), .Y(new_n13278));
  nand_4 g12902(.A(n12044), .B(n8476), .Y(new_n13279));
  xor_3  g12903(.A(new_n13279), .B(new_n13278), .Y(new_n13280));
  nand_4 g12904(.A(n7690), .B(n533), .Y(new_n13281));
  nand_4 g12905(.A(n3616), .B(n1512), .Y(new_n13282));
  xor_3  g12906(.A(new_n13282), .B(new_n13281), .Y(new_n13283));
  xnor_3 g12907(.A(new_n13283), .B(new_n13280), .Y(new_n13284));
  xnor_3 g12908(.A(new_n13284), .B(new_n13277), .Y(new_n13285));
  nand_4 g12909(.A(n5305), .B(n615), .Y(new_n13286));
  not_3  g12910(.A(new_n13286), .Y(new_n13287));
  nand_4 g12911(.A(new_n601), .B(new_n599), .Y(new_n13288));
  nand_4 g12912(.A(new_n610), .B(new_n602), .Y(new_n13289));
  nand_4 g12913(.A(new_n13289), .B(new_n13288), .Y(new_n13290));
  xnor_3 g12914(.A(new_n13290), .B(new_n13287), .Y(new_n13291));
  xnor_3 g12915(.A(new_n13291), .B(new_n13285), .Y(new_n13292));
  xnor_3 g12916(.A(new_n13292), .B(new_n13267), .Y(new_n13293));
  nand_4 g12917(.A(n10848), .B(n5857), .Y(new_n13294));
  nand_4 g12918(.A(n7965), .B(n1906), .Y(new_n13295));
  not_3  g12919(.A(new_n13295), .Y(new_n13296));
  xor_3  g12920(.A(new_n13296), .B(new_n13294), .Y(new_n13297));
  not_3  g12921(.A(new_n467), .Y(new_n13298));
  nor_4  g12922(.A(new_n469), .B(new_n13298), .Y(new_n13299));
  not_3  g12923(.A(new_n466), .Y(new_n13300));
  nor_4  g12924(.A(new_n470), .B(new_n13300), .Y(new_n13301));
  nor_4  g12925(.A(new_n13301), .B(new_n13299), .Y(new_n13302));
  nand_4 g12926(.A(n8028), .B(n45), .Y(new_n13303));
  nand_4 g12927(.A(n12299), .B(n4928), .Y(new_n13304));
  xor_3  g12928(.A(new_n13304), .B(new_n13303), .Y(new_n13305));
  xnor_3 g12929(.A(new_n13305), .B(new_n13302), .Y(new_n13306));
  xnor_3 g12930(.A(new_n13306), .B(new_n13297), .Y(new_n13307));
  nand_4 g12931(.A(new_n973), .B(new_n971), .Y(new_n13308));
  nand_4 g12932(.A(new_n981), .B(new_n974), .Y(new_n13309));
  nand_4 g12933(.A(new_n13309), .B(new_n13308), .Y(new_n13310));
  nand_4 g12934(.A(n8759), .B(n783), .Y(new_n13311));
  nand_4 g12935(.A(n10510), .B(n7500), .Y(new_n13312));
  xor_3  g12936(.A(new_n13312), .B(new_n13311), .Y(new_n13313));
  xnor_3 g12937(.A(new_n13313), .B(new_n13310), .Y(new_n13314));
  xnor_3 g12938(.A(new_n13314), .B(new_n13307), .Y(new_n13315));
  xnor_3 g12939(.A(new_n13315), .B(new_n13293), .Y(new_n13316));
  xnor_3 g12940(.A(new_n13316), .B(new_n13263), .Y(new_n13317));
  xnor_3 g12941(.A(new_n13317), .B(new_n13259), .Y(new_n13318));
  xnor_3 g12942(.A(new_n13318), .B(new_n13220), .Y(new_n13319));
  xnor_3 g12943(.A(new_n13319), .B(new_n13211), .Y(new_n13320));
  xnor_3 g12944(.A(new_n13320), .B(new_n13188), .Y(new_n13321));
  nor_4  g12945(.A(new_n989), .B(new_n955), .Y(new_n13322));
  not_3  g12946(.A(new_n1010), .Y(new_n13323));
  nor_4  g12947(.A(new_n13323), .B(new_n990), .Y(new_n13324));
  nor_4  g12948(.A(new_n13324), .B(new_n13322), .Y(new_n13325));
  nor_4  g12949(.A(new_n774), .B(new_n643), .Y(new_n13326));
  nor_4  g12950(.A(new_n826), .B(new_n775), .Y(new_n13327));
  nor_4  g12951(.A(new_n13327), .B(new_n13326), .Y(new_n13328));
  xnor_3 g12952(.A(new_n13328), .B(new_n13325), .Y(new_n13329));
  xnor_3 g12953(.A(new_n13329), .B(new_n13321), .Y(new_n13330));
  not_3  g12954(.A(new_n513), .Y(new_n13331));
  nand_4 g12955(.A(new_n827), .B(new_n13331), .Y(new_n13332));
  nand_4 g12956(.A(new_n878), .B(new_n828), .Y(new_n13333));
  nand_4 g12957(.A(new_n13333), .B(new_n13332), .Y(new_n13334));
  not_3  g12958(.A(new_n461), .Y(new_n13335));
  nand_4 g12959(.A(new_n492), .B(new_n13335), .Y(new_n13336));
  nand_4 g12960(.A(new_n512), .B(new_n493), .Y(new_n13337));
  nand_4 g12961(.A(new_n13337), .B(new_n13336), .Y(new_n13338));
  nand_4 g12962(.A(n4312), .B(n2585), .Y(new_n13339));
  xor_3  g12963(.A(new_n13339), .B(new_n13338), .Y(new_n13340));
  xnor_3 g12964(.A(new_n13340), .B(new_n13334), .Y(new_n13341));
  not_3  g12965(.A(new_n1065), .Y(new_n13342));
  nand_4 g12966(.A(new_n1066), .B(new_n879), .Y(new_n13343));
  nand_4 g12967(.A(new_n13343), .B(new_n13342), .Y(new_n13344));
  xnor_3 g12968(.A(new_n13344), .B(new_n13341), .Y(new_n13345));
  xnor_3 g12969(.A(new_n13345), .B(new_n13330), .Y(n7966));
  not_3  g12970(.A(new_n12924), .Y(new_n13347));
  nand_4 g12971(.A(new_n12922), .B(new_n12920), .Y(new_n13348));
  xnor_3 g12972(.A(new_n13348), .B(new_n13347), .Y(n7981));
  nand_4 g12973(.A(new_n12530), .B(new_n12512), .Y(new_n13350));
  nand_4 g12974(.A(new_n13350), .B(new_n12511_1), .Y(new_n13351));
  nor_4  g12975(.A(new_n12521), .B(new_n12526), .Y(new_n13352));
  nor_4  g12976(.A(new_n13352), .B(new_n12341), .Y(new_n13353));
  nor_4  g12977(.A(new_n13353), .B(new_n12335), .Y(new_n13354));
  xnor_3 g12978(.A(new_n13353), .B(new_n12335), .Y(new_n13355));
  nor_4  g12979(.A(new_n12507), .B(new_n13355), .Y(new_n13356));
  nor_4  g12980(.A(new_n13356), .B(new_n13354), .Y(new_n13357));
  not_3  g12981(.A(new_n12215), .Y(new_n13358));
  nand_4 g12982(.A(new_n12253), .B(new_n13358), .Y(new_n13359));
  nand_4 g12983(.A(new_n12263), .B(new_n12254), .Y(new_n13360));
  nand_4 g12984(.A(new_n13360), .B(new_n13359), .Y(new_n13361));
  nand_4 g12985(.A(new_n12247_1), .B(new_n12246), .Y(new_n13362));
  nand_4 g12986(.A(new_n12251), .B(new_n13362), .Y(new_n13363));
  nand_4 g12987(.A(n12391), .B(n1353), .Y(new_n13364));
  not_3  g12988(.A(new_n13364), .Y(new_n13365));
  nand_4 g12989(.A(new_n12471), .B(new_n12460), .Y(new_n13366));
  nand_4 g12990(.A(new_n12486), .B(new_n12472), .Y(new_n13367));
  nand_4 g12991(.A(new_n13367), .B(new_n13366), .Y(new_n13368));
  not_3  g12992(.A(new_n12473), .Y(new_n13369));
  nor_4  g12993(.A(new_n12474), .B(new_n13369), .Y(new_n13370));
  nor_4  g12994(.A(new_n12485), .B(new_n12475), .Y(new_n13371));
  nor_4  g12995(.A(new_n13371), .B(new_n13370), .Y(new_n13372));
  nand_4 g12996(.A(n7891), .B(n447), .Y(new_n13373));
  nand_4 g12997(.A(new_n12466), .B(new_n12463), .Y(new_n13374));
  nand_4 g12998(.A(new_n13374), .B(new_n12469), .Y(new_n13375));
  xor_3  g12999(.A(new_n13375), .B(new_n13373), .Y(new_n13376));
  nand_4 g13000(.A(new_n12480), .B(new_n12477), .Y(new_n13377));
  and_4  g13001(.A(new_n13377), .B(new_n12483), .Y(new_n13378));
  nand_4 g13002(.A(n11407), .B(n2087), .Y(new_n13379));
  nand_4 g13003(.A(n6687), .B(n6604), .Y(new_n13380));
  xor_3  g13004(.A(new_n13380), .B(new_n13379), .Y(new_n13381));
  xnor_3 g13005(.A(new_n13381), .B(new_n13378), .Y(new_n13382));
  xnor_3 g13006(.A(new_n13382), .B(new_n13376), .Y(new_n13383));
  xnor_3 g13007(.A(new_n13383), .B(new_n13372), .Y(new_n13384));
  xnor_3 g13008(.A(new_n13384), .B(new_n13368), .Y(new_n13385));
  nand_4 g13009(.A(new_n12428), .B(new_n12421), .Y(new_n13386));
  nand_4 g13010(.A(new_n12439), .B(new_n12429), .Y(new_n13387));
  nand_4 g13011(.A(new_n13387), .B(new_n13386), .Y(new_n13388));
  not_3  g13012(.A(new_n12424), .Y(new_n13389));
  nor_4  g13013(.A(new_n12426), .B(new_n13389), .Y(new_n13390));
  not_3  g13014(.A(new_n12423), .Y(new_n13391));
  nor_4  g13015(.A(new_n12427), .B(new_n13391), .Y(new_n13392));
  nor_4  g13016(.A(new_n13392), .B(new_n13390), .Y(new_n13393));
  xnor_3 g13017(.A(new_n13393), .B(new_n13388), .Y(new_n13394));
  xnor_3 g13018(.A(new_n13394), .B(new_n13385), .Y(new_n13395));
  xnor_3 g13019(.A(new_n13395), .B(new_n13365), .Y(new_n13396));
  not_3  g13020(.A(new_n12431), .Y(new_n13397));
  nand_4 g13021(.A(new_n13397), .B(new_n12430), .Y(new_n13398));
  not_3  g13022(.A(new_n12432), .Y(new_n13399));
  not_3  g13023(.A(new_n12438), .Y(new_n13400));
  nand_4 g13024(.A(new_n13400), .B(new_n13399), .Y(new_n13401));
  nand_4 g13025(.A(new_n13401), .B(new_n13398), .Y(new_n13402));
  nand_4 g13026(.A(n12709), .B(n7523), .Y(new_n13403));
  nand_4 g13027(.A(n12777), .B(n2515), .Y(new_n13404));
  xor_3  g13028(.A(new_n13404), .B(new_n13403), .Y(new_n13405));
  xor_3  g13029(.A(new_n13405), .B(new_n13402), .Y(new_n13406));
  nand_4 g13030(.A(n7159), .B(n1199), .Y(new_n13407));
  nand_4 g13031(.A(n6441), .B(n5314), .Y(new_n13408));
  xor_3  g13032(.A(new_n13408), .B(new_n13407), .Y(new_n13409));
  nand_4 g13033(.A(n11791), .B(n5767), .Y(new_n13410));
  nand_4 g13034(.A(n6254), .B(n4828), .Y(new_n13411));
  xor_3  g13035(.A(new_n13411), .B(new_n13410), .Y(new_n13412));
  xnor_3 g13036(.A(new_n13412), .B(new_n13409), .Y(new_n13413));
  nand_4 g13037(.A(n12069), .B(n4436), .Y(new_n13414));
  nand_4 g13038(.A(n11999), .B(n11153), .Y(new_n13415));
  xor_3  g13039(.A(new_n13415), .B(new_n13414), .Y(new_n13416));
  nand_4 g13040(.A(n12489), .B(n6578), .Y(new_n13417));
  nand_4 g13041(.A(n12947), .B(n996), .Y(new_n13418));
  xor_3  g13042(.A(new_n13418), .B(new_n13417), .Y(new_n13419));
  xnor_3 g13043(.A(new_n13419), .B(new_n13416), .Y(new_n13420));
  xnor_3 g13044(.A(new_n13420), .B(new_n13413), .Y(new_n13421));
  nand_4 g13045(.A(n11967), .B(n7160), .Y(new_n13422));
  not_3  g13046(.A(new_n13422), .Y(new_n13423));
  not_3  g13047(.A(new_n12434), .Y(new_n13424));
  nor_4  g13048(.A(new_n12436), .B(new_n13424), .Y(new_n13425));
  not_3  g13049(.A(new_n12433), .Y(new_n13426));
  nor_4  g13050(.A(new_n12437), .B(new_n13426), .Y(new_n13427));
  nor_4  g13051(.A(new_n13427), .B(new_n13425), .Y(new_n13428));
  xnor_3 g13052(.A(new_n13428), .B(new_n13423), .Y(new_n13429));
  xnor_3 g13053(.A(new_n13429), .B(new_n13421), .Y(new_n13430));
  xnor_3 g13054(.A(new_n13430), .B(new_n13406), .Y(new_n13431));
  xnor_3 g13055(.A(new_n13431), .B(new_n13396), .Y(new_n13432));
  xnor_3 g13056(.A(new_n13432), .B(new_n13363), .Y(new_n13433));
  xnor_3 g13057(.A(new_n13433), .B(new_n13361), .Y(new_n13434));
  not_3  g13058(.A(new_n12304), .Y(new_n13435));
  nand_4 g13059(.A(new_n12333), .B(new_n13435), .Y(new_n13436));
  nand_4 g13060(.A(new_n12334), .B(new_n12303), .Y(new_n13437));
  nand_4 g13061(.A(new_n13437), .B(new_n13436), .Y(new_n13438));
  nor_4  g13062(.A(new_n12221_1), .B(new_n12220), .Y(new_n13439));
  and_4  g13063(.A(new_n12221_1), .B(new_n12220), .Y(new_n13440));
  or_4   g13064(.A(new_n13440), .B(new_n12218), .Y(new_n13441));
  not_3  g13065(.A(new_n13441), .Y(new_n13442));
  nor_4  g13066(.A(new_n13442), .B(new_n13439), .Y(new_n13443));
  nand_4 g13067(.A(n11877), .B(n3627), .Y(new_n13444));
  nand_4 g13068(.A(n8336), .B(n1198), .Y(new_n13445));
  nand_4 g13069(.A(n6770), .B(n5320), .Y(new_n13446));
  xor_3  g13070(.A(new_n13446), .B(new_n13445), .Y(new_n13447));
  xor_3  g13071(.A(new_n13447), .B(new_n13444), .Y(new_n13448));
  xnor_3 g13072(.A(new_n13448), .B(new_n13443), .Y(new_n13449));
  xnor_3 g13073(.A(new_n13449), .B(new_n13438), .Y(new_n13450));
  and_4  g13074(.A(new_n12492), .B(new_n12491), .Y(new_n13451));
  not_3  g13075(.A(new_n12494), .Y(new_n13452));
  nor_4  g13076(.A(new_n13452), .B(new_n12488), .Y(new_n13453));
  nor_4  g13077(.A(new_n13453), .B(new_n13451), .Y(new_n13454));
  nand_4 g13078(.A(new_n12495), .B(new_n12456), .Y(new_n13455));
  nand_4 g13079(.A(new_n12500), .B(new_n12496), .Y(new_n13456));
  nand_4 g13080(.A(new_n13456), .B(new_n13455), .Y(new_n13457));
  xnor_3 g13081(.A(new_n13457), .B(new_n13454), .Y(new_n13458));
  xnor_3 g13082(.A(new_n13458), .B(new_n13450), .Y(new_n13459));
  xnor_3 g13083(.A(new_n13459), .B(new_n13434), .Y(new_n13460));
  not_3  g13084(.A(new_n12501), .Y(new_n13461));
  nand_4 g13085(.A(new_n13461), .B(new_n12453), .Y(new_n13462));
  nand_4 g13086(.A(new_n12506), .B(new_n12502), .Y(new_n13463));
  nand_4 g13087(.A(new_n13463), .B(new_n13462), .Y(new_n13464));
  nand_4 g13088(.A(new_n12447), .B(new_n12371), .Y(new_n13465));
  not_3  g13089(.A(new_n12448), .Y(new_n13466));
  nand_4 g13090(.A(new_n12452), .B(new_n13466), .Y(new_n13467));
  nand_4 g13091(.A(new_n13467), .B(new_n13465), .Y(new_n13468));
  nor_4  g13092(.A(new_n12318), .B(new_n12317), .Y(new_n13469));
  not_3  g13093(.A(new_n12319), .Y(new_n13470));
  nor_4  g13094(.A(new_n12325), .B(new_n13470), .Y(new_n13471));
  nor_4  g13095(.A(new_n13471), .B(new_n13469), .Y(new_n13472));
  nand_4 g13096(.A(n5319), .B(n1478), .Y(new_n13473));
  not_3  g13097(.A(new_n13473), .Y(new_n13474));
  nand_4 g13098(.A(n11728), .B(n7320), .Y(new_n13475));
  nand_4 g13099(.A(n10990), .B(n4817), .Y(new_n13476));
  xor_3  g13100(.A(new_n13476), .B(new_n13475), .Y(new_n13477));
  xnor_3 g13101(.A(new_n13477), .B(new_n13474), .Y(new_n13478));
  not_3  g13102(.A(new_n12310), .Y(new_n13479));
  nor_4  g13103(.A(new_n12312), .B(new_n13479), .Y(new_n13480));
  nor_4  g13104(.A(new_n12313), .B(new_n12309), .Y(new_n13481));
  nor_4  g13105(.A(new_n13481), .B(new_n13480), .Y(new_n13482));
  xnor_3 g13106(.A(new_n13482), .B(new_n13478), .Y(new_n13483));
  nand_4 g13107(.A(n5212), .B(n4516), .Y(new_n13484));
  nand_4 g13108(.A(n12000), .B(n4189), .Y(new_n13485));
  nand_4 g13109(.A(n9725), .B(n2564), .Y(new_n13486));
  xor_3  g13110(.A(new_n13486), .B(new_n13485), .Y(new_n13487));
  xnor_3 g13111(.A(new_n13487), .B(new_n13484), .Y(new_n13488));
  nand_4 g13112(.A(n8819), .B(n1094), .Y(new_n13489));
  nand_4 g13113(.A(n8717), .B(n6986), .Y(new_n13490));
  xor_3  g13114(.A(new_n13490), .B(new_n13489), .Y(new_n13491));
  xnor_3 g13115(.A(new_n13491), .B(new_n13488), .Y(new_n13492));
  xnor_3 g13116(.A(new_n13492), .B(new_n13483), .Y(new_n13493));
  xnor_3 g13117(.A(new_n13493), .B(new_n13472), .Y(new_n13494));
  nand_4 g13118(.A(n2433), .B(n2226), .Y(new_n13495));
  nand_4 g13119(.A(n10678), .B(n6429), .Y(new_n13496));
  xor_3  g13120(.A(new_n13496), .B(new_n13495), .Y(new_n13497));
  not_3  g13121(.A(new_n12321), .Y(new_n13498));
  nor_4  g13122(.A(new_n12323), .B(new_n13498), .Y(new_n13499));
  not_3  g13123(.A(new_n12320), .Y(new_n13500));
  nor_4  g13124(.A(new_n12324), .B(new_n13500), .Y(new_n13501));
  nor_4  g13125(.A(new_n13501), .B(new_n13499), .Y(new_n13502));
  nand_4 g13126(.A(n10928), .B(n7730), .Y(new_n13503));
  xnor_3 g13127(.A(new_n13503), .B(new_n13502), .Y(new_n13504));
  xnor_3 g13128(.A(new_n13504), .B(new_n13497), .Y(new_n13505));
  nand_4 g13129(.A(new_n12227), .B(new_n12225), .Y(new_n13506));
  nand_4 g13130(.A(new_n12237), .B(new_n12228), .Y(new_n13507));
  nand_4 g13131(.A(new_n13507), .B(new_n13506), .Y(new_n13508));
  nand_4 g13132(.A(n9457), .B(n5760), .Y(new_n13509));
  nand_4 g13133(.A(n11222), .B(n10022), .Y(new_n13510));
  xor_3  g13134(.A(new_n13510), .B(new_n13509), .Y(new_n13511));
  xnor_3 g13135(.A(new_n13511), .B(new_n13508), .Y(new_n13512));
  xnor_3 g13136(.A(new_n13512), .B(new_n13505), .Y(new_n13513));
  not_3  g13137(.A(new_n12307), .Y(new_n13514));
  nor_4  g13138(.A(new_n12314), .B(new_n13514), .Y(new_n13515));
  not_3  g13139(.A(new_n12315), .Y(new_n13516));
  nor_4  g13140(.A(new_n12326), .B(new_n13516), .Y(new_n13517));
  nor_4  g13141(.A(new_n13517), .B(new_n13515), .Y(new_n13518));
  xnor_3 g13142(.A(new_n13518), .B(new_n13513), .Y(new_n13519));
  xnor_3 g13143(.A(new_n13519), .B(new_n13494), .Y(new_n13520));
  nand_4 g13144(.A(new_n12444_1), .B(new_n12443), .Y(new_n13521));
  not_3  g13145(.A(new_n12441), .Y(new_n13522));
  nand_4 g13146(.A(new_n12446), .B(new_n13522), .Y(new_n13523));
  nand_4 g13147(.A(new_n13523), .B(new_n13521), .Y(new_n13524));
  nand_4 g13148(.A(new_n12289), .B(new_n12330), .Y(new_n13525));
  not_3  g13149(.A(new_n12327), .Y(new_n13526));
  nand_4 g13150(.A(new_n12332), .B(new_n13526), .Y(new_n13527));
  nand_4 g13151(.A(new_n13527), .B(new_n13525), .Y(new_n13528));
  not_3  g13152(.A(new_n12217), .Y(new_n13529));
  nand_4 g13153(.A(new_n12223), .B(new_n13529), .Y(new_n13530));
  nand_4 g13154(.A(new_n12238), .B(new_n12224), .Y(new_n13531));
  nand_4 g13155(.A(new_n13531), .B(new_n13530), .Y(new_n13532));
  nand_4 g13156(.A(n9920), .B(n4370), .Y(new_n13533));
  not_3  g13157(.A(new_n12229), .Y(new_n13534));
  nand_4 g13158(.A(new_n12232), .B(new_n13534), .Y(new_n13535));
  nand_4 g13159(.A(new_n13535), .B(new_n12235), .Y(new_n13536));
  xor_3  g13160(.A(new_n13536), .B(new_n13533), .Y(new_n13537));
  xnor_3 g13161(.A(new_n13537), .B(new_n13532), .Y(new_n13538));
  xnor_3 g13162(.A(new_n13538), .B(new_n13528), .Y(new_n13539));
  xnor_3 g13163(.A(new_n13539), .B(new_n13524), .Y(new_n13540));
  xnor_3 g13164(.A(new_n13540), .B(new_n13520), .Y(new_n13541));
  xnor_3 g13165(.A(new_n13541), .B(new_n13468), .Y(new_n13542));
  xnor_3 g13166(.A(new_n13542), .B(new_n13464), .Y(new_n13543));
  xnor_3 g13167(.A(new_n13543), .B(new_n13460), .Y(new_n13544));
  xnor_3 g13168(.A(new_n13544), .B(new_n13357), .Y(new_n13545));
  xnor_3 g13169(.A(new_n13545), .B(new_n13351), .Y(n8100));
  not_3  g13170(.A(new_n10018), .Y(new_n13547));
  xor_3  g13171(.A(new_n10019), .B(new_n13547), .Y(n8138));
  not_3  g13172(.A(new_n6278), .Y(new_n13549));
  xor_3  g13173(.A(new_n6280), .B(new_n13549), .Y(n8202));
  xor_3  g13174(.A(new_n3825), .B(new_n3812), .Y(n8303));
  not_3  g13175(.A(new_n3079), .Y(new_n13552));
  xor_3  g13176(.A(new_n3080), .B(new_n13552), .Y(n8398));
  not_3  g13177(.A(new_n4460), .Y(new_n13554));
  xor_3  g13178(.A(new_n4461), .B(new_n13554), .Y(n9137));
  not_3  g13179(.A(new_n7375), .Y(new_n13556));
  xor_3  g13180(.A(new_n13556), .B(new_n7374), .Y(n9387));
  not_3  g13181(.A(new_n11969), .Y(new_n13558));
  xor_3  g13182(.A(new_n13558), .B(new_n11968), .Y(n9571));
  nor_4  g13183(.A(new_n1018), .B(new_n1015), .Y(new_n13560));
  xor_3  g13184(.A(new_n13560), .B(new_n1062), .Y(n9578));
  xor_3  g13185(.A(new_n1212), .B(new_n1209_1), .Y(n9706));
  not_3  g13186(.A(new_n4450), .Y(new_n13563));
  xor_3  g13187(.A(new_n4463), .B(new_n13563), .Y(n9756));
  nand_4 g13188(.A(new_n7039), .B(new_n7015), .Y(new_n13565));
  nand_4 g13189(.A(new_n13565), .B(new_n7018), .Y(new_n13566));
  not_3  g13190(.A(new_n6988), .Y(new_n13567));
  nand_4 g13191(.A(new_n13567), .B(new_n6768), .Y(new_n13568));
  nand_4 g13192(.A(new_n7013), .B(new_n6989), .Y(new_n13569));
  nand_4 g13193(.A(new_n13569), .B(new_n13568), .Y(new_n13570));
  not_3  g13194(.A(new_n6614), .Y(new_n13571));
  nand_4 g13195(.A(new_n6648), .B(new_n13571), .Y(new_n13572));
  nand_4 g13196(.A(new_n6665), .B(new_n6649), .Y(new_n13573));
  nand_4 g13197(.A(new_n13573), .B(new_n13572), .Y(new_n13574));
  nor_4  g13198(.A(new_n6830), .B(new_n6829), .Y(new_n13575));
  not_3  g13199(.A(new_n6831), .Y(new_n13576));
  nor_4  g13200(.A(new_n6837), .B(new_n13576), .Y(new_n13577));
  nor_4  g13201(.A(new_n13577), .B(new_n13575), .Y(new_n13578));
  xnor_3 g13202(.A(new_n13578), .B(new_n13574), .Y(new_n13579));
  not_3  g13203(.A(new_n6947), .Y(new_n13580));
  nand_4 g13204(.A(new_n13580), .B(new_n6912), .Y(new_n13581));
  nand_4 g13205(.A(new_n6962), .B(new_n6948), .Y(new_n13582));
  nand_4 g13206(.A(new_n13582), .B(new_n13581), .Y(new_n13583));
  nor_4  g13207(.A(new_n6733), .B(new_n6732), .Y(new_n13584));
  nor_4  g13208(.A(new_n6741), .B(new_n6735), .Y(new_n13585));
  nor_4  g13209(.A(new_n13585), .B(new_n13584), .Y(new_n13586));
  not_3  g13210(.A(new_n6737), .Y(new_n13587));
  nor_4  g13211(.A(new_n6739), .B(new_n13587), .Y(new_n13588));
  not_3  g13212(.A(new_n6736), .Y(new_n13589));
  nor_4  g13213(.A(new_n6740), .B(new_n13589), .Y(new_n13590));
  nor_4  g13214(.A(new_n13590), .B(new_n13588), .Y(new_n13591));
  nand_4 g13215(.A(n10451), .B(n2226), .Y(new_n13592));
  xnor_3 g13216(.A(new_n13592), .B(new_n13591), .Y(new_n13593));
  xnor_3 g13217(.A(new_n13593), .B(new_n13586), .Y(new_n13594));
  nand_4 g13218(.A(n10278), .B(n6986), .Y(new_n13595));
  nand_4 g13219(.A(n11423), .B(n10928), .Y(new_n13596));
  xor_3  g13220(.A(new_n13596), .B(new_n13595), .Y(new_n13597));
  not_3  g13221(.A(new_n6725), .Y(new_n13598));
  nor_4  g13222(.A(new_n6727), .B(new_n13598), .Y(new_n13599));
  not_3  g13223(.A(new_n6724), .Y(new_n13600));
  nor_4  g13224(.A(new_n6728), .B(new_n13600), .Y(new_n13601));
  nor_4  g13225(.A(new_n13601), .B(new_n13599), .Y(new_n13602));
  nand_4 g13226(.A(n10678), .B(n3022), .Y(new_n13603));
  xnor_3 g13227(.A(new_n13603), .B(new_n13602), .Y(new_n13604));
  xnor_3 g13228(.A(new_n13604), .B(new_n13597), .Y(new_n13605));
  xnor_3 g13229(.A(new_n13605), .B(new_n13594), .Y(new_n13606));
  nand_4 g13230(.A(n10327), .B(n4189), .Y(new_n13607));
  nand_4 g13231(.A(new_n6629), .B(new_n6627), .Y(new_n13608));
  nand_4 g13232(.A(new_n6639), .B(new_n6630), .Y(new_n13609));
  nand_4 g13233(.A(new_n13609), .B(new_n13608), .Y(new_n13610));
  nand_4 g13234(.A(n9583), .B(n2564), .Y(new_n13611));
  not_3  g13235(.A(new_n13611), .Y(new_n13612));
  xnor_3 g13236(.A(new_n13612), .B(new_n13610), .Y(new_n13613));
  xnor_3 g13237(.A(new_n13613), .B(new_n13607), .Y(new_n13614));
  xnor_3 g13238(.A(new_n13614), .B(new_n13606), .Y(new_n13615));
  nand_4 g13239(.A(new_n6729), .B(new_n6722), .Y(new_n13616));
  nand_4 g13240(.A(new_n6742_1), .B(new_n6730), .Y(new_n13617));
  nand_4 g13241(.A(new_n13617), .B(new_n13616), .Y(new_n13618));
  nand_4 g13242(.A(n11023), .B(n1094), .Y(new_n13619));
  nand_4 g13243(.A(n9920), .B(n7456), .Y(new_n13620));
  not_3  g13244(.A(new_n6631), .Y(new_n13621));
  nand_4 g13245(.A(new_n6634), .B(new_n13621), .Y(new_n13622));
  nand_4 g13246(.A(new_n13622), .B(new_n6637), .Y(new_n13623));
  xor_3  g13247(.A(new_n13623), .B(new_n13620), .Y(new_n13624));
  xor_3  g13248(.A(new_n13624), .B(new_n13619), .Y(new_n13625));
  xnor_3 g13249(.A(new_n13625), .B(new_n13618), .Y(new_n13626));
  xnor_3 g13250(.A(new_n13626), .B(new_n13615), .Y(new_n13627));
  xnor_3 g13251(.A(new_n13627), .B(new_n13583), .Y(new_n13628));
  xnor_3 g13252(.A(new_n13628), .B(new_n13579), .Y(new_n13629));
  not_3  g13253(.A(new_n6719), .Y(new_n13630));
  nand_4 g13254(.A(new_n6752), .B(new_n13630), .Y(new_n13631));
  nand_4 g13255(.A(new_n6766), .B(new_n6753), .Y(new_n13632));
  nand_4 g13256(.A(new_n13632), .B(new_n13631), .Y(new_n13633));
  nand_4 g13257(.A(n11662), .B(n6770), .Y(new_n13634));
  nand_4 g13258(.A(new_n6645_1), .B(new_n6644), .Y(new_n13635));
  not_3  g13259(.A(new_n6642), .Y(new_n13636));
  nand_4 g13260(.A(new_n6647), .B(new_n13636), .Y(new_n13637));
  nand_4 g13261(.A(new_n13637), .B(new_n13635), .Y(new_n13638));
  xnor_3 g13262(.A(new_n13638), .B(new_n13634), .Y(new_n13639));
  nand_4 g13263(.A(new_n6625), .B(new_n6618), .Y(new_n13640));
  nand_4 g13264(.A(new_n6640), .B(new_n6626), .Y(new_n13641));
  nand_4 g13265(.A(new_n13641), .B(new_n13640), .Y(new_n13642));
  not_3  g13266(.A(new_n6621), .Y(new_n13643));
  nor_4  g13267(.A(new_n6623), .B(new_n13643), .Y(new_n13644));
  not_3  g13268(.A(new_n6620), .Y(new_n13645));
  nor_4  g13269(.A(new_n6624), .B(new_n13645), .Y(new_n13646));
  nor_4  g13270(.A(new_n13646), .B(new_n13644), .Y(new_n13647));
  nand_4 g13271(.A(n9640), .B(n7320), .Y(new_n13648));
  not_3  g13272(.A(new_n13648), .Y(new_n13649));
  nand_4 g13273(.A(n8336), .B(n2278), .Y(new_n13650));
  nand_4 g13274(.A(n7523), .B(n6703), .Y(new_n13651));
  xor_3  g13275(.A(new_n13651), .B(new_n13650), .Y(new_n13652));
  nand_4 g13276(.A(n12591), .B(n3627), .Y(new_n13653));
  nand_4 g13277(.A(n4516), .B(n3932), .Y(new_n13654));
  xor_3  g13278(.A(new_n13654), .B(new_n13653), .Y(new_n13655));
  xnor_3 g13279(.A(new_n13655), .B(new_n13652), .Y(new_n13656));
  xnor_3 g13280(.A(new_n13656), .B(new_n13649), .Y(new_n13657));
  xnor_3 g13281(.A(new_n13657), .B(new_n13647), .Y(new_n13658));
  xnor_3 g13282(.A(new_n13658), .B(new_n13642), .Y(new_n13659));
  nand_4 g13283(.A(n12247), .B(n11153), .Y(new_n13660));
  not_3  g13284(.A(new_n13660), .Y(new_n13661));
  nor_4  g13285(.A(new_n6835), .B(new_n6834), .Y(new_n13662));
  nand_4 g13286(.A(new_n6835), .B(new_n6834), .Y(new_n13663));
  nand_4 g13287(.A(new_n13663), .B(new_n6833), .Y(new_n13664));
  not_3  g13288(.A(new_n13664), .Y(new_n13665));
  nor_4  g13289(.A(new_n13665), .B(new_n13662), .Y(new_n13666));
  nand_4 g13290(.A(n6687), .B(n753), .Y(new_n13667));
  nand_4 g13291(.A(n2087), .B(n1798), .Y(new_n13668));
  xor_3  g13292(.A(new_n13668), .B(new_n13667), .Y(new_n13669));
  nand_4 g13293(.A(n12826), .B(n7891), .Y(new_n13670));
  nand_4 g13294(.A(n12391), .B(n4094), .Y(new_n13671));
  xor_3  g13295(.A(new_n13671), .B(new_n13670), .Y(new_n13672));
  xnor_3 g13296(.A(new_n13672), .B(new_n13669), .Y(new_n13673));
  xnor_3 g13297(.A(new_n13673), .B(new_n13666), .Y(new_n13674));
  xnor_3 g13298(.A(new_n13674), .B(new_n13661), .Y(new_n13675));
  xnor_3 g13299(.A(new_n13675), .B(new_n13659), .Y(new_n13676));
  nand_4 g13300(.A(new_n6749), .B(new_n6747), .Y(new_n13677));
  nand_4 g13301(.A(new_n6751), .B(new_n6743), .Y(new_n13678));
  nand_4 g13302(.A(new_n13678), .B(new_n13677), .Y(new_n13679));
  nand_4 g13303(.A(new_n6929), .B(new_n6922), .Y(new_n13680));
  nand_4 g13304(.A(new_n6944), .B(new_n6931), .Y(new_n13681));
  nand_4 g13305(.A(new_n13681), .B(new_n13680), .Y(new_n13682));
  xnor_3 g13306(.A(new_n13682), .B(new_n13679), .Y(new_n13683));
  xnor_3 g13307(.A(new_n13683), .B(new_n13676), .Y(new_n13684));
  xnor_3 g13308(.A(new_n13684), .B(new_n13639), .Y(new_n13685));
  xnor_3 g13309(.A(new_n13685), .B(new_n13633), .Y(new_n13686));
  xnor_3 g13310(.A(new_n13686), .B(new_n13629), .Y(new_n13687));
  nand_4 g13311(.A(new_n6986_1), .B(new_n6963), .Y(new_n13688));
  nor_4  g13312(.A(new_n6984), .B(new_n6966), .Y(new_n13689));
  xnor_3 g13313(.A(new_n13689), .B(new_n6963), .Y(new_n13690));
  nand_4 g13314(.A(new_n13690), .B(new_n6863), .Y(new_n13691));
  nand_4 g13315(.A(new_n13691), .B(new_n13688), .Y(new_n13692));
  nand_4 g13316(.A(new_n6847), .B(new_n6815), .Y(new_n13693));
  nand_4 g13317(.A(new_n6862), .B(new_n6848), .Y(new_n13694));
  nand_4 g13318(.A(new_n13694), .B(new_n13693), .Y(new_n13695));
  nand_4 g13319(.A(new_n6934), .B(new_n6932), .Y(new_n13696));
  nand_4 g13320(.A(new_n6943), .B(new_n6935), .Y(new_n13697));
  nand_4 g13321(.A(new_n13697), .B(new_n13696), .Y(new_n13698));
  not_3  g13322(.A(new_n6822_1), .Y(new_n13699));
  nor_4  g13323(.A(new_n6824), .B(new_n13699), .Y(new_n13700));
  not_3  g13324(.A(new_n6821), .Y(new_n13701));
  nor_4  g13325(.A(new_n6825), .B(new_n13701), .Y(new_n13702));
  nor_4  g13326(.A(new_n13702), .B(new_n13700), .Y(new_n13703));
  xnor_3 g13327(.A(new_n13703), .B(new_n13698), .Y(new_n13704));
  nand_4 g13328(.A(n10898), .B(n9457), .Y(new_n13705));
  nand_4 g13329(.A(n12511), .B(n11222), .Y(new_n13706));
  not_3  g13330(.A(new_n13706), .Y(new_n13707));
  xor_3  g13331(.A(new_n13707), .B(new_n13705), .Y(new_n13708));
  nand_4 g13332(.A(n11876), .B(n4817), .Y(new_n13709));
  nand_4 g13333(.A(n5319), .B(n3754), .Y(new_n13710));
  xor_3  g13334(.A(new_n13710), .B(new_n13709), .Y(new_n13711));
  xor_3  g13335(.A(new_n13711), .B(new_n13708), .Y(new_n13712));
  xnor_3 g13336(.A(new_n13712), .B(new_n13704), .Y(new_n13713));
  nand_4 g13337(.A(n12069), .B(n10685), .Y(new_n13714));
  not_3  g13338(.A(new_n13714), .Y(new_n13715));
  not_3  g13339(.A(new_n6925), .Y(new_n13716));
  nor_4  g13340(.A(new_n6927), .B(new_n13716), .Y(new_n13717));
  nor_4  g13341(.A(new_n6928), .B(new_n6924), .Y(new_n13718));
  nor_4  g13342(.A(new_n13718), .B(new_n13717), .Y(new_n13719));
  nand_4 g13343(.A(n6578), .B(n5645), .Y(new_n13720));
  not_3  g13344(.A(new_n13720), .Y(new_n13721));
  xnor_3 g13345(.A(new_n13721), .B(new_n13719), .Y(new_n13722));
  nand_4 g13346(.A(n11922), .B(n4828), .Y(new_n13723));
  nand_4 g13347(.A(n8665), .B(n2515), .Y(new_n13724));
  not_3  g13348(.A(new_n13724), .Y(new_n13725));
  xor_3  g13349(.A(new_n13725), .B(new_n13723), .Y(new_n13726));
  xnor_3 g13350(.A(new_n13726), .B(new_n13722), .Y(new_n13727));
  xnor_3 g13351(.A(new_n13727), .B(new_n13715), .Y(new_n13728));
  xnor_3 g13352(.A(new_n13728), .B(new_n13713), .Y(new_n13729));
  nand_4 g13353(.A(new_n6826_1), .B(new_n6819), .Y(new_n13730));
  not_3  g13354(.A(new_n6838), .Y(new_n13731));
  nand_4 g13355(.A(new_n13731), .B(new_n6827), .Y(new_n13732));
  nand_4 g13356(.A(new_n13732), .B(new_n13730), .Y(new_n13733));
  nand_4 g13357(.A(n996), .B(n159), .Y(new_n13734));
  nand_4 g13358(.A(n5767), .B(n2749), .Y(new_n13735));
  xor_3  g13359(.A(new_n13735), .B(new_n13734), .Y(new_n13736));
  nand_4 g13360(.A(n1199), .B(n1067), .Y(new_n13737));
  nand_4 g13361(.A(n5314), .B(n1510), .Y(new_n13738));
  xor_3  g13362(.A(new_n13738), .B(new_n13737), .Y(new_n13739));
  xor_3  g13363(.A(new_n13739), .B(new_n13736), .Y(new_n13740));
  nand_4 g13364(.A(n7160), .B(n2551), .Y(new_n13741));
  not_3  g13365(.A(new_n6939), .Y(new_n13742));
  nor_4  g13366(.A(new_n6941), .B(new_n13742), .Y(new_n13743));
  nor_4  g13367(.A(new_n6942), .B(new_n6938), .Y(new_n13744));
  nor_4  g13368(.A(new_n13744), .B(new_n13743), .Y(new_n13745));
  xnor_3 g13369(.A(new_n13745), .B(new_n13741), .Y(new_n13746));
  xnor_3 g13370(.A(new_n13746), .B(new_n13740), .Y(new_n13747));
  xnor_3 g13371(.A(new_n13747), .B(new_n13733), .Y(new_n13748));
  xnor_3 g13372(.A(new_n13748), .B(new_n13729), .Y(new_n13749));
  nand_4 g13373(.A(new_n6917), .B(new_n6916), .Y(new_n13750));
  nand_4 g13374(.A(new_n6946), .B(new_n6919), .Y(new_n13751));
  nand_4 g13375(.A(new_n13751), .B(new_n13750), .Y(new_n13752));
  nand_4 g13376(.A(new_n6844), .B(new_n6843), .Y(new_n13753));
  not_3  g13377(.A(new_n6839), .Y(new_n13754));
  nand_4 g13378(.A(new_n6846), .B(new_n13754), .Y(new_n13755));
  nand_4 g13379(.A(new_n13755), .B(new_n13753), .Y(new_n13756));
  xnor_3 g13380(.A(new_n13756), .B(new_n13752), .Y(new_n13757));
  xnor_3 g13381(.A(new_n13757), .B(new_n13749), .Y(new_n13758));
  xnor_3 g13382(.A(new_n13758), .B(new_n13695), .Y(new_n13759));
  xnor_3 g13383(.A(new_n13759), .B(new_n13692), .Y(new_n13760));
  xnor_3 g13384(.A(new_n13760), .B(new_n13687), .Y(new_n13761));
  xnor_3 g13385(.A(new_n13761), .B(new_n13570), .Y(new_n13762));
  xnor_3 g13386(.A(new_n13762), .B(new_n13566), .Y(n9767));
  not_3  g13387(.A(new_n2180), .Y(new_n13764));
  xor_3  g13388(.A(new_n2182), .B(new_n13764), .Y(n9820));
  nand_4 g13389(.A(new_n9990), .B(new_n9989), .Y(new_n13766));
  xnor_3 g13390(.A(new_n13766), .B(new_n10033), .Y(n9938));
  xor_3  g13391(.A(new_n1058), .B(new_n1055), .Y(n10476));
  xor_3  g13392(.A(new_n1052), .B(new_n1041), .Y(n10589));
  not_3  g13393(.A(new_n1205), .Y(new_n13770));
  xor_3  g13394(.A(new_n1207), .B(new_n13770), .Y(n10695));
  not_3  g13395(.A(new_n3842_1), .Y(new_n13772));
  nor_4  g13396(.A(new_n3794), .B(new_n3793), .Y(new_n13773));
  xnor_3 g13397(.A(new_n13773), .B(new_n13772), .Y(n10789));
  xor_3  g13398(.A(new_n3074), .B(new_n3064), .Y(n10851));
  not_3  g13399(.A(new_n5260), .Y(new_n13776));
  xor_3  g13400(.A(new_n5269), .B(new_n13776), .Y(n10913));
  xnor_3 g13401(.A(new_n7512), .B(new_n7379), .Y(n10949));
  xnor_3 g13402(.A(new_n11971), .B(new_n11916), .Y(n11216));
  xor_3  g13403(.A(new_n5261), .B(new_n5251), .Y(n11326));
  not_3  g13404(.A(new_n5571), .Y(new_n13781));
  not_3  g13405(.A(new_n5806), .Y(new_n13782));
  nor_4  g13406(.A(new_n13782), .B(new_n13781), .Y(new_n13783));
  nor_4  g13407(.A(new_n5806), .B(new_n5571), .Y(new_n13784));
  nor_4  g13408(.A(new_n5942), .B(new_n13784), .Y(new_n13785));
  nor_4  g13409(.A(new_n13785), .B(new_n13783), .Y(new_n13786));
  nand_4 g13410(.A(new_n5883), .B(new_n5853), .Y(new_n13787));
  not_3  g13411(.A(new_n5884), .Y(new_n13788));
  nand_4 g13412(.A(new_n5887), .B(new_n13788), .Y(new_n13789));
  nand_4 g13413(.A(new_n13789), .B(new_n13787), .Y(new_n13790));
  nand_4 g13414(.A(n9763), .B(n45), .Y(new_n13791));
  nand_4 g13415(.A(new_n5553), .B(new_n5552), .Y(new_n13792));
  not_3  g13416(.A(new_n5550), .Y(new_n13793));
  nand_4 g13417(.A(new_n5555), .B(new_n13793), .Y(new_n13794));
  nand_4 g13418(.A(new_n13794), .B(new_n13792), .Y(new_n13795));
  xnor_3 g13419(.A(new_n13795), .B(new_n13791), .Y(new_n13796));
  xnor_3 g13420(.A(new_n13796), .B(new_n13790), .Y(new_n13797));
  not_3  g13421(.A(new_n5528), .Y(new_n13798));
  nand_4 g13422(.A(new_n5556), .B(new_n13798), .Y(new_n13799));
  nand_4 g13423(.A(new_n5570), .B(new_n5557), .Y(new_n13800));
  nand_4 g13424(.A(new_n13800), .B(new_n13799), .Y(new_n13801));
  nand_4 g13425(.A(new_n5843), .B(new_n5811), .Y(new_n13802));
  nand_4 g13426(.A(new_n5844), .B(new_n5810), .Y(new_n13803));
  nand_4 g13427(.A(new_n13803), .B(new_n13802), .Y(new_n13804));
  xnor_3 g13428(.A(new_n13804), .B(new_n13801), .Y(new_n13805));
  xnor_3 g13429(.A(new_n13805), .B(new_n13797), .Y(new_n13806));
  nand_4 g13430(.A(new_n5924), .B(new_n5892), .Y(new_n13807));
  nand_4 g13431(.A(new_n5926), .B(new_n5925), .Y(new_n13808));
  nand_4 g13432(.A(new_n13808), .B(new_n13807), .Y(new_n13809));
  nor_4  g13433(.A(new_n5541), .B(new_n5540), .Y(new_n13810));
  not_3  g13434(.A(new_n5542), .Y(new_n13811));
  nor_4  g13435(.A(new_n5548), .B(new_n13811), .Y(new_n13812));
  nor_4  g13436(.A(new_n13812), .B(new_n13810), .Y(new_n13813));
  xnor_3 g13437(.A(new_n13813), .B(new_n13809), .Y(new_n13814));
  not_3  g13438(.A(new_n5814_1), .Y(new_n13815));
  nand_4 g13439(.A(new_n5820), .B(new_n13815), .Y(new_n13816));
  nand_4 g13440(.A(new_n5835), .B(new_n5821), .Y(new_n13817));
  nand_4 g13441(.A(new_n13817), .B(new_n13816), .Y(new_n13818));
  nand_4 g13442(.A(n2253), .B(n1097), .Y(new_n13819));
  not_3  g13443(.A(new_n5816), .Y(new_n13820));
  nor_4  g13444(.A(new_n5818), .B(new_n13820), .Y(new_n13821));
  not_3  g13445(.A(new_n5815), .Y(new_n13822));
  nor_4  g13446(.A(new_n5819), .B(new_n13822), .Y(new_n13823));
  nor_4  g13447(.A(new_n13823), .B(new_n13821), .Y(new_n13824));
  xnor_3 g13448(.A(new_n13824), .B(new_n13819), .Y(new_n13825));
  not_3  g13449(.A(new_n5826), .Y(new_n13826));
  nand_4 g13450(.A(new_n5829), .B(new_n13826), .Y(new_n13827));
  and_4  g13451(.A(new_n13827), .B(new_n5832), .Y(new_n13828));
  nand_4 g13452(.A(n12299), .B(n12221), .Y(new_n13829));
  nand_4 g13453(.A(n9241), .B(n9189), .Y(new_n13830));
  xor_3  g13454(.A(new_n13830), .B(new_n13829), .Y(new_n13831));
  xnor_3 g13455(.A(new_n13831), .B(new_n13828), .Y(new_n13832));
  xnor_3 g13456(.A(new_n13832), .B(new_n13825), .Y(new_n13833));
  nand_4 g13457(.A(n12145), .B(n7436), .Y(new_n13834));
  not_3  g13458(.A(new_n13834), .Y(new_n13835));
  nand_4 g13459(.A(n10217), .B(n6776), .Y(new_n13836));
  nand_4 g13460(.A(n8276), .B(n2522), .Y(new_n13837));
  xor_3  g13461(.A(new_n13837), .B(new_n13836), .Y(new_n13838));
  xnor_3 g13462(.A(new_n13838), .B(new_n13835), .Y(new_n13839));
  nand_4 g13463(.A(new_n5824), .B(new_n5822), .Y(new_n13840));
  nand_4 g13464(.A(new_n5834), .B(new_n5825), .Y(new_n13841));
  nand_4 g13465(.A(new_n13841), .B(new_n13840), .Y(new_n13842));
  xnor_3 g13466(.A(new_n13842), .B(new_n13839), .Y(new_n13843));
  xnor_3 g13467(.A(new_n13843), .B(new_n13833), .Y(new_n13844));
  xnor_3 g13468(.A(new_n13844), .B(new_n13818), .Y(new_n13845));
  nand_4 g13469(.A(new_n5921), .B(new_n5919), .Y(new_n13846));
  nand_4 g13470(.A(new_n5923), .B(new_n5915), .Y(new_n13847));
  nand_4 g13471(.A(new_n13847), .B(new_n13846), .Y(new_n13848));
  not_3  g13472(.A(new_n5544), .Y(new_n13849));
  nor_4  g13473(.A(new_n5546), .B(new_n13849), .Y(new_n13850));
  not_3  g13474(.A(new_n5543), .Y(new_n13851));
  nor_4  g13475(.A(new_n5547), .B(new_n13851), .Y(new_n13852));
  nor_4  g13476(.A(new_n13852), .B(new_n13850), .Y(new_n13853));
  nand_4 g13477(.A(n5964), .B(n3865), .Y(new_n13854));
  nand_4 g13478(.A(n12705), .B(n4634), .Y(new_n13855));
  xor_3  g13479(.A(new_n13855), .B(new_n13854), .Y(new_n13856));
  xor_3  g13480(.A(new_n13856), .B(new_n13853), .Y(new_n13857));
  xnor_3 g13481(.A(new_n13857), .B(new_n13848), .Y(new_n13858));
  xnor_3 g13482(.A(new_n13858), .B(new_n13845), .Y(new_n13859));
  not_3  g13483(.A(new_n5896), .Y(new_n13860));
  nand_4 g13484(.A(new_n5901), .B(new_n13860), .Y(new_n13861));
  nand_4 g13485(.A(new_n5913), .B(new_n5902), .Y(new_n13862));
  nand_4 g13486(.A(new_n13862), .B(new_n13861), .Y(new_n13863));
  not_3  g13487(.A(new_n5904), .Y(new_n13864));
  nand_4 g13488(.A(new_n13864), .B(new_n5903), .Y(new_n13865));
  nand_4 g13489(.A(new_n5911), .B(new_n5905), .Y(new_n13866));
  nand_4 g13490(.A(new_n13866), .B(new_n13865), .Y(new_n13867));
  nand_4 g13491(.A(n3616), .B(n2498), .Y(new_n13868));
  not_3  g13492(.A(new_n13868), .Y(new_n13869));
  nand_4 g13493(.A(n10545), .B(n521), .Y(new_n13870));
  nand_4 g13494(.A(n7690), .B(n5579), .Y(new_n13871));
  xnor_3 g13495(.A(new_n13871), .B(new_n13870), .Y(new_n13872));
  xnor_3 g13496(.A(new_n13872), .B(new_n13869), .Y(new_n13873));
  xnor_3 g13497(.A(new_n13873), .B(new_n13867), .Y(new_n13874));
  and_4  g13498(.A(new_n5899), .B(new_n5898), .Y(new_n13875));
  not_3  g13499(.A(new_n5897), .Y(new_n13876));
  nor_4  g13500(.A(new_n5900), .B(new_n13876), .Y(new_n13877));
  nor_4  g13501(.A(new_n13877), .B(new_n13875), .Y(new_n13878));
  nand_4 g13502(.A(n5860), .B(n806), .Y(new_n13879));
  nand_4 g13503(.A(n4499), .B(n2558), .Y(new_n13880));
  nand_4 g13504(.A(n7270), .B(n2393), .Y(new_n13881));
  xnor_3 g13505(.A(new_n13881), .B(new_n13880), .Y(new_n13882));
  nand_4 g13506(.A(n5331), .B(n1576), .Y(new_n13883));
  nand_4 g13507(.A(n7388), .B(n2507), .Y(new_n13884));
  xnor_3 g13508(.A(new_n13884), .B(new_n13883), .Y(new_n13885));
  xnor_3 g13509(.A(new_n13885), .B(new_n13882), .Y(new_n13886));
  xnor_3 g13510(.A(new_n13886), .B(new_n13879), .Y(new_n13887));
  xnor_3 g13511(.A(new_n13887), .B(new_n13878), .Y(new_n13888));
  xnor_3 g13512(.A(new_n13888), .B(new_n13874), .Y(new_n13889));
  xnor_3 g13513(.A(new_n13889), .B(new_n13863), .Y(new_n13890));
  not_3  g13514(.A(new_n5856), .Y(new_n13891));
  nand_4 g13515(.A(new_n5861), .B(new_n13891), .Y(new_n13892));
  nand_4 g13516(.A(new_n5873), .B(new_n5862), .Y(new_n13893));
  nand_4 g13517(.A(new_n13893), .B(new_n13892), .Y(new_n13894));
  not_3  g13518(.A(new_n5864), .Y(new_n13895));
  nand_4 g13519(.A(new_n13895), .B(new_n5863), .Y(new_n13896));
  nand_4 g13520(.A(new_n5871), .B(new_n5865), .Y(new_n13897));
  nand_4 g13521(.A(new_n13897), .B(new_n13896), .Y(new_n13898));
  and_4  g13522(.A(new_n5869), .B(new_n5868), .Y(new_n13899));
  nor_4  g13523(.A(new_n5870), .B(new_n5867), .Y(new_n13900));
  nor_4  g13524(.A(new_n13900), .B(new_n13899), .Y(new_n13901));
  xnor_3 g13525(.A(new_n13901), .B(new_n13898), .Y(new_n13902));
  nand_4 g13526(.A(n5305), .B(n2512), .Y(new_n13903));
  nand_4 g13527(.A(n12648), .B(n6016), .Y(new_n13904));
  nand_4 g13528(.A(n11892), .B(n5153), .Y(new_n13905));
  xnor_3 g13529(.A(new_n13905), .B(new_n13904), .Y(new_n13906));
  xnor_3 g13530(.A(new_n13906), .B(new_n13903), .Y(new_n13907));
  nor_4  g13531(.A(new_n5859), .B(new_n5858), .Y(new_n13908));
  not_3  g13532(.A(new_n5857_1), .Y(new_n13909));
  nand_4 g13533(.A(new_n5859), .B(new_n5858), .Y(new_n13910));
  nand_4 g13534(.A(new_n13910), .B(new_n13909), .Y(new_n13911));
  not_3  g13535(.A(new_n13911), .Y(new_n13912));
  nor_4  g13536(.A(new_n13912), .B(new_n13908), .Y(new_n13913));
  nand_4 g13537(.A(n5798), .B(n2530), .Y(new_n13914));
  nand_4 g13538(.A(n10547), .B(n7265), .Y(new_n13915));
  nand_4 g13539(.A(n8476), .B(n2347), .Y(new_n13916));
  xnor_3 g13540(.A(new_n13916), .B(new_n13915), .Y(new_n13917));
  xnor_3 g13541(.A(new_n13917), .B(new_n13914), .Y(new_n13918));
  xnor_3 g13542(.A(new_n13918), .B(new_n13913), .Y(new_n13919));
  xnor_3 g13543(.A(new_n13919), .B(new_n13907), .Y(new_n13920));
  xnor_3 g13544(.A(new_n13920), .B(new_n13902), .Y(new_n13921));
  xnor_3 g13545(.A(new_n13921), .B(new_n13894), .Y(new_n13922));
  xnor_3 g13546(.A(new_n13922), .B(new_n13890), .Y(new_n13923));
  nand_4 g13547(.A(n3986), .B(n3342), .Y(new_n13924));
  nand_4 g13548(.A(n11257), .B(n2879), .Y(new_n13925));
  nand_4 g13549(.A(n8759), .B(n7823), .Y(new_n13926));
  xor_3  g13550(.A(new_n13926), .B(new_n13925), .Y(new_n13927));
  xor_3  g13551(.A(new_n13927), .B(new_n13924), .Y(new_n13928));
  xnor_3 g13552(.A(new_n13928), .B(new_n13923), .Y(new_n13929));
  and_4  g13553(.A(new_n5909), .B(new_n5908), .Y(new_n13930));
  nor_4  g13554(.A(new_n5910), .B(new_n5907), .Y(new_n13931));
  nor_4  g13555(.A(new_n13931), .B(new_n13930), .Y(new_n13932));
  nand_4 g13556(.A(new_n5880), .B(new_n5878), .Y(new_n13933));
  nand_4 g13557(.A(new_n5882), .B(new_n5874), .Y(new_n13934));
  nand_4 g13558(.A(new_n13934), .B(new_n13933), .Y(new_n13935));
  xnor_3 g13559(.A(new_n13935), .B(new_n13932), .Y(new_n13936));
  xnor_3 g13560(.A(new_n13936), .B(new_n13929), .Y(new_n13937));
  nand_4 g13561(.A(new_n5839), .B(new_n5838), .Y(new_n13938));
  nand_4 g13562(.A(new_n5841), .B(new_n5836), .Y(new_n13939));
  nand_4 g13563(.A(new_n13939), .B(new_n13938), .Y(new_n13940));
  not_3  g13564(.A(new_n5531), .Y(new_n13941));
  nand_4 g13565(.A(new_n5537), .B(new_n13941), .Y(new_n13942));
  not_3  g13566(.A(new_n5549), .Y(new_n13943));
  nand_4 g13567(.A(new_n13943), .B(new_n5538), .Y(new_n13944));
  nand_4 g13568(.A(new_n13944), .B(new_n13942), .Y(new_n13945));
  not_3  g13569(.A(new_n5533), .Y(new_n13946));
  nor_4  g13570(.A(new_n5535), .B(new_n13946), .Y(new_n13947));
  not_3  g13571(.A(new_n5532), .Y(new_n13948));
  nor_4  g13572(.A(new_n5536), .B(new_n13948), .Y(new_n13949));
  nor_4  g13573(.A(new_n13949), .B(new_n13947), .Y(new_n13950));
  nand_4 g13574(.A(n9195), .B(n4312), .Y(new_n13951));
  nand_4 g13575(.A(n12025), .B(n10223), .Y(new_n13952));
  xor_3  g13576(.A(new_n13952), .B(new_n13951), .Y(new_n13953));
  nand_4 g13577(.A(n10510), .B(n2024), .Y(new_n13954));
  nand_4 g13578(.A(n10644), .B(n7946), .Y(new_n13955));
  xor_3  g13579(.A(new_n13955), .B(new_n13954), .Y(new_n13956));
  xnor_3 g13580(.A(new_n13956), .B(new_n13953), .Y(new_n13957));
  xnor_3 g13581(.A(new_n13957), .B(new_n13950), .Y(new_n13958));
  xnor_3 g13582(.A(new_n13958), .B(new_n13945), .Y(new_n13959));
  xnor_3 g13583(.A(new_n13959), .B(new_n13940), .Y(new_n13960));
  xnor_3 g13584(.A(new_n13960), .B(new_n13937), .Y(new_n13961));
  xnor_3 g13585(.A(new_n13961), .B(new_n13859), .Y(new_n13962));
  xnor_3 g13586(.A(new_n13962), .B(new_n13814), .Y(new_n13963));
  xnor_3 g13587(.A(new_n13963), .B(new_n13806), .Y(new_n13964));
  nand_4 g13588(.A(n9111), .B(n5857), .Y(new_n13965));
  nand_4 g13589(.A(n7965), .B(n6431), .Y(new_n13966));
  xor_3  g13590(.A(new_n13966), .B(new_n13965), .Y(new_n13967));
  not_3  g13591(.A(new_n13967), .Y(new_n13968));
  xnor_3 g13592(.A(new_n13968), .B(new_n13964), .Y(new_n13969));
  not_3  g13593(.A(new_n5845), .Y(new_n13970));
  nand_4 g13594(.A(new_n5849), .B(new_n13970), .Y(new_n13971));
  not_3  g13595(.A(new_n5941), .Y(new_n13972));
  nand_4 g13596(.A(new_n13972), .B(new_n5850), .Y(new_n13973));
  nand_4 g13597(.A(new_n13973), .B(new_n13971), .Y(new_n13974));
  not_3  g13598(.A(new_n5931), .Y(new_n13975));
  not_3  g13599(.A(new_n5938), .Y(new_n13976));
  nand_4 g13600(.A(new_n13976), .B(new_n13975), .Y(new_n13977));
  xnor_3 g13601(.A(new_n13977), .B(new_n13974), .Y(new_n13978));
  xnor_3 g13602(.A(new_n13978), .B(new_n13969), .Y(new_n13979));
  xnor_3 g13603(.A(new_n13979), .B(new_n13786), .Y(n11707));
  not_3  g13604(.A(new_n6521), .Y(new_n13981));
  xor_3  g13605(.A(new_n13981), .B(new_n6520), .Y(n11755));
  xor_3  g13606(.A(new_n3838), .B(new_n3834), .Y(n11780));
  not_3  g13607(.A(new_n10445), .Y(new_n13984));
  xor_3  g13608(.A(new_n10446), .B(new_n13984), .Y(n11919));
  xor_3  g13609(.A(new_n10448), .B(new_n10430), .Y(n12005));
  xnor_3 g13610(.A(new_n10897), .B(new_n10892), .Y(n12014));
  not_3  g13611(.A(new_n9143), .Y(new_n13988));
  xnor_3 g13612(.A(new_n13988), .B(new_n9100), .Y(n12020));
  not_3  g13613(.A(new_n11924), .Y(new_n13990));
  xor_3  g13614(.A(new_n11963), .B(new_n13990), .Y(n12076));
  xnor_3 g13615(.A(new_n12528), .B(new_n12520), .Y(n12111));
  xnor_3 g13616(.A(new_n10899), .B(new_n10883), .Y(n12444));
  nor_4  g13617(.A(new_n5790), .B(new_n5788), .Y(new_n13994));
  xnor_3 g13618(.A(new_n13994), .B(new_n5804), .Y(n12807));
endmodule


