
module top_809568696_809776567_809698999_863110837_1234615 (n74, n203, n271, n394, n411, n427, n462, n498, n650, n656, n666, n674, n702, n730, n737, n760, n844, n977, n1027, n1093, n1222, n1265, n1268, n1347, n1568, n1637, n1702, n1763, n1776, n2048, n2061, n2164, n2166, n2201, n2334, n2454, n2573, n2615, n2674, n2699, n2895, n3130, n3166, n3263, n3367, n3388, n3506, n3532, n3652, n3655, n3673, n3775, n3799, n3804, n3833, n3893, n3910, n3972, n4000, n4022, n4039, n4117, n4131, n4147, n4154, n4172, n4175, n4225, n4282, n4292, n4615, n4659, n4755, n4774, n4785, n4895, n4907, n5009, n5014, n5023, n5033, n5046, n5077, n5184, n5185, n5225, n5430, n5449, n5467, n5502, n5601, n5725, n5786, n5943, n5950, n5960, n6007, n6054, n6114, n6147, n6251, n6258, n6270, n6362, n6436, n6460, n6480, n6517, n6555, n6586, n6680, n6693, n6703, n6758, n6791, n6810, n6873, n6946, n6999, n7104, n7272, n7282, n7354, n7450, n7652, n7667, n7748, n7832, n7941, n7972, n7988, n8002, n8044, n8073, n8204, n8262, n8302, n8315, n8397, n8439, n8463, n8486, n8550, n8552, n8598, n8635, n8649, n8737, n8746, n8780, n8799, n8800, n8873, n8892, n8926, n8997, n9026, n9110, n9154, n9186, n9252, n9314, n9543, n9544, n9555, n9589, n9830, n9893, n9921, n9936, n9977, n10050, n10051, n10061, n10080, n10112, n10147, n10255, n10278, n10283, n10378, n10407, n10426, n10446, n10466, n10470, n10573, n10615, n10630, n10736, n10750, n10765, n10862, n10912, n10945, n11143, n11158, n11269, n11345, n11404, n11529, n11590, n11605, n11666, n11756, n11776, n11842, n11854, n11875, n11902, n11930, n11933, n11961, n12009, n12012, n12025, n12142, n12218, n12270, n12321, n12336, n12573, n12614, n12782, n12829, n12885, n12927, n12976, n13000, n13093, n13102, n13109, n13186, n13224, n13231, n13295, n13363, n13364, n13509, n13511, n13561, n13625, n13636, n13814, n13882, n13890, n13944, n13992, n14072, n14163, n14293, n14303, n14408, n14464, n14475, n14483, n8, n46, n91, n126, n278, n389, n451, n490, n543, n682, n884, n948, n1094, n1122, n1124, n1329, n1545, n1739, n1827, n1900, n1927, n1951, n2027, n2126, n2175, n2223, n2311, n2407, n2556, n2559, n2572, n2672, n2734, n3090, n3242, n3340, n3603, n3854, n3901, n4125, n4279, n4305, n4345, n4437, n4541, n4604, n4672, n4858, n4971, n5479, n5550, n5586, n5806, n5851, n5987, n6012, n6198, n6275, n6314, n6682, n6696, n6786, n6853, n6952, n6979, n7071, n7073, n7132, n7152, n7246, n7265, n7382, n7655, n7771, n7825, n8068, n8085, n8124, n8144, n8215, n8306, n8471, n8604, n8909, n9096, n9342, n9437, n9447, n9570, n9665, n9717, n10515, n10591, n10791, n10802, n10915, n11122, n11393, n11463, n11534, n11627, n11664, n11822, n11847, n12032, n12166, n12232, n12355, n12535, n12989, n13010, n13045, n13114, n13141, n13316, n13577, n13639, n13658, n13693, n13760, n13853, n13870, n13953, n13959, n14289, n14307, n14330, n14399, n14463);
input n74, n203, n271, n394, n411, n427, n462, n498, n650, n656, n666, n674, n702, n730, n737, n760, n844, n977, n1027, n1093, n1222, n1265, n1268, n1347, n1568, n1637, n1702, n1763, n1776, n2048, n2061, n2164, n2166, n2201, n2334, n2454, n2573, n2615, n2674, n2699, n2895, n3130, n3166, n3263, n3367, n3388, n3506, n3532, n3652, n3655, n3673, n3775, n3799, n3804, n3833, n3893, n3910, n3972, n4000, n4022, n4039, n4117, n4131, n4147, n4154, n4172, n4175, n4225, n4282, n4292, n4615, n4659, n4755, n4774, n4785, n4895, n4907, n5009, n5014, n5023, n5033, n5046, n5077, n5184, n5185, n5225, n5430, n5449, n5467, n5502, n5601, n5725, n5786, n5943, n5950, n5960, n6007, n6054, n6114, n6147, n6251, n6258, n6270, n6362, n6436, n6460, n6480, n6517, n6555, n6586, n6680, n6693, n6703, n6758, n6791, n6810, n6873, n6946, n6999, n7104, n7272, n7282, n7354, n7450, n7652, n7667, n7748, n7832, n7941, n7972, n7988, n8002, n8044, n8073, n8204, n8262, n8302, n8315, n8397, n8439, n8463, n8486, n8550, n8552, n8598, n8635, n8649, n8737, n8746, n8780, n8799, n8800, n8873, n8892, n8926, n8997, n9026, n9110, n9154, n9186, n9252, n9314, n9543, n9544, n9555, n9589, n9830, n9893, n9921, n9936, n9977, n10050, n10051, n10061, n10080, n10112, n10147, n10255, n10278, n10283, n10378, n10407, n10426, n10446, n10466, n10470, n10573, n10615, n10630, n10736, n10750, n10765, n10862, n10912, n10945, n11143, n11158, n11269, n11345, n11404, n11529, n11590, n11605, n11666, n11756, n11776, n11842, n11854, n11875, n11902, n11930, n11933, n11961, n12009, n12012, n12025, n12142, n12218, n12270, n12321, n12336, n12573, n12614, n12782, n12829, n12885, n12927, n12976, n13000, n13093, n13102, n13109, n13186, n13224, n13231, n13295, n13363, n13364, n13509, n13511, n13561, n13625, n13636, n13814, n13882, n13890, n13944, n13992, n14072, n14163, n14293, n14303, n14408, n14464, n14475, n14483;
output n8, n46, n91, n126, n278, n389, n451, n490, n543, n682, n884, n948, n1094, n1122, n1124, n1329, n1545, n1739, n1827, n1900, n1927, n1951, n2027, n2126, n2175, n2223, n2311, n2407, n2556, n2559, n2572, n2672, n2734, n3090, n3242, n3340, n3603, n3854, n3901, n4125, n4279, n4305, n4345, n4437, n4541, n4604, n4672, n4858, n4971, n5479, n5550, n5586, n5806, n5851, n5987, n6012, n6198, n6275, n6314, n6682, n6696, n6786, n6853, n6952, n6979, n7071, n7073, n7132, n7152, n7246, n7265, n7382, n7655, n7771, n7825, n8068, n8085, n8124, n8144, n8215, n8306, n8471, n8604, n8909, n9096, n9342, n9437, n9447, n9570, n9665, n9717, n10515, n10591, n10791, n10802, n10915, n11122, n11393, n11463, n11534, n11627, n11664, n11822, n11847, n12032, n12166, n12232, n12355, n12535, n12989, n13010, n13045, n13114, n13141, n13316, n13577, n13639, n13658, n13693, n13760, n13853, n13870, n13953, n13959, n14289, n14307, n14330, n14399, n14463;
wire n0, n1, n2, n3, n4, n5, n6, n7, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n272, n273, n274, n275, n276, n277, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n390, n391, n392, n393, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n491, n492, n493, n494, n495, n496, n497, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n651, n652, n653, n654, n655, n657, n658, n659, n660, n661, n662, n663, n664, n665, n667, n668, n669, n670, n671, n672, n673, n675, n676, n677, n678, n679, n680, n681, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n731, n732, n733, n734, n735, n736, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1123, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1266, n1267, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2165, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2557, n2558, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2673, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3653, n3654, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3800, n3801, n3802, n3803, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4126, n4127, n4128, n4129, n4130, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4148, n4149, n4150, n4151, n4152, n4153, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4173, n4174, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4280, n4281, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5010, n5011, n5012, n5013, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5944, n5945, n5946, n5947, n5948, n5949, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6008, n6009, n6010, n6011, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6252, n6253, n6254, n6255, n6256, n6257, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6271, n6272, n6273, n6274, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6681, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6694, n6695, n6697, n6698, n6699, n6700, n6701, n6702, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6787, n6788, n6789, n6790, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6947, n6948, n6949, n6950, n6951, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7072, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7266, n7267, n7268, n7269, n7270, n7271, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7653, n7654, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7826, n7827, n7828, n7829, n7830, n7831, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8069, n8070, n8071, n8072, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8303, n8304, n8305, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8551, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8599, n8600, n8601, n8602, n8603, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10279, n10280, n10281, n10282, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10467, n10468, n10469, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10913, n10914, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11530, n11531, n11532, n11533, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11665, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11843, n11844, n11845, n11846, n11848, n11849, n11850, n11851, n11852, n11853, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11931, n11932, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12010, n12011, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12026, n12027, n12028, n12029, n12030, n12031, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13103, n13104, n13105, n13106, n13107, n13108, n13110, n13111, n13112, n13113, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13225, n13226, n13227, n13228, n13229, n13230, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13510, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13637, n13638, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13954, n13955, n13956, n13957, n13958, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14290, n14291, n14292, n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14304, n14305, n14306, n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526;
assign n6289 = n9151 | n3294;
assign n7757 = ~(n12807 | n10319);
assign n2651 = ~n13041;
assign n10364 = n12601 | n9558;
assign n1362 = ~n7322;
assign n6140 = n4052 | n8064;
assign n8630 = ~n13734;
assign n14021 = n4289 & n6390;
assign n6317 = n5240 & n5350;
assign n13791 = n4871 | n5786;
assign n178 = n11607 & n9635;
assign n1013 = n12528 | n7972;
assign n5244 = n406 & n40;
assign n2507 = n14188 | n14051;
assign n10110 = ~(n4544 | n11112);
assign n12465 = n13676 & n4145;
assign n2021 = ~n5795;
assign n180 = n4102 & n11811;
assign n5358 = n3986 & n2419;
assign n2530 = ~(n2597 | n7614);
assign n7263 = n7529 & n8354;
assign n9031 = n11687 & n5664;
assign n12876 = ~(n1944 | n5100);
assign n12900 = ~n5725;
assign n13931 = n4300 & n5032;
assign n9422 = ~n1894;
assign n10151 = n4967 | n8596;
assign n10115 = n3271 & n3260;
assign n2332 = n4022 | n11875;
assign n13604 = n5715 | n13570;
assign n10494 = n7116 | n7870;
assign n12899 = n11142 & n12366;
assign n12249 = n10994 & n9776;
assign n1389 = n12918 & n5537;
assign n1944 = ~n11302;
assign n14312 = ~n3287;
assign n11237 = n12870 | n9767;
assign n5724 = ~(n11180 | n2128);
assign n5129 = ~n1243;
assign n7303 = n12020 | n6027;
assign n7754 = n3804 | n7652;
assign n667 = n14373 & n3634;
assign n1675 = ~(n10233 | n7403);
assign n4909 = n4354 & n3671;
assign n3977 = ~n10824;
assign n1030 = n5229 & n8184;
assign n1263 = ~(n9806 | n9496);
assign n10882 = n14042 & n2697;
assign n10974 = n10871 | n12320;
assign n13428 = n11558 | n7538;
assign n7180 = n13103 & n12346;
assign n10950 = n976 | n437;
assign n2889 = ~n13425;
assign n5592 = n4098 & n3065;
assign n10914 = n10808 | n13594;
assign n9665 = n13511 & n9733;
assign n4403 = n8801 & n10549;
assign n13412 = n13083 | n942;
assign n7567 = n14286 & n7644;
assign n781 = ~n7339;
assign n2362 = n3093 | n3943;
assign n6672 = ~n6357;
assign n14005 = n5236 | n11954;
assign n7129 = n13297 & n187;
assign n5481 = n2949 | n9091;
assign n32 = ~(n4913 | n8126);
assign n4943 = n3212 & n4990;
assign n9606 = ~(n1473 | n6423);
assign n6879 = n2177 & n2552;
assign n8081 = ~n4036;
assign n13550 = n10960 | n5342;
assign n3660 = n1137 | n11790;
assign n7712 = n14093 & n5157;
assign n1612 = ~n3572;
assign n8287 = n9229 | n7331;
assign n10768 = n11647 | n1547;
assign n1571 = ~n8357;
assign n10012 = n6383 | n10051;
assign n8432 = ~n8524;
assign n3531 = n8376 | n9589;
assign n114 = n4851 & n14280;
assign n13990 = n13507 | n6436;
assign n1358 = n12401 | n5643;
assign n13163 = ~(n4924 | n5324);
assign n4951 = n4856 & n6884;
assign n4953 = n666 | n13511;
assign n13989 = n4433 & n12947;
assign n6927 = n4422 & n7485;
assign n12632 = n13220 | n7191;
assign n1237 = n10763 & n14040;
assign n11299 = ~(n7011 | n12162);
assign n6595 = ~n5627;
assign n8048 = ~n12014;
assign n1817 = n9375 | n5095;
assign n3861 = ~n2958;
assign n10345 = n5092 & n5407;
assign n10477 = n7421 & n3669;
assign n6283 = n9353 | n11650;
assign n8753 = n13087 | n4518;
assign n7689 = ~n7056;
assign n11411 = ~n4266;
assign n8957 = n14282 | n12902;
assign n3822 = n11345 | n5786;
assign n10518 = n14450 | n10147;
assign n5897 = ~n13967;
assign n2125 = ~(n12904 | n10607);
assign n9733 = ~(n5237 | n8944);
assign n3022 = n6822 & n9199;
assign n13113 = n11710 | n7021;
assign n230 = ~n5178;
assign n2015 = n9140 | n13351;
assign n5150 = n10019 | n6737;
assign n10329 = ~(n13356 | n9372);
assign n14316 = n7219 | n6307;
assign n2931 = n5064 | n4181;
assign n14134 = ~n7940;
assign n3978 = n8950 & n7597;
assign n10926 = n5807 | n12141;
assign n2400 = n8908 | n11465;
assign n3379 = n5064 | n4227;
assign n3473 = n14260 & n4003;
assign n4506 = n1876 & n13713;
assign n1570 = n2878 | n2225;
assign n7120 = ~n9193;
assign n4303 = n14321 & n515;
assign n7496 = ~(n8189 | n12030);
assign n13881 = ~(n906 | n11277);
assign n8378 = ~n409;
assign n10354 = n55 & n876;
assign n671 = n6242 | n10752;
assign n10988 = n14419 | n7643;
assign n9461 = ~n10395;
assign n1521 = n13555 & n5463;
assign n9282 = ~(n4195 | n5747);
assign n923 = n2533 & n872;
assign n475 = n14366 | n43;
assign n10159 = n10461 | n11364;
assign n742 = ~n241;
assign n2487 = n8582 | n4719;
assign n6976 = n2224 & n13663;
assign n11242 = n7957 & n7138;
assign n13973 = n3394 | n13859;
assign n10150 = n14313 & n8116;
assign n6327 = ~(n6672 | n12268);
assign n8613 = n5450 | n6229;
assign n13372 = n12353 | n12385;
assign n4979 = n14213 & n13576;
assign n5403 = n3886 | n13790;
assign n10140 = n10560 | n3600;
assign n7473 = n13297 & n6951;
assign n1260 = n12768 | n8737;
assign n12910 = n2888 | n3360;
assign n11192 = ~(n9795 | n14259);
assign n2440 = n286 & n6562;
assign n9122 = n12100 | n3017;
assign n6330 = n5234 | n9338;
assign n577 = n8412 & n9010;
assign n5991 = n1539 & n8103;
assign n13206 = ~n1813;
assign n3358 = n13698 | n12441;
assign n11824 = ~n730;
assign n8532 = n1431 & n9764;
assign n1239 = n3667 | n7380;
assign n5700 = n6350 | n11949;
assign n9728 = n10589 & n7148;
assign n8319 = n3419 | n13363;
assign n234 = ~n12489;
assign n12215 = n9806 | n3147;
assign n1210 = ~n427;
assign n13229 = n2949 | n12427;
assign n5227 = n13367 & n13687;
assign n5884 = n6016 & n4531;
assign n13142 = ~n3455;
assign n10751 = ~n6989;
assign n4124 = n3025 | n13332;
assign n6783 = n14107 | n1670;
assign n10728 = n3766 & n10226;
assign n12046 = ~n2503;
assign n14459 = n12047 | n3153;
assign n10148 = ~(n13977 | n12002);
assign n225 = ~n13734;
assign n10452 = n5570 | n2786;
assign n4081 = n646 & n12722;
assign n14045 = n1821 | n1663;
assign n6055 = n6937 & n5756;
assign n5661 = n14449 | n13228;
assign n2053 = n390 | n3250;
assign n1666 = ~(n12453 | n1611);
assign n5425 = ~(n5209 | n3973);
assign n7269 = n9297 & n3135;
assign n1247 = ~n4535;
assign n11078 = ~(n12087 | n266);
assign n9429 = ~n11541;
assign n13292 = n163 | n7679;
assign n11582 = ~n9046;
assign n119 = n5139 | n112;
assign n7886 = ~n316;
assign n14368 = ~n9679;
assign n9468 = n12039 & n4393;
assign n10145 = n1520 & n12538;
assign n8413 = n1254 & n176;
assign n7977 = n7391 & n10720;
assign n2850 = ~n1706;
assign n13895 = n3715 & n13290;
assign n5453 = n2901 | n11010;
assign n5577 = ~(n900 | n1159);
assign n3528 = ~(n7551 | n4673);
assign n5191 = n1489 & n3415;
assign n7459 = ~(n13707 | n12055);
assign n4201 = ~(n14058 | n7577);
assign n5876 = ~n14135;
assign n132 = n12820 | n12260;
assign n6384 = ~(n13361 | n1887);
assign n12909 = n2608 | n6270;
assign n4115 = n6649 & n1186;
assign n6694 = n1051 | n13427;
assign n7923 = n12335 & n566;
assign n9196 = n3424 & n13690;
assign n9257 = n7961 & n14348;
assign n3378 = n14063 & n1429;
assign n904 = ~n5675;
assign n7591 = n12994 | n4852;
assign n3557 = ~(n2417 | n5339);
assign n3007 = n9041 & n53;
assign n13692 = n9375 | n292;
assign n11829 = n9218 | n1730;
assign n9459 = n747 | n14064;
assign n12492 = ~(n14216 | n11505);
assign n7739 = ~n12846;
assign n2077 = n10089 | n4450;
assign n599 = n2055 | n3975;
assign n621 = n3134 | n11268;
assign n6340 = n12759 | n14415;
assign n2958 = ~n744;
assign n9993 = n13718 | n2296;
assign n8041 = n1662 & n9420;
assign n13836 = n1480 | n8774;
assign n9379 = n12721 & n6215;
assign n10898 = n6649 & n7074;
assign n2692 = ~n2520;
assign n5328 = n28 | n1759;
assign n7005 = n1071 & n8665;
assign n2054 = ~(n10535 | n11034);
assign n5117 = n2067 & n6643;
assign n5794 = n1140 & n4191;
assign n5551 = n839 | n3185;
assign n3416 = n9920 & n11878;
assign n11617 = n2608 & n12132;
assign n5873 = ~n4022;
assign n14485 = ~(n4092 | n5385);
assign n14203 = n14227 & n13897;
assign n8222 = n392 & n11789;
assign n2784 = ~n7086;
assign n7805 = n3047 | n5590;
assign n8401 = ~n7275;
assign n9719 = n9564 & n1104;
assign n10930 = ~n14075;
assign n7762 = n8025 & n12129;
assign n4832 = n5800 | n9845;
assign n10338 = ~n3577;
assign n4103 = n6891 | n12575;
assign n13822 = n3952 & n10487;
assign n4028 = n12460 & n5859;
assign n4453 = n1339 & n7868;
assign n8514 = n13103 & n7290;
assign n12004 = n850 | n12983;
assign n3182 = ~n14164;
assign n11464 = n13952 & n12180;
assign n12070 = n2597 | n2062;
assign n6184 = ~(n3034 | n6131);
assign n9658 = n13650 & n1748;
assign n10730 = ~n13158;
assign n11610 = n8431 & n11351;
assign n14151 = n4844 & n2140;
assign n9814 = n13675 | n13972;
assign n1947 = n5084 | n8260;
assign n13399 = ~n2409;
assign n11778 = n12808 & n11452;
assign n5800 = ~n5242;
assign n12124 = n11048 | n9473;
assign n5432 = ~n13752;
assign n356 = n679 & n11927;
assign n10349 = ~(n9810 | n1469);
assign n6119 = ~n7533;
assign n6187 = n2985 & n11919;
assign n12032 = n8550 & n11192;
assign n8367 = n6109 | n2070;
assign n7808 = ~n10603;
assign n3524 = ~(n9124 | n1323);
assign n10771 = n12023 | n9312;
assign n7945 = n5587 | n4516;
assign n4219 = n8638 | n829;
assign n6543 = n7250 | n9003;
assign n3081 = n11411 & n3788;
assign n3507 = n11048 | n14513;
assign n5701 = n13535 & n1630;
assign n11650 = n406 & n2019;
assign n10677 = n7011 | n8863;
assign n11094 = ~n11415;
assign n1128 = n2897 | n12487;
assign n1493 = n1051 | n13543;
assign n4856 = ~n2744;
assign n5692 = n3607 & n10293;
assign n12075 = ~n11152;
assign n6194 = ~(n12087 | n3436);
assign n2761 = ~n1676;
assign n807 = n1844 | n14232;
assign n11565 = n10300 | n5433;
assign n3945 = n6822 & n2377;
assign n4966 = n8252 & n12430;
assign n12554 = n283 | n7190;
assign n7001 = n12353 | n1384;
assign n9647 = n2985 & n3283;
assign n563 = n2857 | n7982;
assign n7089 = n406 & n13;
assign n9258 = n10331 | n8968;
assign n1697 = ~n1220;
assign n10039 = n11028 & n7268;
assign n7919 = ~n13437;
assign n2773 = n11011 | n3246;
assign n12803 = n2790 | n11480;
assign n11048 = ~n11152;
assign n14245 = ~n12336;
assign n13564 = n889 & n2585;
assign n11789 = n6730 | n3299;
assign n6081 = ~(n12693 | n1782);
assign n13036 = n10351 | n7918;
assign n693 = n6854 & n13957;
assign n13901 = n1161 & n13128;
assign n5877 = n10134 & n4955;
assign n3982 = n4978 | n7155;
assign n6574 = n7122 | n6722;
assign n6648 = n11036 | n11273;
assign n6849 = ~n10466;
assign n8064 = n13236 & n13216;
assign n7519 = ~n11792;
assign n3555 = n7862 | n10379;
assign n4229 = n2510 | n3878;
assign n9680 = n4880 & n10324;
assign n3836 = n13446 | n7487;
assign n2578 = n13952 & n9827;
assign n13748 = n10072 & n11126;
assign n11639 = n2682 & n9993;
assign n4865 = ~n3542;
assign n2712 = n7003 | n1270;
assign n2643 = ~n11715;
assign n4834 = n13806 | n10935;
assign n3433 = n13656 & n9333;
assign n8535 = n3635 & n1216;
assign n5541 = n13877 & n10725;
assign n13660 = n11569 & n9112;
assign n1528 = n13555 & n9034;
assign n6880 = n8908 | n2496;
assign n1930 = n13433 & n11344;
assign n6822 = ~n6559;
assign n5349 = n3193 | n3142;
assign n8956 = n11360 | n12596;
assign n6526 = n10710 & n5965;
assign n766 = ~n4317;
assign n3026 = n1339 & n8846;
assign n7575 = ~n8565;
assign n6109 = ~n4606;
assign n12245 = n2983 & n8614;
assign n5293 = n11867 & n2411;
assign n2093 = n3800 | n8935;
assign n7238 = ~n11071;
assign n10169 = n10032 & n3656;
assign n3716 = ~(n12934 | n3464);
assign n5013 = n14404 | n9774;
assign n3422 = n6781 | n13546;
assign n1624 = n13069 & n8837;
assign n9847 = ~(n1697 | n8720);
assign n13517 = n6288 | n14169;
assign n12662 = n4407 | n10223;
assign n164 = ~(n8378 | n3964);
assign n7866 = n2099 & n14226;
assign n7440 = n8630 & n140;
assign n4434 = n12013 & n8017;
assign n4669 = n511 | n6553;
assign n3190 = n8066 & n1913;
assign n5256 = n7612 | n12573;
assign n97 = n1876 & n14338;
assign n469 = n10224 | n12365;
assign n10299 = n80 & n11237;
assign n8893 = n8427 & n3178;
assign n2447 = n5999 & n13452;
assign n2106 = n12278 | n7466;
assign n464 = n838 | n9489;
assign n11193 = n10960 | n12073;
assign n2723 = n4573 & n11068;
assign n11344 = n4180 | n9316;
assign n4244 = ~n7681;
assign n4477 = ~(n10323 | n2988);
assign n8706 = n10846 | n14408;
assign n7036 = n7354 | n13363;
assign n11846 = n1147 | n5771;
assign n1824 = n1489 & n863;
assign n4554 = ~n4135;
assign n3256 = n2724 & n11973;
assign n14179 = n7627 & n6188;
assign n7260 = n5603 | n3385;
assign n6220 = n10072 & n12861;
assign n7201 = n6389 & n10895;
assign n10990 = n4468 | n13479;
assign n2608 = ~n9830;
assign n8897 = ~n8148;
assign n4074 = n12428 | n14142;
assign n11295 = n4033 | n12341;
assign n8394 = n8045 | n9419;
assign n1025 = n1047 & n1208;
assign n3373 = n2587 & n7554;
assign n5161 = n5279 & n267;
assign n9966 = n3491 & n4649;
assign n12998 = ~n5268;
assign n9487 = n2098 | n1314;
assign n2385 = n3268 & n1503;
assign n2683 = n3559 | n4351;
assign n10172 = n14286 & n10157;
assign n2944 = n10035 | n5555;
assign n8826 = n769 | n7520;
assign n11318 = n69 | n4870;
assign n1403 = ~(n2889 | n606);
assign n1719 = n405 & n6165;
assign n12980 = n776 & n3930;
assign n8924 = n3320 | n14340;
assign n12466 = n5459 & n7869;
assign n4603 = n12092 & n14361;
assign n1478 = ~n10047;
assign n873 = ~n5153;
assign n1193 = ~n13003;
assign n9554 = n10834 | n941;
assign n14229 = n14450 & n13415;
assign n3295 = n12460 & n13188;
assign n8617 = ~(n9601 | n1954);
assign n14226 = n10019 | n10727;
assign n6709 = n405 & n4701;
assign n1914 = ~n13901;
assign n12916 = n5825 & n8525;
assign n4875 = n11048 | n13872;
assign n9166 = n10136 | n4505;
assign n10531 = n5252 & n9116;
assign n10629 = n752 & n9465;
assign n12777 = n12820 | n13918;
assign n8934 = n2587 & n7878;
assign n12734 = n9972 & n764;
assign n412 = ~n3357;
assign n6291 = n5472 | n756;
assign n3421 = ~(n4877 | n3997);
assign n2640 = n5458 & n9397;
assign n527 = ~(n7886 | n8388);
assign n8554 = n1924 & n13923;
assign n12658 = n848 | n9936;
assign n13493 = n5317 & n6890;
assign n11181 = n8332 | n72;
assign n11082 = n28 | n7947;
assign n9757 = n350 & n8365;
assign n7119 = n12543 | n4040;
assign n6981 = ~n977;
assign n1279 = n4923 | n13750;
assign n12954 = n8747 | n6571;
assign n6841 = ~(n9305 | n13053);
assign n6115 = n6350 | n1968;
assign n11399 = n5236 | n11899;
assign n8526 = n1137 | n10910;
assign n6288 = ~n9959;
assign n2909 = n7768 & n3127;
assign n9318 = ~(n11697 | n4975);
assign n1395 = n7171 & n2627;
assign n5958 = ~(n4978 | n2189);
assign n14037 = n4790 & n3993;
assign n145 = n904 & n14224;
assign n12196 = n2783 & n9599;
assign n5376 = ~(n1127 | n725);
assign n9613 = ~n2816;
assign n6048 = ~(n1771 | n4696);
assign n10667 = n11176 | n2551;
assign n10802 = n13186 & n6448;
assign n1499 = n4128 | n10292;
assign n5924 = n5450 | n14448;
assign n12188 = n6649 & n3300;
assign n4694 = ~(n13875 | n7606);
assign n6928 = n400 & n10231;
assign n3086 = n14319 | n11596;
assign n7404 = n11654 & n6742;
assign n7811 = n10660 & n8706;
assign n11502 = n1660 | n167;
assign n3392 = n6206 | n5604;
assign n13934 = n7717 & n7218;
assign n6701 = n5048 & n9957;
assign n9444 = ~(n13283 | n2522);
assign n12115 = n5493 | n2632;
assign n13161 = n12039 & n4141;
assign n5043 = n8247 & n4964;
assign n3729 = n14430 | n13320;
assign n6434 = ~n10529;
assign n12313 = n13404 & n9528;
assign n14182 = n11576 | n10594;
assign n8745 = n432 & n10504;
assign n1489 = ~n5525;
assign n13479 = n7691 & n7504;
assign n12168 = n9206 | n5449;
assign n13337 = ~(n12922 | n5654);
assign n13009 = ~(n4144 | n12878);
assign n8794 = n3419 & n6144;
assign n7745 = ~n3926;
assign n13317 = ~n12909;
assign n1618 = n10408 & n5903;
assign n12128 = n9232 & n6621;
assign n12713 = n7898 | n8776;
assign n5423 = n7392 & n8292;
assign n10167 = n13700 & n12108;
assign n2516 = n7208 & n10836;
assign n3726 = ~(n6266 | n2854);
assign n8786 = ~n230;
assign n4312 = n2904 & n5506;
assign n11146 = n7708 | n8302;
assign n8570 = n13854 | n8954;
assign n5597 = ~(n1713 | n10604);
assign n12043 = n4788 & n1923;
assign n13601 = n12620 & n6983;
assign n2728 = n10458 & n7110;
assign n7283 = n5948 & n10778;
assign n7841 = ~(n12403 | n11898);
assign n11676 = ~n8598;
assign n2223 = n4175 & n6721;
assign n3571 = n2461 & n2526;
assign n382 = n2788 & n12304;
assign n104 = n13074 | n7797;
assign n11861 = ~n11195;
assign n8652 = n7887 | n4387;
assign n1492 = ~(n5762 | n7582);
assign n9984 = ~n1267;
assign n1910 = ~(n3768 | n13378);
assign n324 = n4195 | n1732;
assign n11500 = n10855 & n4680;
assign n10373 = ~(n12075 | n8143);
assign n7205 = n8358 & n14184;
assign n404 = n12057 & n13773;
assign n8943 = ~(n4877 | n11260);
assign n3668 = n8816 | n4916;
assign n11187 = n3370 & n5682;
assign n7543 = n965 & n2105;
assign n2836 = n747 | n12867;
assign n14526 = ~(n4829 | n13632);
assign n4737 = n2224 & n10514;
assign n2009 = n8799 | n12614;
assign n9795 = ~n2772;
assign n1813 = ~n2371;
assign n11691 = n8581 | n11461;
assign n10794 = n12292 | n6440;
assign n13689 = n6205 | n9237;
assign n11061 = n6046 | n9434;
assign n2844 = ~(n8301 | n7105);
assign n5266 = ~n5901;
assign n10835 = n2330 & n6599;
assign n5464 = n1061 | n8585;
assign n10117 = n11303 | n2078;
assign n9961 = n6192 & n269;
assign n5173 = n4098 & n12914;
assign n4495 = n8986 | n4768;
assign n7013 = ~(n11094 | n8982);
assign n10777 = n2149 | n3295;
assign n4613 = n6016 & n8254;
assign n5629 = n3405 & n9298;
assign n10739 = ~(n12705 | n10235);
assign n1132 = n286 & n4190;
assign n1698 = n4908 | n6550;
assign n8030 = n8393 & n5346;
assign n2565 = n4407 | n6591;
assign n17 = n11679 & n7635;
assign n3314 = n1266 & n4411;
assign n1673 = n4394 & n11528;
assign n3937 = ~(n8663 | n10952);
assign n5409 = ~n1833;
assign n1191 = n228 | n10137;
assign n6861 = n9819 | n1093;
assign n5270 = n4435 | n11855;
assign n3240 = n11157 & n3690;
assign n6921 = n10338 & n8915;
assign n3711 = n11724 | n136;
assign n7592 = n687 & n3379;
assign n10979 = n14351 & n12137;
assign n13577 = n9110 & n467;
assign n4332 = n8702 & n10389;
assign n2472 = n3233 & n11617;
assign n4505 = n4095 & n10545;
assign n4079 = ~(n7904 | n12430);
assign n3855 = n12335 & n9676;
assign n7836 = n2942 & n5452;
assign n12547 = n976 | n6924;
assign n10698 = n14404 | n9222;
assign n3714 = n8250 & n9777;
assign n10702 = n13847 | n9860;
assign n2120 = n4574 & n14185;
assign n896 = n2179 | n4587;
assign n115 = n14210 & n10000;
assign n8297 = n7462 | n5215;
assign n12516 = n12015 & n2392;
assign n3361 = ~n13983;
assign n661 = n13991 | n14444;
assign n3640 = ~n8899;
assign n14019 = ~(n3822 | n11763);
assign n6975 = ~n2011;
assign n14493 = n10855 & n12796;
assign n11750 = n9807 | n7713;
assign n8582 = ~n2918;
assign n4871 = ~n3532;
assign n10850 = n2229 | n8077;
assign n4011 = n12226 & n1510;
assign n7341 = n11722 | n10826;
assign n13559 = n8043 & n13280;
assign n3514 = n1854 & n2839;
assign n12177 = n501 & n4192;
assign n2169 = n2064 & n13292;
assign n5172 = ~n521;
assign n9895 = n2587 & n1067;
assign n4387 = n406 & n10926;
assign n14390 = ~(n882 | n11671);
assign n5663 = n4382 & n7758;
assign n6100 = n7914 | n1146;
assign n5468 = ~n3007;
assign n12578 = n6373 | n8588;
assign n7418 = ~n11456;
assign n9810 = n4147 | n10378;
assign n5121 = n5570 | n6800;
assign n4 = ~(n6797 | n8449);
assign n11709 = ~(n5365 | n4645);
assign n11796 = ~(n1480 | n6646);
assign n2777 = n1354 & n14105;
assign n10554 = ~(n13201 | n10900);
assign n260 = n4422 & n7330;
assign n12092 = ~n13383;
assign n12444 = n6536 & n510;
assign n6094 = ~(n14370 | n6918);
assign n320 = ~n5950;
assign n6502 = ~(n8592 | n13214);
assign n10738 = n12092 & n8725;
assign n4498 = ~n12249;
assign n3108 = n2747 | n9173;
assign n2205 = n172 | n1704;
assign n5272 = n2330 & n9857;
assign n3380 = ~(n11998 | n10655);
assign n3218 = n6271 | n6748;
assign n7678 = ~n238;
assign n12918 = ~n13219;
assign n5167 = n6128 & n9161;
assign n4233 = ~n4465;
assign n1087 = n9724 & n1516;
assign n3860 = n9442 | n12550;
assign n11390 = n13107 & n677;
assign n3099 = ~n5974;
assign n12309 = n12229 & n5988;
assign n4707 = n5507 | n12775;
assign n149 = n7003 | n5746;
assign n12386 = n7779 & n372;
assign n4198 = n7203 & n14445;
assign n12383 = n6135 & n12788;
assign n6754 = ~n11975;
assign n3848 = ~(n11325 | n11999);
assign n12816 = n11576 | n5367;
assign n1954 = ~(n9035 | n7143);
assign n8115 = ~n6074;
assign n5872 = n348 & n13207;
assign n6071 = n1427 & n6005;
assign n842 = n7826 & n12497;
assign n9884 = n11951 | n5136;
assign n8411 = n5936 | n485;
assign n2210 = n4757 & n13143;
assign n4396 = ~(n5780 | n14243);
assign n721 = n4581 & n1008;
assign n4441 = n11804 | n4436;
assign n3597 = n2643 & n9761;
assign n2273 = n7826 & n9538;
assign n12792 = n6109 | n10060;
assign n1785 = n12549 | n13614;
assign n12933 = ~n12321;
assign n1588 = ~n8656;
assign n13273 = ~(n5468 | n4063);
assign n4370 = n3161 | n531;
assign n214 = n5800 | n1877;
assign n3055 = n8300 & n3570;
assign n10463 = n3405 & n2013;
assign n2808 = ~n4510;
assign n2502 = n1117 & n3617;
assign n13159 = ~(n3546 | n2345);
assign n12991 = n2315 | n2196;
assign n10037 = n7898 | n2388;
assign n5882 = n1904 & n9221;
assign n7419 = ~n1478;
assign n12304 = ~n13714;
assign n9271 = n12759 | n7730;
assign n2364 = n4347 & n14462;
assign n9120 = n4340 | n3391;
assign n190 = n1362 | n13031;
assign n9867 = n14351 & n10891;
assign n12272 = n6848 & n1165;
assign n7026 = ~n6559;
assign n11371 = ~(n11259 | n5199);
assign n3220 = n14465 & n6775;
assign n1422 = n13155 | n10526;
assign n7809 = ~n9231;
assign n3312 = n10595 & n4616;
assign n12432 = n8096 | n8955;
assign n7044 = n116 | n8634;
assign n7430 = ~n11331;
assign n1835 = n8396 | n1078;
assign n13823 = ~n4928;
assign n9264 = n7430 | n12418;
assign n5021 = n900 | n7746;
assign n14110 = ~n12687;
assign n2732 = n3826 | n12234;
assign n12602 = n1261 | n3448;
assign n3297 = n904 & n6876;
assign n8150 = n5406 | n1931;
assign n4026 = n850 | n7964;
assign n6848 = ~n4292;
assign n4817 = n5493 | n10948;
assign n3481 = n12013 & n8788;
assign n13315 = n10357 & n14140;
assign n4676 = n12625 | n1963;
assign n471 = n6753 & n7119;
assign n6557 = n3405 & n4420;
assign n14138 = n7358 | n8281;
assign n6107 = n2315 | n8808;
assign n877 = n3942 & n9346;
assign n4830 = n11676 & n6408;
assign n14377 = ~n9721;
assign n6262 = n12185 & n6717;
assign n5723 = n3169 & n5211;
assign n12026 = n13362 & n12597;
assign n12285 = n4908 | n471;
assign n8874 = ~(n11580 | n6191);
assign n7391 = ~n11369;
assign n5088 = ~n1639;
assign n9143 = n10933 | n9823;
assign n13929 = n3672 & n8842;
assign n9033 = ~(n4092 | n13984);
assign n8173 = n1821 | n9663;
assign n1846 = n7156 | n1113;
assign n11171 = ~n2970;
assign n5834 = n1348 | n1706;
assign n4888 = n4544 | n3378;
assign n8847 = n13867 | n10061;
assign n8891 = n9211 | n8832;
assign n10280 = ~n5738;
assign n12434 = n1729 & n4087;
assign n5137 = ~n6657;
assign n7744 = n6344 | n12819;
assign n4698 = ~n6362;
assign n13079 = n10523 | n5681;
assign n10928 = n3047 | n8024;
assign n10868 = n817 | n577;
assign n575 = n5553 & n2968;
assign n3828 = n6343 & n6901;
assign n10276 = ~n2428;
assign n3767 = n3986 & n7260;
assign n8604 = n5786 & n2183;
assign n12119 = ~(n8277 | n5676);
assign n2095 = n12858 & n9098;
assign n8491 = n820 | n13302;
assign n285 = n4690 & n11663;
assign n2018 = n6625 & n3599;
assign n697 = n781 | n10546;
assign n1432 = ~(n1844 | n10823);
assign n3203 = n678 & n6453;
assign n5549 = n7433 & n13132;
assign n6121 = ~(n7754 | n6948);
assign n10829 = n1623 | n7763;
assign n13883 = n7122 | n8264;
assign n4337 = ~(n1628 | n13070);
assign n7147 = n1708 & n14323;
assign n4161 = n1937 & n13293;
assign n9949 = n10247 & n6286;
assign n3981 = n6486 & n798;
assign n6491 = n5062 & n520;
assign n5101 = n11803 & n14308;
assign n2947 = ~(n5986 | n1762);
assign n4363 = ~(n10179 | n11964);
assign n2078 = n4244 & n10404;
assign n1194 = ~(n919 | n11685);
assign n8698 = n1788 & n9077;
assign n9195 = n9541 | n7080;
assign n11703 = n8897 | n2083;
assign n326 = n55 & n11256;
assign n13120 = n13978 | n468;
assign n11742 = n12633 | n8678;
assign n13115 = n3219 | n8625;
assign n3407 = n8950 & n2954;
assign n4678 = n2527 & n3329;
assign n4072 = n14376 | n13364;
assign n10010 = n12023 | n2771;
assign n10929 = ~n8131;
assign n8165 = n14091 & n5087;
assign n4491 = ~n2470;
assign n7359 = ~n8272;
assign n5178 = n4871 & n11763;
assign n8898 = n9289 | n2825;
assign n2810 = n10781 | n2247;
assign n36 = n748 & n7950;
assign n3044 = n12820 | n2321;
assign n13764 = n12994 | n8931;
assign n4779 = n225 & n3205;
assign n9093 = n2378 & n8491;
assign n12090 = n12149 | n7836;
assign n8172 = ~n565;
assign n11555 = n13676 & n2842;
assign n4148 = n7970 & n4689;
assign n7533 = n10660 & n7087;
assign n8481 = ~(n1425 | n13400);
assign n11176 = ~n1060;
assign n996 = n10024 | n9421;
assign n6028 = ~(n2086 | n9785);
assign n8191 = n11580 | n6736;
assign n9568 = n3932 & n5707;
assign n10383 = ~n12687;
assign n3953 = n10960 | n10113;
assign n2807 = ~(n14238 | n8201);
assign n8054 = n6343 & n8387;
assign n2716 = n8692 & n12291;
assign n10880 = n2067 & n8472;
assign n6212 = n5188 & n11778;
assign n9168 = n791 | n9870;
assign n2085 = n2177 & n4459;
assign n9412 = n14282 | n4909;
assign n9741 = n14150 & n853;
assign n13683 = n4581 & n8731;
assign n7780 = n647 | n6846;
assign n8546 = n222 & n174;
assign n10684 = n14260 & n5911;
assign n39 = n9232 & n12134;
assign n6453 = n3527 | n5272;
assign n10421 = n5335 & n8344;
assign n4319 = n11379 | n1155;
assign n11734 = n2857 | n6526;
assign n3350 = n1660 | n2299;
assign n11332 = ~(n9216 | n4469);
assign n5578 = n432 & n464;
assign n13116 = n13209 & n6569;
assign n8708 = n8300 & n899;
assign n596 = n3365 & n9621;
assign n9906 = n10534 | n5953;
assign n8445 = n6781 | n9919;
assign n2476 = n2998 & n6973;
assign n4239 = ~n9354;
assign n7677 = ~n8168;
assign n11702 = ~n3313;
assign n7439 = ~(n10309 | n11755);
assign n14435 = ~n4939;
assign n10131 = n10383 | n0;
assign n4016 = n8232 & n6880;
assign n11337 = n10637 | n12356;
assign n8797 = n555 | n1743;
assign n291 = n172 | n12502;
assign n45 = n6609 & n9598;
assign n10651 = ~n5905;
assign n11042 = n10566 & n3253;
assign n5203 = n8801 & n5284;
assign n11785 = n9422 | n6465;
assign n1609 = n13112 | n5656;
assign n13839 = ~(n13190 | n12467);
assign n7483 = n14198 | n5530;
assign n4447 = ~n6586;
assign n7431 = ~(n9546 | n9203);
assign n14375 = n10197 & n1336;
assign n497 = n13745 & n2366;
assign n12626 = ~(n12311 | n491);
assign n8521 = n12992 | n656;
assign n4489 = n13342 & n6523;
assign n8049 = n2804 & n6640;
assign n9094 = ~(n2218 | n4664);
assign n5242 = n4047 & n10236;
assign n692 = n4123 | n10862;
assign n47 = ~(n4608 | n4507);
assign n251 = ~n14354;
assign n7505 = n8980 | n1942;
assign n1726 = n11406 & n4780;
assign n10650 = ~n8345;
assign n4425 = n9972 & n11029;
assign n6380 = n536 & n9085;
assign n12404 = ~n11547;
assign n10947 = n4655 & n4339;
assign n9745 = ~n3356;
assign n87 = n3076 | n12608;
assign n8139 = ~(n11094 | n9498);
assign n5766 = n9806 | n9457;
assign n9519 = ~(n11580 | n2350);
assign n4428 = n6891 | n943;
assign n9426 = n1788 & n14014;
assign n6681 = n12651 | n11984;
assign n4334 = n14465 & n3684;
assign n7064 = n5980 & n7077;
assign n3184 = n4602 | n7316;
assign n3189 = n2961 & n11522;
assign n9675 = ~(n13248 | n5714);
assign n1164 = n13421 & n10227;
assign n400 = ~n7652;
assign n1782 = n2758 & n10442;
assign n8782 = n1628 | n11242;
assign n11407 = n1857 & n9828;
assign n2475 = n3762 & n4067;
assign n9245 = ~n13231;
assign n11072 = n10871 | n7854;
assign n10404 = n10449 | n10365;
assign n9175 = n1840 | n1721;
assign n9403 = ~n7064;
assign n6623 = n12968 | n9256;
assign n11432 = ~(n10977 | n11802);
assign n6933 = ~n9377;
assign n5883 = ~(n13981 | n2122);
assign n2404 = n4562 | n4032;
assign n1497 = n7768 & n12908;
assign n1486 = ~(n6039 | n11926);
assign n8936 = n9191 & n12350;
assign n10144 = n10197 & n2993;
assign n8273 = n12494 | n4122;
assign n7170 = ~(n329 | n6172);
assign n6403 = ~(n1617 | n2879);
assign n1276 = n12934 | n1467;
assign n8692 = ~n4824;
assign n8255 = n1535 | n3240;
assign n7662 = ~n4835;
assign n10293 = n227 | n3081;
assign n7985 = ~(n300 | n11246);
assign n10833 = n12147 & n2840;
assign n11838 = ~n8451;
assign n2618 = n10458 & n13245;
assign n12707 = n4340 | n14131;
assign n4168 = n7888 | n8514;
assign n4474 = n3093 | n2144;
assign n6961 = n11953 | n12125;
assign n2662 = n6544 | n2808;
assign n10670 = n12414 | n5877;
assign n1682 = ~(n4877 | n701);
assign n9833 = n8986 | n9240;
assign n11207 = n706 & n277;
assign n13014 = n1711 | n8010;
assign n12083 = n1602 | n13504;
assign n11620 = ~n4465;
assign n9192 = ~(n7720 | n5982);
assign n4815 = n7068 & n10983;
assign n10787 = n5975 & n987;
assign n10639 = n619 | n5051;
assign n1708 = ~n7052;
assign n8534 = ~(n8015 | n11434);
assign n13838 = n13706 | n4025;
assign n10954 = n769 | n27;
assign n6678 = n4092 | n699;
assign n14080 = ~(n10715 | n5075);
assign n8933 = n6157 & n6468;
assign n1438 = n4822 | n683;
assign n14340 = n13676 & n12686;
assign n5450 = ~n630;
assign n12634 = n13367 & n12223;
assign n8216 = ~n8750;
assign n715 = n1391 | n1408;
assign n7256 = n13227 & n1590;
assign n11423 = n14227 & n10771;
assign n10617 = ~n1178;
assign n6971 = ~n2918;
assign n7055 = n5406 | n9370;
assign n3309 = ~n6308;
assign n8077 = n6051 & n3399;
assign n1314 = n5279 & n13077;
assign n13198 = n3667 | n8265;
assign n3034 = ~n1161;
assign n5679 = n12521 & n3938;
assign n6626 = n7060 & n4031;
assign n7478 = n6654 | n10252;
assign n13752 = n11852 & n9142;
assign n6503 = n1198 | n758;
assign n3803 = n13626 & n6104;
assign n9408 = ~(n8825 | n9901);
assign n2560 = n2055 | n6882;
assign n7563 = n3813 & n12744;
assign n4944 = ~(n10189 | n1777);
assign n9952 = ~n14011;
assign n6862 = n5493 | n2722;
assign n6338 = n7971 | n14423;
assign n9221 = n1538 | n6769;
assign n7932 = n10731 | n7361;
assign n767 = n12404 & n13157;
assign n4381 = n8147 & n9682;
assign n2538 = n1489 & n444;
assign n7414 = n6754 & n1244;
assign n10563 = n3445 | n4997;
assign n3223 = n4932 & n1052;
assign n12883 = n5948 & n7213;
assign n3023 = n10245 | n2634;
assign n2211 = n1821 | n6976;
assign n12891 = ~(n4270 | n1790);
assign n13613 = n6507 & n3425;
assign n12895 = n4102 & n11604;
assign n3522 = n5940 & n10429;
assign n13789 = n8980 | n9883;
assign n1005 = n5715 | n2777;
assign n8643 = ~(n31 | n9253);
assign n5799 = n11674 & n1296;
assign n10053 = n11620 | n6204;
assign n5393 = n1728 | n8587;
assign n7460 = n2820 & n5900;
assign n8887 = n9589 | n11404;
assign n8466 = ~(n7919 | n9150);
assign n915 = n1202 | n8919;
assign n6545 = n6316 & n4116;
assign n14006 = ~n4615;
assign n3995 = n12764 | n127;
assign n11733 = n4102 & n13019;
assign n12512 = n10457 & n10964;
assign n6959 = n7700 | n11053;
assign n13059 = n8714 | n11586;
assign n8042 = n6706 | n11370;
assign n3145 = ~(n3443 | n3581);
assign n9165 = n954 | n9515;
assign n3498 = n7779 & n3793;
assign n4044 = n13142 | n10616;
assign n7469 = n6486 & n5274;
assign n3832 = n1613 | n10027;
assign n9930 = n4690 & n14082;
assign n13003 = ~n11120;
assign n5733 = n10822 & n9561;
assign n3242 = n6147 & n685;
assign n4850 = n12741 & n13731;
assign n10194 = n286 & n2439;
assign n6419 = ~(n7375 | n5611);
assign n3405 = ~n1911;
assign n2654 = n6744 & n10474;
assign n10344 = ~(n11285 | n7555);
assign n6169 = n14466 | n8089;
assign n3854 = n3799 & n10776;
assign n390 = ~n10204;
assign n10089 = ~n6123;
assign n8969 = ~n1894;
assign n388 = n3586 & n4170;
assign n1728 = ~n2484;
assign n4948 = n4276 & n14148;
assign n3829 = n13367 & n9540;
assign n10008 = n6354 & n6814;
assign n3677 = ~(n12288 | n731);
assign n13606 = n3536 & n13928;
assign n4894 = n12391 | n8550;
assign n10075 = n12461 & n2737;
assign n7565 = n2878 | n6355;
assign n12384 = n4913 | n6231;
assign n1399 = n8386 & n8194;
assign n4256 = n4614 & n8039;
assign n13353 = ~(n1417 | n4730);
assign n885 = n5634 & n2524;
assign n5111 = n13083 | n13478;
assign n10445 = n11935 | n6152;
assign n11786 = n5732 | n8845;
assign n4364 = n2322 & n8772;
assign n12822 = n8372 & n13692;
assign n1745 = n8386 & n275;
assign n7107 = n5229 & n1134;
assign n9171 = n11329 & n2348;
assign n13396 = n13978 | n9649;
assign n8713 = n8747 | n5968;
assign n4086 = ~(n12568 | n5323);
assign n12385 = n8238 & n1396;
assign n8690 = n10857 | n9693;
assign n2872 = n1051 | n4706;
assign n1952 = n13535 & n8340;
assign n689 = n1031 | n8785;
assign n8574 = n8209 | n13688;
assign n9824 = ~n4050;
assign n4916 = ~(n8543 | n2483);
assign n6736 = ~(n9176 | n244);
assign n1369 = n8855 & n12094;
assign n13387 = ~(n8223 | n3413);
assign n1354 = ~n442;
assign n4917 = ~(n11584 | n4763);
assign n8998 = n5891 | n8128;
assign n9886 = n7057 & n7498;
assign n5429 = ~n13765;
assign n1866 = n3332 & n5776;
assign n2668 = n2445 & n13348;
assign n4639 = ~n7518;
assign n13897 = n8748 | n2376;
assign n1551 = n2465 & n35;
assign n5483 = ~n12249;
assign n13240 = ~n2744;
assign n1255 = ~n13154;
assign n9217 = n7481 | n1896;
assign n820 = ~n13901;
assign n12720 = n13078 & n353;
assign n6070 = ~(n8378 | n13377);
assign n8761 = n2961 & n11389;
assign n12556 = n4925 | n6056;
assign n12767 = n172 | n2059;
assign n953 = n9422 | n11081;
assign n9035 = ~n8595;
assign n1505 = n1414 & n12484;
assign n6950 = n14449 | n11649;
assign n1545 = n4117 & n9840;
assign n3211 = ~n4533;
assign n12239 = n12211 | n8522;
assign n3669 = n13016 | n6825;
assign n2513 = n12112 | n8621;
assign n8067 = n5088 & n10411;
assign n5881 = n9353 | n12845;
assign n1892 = n12712 | n3750;
assign n13610 = n7971 | n11560;
assign n12108 = n194 | n4552;
assign n5386 = n7670 & n1504;
assign n13802 = n7429 & n1523;
assign n12213 = n9140 | n13741;
assign n3519 = n5825 & n4762;
assign n8467 = ~(n9035 | n1869);
assign n422 = n791 | n12817;
assign n1557 = n6556 | n10736;
assign n1590 = n100 | n869;
assign n5602 = n5279 & n10860;
assign n12276 = n11142 & n8062;
assign n13510 = n838 | n10194;
assign n3650 = n3076 | n12359;
assign n8379 = n10134 & n2754;
assign n7555 = ~(n1218 | n3302);
assign n11129 = ~n2094;
assign n7268 = n13978 | n3695;
assign n12981 = n3120 | n4288;
assign n3225 = ~(n13310 | n6513);
assign n772 = ~n12323;
assign n2964 = n6607 | n6985;
assign n8880 = ~(n4195 | n12275);
assign n1234 = ~(n4988 | n6403);
assign n1038 = n3125 | n138;
assign n8455 = n1414 & n5740;
assign n2353 = n10084 & n6398;
assign n9343 = n13847 | n9279;
assign n2417 = ~n6451;
assign n10222 = n13626 & n8946;
assign n8909 = n9589 & n1196;
assign n1861 = n7997 & n7925;
assign n2955 = n7364 | n9283;
assign n4232 = n791 | n10116;
assign n14352 = ~(n10803 | n14019);
assign n10437 = n3942 & n6958;
assign n866 = n234 | n1439;
assign n3290 = ~n1312;
assign n13685 = n2089 | n11471;
assign n3074 = n11542 | n2285;
assign n8701 = ~n2484;
assign n8837 = n8881 | n7544;
assign n6786 = n11875 & n4247;
assign n3890 = ~(n12294 | n10002);
assign n2768 = ~(n8462 | n12454);
assign n6247 = n4104 & n3687;
assign n5927 = n12953 & n14189;
assign n2896 = n7011 | n8418;
assign n4336 = n6016 & n8675;
assign n6552 = n8983 | n5205;
assign n12972 = n412 | n10132;
assign n13291 = n12019 | n2582;
assign n2122 = ~(n4561 | n7879);
assign n11044 = ~(n13276 | n12539);
assign n12476 = n7812 | n10430;
assign n14424 = n7530 | n10986;
assign n12681 = ~(n11047 | n10390);
assign n6325 = ~(n9414 | n14236);
assign n5433 = n1804 & n3149;
assign n3638 = ~(n425 | n4301);
assign n1754 = n5825 & n4021;
assign n7155 = n2021 & n1211;
assign n8735 = n14016 & n4963;
assign n2220 = n1610 & n8973;
assign n13788 = n2445 & n4878;
assign n10944 = n11950 & n1856;
assign n8723 = n5695 | n6033;
assign n12619 = n5062 & n11386;
assign n9916 = n7284 & n1566;
assign n2124 = n3088 | n12381;
assign n11720 = n11097 | n4401;
assign n6547 = n492 | n12374;
assign n13767 = n4052 | n12059;
assign n13506 = n7803 | n3328;
assign n12967 = n12292 | n9030;
assign n274 = n12018 & n2553;
assign n5910 = n3099 | n743;
assign n9261 = n12428 | n9013;
assign n8813 = n692 & n8349;
assign n14386 = n5409 | n589;
assign n1953 = ~(n14370 | n11767);
assign n11569 = ~n11547;
assign n3906 = ~(n7364 | n14052);
assign n3513 = n13362 & n1828;
assign n5205 = n11142 & n10669;
assign n13937 = ~n11574;
assign n9432 = ~(n8197 | n6864);
assign n9280 = ~n10765;
assign n330 = ~(n10402 | n14070);
assign n8227 = n9972 & n3636;
assign n4796 = n11171 | n5422;
assign n4310 = n11621 | n8317;
assign n2687 = n2790 | n7093;
assign n9634 = ~(n9550 | n12111);
assign n1701 = ~n10775;
assign n12137 = n12023 | n3563;
assign n4575 = ~(n6672 | n12988);
assign n5052 = n13806 | n4513;
assign n4329 = n200 & n14509;
assign n4940 = n2272 | n13534;
assign n7094 = ~(n13050 | n10959);
assign n3624 = n8047 & n479;
assign n12462 = n10781 | n1456;
assign n3326 = n11422 & n3555;
assign n13250 = n5362 | n11349;
assign n12053 = n2783 & n8889;
assign n6692 = n4498 | n11645;
assign n13541 = n14260 & n3001;
assign n4459 = n5064 | n2167;
assign n5029 = n14200 | n9026;
assign n7211 = ~n2432;
assign n10633 = n7187 & n1737;
assign n3360 = n12449 & n6347;
assign n3679 = n9541 | n3407;
assign n13567 = n7419 & n8764;
assign n6685 = n7914 | n6597;
assign n2815 = n100 | n14441;
assign n2342 = n11572 | n12574;
assign n3974 = n8983 | n1288;
assign n8383 = n8452 | n4712;
assign n7324 = n13147 & n4625;
assign n13753 = ~(n9806 | n14297);
assign n11527 = n4205 | n12916;
assign n8626 = n10516 & n110;
assign n9449 = n4205 | n3291;
assign n11928 = ~(n8209 | n7160);
assign n13047 = n7618 & n1959;
assign n14518 = n9509 & n6662;
assign n2422 = ~n13447;
assign n7497 = n1189 | n7821;
assign n3091 = n5936 | n4569;
assign n12896 = n4033 | n9310;
assign n1751 = n776 & n12392;
assign n52 = n14038 & n2379;
assign n6090 = ~n12394;
assign n7384 = n10637 | n14344;
assign n264 = ~n9388;
assign n4169 = n6537 & n13858;
assign n9937 = n6206 | n13647;
assign n13795 = n14213 & n13256;
assign n256 = n6323 | n5027;
assign n1151 = n1431 & n3122;
assign n13719 = n3286 & n10049;
assign n1858 = ~(n13941 | n9820);
assign n12018 = ~n7621;
assign n7761 = n13464 & n14451;
assign n2963 = n7963 | n4147;
assign n11592 = n6654 | n13161;
assign n12470 = n2412 | n9259;
assign n13338 = ~n9865;
assign n1019 = ~(n1685 | n10065);
assign n11416 = n8630 & n8362;
assign n544 = n3097 & n13666;
assign n2548 = ~n3822;
assign n4432 = n7122 | n12514;
assign n11211 = n13359 & n12742;
assign n10412 = n3667 | n693;
assign n11392 = ~n13186;
assign n7040 = n14351 & n11907;
assign n6029 = n10854 & n3574;
assign n5074 = n11213 & n8314;
assign n7671 = n12020 | n11825;
assign n9348 = n7079 & n12080;
assign n6062 = ~n10897;
assign n9556 = n1202 | n5767;
assign n5451 = n194 | n6269;
assign n4626 = n2098 | n7164;
assign n6962 = n11839 | n1072;
assign n6770 = n4128 | n13493;
assign n10986 = n12521 & n8987;
assign n7951 = n2985 & n1135;
assign n2443 = ~(n6424 | n1055);
assign n2465 = ~n6905;
assign n5166 = n8721 & n6984;
assign n13392 = n5625 | n7374;
assign n2610 = ~(n13875 | n206);
assign n5460 = ~n834;
assign n2616 = n7852 & n1236;
assign n5755 = n8786 & n12221;
assign n13820 = n9571 & n9603;
assign n1674 = n6157 & n11521;
assign n11185 = n6013 & n5667;
assign n7039 = n5459 & n9438;
assign n7680 = n6830 & n3698;
assign n2984 = n12601 | n4943;
assign n4776 = n12821 | n8627;
assign n2012 = ~n12976;
assign n3161 = ~n9959;
assign n12067 = n11867 & n13618;
assign n13565 = n3401 & n12488;
assign n11754 = n10713 | n10145;
assign n11249 = n480 | n4198;
assign n11929 = ~(n4092 | n9207);
assign n6265 = n11093 & n7332;
assign n7672 = n10449 | n10553;
assign n5818 = n2367 & n9391;
assign n10643 = n6525 & n10435;
assign n8112 = ~n13109;
assign n2174 = n4741 | n10114;
assign n1461 = n8605 & n6815;
assign n7417 = n5240 & n7189;
assign n6011 = n3799 | n8746;
assign n6889 = ~(n600 | n2646);
assign n14205 = n9174 | n8988;
assign n7839 = n8304 | n2151;
assign n9621 = n12149 | n5060;
assign n3919 = n13755 & n5372;
assign n9074 = n11484 & n5993;
assign n935 = n12147 & n9247;
assign n7706 = n14366 | n9715;
assign n8124 = n9154 & n8991;
assign n11144 = n5434 & n9146;
assign n11548 = ~n11324;
assign n7539 = n8020 & n7303;
assign n6211 = ~n12086;
assign n4075 = n9269 | n2372;
assign n3709 = ~n6054;
assign n342 = n3546 | n10071;
assign n14388 = ~n11474;
assign n4571 = n1044 | n447;
assign n4809 = n11240 & n12237;
assign n1525 = n5587 | n232;
assign n6902 = n1678 & n3392;
assign n4898 = ~n10985;
assign n2007 = n687 & n7286;
assign n931 = ~n2355;
assign n14017 = ~(n5429 | n4409);
assign n9355 = n6957 & n7975;
assign n2771 = n12592 & n12554;
assign n7992 = n2564 & n2931;
assign n7864 = n12265 & n125;
assign n4091 = ~n8288;
assign n8410 = n986 & n5295;
assign n1951 = n10050 & n11088;
assign n6278 = ~(n10136 | n10041);
assign n11757 = ~(n4518 | n220);
assign n2307 = n9856 | n3522;
assign n10795 = n9403 | n2905;
assign n12649 = n10710 & n2793;
assign n3990 = ~(n8458 | n2990);
assign n11887 = n6629 | n8839;
assign n668 = n13362 & n4488;
assign n5851 = n13944 & n4183;
assign n11050 = ~(n9423 | n2010);
assign n4452 = n3394 | n6608;
assign n14089 = n7221 & n161;
assign n982 = n4619 & n12723;
assign n7623 = n11336 & n4073;
assign n3665 = n11510 | n10251;
assign n13558 = n13860 & n4452;
assign n9590 = ~(n10036 | n9309);
assign n9953 = ~n8650;
assign n13191 = n2784 | n2701;
assign n7845 = n9864 | n1237;
assign n2115 = ~(n4284 | n11916);
assign n8929 = ~(n1760 | n5208);
assign n11562 = ~(n48 | n3894);
assign n13091 = n815 | n10615;
assign n10487 = n8452 | n10070;
assign n7137 = n12149 | n1994;
assign n3556 = n6898 & n8687;
assign n3810 = n9191 & n4229;
assign n3365 = ~n1571;
assign n13829 = ~(n900 | n12706);
assign n235 = ~n11901;
assign n8242 = ~n7339;
assign n10939 = n2387 | n9958;
assign n4078 = n9297 & n8659;
assign n12449 = ~n8524;
assign n5342 = n1904 & n10146;
assign n9717 = n6873 & n1241;
assign n8720 = ~(n13327 | n9799);
assign n4521 = n428 & n1038;
assign n654 = n2533 & n9165;
assign n2785 = n11121 | n4920;
assign n5100 = ~(n163 | n8590);
assign n1850 = ~n4175;
assign n13647 = n7203 & n10543;
assign n5307 = n12445 & n2124;
assign n6544 = ~n2609;
assign n13806 = ~n7086;
assign n11374 = n4581 & n2887;
assign n6901 = n11909 | n7103;
assign n12731 = n12986 & n7449;
assign n12592 = ~n1724;
assign n13314 = n11300 & n12289;
assign n11000 = ~(n2780 | n12654);
assign n3122 = n648 | n4628;
assign n4803 = ~n9416;
assign n13574 = n8111 & n4460;
assign n1023 = ~n3054;
assign n10619 = ~n9543;
assign n7854 = n11636 & n5829;
assign n1131 = n766 | n2464;
assign n5229 = ~n9450;
assign n9891 = n8630 & n1570;
assign n4634 = ~n7200;
assign n92 = n4239 | n5802;
assign n5801 = n3724 & n5931;
assign n557 = n986 & n7078;
assign n2983 = ~n13734;
assign n7317 = n4244 & n1750;
assign n9975 = n7358 | n13649;
assign n13812 = n3923 & n9424;
assign n6468 = n11951 | n7385;
assign n13693 = n74 & n7669;
assign n13234 = n11066 & n4510;
assign n994 = n12324 | n1918;
assign n2532 = n4898 | n10437;
assign n8710 = n14110 | n7482;
assign n8648 = n7057 & n13886;
assign n12830 = n10781 | n13262;
assign n8764 = n77 | n2476;
assign n11222 = n8527 | n13322;
assign n3398 = n4045 | n1369;
assign n3013 = n13016 | n7199;
assign n1208 = n13806 | n4833;
assign n4053 = n7208 & n13150;
assign n1424 = n13875 | n12067;
assign n8705 = n6527 & n7396;
assign n5588 = n8965 & n4220;
assign n8348 = n5575 | n13782;
assign n4662 = n5053 & n8803;
assign n6294 = n5315 | n12778;
assign n11716 = n12019 | n7369;
assign n7110 = n1538 | n6626;
assign n13452 = n555 | n10744;
assign n8303 = n9297 & n4872;
assign n6389 = ~n5990;
assign n14129 = n1937 & n12393;
assign n12818 = n11420 | n2633;
assign n12508 = ~(n3944 | n2052);
assign n3605 = n200 & n11298;
assign n3664 = n820 | n4660;
assign n3456 = n11220 & n10126;
assign n2325 = n13781 & n2260;
assign n4537 = n2843 | n1364;
assign n1538 = ~n777;
assign n6537 = ~n3775;
assign n9912 = n387 | n9517;
assign n11783 = n6822 & n11229;
assign n11532 = n12858 & n7694;
assign n5212 = n2098 | n2749;
assign n4116 = n9429 | n14359;
assign n1387 = n12601 | n3157;
assign n5235 = n3536 & n13335;
assign n6483 = n5275 & n10993;
assign n11645 = n8025 & n11890;
assign n2564 = ~n12503;
assign n12761 = ~(n3165 | n4912);
assign n10703 = n6595 | n14482;
assign n14396 = n10072 & n7051;
assign n2917 = ~(n1914 | n2113);
assign n1597 = n2025 | n1624;
assign n5839 = ~n10837;
assign n6972 = ~(n7227 | n10938);
assign n8012 = n3011 | n11064;
assign n2922 = n7419 & n13691;
assign n4065 = ~n2934;
assign n255 = n1117 & n9072;
assign n7768 = ~n1955;
assign n8322 = n13252 & n1181;
assign n7624 = ~n13476;
assign n4572 = ~n11582;
assign n5124 = n6857 | n3883;
assign n12159 = ~n448;
assign n6781 = ~n3681;
assign n2428 = n12025 | n3673;
assign n7471 = n13404 & n847;
assign n5524 = n10357 & n9195;
assign n10267 = n8332 | n7960;
assign n11849 = n317 | n9576;
assign n2083 = n11093 & n10163;
assign n10252 = n1489 & n11137;
assign n11558 = ~n8813;
assign n2736 = n13860 & n8779;
assign n1388 = n6556 & n8795;
assign n4421 = n5762 | n12882;
assign n7963 = ~n6251;
assign n12365 = n2942 & n3903;
assign n6414 = n5997 | n12638;
assign n5309 = n7678 | n12570;
assign n6519 = ~n7086;
assign n12665 = n12802 & n9906;
assign n12289 = n3168 | n721;
assign n2939 = n225 & n9356;
assign n11284 = n2181 | n8308;
assign n5999 = ~n3361;
assign n617 = n8697 & n14094;
assign n4589 = ~n6855;
assign n2252 = n2908 | n2391;
assign n4720 = n7710 & n12886;
assign n9915 = n4357 | n2447;
assign n10385 = n4739 | n14469;
assign n11251 = ~n1932;
assign n1042 = ~(n11714 | n2611);
assign n4160 = n10302 & n9374;
assign n10213 = n9174 | n4643;
assign n3210 = ~n10314;
assign n9792 = ~n11158;
assign n13516 = ~n5242;
assign n13525 = ~n6787;
assign n3138 = n9289 | n13620;
assign n8505 = n11440 | n14265;
assign n592 = ~(n3132 | n2703);
assign n2199 = ~(n12968 | n8276);
assign n9718 = ~n13429;
assign n5186 = n5857 & n672;
assign n7116 = ~n2970;
assign n4513 = n3724 & n11957;
assign n1603 = n327 & n3152;
assign n5213 = n12542 & n13329;
assign n11755 = ~(n13324 | n10308);
assign n6063 = n4790 & n2966;
assign n7488 = n4233 | n9178;
assign n8915 = n5562 | n5474;
assign n10676 = n8769 & n8509;
assign n9386 = n12953 & n193;
assign n11945 = ~(n473 | n933);
assign n13720 = ~n6460;
assign n6738 = n2583 & n1491;
assign n8999 = ~(n1820 | n14352);
assign n2622 = n11470 & n5652;
assign n5916 = ~(n5919 | n9787);
assign n947 = n8877 | n3654;
assign n3400 = ~n13084;
assign n7074 = n2694 | n13152;
assign n11184 = ~(n1681 | n9205);
assign n571 = n1028 | n5970;
assign n503 = n4925 | n10366;
assign n9055 = n10351 | n10598;
assign n3323 = n4880 & n4640;
assign n8331 = n7678 | n1592;
assign n11584 = ~n12358;
assign n11262 = ~n9252;
assign n6779 = n1198 | n10007;
assign n4290 = n9226 | n9712;
assign n12079 = ~n513;
assign n12335 = ~n12970;
assign n584 = ~n11788;
assign n11572 = ~n7064;
assign n4941 = n7229 | n3721;
assign n14259 = n225 & n12690;
assign n6978 = n10384 & n5905;
assign n6892 = n10062 | n10093;
assign n3963 = ~(n9046 | n7714);
assign n3530 = ~n10012;
assign n3544 = n8376 & n2854;
assign n9135 = n7221 & n11974;
assign n12524 = n13854 | n8054;
assign n14427 = n5926 & n6633;
assign n882 = ~n3054;
assign n5829 = n4807 | n12150;
assign n3097 = ~n5613;
assign n9062 = n12445 & n12297;
assign n1410 = n10019 | n96;
assign n12712 = ~n7600;
assign n12622 = ~n11541;
assign n6528 = n1189 | n7733;
assign n5381 = n222 & n757;
assign n10983 = n12622 | n14037;
assign n5721 = n5409 | n6539;
assign n2228 = n7429 & n9001;
assign n14439 = n1711 | n4138;
assign n9331 = n6090 | n11758;
assign n2977 = n10019 | n11517;
assign n5416 = n5855 | n4907;
assign n12167 = ~n3833;
assign n6796 = n3093 | n8239;
assign n2711 = n329 | n7991;
assign n7760 = n5489 & n8886;
assign n1152 = ~n4769;
assign n4141 = n3569 | n19;
assign n10271 = ~(n6765 | n2323);
assign n11121 = ~n14412;
assign n107 = n6311 & n280;
assign n5843 = n9345 & n135;
assign n3005 = n4207 | n10869;
assign n279 = n10815 & n4038;
assign n3942 = ~n3440;
assign n8187 = n13016 | n10371;
assign n5708 = n12858 & n7114;
assign n790 = n2318 | n10941;
assign n4667 = n8034 | n10477;
assign n4578 = n11105 | n7232;
assign n5639 = n6288 | n1993;
assign n7024 = ~(n5919 | n3749);
assign n10981 = n1480 | n13494;
assign n13076 = n1962 & n7270;
assign n2113 = ~(n8856 | n3769);
assign n315 = n12475 & n11782;
assign n4790 = ~n9450;
assign n11108 = n1223 | n14440;
assign n10134 = ~n6139;
assign n3490 = n8015 | n12655;
assign n9401 = n231 & n12532;
assign n11090 = ~n10629;
assign n12001 = n11679 & n11725;
assign n9632 = n5434 & n4993;
assign n10559 = n10154 | n5515;
assign n10204 = n4533 & n2848;
assign n8803 = n1189 | n3962;
assign n10612 = n4435 | n8615;
assign n683 = n4394 & n10640;
assign n4822 = ~n9580;
assign n3281 = n2750 | n12656;
assign n13590 = n317 | n11074;
assign n13612 = n11935 | n12875;
assign n1074 = ~n1639;
assign n2177 = ~n12503;
assign n5538 = n14093 & n13254;
assign n9701 = ~(n11305 | n66);
assign n8751 = ~(n4233 | n7244);
assign n13803 = n5977 | n10013;
assign n4722 = ~n8451;
assign n11914 = n3320 | n5499;
assign n10263 = ~(n5986 | n6047);
assign n10171 = n14093 & n4635;
assign n4087 = n8209 | n2498;
assign n11356 = n2750 | n11639;
assign n14323 = n4180 | n14431;
assign n3486 = n9705 & n324;
assign n9184 = n12576 | n156;
assign n10621 = n10331 | n4053;
assign n4439 = ~n2069;
assign n2740 = n4033 | n12523;
assign n5975 = ~n5449;
assign n2466 = n11405 | n9999;
assign n12716 = n627 & n8408;
assign n1607 = n8412 & n13215;
assign n13797 = n234 | n9667;
assign n3274 = n4546 & n7425;
assign n10202 = n8986 | n4732;
assign n13265 = ~(n11765 | n11054);
assign n707 = n6130 & n7366;
assign n9380 = ~(n10312 | n6284);
assign n8770 = n14091 & n3358;
assign n2669 = ~n6829;
assign n2566 = ~n13983;
assign n11732 = ~(n13324 | n8072);
assign n243 = n1660 | n7102;
assign n13935 = n11360 | n9624;
assign n6576 = n390 | n8356;
assign n4778 = n14088 | n10361;
assign n3288 = n1258 | n10605;
assign n7898 = ~n13696;
assign n1981 = n11303 | n601;
assign n7276 = n12250 & n14159;
assign n1284 = n14282 | n2751;
assign n12520 = n11838 & n6934;
assign n2685 = n6288 | n5609;
assign n5339 = ~(n11285 | n10109);
assign n6279 = ~(n2017 | n14017);
assign n5714 = ~(n194 | n11184);
assign n6632 = n8172 | n12734;
assign n10512 = ~n10912;
assign n7586 = n7736 | n579;
assign n13177 = n1669 | n9699;
assign n12027 = n9275 & n6970;
assign n7649 = n4741 | n8110;
assign n13195 = n7997 | n6517;
assign n10521 = n10015 & n8187;
assign n9652 = ~(n329 | n8902);
assign n12892 = n541 & n12173;
assign n11952 = n13675 | n3488;
assign n10405 = n11867 & n13736;
assign n1464 = n13252 & n9691;
assign n12607 = n6527 & n2767;
assign n8230 = n1535 | n13251;
assign n6 = ~(n6953 | n12456);
assign n9557 = ~n13784;
assign n12326 = n4790 & n3238;
assign n7188 = ~n12397;
assign n3346 = n9211 | n916;
assign n2355 = n3910 | n5467;
assign n2150 = ~(n14466 | n8186);
assign n4140 = n11459 | n1305;
assign n11937 = n13718 | n12333;
assign n2111 = ~n7441;
assign n5288 = ~n13593;
assign n1724 = ~n4595;
assign n2991 = n1261 | n3426;
assign n346 = n4468 | n4381;
assign n3195 = n2564 & n6575;
assign n6951 = n12712 | n12140;
assign n8161 = n2669 & n6594;
assign n8661 = n930 | n13583;
assign n14074 = ~n10446;
assign n1826 = n11542 | n12648;
assign n9373 = n9819 & n8309;
assign n7545 = n10136 | n13768;
assign n8559 = n13484 & n12372;
assign n7844 = n9952 & n11391;
assign n5488 = ~n10282;
assign n10462 = ~(n11680 | n1399);
assign n3984 = n12400 | n10074;
assign n9194 = n14401 | n6068;
assign n11253 = n7736 | n7864;
assign n14157 = ~n9197;
assign n11836 = n839 | n3496;
assign n4291 = n13078 & n861;
assign n14487 = n14042 & n7083;
assign n615 = n5315 | n13909;
assign n14164 = n2080 | n10278;
assign n8886 = n820 | n8705;
assign n2860 = n13520 & n6757;
assign n14249 = ~n14303;
assign n4094 = n12412 & n5984;
assign n568 = ~n3007;
assign n12558 = n14337 | n11905;
assign n4649 = n6711 | n3297;
assign n1287 = n12542 & n922;
assign n8596 = n13641 & n1394;
assign n11833 = n9564 & n2410;
assign n638 = ~n1843;
assign n12396 = ~(n163 | n8612);
assign n28 = ~n4203;
assign n10310 = ~n3655;
assign n1067 = n2229 | n2101;
assign n1558 = n6318 & n14242;
assign n1267 = n8500 & n13752;
assign n9123 = n9191 & n13483;
assign n11081 = n873 & n10158;
assign n5452 = n9218 | n8494;
assign n12738 = n13017 | n5185;
assign n13926 = n12633 | n2517;
assign n7904 = n8800 | n203;
assign n9189 = n3485 & n7274;
assign n14393 = n4095 & n6956;
assign n825 = n2694 | n2351;
assign n6151 = n13464 & n243;
assign n655 = n3097 & n10246;
assign n6126 = n4018 & n6912;
assign n2489 = n4544 | n3198;
assign n3587 = ~n2405;
assign n7612 = ~n4131;
assign n7498 = n10834 | n5146;
assign n6890 = n8881 | n9636;
assign n12367 = n12229 & n3869;
assign n1994 = n2422 & n5397;
assign n6656 = n12038 & n2602;
assign n7822 = n12303 | n8262;
assign n71 = n5483 | n11934;
assign n12247 = n14466 | n6395;
assign n3924 = ~(n7683 | n12451);
assign n900 = ~n426;
assign n12612 = ~(n3255 | n7386);
assign n8788 = n12428 | n9426;
assign n14064 = n2158 & n10667;
assign n14468 = n12986 & n4956;
assign n2695 = ~(n12292 | n7709);
assign n5889 = n13516 | n12577;
assign n13017 = ~n7988;
assign n8473 = ~(n11492 | n3771);
assign n7481 = ~n9453;
assign n4345 = n2615 & n5893;
assign n1535 = ~n9580;
assign n2250 = n1136 & n6298;
assign n559 = n3093 | n13133;
assign n1934 = n1728 | n1310;
assign n12925 = n673 & n13371;
assign n13012 = n1332 | n11269;
assign n5552 = n13485 | n4511;
assign n9970 = n7418 | n10370;
assign n10312 = ~n2451;
assign n6931 = n11503 & n3955;
assign n4625 = n10637 | n9133;
assign n9849 = n1576 | n4427;
assign n13503 = n4095 & n5979;
assign n1174 = ~(n13522 | n6094);
assign n8342 = n5279 & n9638;
assign n5612 = n5048 & n2282;
assign n14385 = ~(n10620 | n6416);
assign n13782 = n11484 & n6510;
assign n6512 = ~(n13759 | n4096);
assign n3949 = n14481 | n5281;
assign n8906 = n12445 & n1230;
assign n1706 = n13102 | n7354;
assign n5295 = n14188 | n8436;
assign n3508 = n4913 | n11191;
assign n1798 = ~(n5848 | n10737);
assign n2845 = ~n12614;
assign n4585 = n6486 & n1598;
assign n10272 = n13823 & n3137;
assign n4555 = n6957 & n307;
assign n12293 = n4614 & n10237;
assign n791 = ~n10985;
assign n508 = n85 | n9469;
assign n2742 = ~n316;
assign n8113 = n7779 & n9597;
assign n3270 = n13155 | n1511;
assign n11545 = n8582 | n1123;
assign n12699 = n3424 & n13039;
assign n9698 = n5834 | n2106;
assign n2992 = n6471 | n7186;
assign n2314 = ~(n7052 | n2795);
assign n1840 = ~n1041;
assign n13249 = ~(n584 | n4663);
assign n2190 = n7673 & n2274;
assign n11509 = n13501 | n6795;
assign n9578 = n12412 & n5473;
assign n11675 = n7767 & n9713;
assign n12227 = n5132 | n686;
assign n6788 = ~n6254;
assign n9603 = n4357 | n1907;
assign n8656 = ~n11195;
assign n11147 = ~(n8529 | n6966);
assign n12366 = n6629 | n4982;
assign n2366 = n8480 | n5031;
assign n3765 = n10238 | n10750;
assign n5954 = n10383 | n6336;
assign n4088 = n13952 & n10748;
assign n7318 = n1136 | n3799;
assign n12179 = ~n5416;
assign n5780 = ~n2369;
assign n13835 = ~n12096;
assign n1662 = ~n14525;
assign n2856 = ~(n12040 | n8677);
assign n7704 = ~n11870;
assign n3154 = n12015 & n4816;
assign n5292 = n9509 & n13917;
assign n4388 = n2908 | n5588;
assign n215 = n13359 & n715;
assign n4655 = ~n14525;
assign n1117 = ~n9450;
assign n3626 = n5236 | n4853;
assign n10107 = n2669 & n10761;
assign n13597 = ~n1769;
assign n4870 = n13421 & n2818;
assign n13204 = n10461 | n2675;
assign n8038 = n11620 | n10230;
assign n9716 = ~n13668;
assign n1186 = n7438 | n10882;
assign n7938 = ~n8892;
assign n155 = n2669 & n7166;
assign n13145 = ~(n6041 | n6246);
assign n11388 = n3435 & n5673;
assign n12147 = ~n9950;
assign n8675 = n5472 | n7062;
assign n1318 = n13575 & n5320;
assign n1941 = n7043 & n12884;
assign n8567 = n9931 | n2361;
assign n13236 = ~n8122;
assign n12451 = ~(n1127 | n13753);
assign n13760 = n9921 & n2443;
assign n420 = n13485 | n3547;
assign n11818 = n11901 | n6011;
assign n7115 = n12336 | n12782;
assign n9957 = n2843 | n2693;
assign n8750 = n1210 & n13912;
assign n13779 = ~n10368;
assign n13239 = n10781 | n495;
assign n7862 = ~n13901;
assign n9418 = n2527 & n3045;
assign n5880 = n14091 & n11059;
assign n3143 = n8692 & n8470;
assign n7609 = ~n8349;
assign n11479 = ~n8800;
assign n5730 = n1520 & n5135;
assign n9360 = n14401 | n12784;
assign n11643 = n28 | n8328;
assign n11321 = n4684 | n11648;
assign n10130 = n11704 | n4658;
assign n9644 = n1339 & n6925;
assign n13891 = n3607 & n14291;
assign n2181 = ~n1220;
assign n11428 = ~n5257;
assign n10015 = ~n10975;
assign n10800 = n5823 & n1175;
assign n9044 = n9442 | n5850;
assign n3284 = n11793 & n6638;
assign n14215 = n10969 & n9392;
assign n5513 = ~(n13365 | n8407);
assign n1307 = n3675 & n11146;
assign n7846 = n9654 | n8204;
assign n10319 = n5779 & n4969;
assign n9596 = n8814 & n9718;
assign n8171 = n13142 | n4235;
assign n14188 = ~n7404;
assign n964 = ~(n5897 | n13505);
assign n1504 = n13698 | n10463;
assign n10124 = n965 & n338;
assign n4787 = n9140 | n14087;
assign n8622 = n4614 & n3216;
assign n1000 = n13518 | n12511;
assign n11867 = ~n9613;
assign n11677 = n9972 & n11787;
assign n9482 = ~(n13835 | n13569);
assign n10815 = ~n14501;
assign n9901 = ~(n7575 | n2881);
assign n2155 = n3800 | n3459;
assign n4637 = ~n2470;
assign n11621 = ~n7289;
assign n12652 = n1356 | n9139;
assign n6064 = n4791 | n10867;
assign n10562 = ~n9592;
assign n123 = ~(n5486 | n11798);
assign n9873 = n6486 & n697;
assign n9760 = n5459 & n9549;
assign n11570 = n2401 | n5874;
assign n13433 = ~n11425;
assign n7444 = ~(n6428 | n7801);
assign n13136 = n13885 | n197;
assign n9743 = ~n11511;
assign n3116 = n8768 & n9833;
assign n5251 = n1071 & n14383;
assign n241 = n10760 & n14057;
assign n4467 = n4657 & n7096;
assign n410 = n5234 | n1600;
assign n6956 = n11094 | n3323;
assign n9600 = n2709 & n8949;
assign n5673 = n5266 | n11865;
assign n2335 = n11121 | n13331;
assign n11549 = n7700 | n11266;
assign n5253 = ~n3007;
assign n11186 = n4684 | n1459;
assign n8108 = n12531 & n10445;
assign n11219 = n5092 & n2453;
assign n479 = n10394 | n5235;
assign n1765 = n3709 & n8319;
assign n7446 = n10731 | n8739;
assign n2556 = n8799 & n7638;
assign n10250 = n2510 | n12621;
assign n10058 = n11739 | n5884;
assign n12412 = ~n12403;
assign n761 = n3871 | n6738;
assign n9012 = n1223 | n2716;
assign n12199 = n13718 | n2860;
assign n13946 = n1125 & n5923;
assign n7428 = n4840 | n6577;
assign n270 = n4828 | n3470;
assign n7837 = n1729 & n12205;
assign n6337 = n14430 | n3048;
assign n3029 = n8630 & n217;
assign n12378 = n10032 & n12081;
assign n5180 = ~n8813;
assign n12178 = n478 | n3556;
assign n7339 = n5218 & n7689;
assign n5152 = n8605 & n546;
assign n6005 = n8277 | n11986;
assign n1699 = ~n4824;
assign n6715 = ~(n2822 | n6217);
assign n4960 = ~(n8209 | n2811);
assign n4786 = n6640 | n5601;
assign n3165 = ~n5734;
assign n1974 = n1834 | n7926;
assign n8730 = ~(n13327 | n11046);
assign n2914 = n10622 & n3060;
assign n8651 = n3777 | n4069;
assign n158 = n873 & n4749;
assign n9133 = n2527 & n1420;
assign n13312 = n8527 | n265;
assign n3121 = n7187 & n8339;
assign n12680 = n12821 | n11858;
assign n10047 = n320 & n115;
assign n7113 = n14449 | n8606;
assign n3267 = n5335 & n14195;
assign n93 = ~n12872;
assign n11405 = ~n4606;
assign n5198 = n10089 | n2452;
assign n13383 = ~n4835;
assign n6884 = n13718 | n13480;
assign n8444 = n10516 & n14514;
assign n9845 = n12445 & n3659;
assign n4123 = ~n6999;
assign n881 = n6527 & n10364;
assign n14450 = ~n11930;
assign n3485 = ~n7275;
assign n5174 = n6753 & n7001;
assign n11510 = ~n8595;
assign n13280 = n13413 | n3438;
assign n5232 = n8210 | n3981;
assign n12944 = n5315 | n1087;
assign n2972 = n12445 & n6026;
assign n12808 = ~n1347;
assign n11552 = n5434 & n11399;
assign n6179 = n4498 | n13099;
assign n8979 = n103 & n7585;
assign n4413 = n9953 & n5677;
assign n8716 = n4156 & n4071;
assign n13742 = n1356 | n4551;
assign n2897 = ~n11456;
assign n5750 = n11607 & n4710;
assign n4561 = n10615 | n9830;
assign n1642 = n1138 & n5379;
assign n4690 = ~n13447;
assign n758 = n9232 & n9814;
assign n8842 = n10083 | n713;
assign n5119 = n2521 & n6059;
assign n6934 = n8034 | n4478;
assign n7776 = n791 | n5190;
assign n8275 = n6013 & n1829;
assign n5093 = n9375 | n9772;
assign n2045 = n12521 & n8026;
assign n11258 = n10516 & n6259;
assign n10955 = n116 | n1352;
assign n618 = ~(n3394 | n9092);
assign n604 = n5275 & n1803;
assign n7433 = ~n13890;
assign n12325 = n2897 | n2927;
assign n3526 = ~n1784;
assign n769 = ~n1966;
assign n11084 = n9375 | n13929;
assign n4012 = n13080 | n10405;
assign n11391 = n5007 | n5213;
assign n13458 = ~n14406;
assign n11054 = ~(n5271 | n11190);
assign n2255 = ~(n955 | n7514);
assign n679 = ~n9314;
assign n8615 = n10668 & n7468;
assign n53 = n4887 & n2505;
assign n6676 = n5493 | n5448;
assign n10449 = ~n1214;
assign n11904 = n13083 | n6991;
assign n451 = n11842 & n8518;
assign n9083 = n11935 | n3035;
assign n4843 = n5475 & n2279;
assign n606 = ~(n11581 | n5015);
assign n6827 = n480 | n13271;
assign n7306 = n6606 & n3106;
assign n7487 = n3923 & n3095;
assign n6320 = n3766 & n4254;
assign n7758 = n673 | n11875;
assign n13054 = n9102 & n12384;
assign n7622 = n5825 & n12552;
assign n12826 = ~(n7662 | n1337);
assign n5804 = n13112 | n4263;
assign n7061 = n6192 & n12519;
assign n11539 = n9571 & n10954;
assign n3179 = n1662 & n9607;
assign n5599 = ~(n2405 | n4471);
assign n9608 = n14521 & n13989;
assign n7146 = ~n3493;
assign n1096 = n1821 | n2796;
assign n3411 = n5507 | n3511;
assign n8728 = n3286 & n10955;
assign n4913 = ~n13165;
assign n6536 = n2505 | n12009;
assign n6077 = n12428 | n3520;
assign n329 = ~n5974;
assign n5638 = n12421 & n6080;
assign n3518 = n12147 & n11913;
assign n9563 = ~n4169;
assign n4450 = n14358 & n6892;
assign n6851 = n15 & n4083;
assign n9285 = ~n1833;
assign n532 = ~(n4210 | n6723);
assign n8285 = n4233 | n3831;
assign n13491 = n12353 | n5845;
assign n4200 = ~n3094;
assign n9565 = n1117 & n7839;
assign n12429 = n14088 | n10531;
assign n262 = n9780 | n10103;
assign n10505 = n9806 | n10022;
assign n2805 = n4739 | n7299;
assign n8268 = n2758 & n6968;
assign n1842 = n13367 & n10572;
assign n2762 = n8047 & n6718;
assign n2650 = n1854 & n13686;
assign n9822 = n2521 & n9061;
assign n3032 = ~(n12292 | n9590);
assign n719 = n8432 & n7037;
assign n9731 = n12695 | n5610;
assign n11442 = n12857 & n3646;
assign n1471 = n6607 | n793;
assign n3688 = n2272 | n2239;
assign n5772 = n5825 & n13071;
assign n2527 = ~n9583;
assign n4341 = n177 | n13295;
assign n1083 = n8432 & n10621;
assign n12334 = ~n9329;
assign n13082 = n3888 | n5500;
assign n9406 = n13682 & n2002;
assign n8492 = n412 | n10176;
assign n12260 = n1937 & n12342;
assign n3934 = ~(n1425 | n1283);
assign n3404 = n6867 | n5772;
assign n445 = n2527 & n3005;
assign n8947 = n3724 & n925;
assign n8940 = n13531 | n8579;
assign n12269 = ~(n8592 | n2234);
assign n11469 = ~(n1628 | n4756);
assign n4711 = ~n355;
assign n8592 = ~n81;
assign n3631 = n638 & n8681;
assign n6296 = n12953 & n11318;
assign n1999 = n14337 | n10762;
assign n10054 = n13547 | n1764;
assign n580 = ~(n14377 | n6158);
assign n1230 = n11223 | n12600;
assign n13954 = n2111 | n7248;
assign n12028 = ~(n619 | n2195);
assign n3907 = ~n9778;
assign n1291 = n1074 & n6481;
assign n5836 = n7438 | n4111;
assign n1917 = n9422 | n7508;
assign n11685 = n9853 & n12763;
assign n14437 = n11329 & n8609;
assign n12790 = ~(n11455 | n10222);
assign n9836 = n4876 | n2397;
assign n12902 = n4354 & n519;
assign n2075 = n12592 & n12206;
assign n14406 = n13728 & n6482;
assign n10610 = n6609 & n12510;
assign n5603 = ~n12106;
assign n2286 = n6263 | n13568;
assign n7063 = ~n6807;
assign n12990 = ~n14501;
assign n11546 = ~n7455;
assign n4661 = n9323 & n7489;
assign n8586 = ~(n4978 | n5635);
assign n7296 = n13860 & n8059;
assign n9978 = n2843 | n12634;
assign n5298 = n163 | n1642;
assign n3754 = n2486 & n6908;
assign n10726 = n8247 & n11234;
assign n13351 = n11422 & n3892;
assign n12532 = n7481 | n3416;
assign n9881 = n1857 & n12222;
assign n10671 = n4468 | n7647;
assign n11178 = n8401 & n4905;
assign n5631 = n7171 & n9017;
assign n7694 = n5562 | n9401;
assign n5558 = ~n1985;
assign n7771 = n1763 & n2488;
assign n2606 = n8452 | n13001;
assign n2529 = ~n6873;
assign n4284 = ~n8027;
assign n9330 = n10367 & n10076;
assign n561 = n555 | n2353;
assign n4753 = n79 & n2471;
assign n3551 = n2006 & n12469;
assign n4801 = n2089 | n4584;
assign n5769 = n747 | n972;
assign n6750 = n9111 | n9951;
assign n2783 = ~n10303;
assign n3001 = n1006 | n8293;
assign n10196 = n15 & n5793;
assign n4007 = ~n12765;
assign n5611 = ~(n5762 | n11791);
assign n14067 = n116 | n4812;
assign n5427 = ~n4169;
assign n6755 = n10922 & n5706;
assign n8747 = ~n2320;
assign n2930 = n7826 & n8658;
assign n7861 = n4065 | n6627;
assign n3173 = n7768 & n11394;
assign n14197 = n7481 | n9386;
assign n8058 = ~(n700 | n1793);
assign n13924 = ~(n1929 | n8459);
assign n7581 = n8692 & n3342;
assign n5790 = n11020 & n9934;
assign n11360 = ~n13668;
assign n1085 = n13978 | n10138;
assign n14 = n1904 & n2200;
assign n7659 = n5857 & n11128;
assign n3723 = n13656 & n1131;
assign n10820 = ~n11548;
assign n627 = ~n5182;
assign n1517 = n4574 & n13403;
assign n12489 = n9156 & n3583;
assign n2788 = n11328 | n3532;
assign n14092 = n49 | n664;
assign n12405 = n3365 & n2974;
assign n11128 = n283 | n3447;
assign n13514 = n7063 & n12070;
assign n9008 = ~n13509;
assign n12962 = n1741 | n7470;
assign n12579 = n553 | n439;
assign n11606 = n4123 & n848;
assign n10574 = n12131 | n11960;
assign n12379 = n3569 | n13029;
assign n14000 = n808 & n5680;
assign n1299 = ~n5595;
assign n10400 = ~n12925;
assign n3076 = ~n13234;
assign n2913 = n14327 & n13935;
assign n9686 = n9329 & n14312;
assign n12315 = ~(n1086 | n10565);
assign n8100 = n6603 | n11714;
assign n6665 = n6389 & n5554;
assign n2612 = n8801 & n12415;
assign n8024 = n9321 & n2800;
assign n11384 = ~n2166;
assign n14270 = n12057 & n8914;
assign n11109 = n1339 & n10946;
assign n11074 = n11240 & n3194;
assign n1241 = ~(n13467 | n4237);
assign n5635 = ~(n4135 | n1321);
assign n12751 = n7068 & n8385;
assign n12266 = n11438 | n2852;
assign n5531 = n12226 & n8142;
assign n10105 = n12265 & n6337;
assign n3971 = ~(n13811 | n9170);
assign n14502 = n7957 & n5068;
assign n8418 = n4018 & n12213;
assign n1012 = ~(n4050 | n11418);
assign n14152 = n769 | n2770;
assign n5146 = n4095 & n418;
assign n1135 = n2179 | n9706;
assign n3693 = n10933 | n8716;
assign n2046 = n8582 | n11613;
assign n11400 = n1339 & n8338;
assign n13094 = n10383 | n5152;
assign n2852 = n3635 & n11594;
assign n9193 = n12808 & n5183;
assign n5764 = ~n304;
assign n10502 = n5038 & n6425;
assign n8489 = n14370 | n7844;
assign n11149 = n782 | n10654;
assign n5532 = n6838 & n12642;
assign n6128 = ~n261;
assign n13591 = n6192 & n10261;
assign n6768 = ~n2503;
assign n6358 = ~(n1697 | n964);
assign n9819 = ~n10862;
assign n13415 = n12636 | n7667;
assign n9939 = n7081 & n11777;
assign n2096 = n7530 | n5231;
assign n5716 = n1391 | n564;
assign n9509 = ~n2906;
assign n2441 = n14481 | n10753;
assign n11678 = ~(n4741 | n4109);
assign n4771 = ~n2370;
assign n4746 = n5362 | n10582;
assign n3946 = n12933 & n13466;
assign n10841 = n11171 | n14003;
assign n4949 = n5591 | n13186;
assign n2161 = n13516 | n1324;
assign n9262 = n7462 | n12815;
assign n11319 = n9442 | n5194;
assign n14269 = n1125 & n5967;
assign n9203 = ~(n7036 | n11);
assign n6033 = n13246 & n4483;
assign n11523 = n1100 & n402;
assign n2690 = ~(n4865 | n13416);
assign n13321 = n11123 | n4361;
assign n8685 = n11739 | n12795;
assign n11738 = ~n9936;
assign n12051 = n12131 | n12058;
assign n5025 = n13220 | n9101;
assign n1360 = n9111 | n4577;
assign n12711 = n5628 & n1974;
assign n12668 = n4180 | n7319;
assign n869 = n12953 & n11241;
assign n9575 = n1258 | n10918;
assign n11625 = n4807 | n5711;
assign n9947 = n7081 & n8553;
assign n12789 = n13103 & n12485;
assign n505 = n2983 & n248;
assign n318 = n5071 & n14147;
assign n4080 = n13107 & n5662;
assign n12499 = n10396 | n12871;
assign n10830 = n673 & n63;
assign n6575 = n4205 | n8113;
assign n10761 = n2318 | n770;
assign n13999 = n3608 & n14076;
assign n888 = ~n12573;
assign n2460 = n10556 & n9393;
assign n13221 = n6389 & n9202;
assign n6252 = n13446 | n7630;
assign n5574 = ~n462;
assign n12621 = n2564 & n13902;
assign n2795 = ~(n3230 | n5166);
assign n4243 = n541 & n13263;
assign n5622 = n10678 & n13120;
assign n12109 = n8983 | n8715;
assign n11631 = n14213 & n2487;
assign n4802 = n11303 | n5783;
assign n5340 = n1678 & n6338;
assign n7067 = n8969 | n10799;
assign n5321 = n1409 | n271;
assign n9352 = ~(n1417 | n2030);
assign n1205 = n89 | n4996;
assign n1986 = n4357 | n1842;
assign n5230 = n6090 | n5880;
assign n11393 = n7748 & n9595;
assign n11932 = n11090 | n802;
assign n8384 = n3134 | n11361;
assign n4014 = n13555 & n3057;
assign n6748 = n10084 & n170;
assign n5066 = n9211 | n9501;
assign n1501 = ~(n8337 | n4687);
assign n1338 = ~(n5504 | n6199);
assign n3159 = n13781 & n12481;
assign n5823 = ~n3926;
assign n6850 = n7208 & n465;
assign n1636 = n2330 & n8313;
assign n9339 = n7245 | n4854;
assign n2118 = ~(n6888 | n13406);
assign n358 = n5587 | n14214;
assign n9934 = n11097 | n796;
assign n2313 = n5053 & n2976;
assign n361 = ~n4606;
assign n3139 = ~(n5621 | n4797);
assign n4795 = ~(n600 | n2554);
assign n143 = n13875 | n13513;
assign n1457 = n5936 | n5733;
assign n9024 = n9952 & n2155;
assign n9163 = n1202 | n13600;
assign n8223 = ~n8224;
assign n6152 = n3710 & n1239;
assign n14490 = n11814 & n4733;
assign n2554 = ~(n7887 | n4718);
assign n8950 = ~n13908;
assign n8420 = ~(n1577 | n4196);
assign n10588 = ~(n4333 | n13709);
assign n14172 = n13877 & n14113;
assign n2462 = n2615 | n8737;
assign n9525 = ~n6928;
assign n4367 = n3273 | n1183;
assign n7162 = n1125 & n6484;
assign n5875 = n6672 | n6145;
assign n7873 = n1494 | n4115;
assign n1509 = ~(n4091 | n4458);
assign n12112 = ~n11331;
assign n1540 = n428 & n2047;
assign n1428 = ~n5153;
assign n2743 = n7670 & n10773;
assign n4965 = n1112 | n11235;
assign n10468 = n13745 & n2542;
assign n5626 = ~(n12651 | n4383);
assign n10790 = n10871 | n9109;
assign n9345 = ~n10469;
assign n11005 = n14145 & n5533;
assign n9377 = ~n2468;
assign n8059 = n11097 | n12011;
assign n5879 = ~(n13050 | n10878);
assign n8008 = ~n12675;
assign n14165 = n3536 & n3585;
assign n4136 = n1772 & n10701;
assign n4058 = n8301 | n11764;
assign n6104 = n14166 | n3408;
assign n7490 = n1623 | n8395;
assign n4174 = ~n10714;
assign n6546 = n14376 & n2537;
assign n7504 = n1061 | n3834;
assign n10949 = n10815 & n10866;
assign n11900 = n5137 & n14115;
assign n2051 = n8980 | n4403;
assign n7617 = ~(n478 | n9862);
assign n9748 = n9885 & n2304;
assign n4469 = n11814 & n10188;
assign n2980 = n6711 | n8535;
assign n9072 = n5234 | n6472;
assign n7244 = ~(n10368 | n9586);
assign n4277 = n10408 & n13510;
assign n10350 = n9429 | n2414;
assign n425 = ~n692;
assign n11559 = n1904 & n13940;
assign n681 = ~(n2241 | n3171);
assign n11173 = n3120 | n6900;
assign n6019 = n9571 & n9002;
assign n13962 = n6373 | n1291;
assign n1596 = n5977 | n3612;
assign n5520 = n627 & n9759;
assign n12616 = n5625 | n4641;
assign n8498 = n2474 | n11158;
assign n5380 = n6206 | n6015;
assign n13697 = n1588 & n11378;
assign n3785 = ~n10368;
assign n10826 = n9113 & n1691;
assign n10011 = n1356 | n1731;
assign n12066 = n8378 | n1106;
assign n10816 = n9078 | n12987;
assign n4691 = n9650 & n7633;
assign n9392 = n10035 | n9071;
assign n484 = n10062 | n9641;
assign n752 = n7433 | n6258;
assign n4476 = n11572 | n14504;
assign n276 = n7826 & n6688;
assign n3838 = n13074 | n4184;
assign n11060 = n7391 & n5273;
assign n10797 = n13078 & n420;
assign n7340 = ~(n9525 | n9138);
assign n169 = n6891 | n4410;
assign n108 = n4156 & n11836;
assign n10163 = n5468 | n1162;
assign n1601 = n1804 & n3042;
assign n13046 = n11702 & n13705;
assign n328 = n6316 & n7416;
assign n8682 = n9654 & n11479;
assign n12879 = ~(n1575 | n454);
assign n5216 = ~(n2087 | n6444);
assign n1631 = n8726 | n12417;
assign n7729 = n6525 & n9441;
assign n10523 = ~n7289;
assign n7994 = n627 & n2691;
assign n11993 = ~(n1914 | n14044);
assign n11370 = n13641 & n7228;
assign n1187 = n12543 | n12219;
assign n3779 = ~(n1742 | n11929);
assign n9853 = ~n8650;
assign n344 = ~(n13981 | n5041);
assign n1943 = n13877 & n4860;
assign n8009 = n5918 & n9574;
assign n3880 = n8789 & n13386;
assign n9861 = n4562 | n13495;
assign n8497 = n4346 & n12893;
assign n14362 = ~(n3333 | n4524);
assign n14409 = n8747 | n10661;
assign n13961 = n2422 & n7410;
assign n12113 = n5926 & n562;
assign n672 = n5815 | n13225;
assign n8807 = n2531 | n2705;
assign n12268 = ~(n14524 | n3225);
assign n13262 = n8358 & n8741;
assign n12882 = n10134 & n4372;
assign n6395 = ~(n13081 | n3702);
assign n1926 = n8726 | n8166;
assign n1716 = n14321 & n11742;
assign n11106 = n13676 & n10991;
assign n1116 = n13220 | n10478;
assign n6659 = n7079 & n9428;
assign n10508 = n8580 | n12823;
assign n13640 = ~(n1638 | n11993);
assign n1212 = n5454 | n3961;
assign n12169 = ~n11055;
assign n2641 = n11614 & n10951;
assign n11782 = n1838 | n3859;
assign n6904 = n4967 | n11466;
assign n8974 = n11008 & n1271;
assign n12486 = n13991 | n13533;
assign n12611 = ~n6807;
assign n12350 = n5450 | n11635;
assign n3654 = n11702 & n3727;
assign n12715 = n10247 & n8489;
assign n3596 = n11953 | n9145;
assign n9767 = n6838 & n6112;
assign n7486 = n9953 & n14363;
assign n14309 = n2378 & n10559;
assign n3463 = n8638 | n13609;
assign n4565 = n12229 & n3615;
assign n917 = n28 | n7642;
assign n12181 = n889 & n12562;
assign n8553 = n12400 | n5085;
assign n5740 = n13083 | n9642;
assign n6242 = ~n10346;
assign n84 = n7673 & n11431;
assign n8214 = ~(n727 | n5116);
assign n5744 = n7957 & n3228;
assign n2240 = n678 & n12898;
assign n11761 = ~n14118;
assign n7835 = n865 & n14217;
assign n11157 = ~n8963;
assign n196 = n14120 & n10291;
assign n11183 = ~n12331;
assign n11689 = n9198 & n5808;
assign n1111 = ~(n7091 | n7954);
assign n2399 = n12821 | n5708;
assign n5202 = n5139 | n2588;
assign n2948 = ~(n2016 | n10441);
assign n161 = n13547 | n2492;
assign n10301 = n12351 | n11537;
assign n3101 = ~(n4589 | n4079);
assign n3956 = n4498 | n6138;
assign n5010 = n9811 & n10100;
assign n3028 = ~n13365;
assign n9351 = n7267 & n12717;
assign n9240 = n13489 & n755;
assign n8850 = n2177 & n8055;
assign n14241 = n1805 | n4568;
assign n6437 = n10960 | n9645;
assign n10824 = n8737 | n4615;
assign n9592 = ~n7931;
assign n160 = n13310 | n3908;
assign n8968 = n3268 & n2297;
assign n7332 = n568 | n9508;
assign n4576 = n12414 | n12635;
assign n496 = ~n2932;
assign n7685 = n6311 & n10988;
assign n12114 = n2246 | n11783;
assign n10961 = n5570 | n624;
assign n4675 = n13520 & n6552;
assign n2056 = n3120 | n6863;
assign n1430 = n3168 | n13261;
assign n7261 = n12821 | n1687;
assign n2724 = ~n13181;
assign n2276 = ~(n13875 | n1149);
assign n12904 = ~n4379;
assign n1833 = n11511 & n12243;
assign n12855 = n2021 & n12579;
assign n11613 = n6609 & n2570;
assign n7816 = n9941 | n10765;
assign n5672 = n12425 & n8723;
assign n2539 = n5092 & n12262;
assign n2851 = ~(n8404 | n6324);
assign n12005 = ~(n9078 | n7890);
assign n7991 = n12611 & n6427;
assign n4867 = n13246 & n2902;
assign n10625 = ~(n14166 | n13124);
assign n1185 = ~(n11765 | n11125);
assign n2627 = n11688 | n10050;
assign n10238 = ~n9589;
assign n1321 = ~(n13875 | n11131);
assign n4725 = n5825 & n2719;
assign n3289 = n9571 & n13095;
assign n3066 = n4844 & n11397;
assign n8199 = ~(n11870 | n10287);
assign n4709 = n3212 & n2885;
assign n1629 = n13781 & n4802;
assign n4510 = n9792 & n6383;
assign n4896 = n1431 & n7108;
assign n8247 = ~n5108;
assign n5987 = n4659 & n12912;
assign n11268 = n13407 & n9166;
assign n9054 = n5139 | n7989;
assign n13218 = n5641 | n6034;
assign n8961 = n1031 | n5163;
assign n8795 = n2067 | n6555;
assign n309 = ~n5118;
assign n332 = n5236 | n7613;
assign n8888 = n14358 & n6267;
assign n8488 = n5483 | n12501;
assign n2283 = n2587 & n7055;
assign n9776 = ~n6520;
assign n1938 = n679 & n7397;
assign n6614 = ~n99;
assign n6310 = n11422 & n14049;
assign n3993 = n13142 | n6309;
assign n2816 = n5591 & n5645;
assign n14105 = n2179 | n1195;
assign n319 = n6957 & n11585;
assign n12676 = n2908 | n7610;
assign n5779 = ~n1495;
assign n10227 = n2089 | n477;
assign n166 = n2422 & n7038;
assign n7289 = n461 & n6614;
assign n11649 = n5071 & n11879;
assign n88 = n838 | n9407;
assign n2179 = ~n238;
assign n13327 = ~n13967;
assign n12288 = ~n3742;
assign n5542 = ~(n8816 | n10082);
assign n13222 = n687 & n4304;
assign n1978 = n10408 & n528;
assign n2698 = n11909 | n5692;
assign n7764 = n10332 & n1967;
assign n5226 = ~n7832;
assign n7928 = n446 & n11603;
assign n8043 = ~n6119;
assign n6238 = n4988 | n4622;
assign n4970 = n1047 & n2960;
assign n587 = n3755 & n13824;
assign n6172 = ~(n5852 | n8370);
assign n13799 = n12998 & n9532;
assign n8527 = ~n9686;
assign n6268 = n320 & n3549;
assign n10708 = n7768 & n7181;
assign n13463 = n6016 & n5498;
assign n13451 = n4684 | n6009;
assign n9504 = n7691 & n8087;
assign n14159 = n2229 | n12665;
assign n13871 = n12335 & n11989;
assign n8769 = ~n5427;
assign n4972 = n10534 | n8379;
assign n6025 = n13103 & n5828;
assign n13918 = n8025 & n12375;
assign n10638 = ~n7518;
assign n14096 = ~(n799 | n5043);
assign n6487 = n965 & n12138;
assign n94 = n7427 & n14497;
assign n13371 = n5975 & n11385;
assign n7329 = n5857 & n10450;
assign n6031 = n12802 & n12669;
assign n282 = n9015 & n629;
assign n8086 = ~(n2017 | n8939);
assign n2861 = n7768 & n41;
assign n13028 = n1140 & n905;
assign n9117 = n14472 | n10156;
assign n8921 = n1844 | n8178;
assign n8510 = n6672 | n3061;
assign n10387 = ~(n13675 | n10719);
assign n5195 = ~n5852;
assign n10288 = n1147 | n3784;
assign n10474 = n14107 | n8523;
assign n10184 = n8969 | n5566;
assign n4706 = n4104 & n1410;
assign n1992 = n13537 | n1928;
assign n5500 = n4358 & n5233;
assign n7245 = ~n9596;
assign n6464 = n7683 | n9246;
assign n741 = n4156 & n5551;
assign n2092 = n7970 & n10670;
assign n12631 = n5732 | n4904;
assign n12796 = n4255 | n509;
assign n7075 = ~n13408;
assign n12265 = ~n9197;
assign n4782 = ~(n13458 | n5649);
assign n3264 = n8726 | n8182;
assign n8128 = n13227 & n11095;
assign n11348 = n1362 | n8602;
assign n2386 = n7212 | n3163;
assign n9635 = n10825 | n9605;
assign n11359 = n2149 | n6237;
assign n5497 = ~(n13310 | n2807);
assign n5537 = n4807 | n14103;
assign n6533 = n9864 | n6780;
assign n9991 = n12870 | n5532;
assign n11076 = n9315 & n13082;
assign n9049 = n9724 & n2965;
assign n11909 = ~n14354;
assign n11456 = n9679 & n5959;
assign n4217 = n12712 | n9755;
assign n7140 = n12229 & n4062;
assign n13205 = n7221 & n7135;
assign n13602 = n10784 | n10262;
assign n7383 = n8247 & n3839;
assign n3815 = ~n5901;
assign n5337 = n9111 | n2280;
assign n11811 = n11123 | n6573;
assign n13972 = n11614 & n978;
assign n1684 = n4562 | n4674;
assign n1791 = ~(n6768 | n5006);
assign n13245 = n1538 | n1242;
assign n10778 = n2645 | n14468;
assign n11863 = n12601 | n11252;
assign n8168 = ~n14181;
assign n7604 = n5491 | n11753;
assign n9191 = ~n5460;
assign n11938 = ~n4342;
assign n5145 = n11935 | n9472;
assign n5051 = ~(n11481 | n11073);
assign n4001 = n5940 & n8811;
assign n14433 = ~n6743;
assign n8949 = n11704 | n11939;
assign n920 = ~n4715;
assign n5734 = n2090 | n9314;
assign n10067 = n6898 & n4395;
assign n6474 = ~(n3003 | n6729);
assign n13963 = n678 & n13762;
assign n10334 = n9297 & n6962;
assign n535 = n55 & n7150;
assign n4879 = n10731 | n4994;
assign n10578 = n8512 & n10623;
assign n7050 = ~n4518;
assign n9489 = n10367 & n4594;
assign n8577 = ~(n14196 | n5210);
assign n811 = n1031 | n1874;
assign n11220 = ~n3356;
assign n5508 = n3777 | n864;
assign n1071 = ~n11715;
assign n2023 = n2901 | n11686;
assign n10931 = n747 | n7347;
assign n590 = n9507 | n4166;
assign n986 = ~n5951;
assign n14225 = n12015 & n5766;
assign n4596 = n13854 | n9385;
assign n9791 = n8096 | n5016;
assign n1439 = n11033 & n8297;
assign n4057 = n13626 & n8790;
assign n8389 = ~(n450 | n5542);
assign n13736 = n9541 | n3978;
assign n4609 = n4146 & n5131;
assign n5627 = n7846 & n2738;
assign n2329 = n14472 | n2569;
assign n7399 = n4923 | n404;
assign n3827 = n7462 | n5019;
assign n6707 = n7683 | n5376;
assign n4326 = n10367 & n14515;
assign n11325 = ~n2202;
assign n4499 = n4923 | n4413;
assign n1663 = n4354 & n8981;
assign n8374 = ~(n10609 | n11178);
assign n13996 = ~(n5833 | n5669);
assign n4740 = n3813 & n6812;
assign n8083 = n1904 & n4495;
assign n1955 = ~n6305;
assign n6986 = n6781 | n13046;
assign n9793 = ~n7036;
assign n12858 = ~n6113;
assign n7320 = n6697 & n13123;
assign n11609 = ~(n9807 | n12920);
assign n12152 = n10458 & n7300;
assign n7114 = n5891 | n13127;
assign n5996 = n1061 | n4621;
assign n10711 = n103 & n7572;
assign n9965 = n2904 & n6064;
assign n5443 = n9716 | n1978;
assign n2575 = ~n3233;
assign n4064 = ~(n6520 | n6482);
assign n7936 = n14093 & n660;
assign n277 = n9716 | n3227;
assign n4492 = n14157 & n11592;
assign n188 = n7187 & n2869;
assign n1463 = ~(n6883 | n13244);
assign n14263 = n11094 | n4014;
assign n4468 = ~n3616;
assign n9562 = ~n3673;
assign n13471 = ~(n7245 | n13573);
assign n3697 = n12568 | n4330;
assign n9852 = n5553 & n8637;
assign n2858 = n8980 | n7254;
assign n14371 = n5997 | n5008;
assign n11346 = n2597 | n8698;
assign n5442 = n12542 & n8771;
assign n13532 = n12169 | n1176;
assign n10486 = n11803 & n8905;
assign n10258 = n2016 | n8289;
assign n9047 = ~(n8081 | n2085);
assign n162 = ~n13900;
assign n2102 = n11704 | n13961;
assign n7915 = n13650 & n10002;
assign n11105 = ~n14154;
assign n4145 = n5936 | n6148;
assign n8237 = n8881 | n11063;
assign n7853 = n3536 & n3261;
assign n8221 = n12615 & n475;
assign n7057 = ~n8555;
assign n14012 = n2724 & n11963;
assign n13586 = ~(n3210 | n1682);
assign n11053 = n13863 & n1774;
assign n6000 = ~n12691;
assign n7926 = n7391 & n6003;
assign n3612 = n7767 & n13043;
assign n6790 = ~(n12548 | n10475);
assign n9394 = n13706 | n810;
assign n5901 = n1506 & n3704;
assign n13390 = n8507 | n9154;
assign n3020 = n3169 & n3665;
assign n11468 = n1051 | n4789;
assign n4257 = n12042 & n10081;
assign n2522 = n2521 & n11941;
assign n11794 = n14088 | n5624;
assign n4928 = ~n12975;
assign n11071 = ~n2241;
assign n4627 = ~n6113;
assign n11739 = ~n10108;
assign n12190 = n3062 | n5340;
assign n3645 = ~(n3428 | n3927);
assign n7322 = n8884 & n11882;
assign n6214 = n13537 | n5332;
assign n8738 = n13112 | n9946;
assign n11835 = n9856 | n1301;
assign n14308 = n13108 | n816;
assign n6307 = n5011 & n1885;
assign n11250 = n4851 & n13766;
assign n2786 = n9944 & n6084;
assign n6831 = n2942 & n11982;
assign n3168 = ~n777;
assign n10168 = n12844 | n3292;
assign n12501 = n10930 & n14262;
assign n7544 = n11838 & n7974;
assign n1766 = n4486 & n4864;
assign n12703 = n13941 | n13646;
assign n12500 = ~n11152;
assign n2536 = n13362 & n6473;
assign n7323 = n6781 | n13558;
assign n10840 = n10539 | n42;
assign n6117 = ~(n4637 | n6089);
assign n4947 = n1137 | n1830;
assign n12198 = ~(n7245 | n7658);
assign n1519 = ~(n3132 | n6048);
assign n5860 = ~(n588 | n575);
assign n8427 = ~n9197;
assign n11912 = n12042 & n8722;
assign n14258 = n3268 & n10452;
assign n170 = n9403 | n8622;
assign n11594 = n11710 | n7276;
assign n9720 = n5275 & n5887;
assign n11905 = n5252 & n11228;
assign n13178 = n8332 | n4843;
assign n12406 = n8513 | n8410;
assign n6601 = n1489 & n9209;
assign n14015 = n3755 & n14281;
assign n7435 = n7436 | n4238;
assign n11968 = n457 & n6871;
assign n6452 = n10154 | n4935;
assign n14039 = ~n6480;
assign n12800 = ~n6554;
assign n12387 = n2082 & n13930;
assign n10924 = ~(n2790 | n12530);
assign n14102 = n361 | n1646;
assign n9614 = ~(n12522 | n7500);
assign n2074 = n781 | n1783;
assign n12074 = n10767 & n1325;
assign n5343 = ~(n6313 | n13422);
assign n298 = ~n13356;
assign n8938 = n3125 | n3431;
assign n13052 = n1356 | n13042;
assign n1979 = n3492 & n11190;
assign n13130 = ~n3046;
assign n11507 = n12105 & n12830;
assign n2827 = n392 & n3429;
assign n13469 = n7914 | n141;
assign n122 = n3491 & n8941;
assign n14108 = n11459 | n6372;
assign n4261 = ~n8555;
assign n9129 = n4856 & n9940;
assign n9419 = n1427 & n2785;
assign n13817 = n14198 | n13440;
assign n9254 = n8238 & n4076;
assign n14065 = ~n6946;
assign n14120 = ~n1120;
assign n12416 = n13706 | n2097;
assign n13687 = n1044 | n14328;
assign n11032 = n12389 & n11716;
assign n8684 = n838 | n11800;
assign n10672 = n1802 | n10080;
assign n8638 = ~n8813;
assign n5667 = n5144 | n1213;
assign n2686 = ~n11788;
assign n367 = n3445 | n10421;
assign n418 = n8480 | n11553;
assign n13294 = n8923 & n924;
assign n14195 = n14058 | n4016;
assign n8529 = ~n1997;
assign n7934 = ~n13625;
assign n9378 = ~(n4544 | n2398);
assign n1744 = ~(n3444 | n6447);
assign n3201 = n7779 & n13843;
assign n8026 = n2055 | n4268;
assign n12757 = ~n10965;
assign n1841 = n8965 & n9114;
assign n1062 = n4698 & n10198;
assign n6058 = n11687 & n220;
assign n7882 = n14029 | n2926;
assign n4781 = n12259 & n728;
assign n9656 = n5628 & n1565;
assign n8762 = ~(n8877 | n13063);
assign n3935 = n13155 | n10879;
assign n8561 = n7364 | n13603;
assign n6522 = n7419 & n8129;
assign n9383 = n3 & n1292;
assign n11415 = n11218 & n5782;
assign n8548 = ~(n7359 | n8389);
assign n7773 = n361 | n124;
assign n2455 = n49 | n2648;
assign n5831 = n11704 | n2278;
assign n9396 = ~(n5391 | n5585);
assign n4982 = n9811 & n1950;
assign n9897 = n9617 & n11140;
assign n10343 = n5406 | n10686;
assign n10895 = n9229 | n6126;
assign n7499 = n4300 & n14470;
assign n6438 = n6654 | n10424;
assign n5665 = ~n11347;
assign n4859 = n1203 & n9008;
assign n9322 = n1339 & n10003;
assign n9421 = n10408 & n383;
assign n9411 = n11121 | n12398;
assign n4025 = n11674 & n3763;
assign n6679 = ~n2996;
assign n2357 = n13209 | n3910;
assign n11474 = ~n6212;
assign n2581 = n13535 & n3956;
assign n2229 = ~n4609;
assign n7924 = n6730 | n6216;
assign n6469 = n1669 | n13423;
assign n12781 = n9984 | n7195;
assign n1935 = n5104 & n2898;
assign n6359 = n10589 & n12261;
assign n8501 = n7530 | n11419;
assign n13275 = n6607 | n1345;
assign n1415 = n480 | n13922;
assign n7342 = n13155 | n8400;
assign n12192 = ~n2332;
assign n7695 = ~(n5480 | n1092);
assign n11280 = ~(n8361 | n3582);
assign n11467 = n1588 & n538;
assign n236 = n3512 | n8283;
assign n3979 = n13718 | n2490;
assign n3423 = n13379 & n4012;
assign n6935 = n14145 & n7085;
assign n11462 = n4876 | n8967;
assign n3246 = n5628 & n3036;
assign n2892 = ~(n3802 | n6150);
assign n3511 = n13952 & n6032;
assign n8686 = n11048 | n4408;
assign n6729 = ~(n10136 | n8481);
assign n2752 = ~n10861;
assign n1356 = ~n7819;
assign n4593 = n5800 | n2373;
assign n11039 = n6311 & n10875;
assign n483 = ~(n13435 | n13939);
assign n14069 = n1840 | n7185;
assign n392 = ~n14525;
assign n3856 = n5064 | n3519;
assign n7239 = n12721 & n9262;
assign n13193 = ~(n11706 | n5196);
assign n6433 = n2158 & n8530;
assign n5572 = n4052 | n11013;
assign n5254 = n14481 | n12387;
assign n12038 = ~n5153;
assign n3348 = n10331 | n4813;
assign n10799 = n12038 & n1884;
assign n2426 = n9920 & n6045;
assign n798 = n8242 | n10313;
assign n6633 = n2843 | n14022;
assign n8424 = ~n5761;
assign n4756 = ~(n6326 | n11911);
assign n5830 = n11440 | n13552;
assign n7167 = n11220 & n8510;
assign n3955 = n14404 | n2715;
assign n7610 = n8965 & n8448;
assign n3793 = n6607 | n13232;
assign n10104 = n9423 | n4570;
assign n8005 = n446 & n14237;
assign n9106 = n12990 & n547;
assign n6006 = n898 & n10950;
assign n3567 = n11411 & n1286;
assign n7576 = n12622 | n2502;
assign n5961 = n8789 & n518;
assign n13408 = ~n12069;
assign n9844 = n11953 | n10711;
assign n13593 = n12852 & n5398;
assign n6446 = n4913 | n12376;
assign n11893 = n11702 & n7360;
assign n1122 = n12270 & n6384;
assign n6723 = ~(n4082 | n356);
assign n10433 = n3276 & n5249;
assign n6922 = n11737 & n1785;
assign n3894 = ~(n13213 | n14183);
assign n9628 = n1660 | n205;
assign n4374 = n5553 & n5456;
assign n2320 = n5678 & n6099;
assign n3355 = ~(n10637 | n13776);
assign n5621 = ~n11350;
assign n482 = ~n2462;
assign n219 = n13991 | n4492;
assign n4265 = n9238 & n5204;
assign n8154 = ~(n12888 | n11566);
assign n10197 = ~n9583;
assign n12506 = n10360 | n7272;
assign n1161 = n2924 | n6362;
assign n9649 = n13863 & n13336;
assign n2770 = n12421 & n3218;
assign n1516 = n5406 | n4148;
assign n116 = ~n14412;
assign n10532 = n1261 | n10256;
assign n9346 = n6706 | n6001;
assign n5243 = ~(n5505 | n5497);
assign n11823 = n4973 & n13619;
assign n5982 = ~(n2057 | n3487);
assign n6125 = ~(n10649 | n386);
assign n11239 = n10289 | n13492;
assign n7899 = n12651 | n2929;
assign n222 = ~n1639;
assign n9877 = n14282 | n7765;
assign n10854 = ~n12450;
assign n5436 = n5926 & n9915;
assign n10781 = ~n5627;
assign n11342 = n7911 & n5327;
assign n9866 = n7970 & n4576;
assign n14140 = n9541 | n4466;
assign n5028 = n12521 & n357;
assign n11224 = n3715 & n12212;
assign n12221 = n6111 | n12184;
assign n13967 = ~n7091;
assign n7197 = ~(n2098 | n5938);
assign n6098 = n9211 | n24;
assign n7823 = n12105 & n11098;
assign n2629 = n7898 | n13571;
assign n11414 = n103 & n5670;
assign n7637 = n2888 | n10870;
assign n13257 = n12779 & n1210;
assign n6236 = n4821 | n3707;
assign n14382 = n2330 & n3335;
assign n2544 = ~(n7359 | n7692);
assign n10230 = n3785 & n694;
assign n1215 = n9617 & n7198;
assign n11986 = n10374 & n7607;
assign n12166 = n7354 & n3734;
assign n12080 = n3667 | n6604;
assign n980 = n12139 | n812;
assign n12331 = n8446 & n8131;
assign n10992 = n900 | n11038;
assign n14462 = n12131 | n12118;
assign n6023 = ~n1568;
assign n3784 = n2961 & n9522;
assign n1690 = n584 | n5074;
assign n5419 = n12953 & n9851;
assign n4093 = ~(n8701 | n2515);
assign n2959 = n9742 | n4005;
assign n9481 = n3536 & n371;
assign n3320 = ~n8148;
assign n1058 = n11542 | n4543;
assign n5168 = n2461 & n12854;
assign n12200 = ~n5678;
assign n7131 = n8849 & n11022;
assign n1450 = n9080 & n7648;
assign n1218 = ~n2577;
assign n11660 = n7938 | n1268;
assign n10746 = ~(n8015 | n14104);
assign n12441 = n3405 & n8406;
assign n4449 = n11737 & n652;
assign n11375 = n13867 & n5663;
assign n13774 = n6163 | n8753;
assign n7910 = n5007 | n5442;
assign n12057 = ~n8650;
assign n5461 = n5815 | n2590;
assign n3186 = n2422 & n2300;
assign n11953 = ~n4317;
assign n7865 = n13484 & n11202;
assign n8149 = n9422 | n10207;
assign n959 = n1804 & n671;
assign n13572 = ~n3870;
assign n3959 = ~n13476;
assign n12337 = n5406 | n2092;
assign n1526 = ~n13213;
assign n12999 = ~n14320;
assign n10374 = ~n8451;
assign n6548 = n11620 | n13606;
assign n9278 = n9742 | n6522;
assign n4106 = n2086 | n5822;
assign n3536 = ~n5460;
assign n13397 = n8183 & n7807;
assign n11472 = ~n3616;
assign n1799 = n3424 & n1998;
assign n11840 = n9353 | n2823;
assign n5313 = n8393 & n11972;
assign n4286 = n13518 | n3012;
assign n8500 = n1850 | n10446;
assign n7008 = ~(n6765 | n13313);
assign n5466 = n766 | n2576;
assign n5992 = n405 & n10143;
assign n701 = ~(n11975 | n2424);
assign n13447 = ~n6714;
assign n2987 = n1452 & n499;
assign n10526 = n8412 & n14069;
assign n10242 = n2983 & n12476;
assign n6668 = n8453 & n5863;
assign n1199 = n11839 | n7040;
assign n8948 = n11153 & n11750;
assign n9327 = n11558 | n14264;
assign n457 = ~n12450;
assign n7062 = n2904 & n2836;
assign n4307 = ~(n9529 | n7371);
assign n6720 = n7530 | n1320;
assign n10251 = n8630 & n1683;
assign n13209 = ~n8873;
assign n237 = ~(n2799 | n9039);
assign n5793 = n10784 | n7977;
assign n13733 = n9490 | n4700;
assign n9283 = n7053 & n10839;
assign n13208 = ~(n3248 | n13858);
assign n7112 = n3286 & n11217;
assign n11127 = n7370 & n13932;
assign n12642 = n2761 | n5983;
assign n6711 = ~n10346;
assign n14070 = ~(n1112 | n4848);
assign n13907 = n13641 & n10805;
assign n768 = n3815 | n11311;
assign n6130 = ~n5606;
assign n14281 = n4033 | n12892;
assign n4483 = n10523 | n11230;
assign n11159 = n5807 | n10129;
assign n9689 = n6039 | n1372;
assign n1777 = ~(n8877 | n13670);
assign n13737 = n3768 | n5826;
assign n2069 = ~n1760;
assign n4171 = n13226 | n9696;
assign n11805 = ~(n5605 | n36);
assign n6817 = ~(n584 | n6590);
assign n5019 = n8183 & n5036;
assign n3702 = ~(n7011 | n5410);
assign n13421 = ~n6657;
assign n6334 = n10624 | n617;
assign n2837 = n4898 | n6110;
assign n13298 = ~n3230;
assign n1329 = n1268 & n2255;
assign n13308 = n5471 & n11693;
assign n13513 = n4619 & n11600;
assign n12948 = n8692 & n7668;
assign n13050 = ~n13158;
assign n10605 = n1610 & n10123;
assign n10484 = n7267 & n8256;
assign n7461 = n5317 & n8237;
assign n5994 = n5997 | n4223;
assign n11236 = n8513 | n753;
assign n9813 = n5926 & n13933;
assign n4857 = n8969 | n6429;
assign n12869 = n9111 | n8094;
assign n7981 = ~(n448 | n3726);
assign n7946 = ~(n3577 | n1063);
assign n11641 = ~(n10241 | n2612);
assign n10153 = n8697 & n7944;
assign n1712 = ~(n10312 | n13148);
assign n5479 = n14072 & n5728;
assign n9438 = n14107 | n595;
assign n763 = n4065 | n14015;
assign n7111 = n8476 | n6411;
assign n9979 = n11569 & n2436;
assign n10490 = n4261 & n13305;
assign n14167 = n2518 | n1867;
assign n14171 = n13535 & n14345;
assign n11873 = n2878 | n7042;
assign n1351 = n1044 | n6919;
assign n4407 = ~n1833;
assign n500 = ~n4634;
assign n6719 = n6724 & n8589;
assign n259 = n7862 | n13732;
assign n8588 = n222 & n14494;
assign n6917 = n3545 | n8100;
assign n10978 = n11123 | n5630;
assign n2956 = n5071 & n6452;
assign n5140 = n12460 & n7796;
assign n2094 = n10050 | n5046;
assign n5893 = ~(n7755 | n4662);
assign n10023 = n1172 | n805;
assign n12588 = n13756 & n3037;
assign n13535 = ~n10322;
assign n13498 = ~(n11428 | n8727);
assign n8791 = n14327 & n5329;
assign n3909 = ~(n2094 | n9017);
assign n1600 = n11329 & n7517;
assign n2192 = n14446 & n12682;
assign n2055 = ~n4777;
assign n2430 = n5647 | n6262;
assign n10595 = ~n14332;
assign n1630 = n5483 | n8342;
assign n9765 = ~(n11667 | n6877);
assign n12778 = n2587 & n2657;
assign n6375 = n3168 | n12373;
assign n6567 = ~(n2923 | n8134);
assign n1035 = n1258 | n7531;
assign n1482 = n13863 & n10831;
assign n4327 = n1189 | n8343;
assign n5246 = n2998 & n6464;
assign n12380 = ~(n8752 | n10326);
assign n11306 = n5458 & n10939;
assign n3830 = n11411 & n14045;
assign n2635 = n3724 & n4697;
assign n6911 = n7116 | n7417;
assign n5553 = ~n2619;
assign n8376 = ~n1637;
assign n14506 = n13675 | n12883;
assign n11303 = ~n11456;
assign n5035 = ~n56;
assign n2128 = ~(n5833 | n11376);
assign n7711 = n6609 & n6548;
assign n11812 = ~(n7227 | n1675);
assign n2180 = ~n9546;
assign n14094 = n12633 | n9196;
assign n9204 = n9269 | n1696;
assign n2248 = n5800 | n2972;
assign n6451 = n14210 & n12964;
assign n8072 = ~(n1914 | n5912);
assign n10308 = ~(n1914 | n13637);
assign n6550 = n6753 & n7903;
assign n3758 = n14058 | n6644;
assign n10742 = n10072 & n1232;
assign n7321 = n873 & n1015;
assign n3000 = n4394 & n3050;
assign n13356 = n5467 | n7282;
assign n8037 = n9151 | n11494;
assign n9474 = n13780 & n586;
assign n3071 = n13847 | n8119;
assign n5264 = n7053 & n10794;
assign n7159 = n10909 & n6802;
assign n7429 = ~n8168;
assign n12014 = n8450 & n1469;
assign n1337 = ~(n3427 | n10697);
assign n611 = n3009 | n3609;
assign n339 = n5948 & n13898;
assign n11583 = n2367 & n13783;
assign n2184 = n13236 & n14095;
assign n4424 = ~n12189;
assign n9089 = n11097 | n2325;
assign n10027 = n4546 & n12729;
assign n11669 = n14400 | n10684;
assign n7154 = n6609 & n10053;
assign n3271 = ~n4774;
assign n10823 = ~(n10186 | n6476);
assign n2821 = n1728 | n5179;
assign n12029 = n7358 | n14278;
assign n2562 = ~n14354;
assign n9335 = n12500 | n2909;
assign n12821 = ~n8272;
assign n3213 = n14472 | n9464;
assign n7174 = n3219 | n7283;
assign n3282 = n2750 | n11958;
assign n13406 = ~(n12568 | n12170);
assign n10791 = n10378 & n2014;
assign n608 = n9190 & n3783;
assign n7031 = n8932 & n6619;
assign n10701 = n2086 | n2647;
assign n10704 = n5899 & n6136;
assign n13813 = n10300 | n5796;
assign n8509 = n1834 | n331;
assign n5969 = n2761 | n5462;
assign n1053 = n7476 | n5943;
assign n11844 = n10562 & n12;
assign n1878 = n898 & n3275;
assign n512 = ~n8162;
assign n2906 = ~n6855;
assign n10113 = n8768 & n10409;
assign n10755 = n9232 & n13115;
assign n5606 = ~n8927;
assign n11020 = ~n3313;
assign n8170 = n5507 | n11464;
assign n3563 = n6525 & n8373;
assign n2221 = n9705 & n5200;
assign n5548 = ~n630;
assign n11021 = n11867 & n12639;
assign n13875 = ~n4325;
assign n12783 = n7678 | n596;
assign n14428 = n251 | n12448;
assign n6368 = n4484 & n7318;
assign n10161 = n7898 | n12584;
assign n5659 = n7250 | n8601;
assign n3948 = n14120 & n2748;
assign n4619 = ~n3922;
assign n2506 = n9403 | n5991;
assign n2725 = n13107 & n1658;
assign n7337 = n553 | n13315;
assign n11293 = n7684 | n8918;
assign n10503 = n3635 & n14277;
assign n6432 = n10589 & n859;
assign n11139 = n1741 | n3409;
assign n7589 = ~n2354;
assign n12197 = ~n13084;
assign n11450 = n781 | n2215;
assign n8119 = n9069 & n4314;
assign n10673 = n1266 & n11626;
assign n9755 = n11748 & n12344;
assign n12296 = n12013 & n11845;
assign n731 = ~(n12968 | n4118);
assign n8766 = n77 | n4902;
assign n3720 = n8431 & n7560;
assign n4805 = n4095 & n7833;
assign n1653 = n10224 | n13729;
assign n7784 = n2998 & n5878;
assign n10900 = n3736 & n13195;
assign n10314 = ~n1769;
assign n3318 = n1623 | n535;
assign n8905 = n13155 | n1607;
assign n12945 = n4657 & n1597;
assign n13382 = n14358 & n5443;
assign n8446 = n6256 | n6946;
assign n8714 = ~n7322;
assign n10325 = n8015 | n7020;
assign n12454 = n7852 & n13889;
assign n4515 = n4382 | n4117;
assign n10127 = n10539 | n7338;
assign n1544 = n11384 & n12310;
assign n602 = ~(n1838 | n12513);
assign n4415 = ~n8223;
assign n13649 = n231 & n12770;
assign n2667 = n1193 & n4494;
assign n11557 = n9188 & n4487;
assign n10355 = ~(n8487 | n6368);
assign n14278 = n13227 & n2591;
assign n148 = n12229 & n13532;
assign n12008 = ~(n7227 | n9137);
assign n2253 = n11105 | n14299;
assign n1654 = n3569 | n6101;
assign n130 = n1031 | n9074;
assign n8464 = ~(n2875 | n7617);
assign n14394 = n8393 & n9382;
assign n10347 = ~(n6888 | n3863);
assign n7616 = n8412 & n4947;
assign n1147 = ~n2934;
assign n541 = ~n8650;
assign n5530 = n10622 & n3013;
assign n11495 = ~n14525;
assign n6157 = ~n5427;
assign n8360 = ~(n8209 | n9875);
assign n10241 = ~n5788;
assign n6611 = n4065 | n587;
assign n12992 = ~n2615;
assign n12360 = n14481 | n8664;
assign n884 = n13224 & n5860;
assign n13402 = n8401 & n6283;
assign n5018 = ~n5921;
assign n11719 = n10913 | n11250;
assign n9774 = n4574 & n1667;
assign n6440 = ~(n4046 | n6028);
assign n12329 = n5180 | n12442;
assign n2403 = n8950 & n13610;
assign n13179 = n13850 & n8844;
assign n2919 = ~n381;
assign n8841 = n12611 & n3627;
assign n10450 = n283 | n5930;
assign n5361 = ~(n1838 | n6512);
assign n5284 = n2790 | n2148;
assign n12561 = n4300 & n11869;
assign n12131 = ~n6332;
assign n6204 = n3370 & n10240;
assign n2416 = n12401 | n1256;
assign n3443 = ~n3812;
assign n11099 = n3766 & n6214;
assign n5400 = ~(n619 | n9066);
assign n8403 = n6690 | n11127;
assign n2999 = ~(n2742 | n7170);
assign n246 = n7122 | n6885;
assign n10697 = n7618 & n13819;
assign n10544 = n8513 | n4612;
assign n6700 = ~n13756;
assign n1560 = n14449 | n7760;
assign n3682 = n11123 | n6739;
assign n3899 = ~(n2086 | n5724);
assign n8731 = n10383 | n8974;
assign n7184 = n8450 & n2963;
assign n4908 = ~n7064;
assign n1466 = n11406 & n3860;
assign n3231 = n783 & n1695;
assign n9740 = ~n1417;
assign n567 = n13433 & n8928;
assign n7058 = n6109 | n8711;
assign n1397 = n12425 & n5201;
assign n6535 = n14029 | n12945;
assign n6765 = ~n1984;
assign n992 = n5315 | n7348;
assign n2609 = n4320 & n13682;
assign n5547 = n10834 | n4805;
assign n2149 = ~n3284;
assign n3483 = n4803 & n1541;
assign n11901 = n271 | n3367;
assign n3648 = n9345 & n3968;
assign n13435 = ~n4415;
assign n6367 = n1354 & n12547;
assign n10100 = n194 | n12661;
assign n6751 = ~(n1812 | n13585);
assign n11907 = n11183 | n11552;
assign n448 = ~n7258;
assign n85 = ~n1894;
assign n9605 = n9188 & n10683;
assign n9705 = ~n10376;
assign n13828 = n4880 & n9708;
assign n3169 = ~n9592;
assign n11124 = n8232 & n8125;
assign n5922 = n10909 & n10832;
assign n3573 = n1937 & n6801;
assign n10906 = n10909 & n3108;
assign n5445 = n11231 | n12856;
assign n6445 = n2682 & n11091;
assign n1739 = n12336 & n9432;
assign n4262 = n9705 & n10795;
assign n5709 = n6724 & n8435;
assign n13725 = n5640 & n3760;
assign n3212 = ~n1478;
assign n6404 = ~(n10136 | n3934);
assign n13431 = n6471 | n14473;
assign n1123 = n6609 & n966;
assign n10718 = n6649 & n825;
assign n14431 = n10562 & n4945;
assign n13723 = ~n1938;
assign n3412 = n13626 & n8240;
assign n5715 = ~n6332;
assign n12277 = n11240 & n8962;
assign n491 = ~(n573 | n8688);
assign n12799 = n185 | n6987;
assign n13732 = n6527 & n10098;
assign n476 = n3427 | n4248;
assign n6642 = n6854 & n10914;
assign n91 = n3833 & n12664;
assign n8234 = n2761 | n10724;
assign n2568 = n14063 & n8053;
assign n8490 = ~n10204;
assign n4440 = n9345 & n3550;
assign n7072 = ~(n6743 | n6228);
assign n13635 = n12047 | n813;
assign n9983 = n1061 | n9128;
assign n7828 = n13108 | n3117;
assign n7955 = ~(n4742 | n12028);
assign n9919 = n13860 & n13689;
assign n1167 = n13555 & n2306;
assign n11057 = n4899 | n255;
assign n9182 = n13968 | n11605;
assign n2541 = ~(n11980 | n2118);
assign n375 = n10449 | n5985;
assign n44 = n12047 | n9943;
assign n2501 = n8172 | n6061;
assign n13043 = n9507 | n1098;
assign n6450 = n7421 & n8014;
assign n12733 = n13755 & n9892;
assign n13117 = n2149 | n10796;
assign n2718 = n4692 & n1295;
assign n13025 = n7943 & n4155;
assign n405 = ~n5613;
assign n10938 = ~(n5278 | n4307);
assign n11834 = n11710 | n9773;
assign n7699 = n776 & n14304;
assign n2710 = n2367 & n14459;
assign n7004 = ~n8163;
assign n11976 = n13484 & n4767;
assign n14471 = n7684 | n13796;
assign n3850 = n14213 & n9945;
assign n11357 = n98 & n2386;
assign n3548 = n7961 & n5636;
assign n9546 = ~n8903;
assign n1010 = n3442 & n11129;
assign n4752 = n9198 & n3307;
assign n13659 = n10824 | n3822;
assign n1320 = n12521 & n3258;
assign n10321 = ~(n1844 | n12923);
assign n13695 = n1414 & n8200;
assign n9017 = n11688 & n4311;
assign n1898 = n13656 & n12368;
assign n2005 = ~n4906;
assign n2088 = n2901 | n12958;
assign n13087 = ~n1045;
assign n10686 = n12741 & n4861;
assign n8391 = n7803 | n5090;
assign n3819 = n3871 | n6049;
assign n6429 = n1428 & n13281;
assign n12479 = n12759 | n7456;
assign n9910 = n7392 & n1048;
assign n9105 = n12521 & n3053;
assign n1923 = n3219 | n1794;
assign n9131 = n1427 & n5322;
assign n9630 = ~(n10593 | n6132);
assign n1573 = n1662 & n7924;
assign n10962 = n5450 | n1943;
assign n5320 = n77 | n5246;
assign n3093 = ~n6804;
assign n2744 = ~n5151;
assign n6379 = n511 | n6617;
assign n9229 = ~n7289;
assign n12766 = ~(n4464 | n3278);
assign n13319 = n4098 & n4232;
assign n2336 = n9052 & n801;
assign n9063 = n13525 & n7753;
assign n6756 = n13847 | n8282;
assign n13966 = n4901 & n2448;
assign n12382 = n12414 | n4555;
assign n870 = n5362 | n688;
assign n8781 = n14430 | n13166;
assign n10620 = ~n7007;
assign n12627 = ~(n12727 | n14123);
assign n5526 = n13518 | n5674;
assign n7134 = n8849 & n4857;
assign n8177 = n12592 & n3626;
assign n2089 = ~n6332;
assign n7336 = n957 & n8975;
assign n3125 = ~n11308;
assign n4043 = n10035 | n11556;
assign n184 = n14321 & n5846;
assign n4033 = ~n9596;
assign n5539 = n11495 & n822;
assign n14481 = ~n11456;
assign n2025 = ~n3046;
assign n14289 = n14303 & n6630;
assign n3961 = n79 & n4428;
assign n2855 = n7911 & n7723;
assign n1077 = n850 | n940;
assign n1380 = n568 | n14171;
assign n13264 = n3401 & n11640;
assign n9297 = ~n12450;
assign n727 = ~n11793;
assign n2420 = ~(n10568 | n1765);
assign n623 = n5312 & n3596;
assign n9907 = ~(n2566 | n9065);
assign n11879 = n13118 | n9748;
assign n4860 = n5064 | n8035;
assign n13135 = n1361 & n9138;
assign n6865 = n2006 & n10881;
assign n12230 = n9824 & n11297;
assign n9627 = n11300 & n1248;
assign n8964 = ~n12444;
assign n4789 = n1857 & n934;
assign n13526 = ~(n14455 | n5058);
assign n4151 = n4821 | n5344;
assign n14254 = ~(n6603 | n9611);
assign n10118 = n2694 | n4679;
assign n14132 = n13676 & n824;
assign n3444 = ~n11052;
assign n8046 = n10166 & n13014;
assign n6991 = n5899 & n14499;
assign n10758 = n12721 & n10352;
assign n5845 = n8238 & n996;
assign n9908 = n6899 & n1679;
assign n11065 = n2790 | n12220;
assign n9237 = n12335 & n1981;
assign n12123 = n11220 & n9311;
assign n6234 = n7208 & n12524;
assign n7902 = ~n8903;
assign n13913 = n5926 & n8858;
assign n5569 = ~n1060;
assign n8763 = n5062 & n10707;
assign n3895 = ~n3799;
assign n9390 = ~(n5762 | n558);
assign n3333 = ~n14512;
assign n11843 = n2901 | n13375;
assign n7489 = n11223 | n3764;
assign n8779 = n11097 | n11043;
assign n6834 = n2750 | n11908;
assign n14463 = n11776 & n3450;
assign n9311 = n7436 | n13904;
assign n9236 = ~n3428;
assign n9532 = n12112 | n9910;
assign n3807 = n12960 & n12201;
assign n8 = n13509 & n1714;
assign n2583 = ~n12930;
assign n12183 = n12858 & n690;
assign n5968 = n12404 & n13605;
assign n6365 = ~(n8404 | n11116);
assign n981 = n3370 & n571;
assign n6579 = n12147 & n2605;
assign n10757 = n8714 | n12459;
assign n1425 = ~n12846;
assign n6409 = n5084 | n10628;
assign n72 = n8393 & n1700;
assign n9064 = n5279 & n8469;
assign n11 = n10760 & n7309;
assign n5455 = n11403 & n7048;
assign n6015 = n4655 & n3953;
assign n548 = n5548 | n6879;
assign n13020 = n7677 & n376;
assign n8564 = n6625 & n5477;
assign n9152 = n98 & n5658;
assign n10936 = ~n3284;
assign n9104 = n533 & n12452;
assign n5252 = ~n5606;
assign n8655 = ~n6436;
assign n9486 = n7156 | n10657;
assign n10972 = n7529 & n5713;
assign n861 = n12576 | n1521;
assign n10517 = n5807 | n11200;
assign n11247 = n5833 | n3644;
assign n11775 = n5234 | n2667;
assign n1689 = n14120 & n13662;
assign n12398 = n7443 & n11348;
assign n12023 = ~n12331;
assign n8870 = n185 | n3368;
assign n13044 = n2888 | n6177;
assign n8143 = ~(n7200 | n13551);
assign n12305 = n283 | n10780;
assign n2649 = n8748 | n12959;
assign n6980 = n541 & n14349;
assign n3845 = ~n7822;
assign n11297 = n504 | n3029;
assign n9176 = ~n10358;
assign n1527 = ~(n9563 | n12390);
assign n1644 = n10713 | n2141;
assign n10234 = ~n7875;
assign n1180 = ~(n12673 | n9737);
assign n3408 = n7327 & n4153;
assign n3986 = ~n5618;
assign n9040 = n10458 & n13411;
assign n4628 = n12592 & n12371;
assign n7759 = ~n12924;
assign n10566 = ~n355;
assign n9090 = ~(n4213 | n12966);
assign n12599 = n14400 | n3293;
assign n5728 = ~(n12827 | n4256);
assign n2 = n9230 | n2519;
assign n14146 = n12542 & n13549;
assign n1031 = ~n11308;
assign n3960 = n251 | n988;
assign n7896 = n6606 & n11815;
assign n8916 = n12500 | n1497;
assign n3704 = n7216 & n9654;
assign n8310 = n2177 & n7829;
assign n9887 = n12414 | n5531;
assign n3102 = n11621 | n12931;
assign n8359 = ~(n8529 | n8633);
assign n2294 = n10922 & n11891;
assign n10911 = n12131 | n7237;
assign n13842 = ~(n8576 | n5183);
assign n7522 = n3126 | n6201;
assign n9457 = n5876 & n11652;
assign n1932 = n10248 | n13561;
assign n5896 = n11839 | n10979;
assign n13979 = ~n11350;
assign n11860 = n5800 | n5307;
assign n4769 = n8975 & n1640;
assign n6377 = n6318 & n4922;
assign n7406 = n2111 | n11920;
assign n13238 = ~(n2218 | n3101);
assign n3539 = n10668 & n9843;
assign n2080 = ~n7748;
assign n12191 = ~n10406;
assign n14321 = ~n9583;
assign n7638 = ~(n9743 | n6057);
assign n2940 = n12185 & n10618;
assign n10461 = ~n4203;
assign n13346 = n12968 | n14285;
assign n7468 = n12047 | n7550;
assign n7800 = n14358 & n13925;
assign n5350 = n3164 | n1182;
assign n3983 = n533 & n9692;
assign n3545 = n8607 | n3457;
assign n6397 = ~n12675;
assign n4463 = ~(n3445 | n13085);
assign n13519 = ~(n6020 | n6972);
assign n7221 = ~n2932;
assign n10485 = n9803 & n7879;
assign n1507 = n3527 | n11225;
assign n10048 = n2783 & n1870;
assign n6859 = n873 & n6261;
assign n1556 = n13706 | n10107;
assign n11974 = n14366 | n6585;
assign n56 = n10953 | n11961;
assign n6490 = n4180 | n8945;
assign n4038 = n8877 | n7296;
assign n12490 = n1481 & n8093;
assign n12421 = ~n3361;
assign n11815 = n4340 | n5360;
assign n10219 = n636 & n723;
assign n486 = n6753 & n12082;
assign n2595 = n5409 | n2654;
assign n6207 = n1708 & n616;
assign n13011 = ~(n5042 | n2395);
assign n37 = n5454 | n11132;
assign n3382 = n5507 | n785;
assign n13106 = n706 & n2994;
assign n7037 = n10539 | n7511;
assign n11505 = ~(n3871 | n9690);
assign n5732 = ~n9354;
assign n4750 = n14404 | n12797;
assign n4478 = n10229 & n7873;
assign n11991 = n14446 & n132;
assign n3579 = n13413 | n2555;
assign n8416 = n10191 | n14287;
assign n10603 = n9673 & n379;
assign n11194 = n9885 & n729;
assign n7962 = ~(n10254 | n1615);
assign n4841 = n4790 & n11775;
assign n2576 = n986 & n1883;
assign n5248 = n2017 | n7315;
assign n5112 = ~(n9107 | n9658);
assign n5384 = n10822 & n3044;
assign n2962 = n2682 & n13192;
assign n2571 = ~n12102;
assign n14234 = n13525 & n4286;
assign n2312 = ~(n14370 | n2024);
assign n6044 = ~n359;
assign n9404 = ~n10714;
assign n991 = n4445 & n12602;
assign n3409 = n8769 & n1306;
assign n9943 = n13656 & n10267;
assign n3413 = ~(n4988 | n4808);
assign n11563 = n11702 & n8958;
assign n1582 = ~n6357;
assign n12031 = n6471 | n9568;
assign n10248 = ~n8737;
assign n714 = n10589 & n3808;
assign n8029 = n14465 & n9800;
assign n4191 = n3164 | n9664;
assign n10146 = n3168 | n13233;
assign n12875 = n7079 & n13196;
assign n12318 = n5999 & n10919;
assign n5412 = ~n8647;
assign n10093 = n8401 & n7493;
assign n12149 = ~n8735;
assign n8200 = n2686 | n16;
assign n11869 = n11438 | n13173;
assign n8572 = ~n13458;
assign n8960 = n12475 & n1653;
assign n13171 = n12953 & n2817;
assign n11600 = n10933 | n13189;
assign n9060 = n11838 & n13817;
assign n2279 = n11011 | n10196;
assign n1869 = ~(n13979 | n7035);
assign n9674 = n8476 | n14375;
assign n13199 = n12400 | n10135;
assign n3515 = n2784 | n9826;
assign n2637 = n12542 & n8445;
assign n5078 = n1202 | n13223;
assign n11982 = n9218 | n13020;
assign n118 = n850 | n9530;
assign n183 = ~n8179;
assign n10719 = ~(n12957 | n13829);
assign n13754 = n13774 | n10339;
assign n6571 = n6899 & n13887;
assign n9157 = n10969 & n4522;
assign n206 = ~(n9291 | n1806);
assign n6479 = n7081 & n13199;
assign n6299 = n10191 | n6029;
assign n11497 = n4913 | n6302;
assign n10592 = n11950 & n8830;
assign n4682 = ~n8341;
assign n223 = n11576 | n2962;
assign n5510 = n7219 | n1956;
assign n6175 = n8964 | n2394;
assign n2038 = n13952 & n12726;
assign n8251 = n7898 | n3353;
assign n11918 = n8452 | n8520;
assign n12 = n11510 | n12349;
assign n10072 = ~n9950;
assign n2014 = ~(n5488 | n2418);
assign n7669 = ~(n12079 | n843);
assign n744 = n1855 & n9317;
assign n4697 = n13537 | n11015;
assign n11141 = n7768 & n5285;
assign n3681 = n1365 & n9214;
assign n6441 = n10357 & n2238;
assign n8995 = n4394 & n3832;
assign n12477 = n4806 & n14054;
assign n12940 = n13850 & n1961;
assign n13707 = ~n3616;
assign n6416 = ~(n12292 | n6194);
assign n11439 = ~(n6074 | n2475);
assign n10052 = n11123 | n14522;
assign n10333 = n10245 | n12833;
assign n4872 = n492 | n14203;
assign n9775 = n9742 | n6002;
assign n11465 = n1140 & n1912;
assign n6396 = n10015 & n11239;
assign n10839 = n5603 | n9816;
assign n10149 = n12870 | n211;
assign n1576 = ~n11541;
assign n6631 = n7081 & n3984;
assign n1204 = n7392 & n6497;
assign n13936 = n1613 | n14407;
assign n5091 = n457 & n1532;
assign n10879 = n1074 & n11871;
assign n13653 = n2387 | n4977;
assign n13691 = n5625 | n8778;
assign n7967 = n10374 & n13349;
assign n5188 = ~n6258;
assign n12201 = n3320 | n6713;
assign n1300 = n2669 & n11985;
assign n8309 = n3736 | n6999;
assign n8542 = n9806 | n6239;
assign n2677 = ~n11066;
assign n13927 = n2236 | n281;
assign n875 = n12633 | n1650;
assign n11963 = n6263 | n3543;
assign n6344 = n10508 | n10201;
assign n948 = n2674 & n10462;
assign n10086 = n4791 | n5629;
assign n4356 = n1805 | n7916;
assign n8125 = n11171 | n337;
assign n647 = ~n12331;
assign n7203 = ~n7940;
assign n13228 = n5489 & n1366;
assign n13335 = n1875 | n12332;
assign n221 = n11094 | n13487;
assign n2826 = n9265 & n11287;
assign n11110 = n5409 | n12466;
assign n6222 = n3586 & n12707;
assign n6080 = n9211 | n9809;
assign n349 = n10922 & n4331;
assign n11626 = n8332 | n11080;
assign n12279 = n1401 & n957;
assign n6016 = ~n4618;
assign n3616 = n1109 & n2343;
assign n1500 = n11438 | n8246;
assign n6874 = ~n7023;
assign n3521 = ~n9377;
assign n3170 = ~(n5762 | n1426);
assign n4995 = n4821 | n6378;
assign n11624 = ~(n5432 | n12932);
assign n7976 = n2897 | n6086;
assign n13619 = n11472 | n1823;
assign n9707 = n7068 & n13671;
assign n10376 = ~n746;
assign n8939 = ~(n5429 | n14136);
assign n13884 = n5234 | n6940;
assign n6020 = ~n7455;
assign n2379 = n2878 | n11224;
assign n3741 = n8517 | n70;
assign n3384 = n7909 & n2501;
assign n5586 = n8552 & n8547;
assign n8224 = n10846 & n11291;
assign n10467 = n7358 | n6818;
assign n9041 = n7255 | n2573;
assign n9742 = ~n13165;
assign n8917 = n12092 & n13813;
assign n9925 = n9422 | n14402;
assign n9009 = n2486 & n3091;
assign n5536 = ~(n6211 | n1319);
assign n9082 = n5695 | n9084;
assign n1090 = ~(n1383 | n14416);
assign n9333 = n766 | n7640;
assign n12540 = n8638 | n3383;
assign n6775 = n11405 | n2812;
assign n528 = n838 | n9330;
assign n11693 = n817 | n967;
assign n9624 = n3485 & n8684;
assign n4618 = ~n11343;
assign n3042 = n6711 | n534;
assign n8167 = n4546 & n7899;
assign n1373 = n8923 & n6811;
assign n10937 = n10032 & n13355;
assign n4158 = n6323 | n8181;
assign n10135 = n8043 & n3390;
assign n9826 = n12259 & n11754;
assign n13303 = n5999 & n2326;
assign n10459 = ~(n8065 | n13958);
assign n9835 = n4486 & n5694;
assign n10188 = n13485 | n3480;
assign n7578 = n695 | n10541;
assign n11740 = n1804 & n563;
assign n3678 = n7812 | n1455;
assign n2590 = n4554 & n9986;
assign n846 = n11176 | n13397;
assign n9973 = n5144 | n1930;
assign n6923 = n3815 | n14012;
assign n11322 = n10408 & n2732;
assign n14218 = n3435 & n4024;
assign n1280 = ~(n6062 | n2880);
assign n4542 = ~(n10936 | n1839);
assign n1756 = n428 & n8961;
assign n6224 = n9345 & n5063;
assign n9112 = n5575 | n3406;
assign n13598 = n7212 | n4355;
assign n5619 = n4156 & n4810;
assign n4704 = n7798 & n10497;
assign n2986 = n781 | n7157;
assign n2597 = ~n8148;
assign n7752 = n12475 & n6213;
assign n10138 = n11020 & n9089;
assign n4692 = ~n3443;
assign n2709 = ~n1571;
assign n11920 = n10134 & n640;
assign n4885 = n5764 & n1815;
assign n11951 = ~n3070;
assign n5589 = n900 | n12868;
assign n13309 = n13525 & n3778;
assign n12484 = n584 | n10704;
assign n1055 = n8769 & n12362;
assign n429 = n9275 & n2056;
assign n3135 = n492 | n8532;
assign n12836 = n11636 & n2867;
assign n13533 = n8427 & n4085;
assign n11913 = n2645 | n9294;
assign n7415 = n14120 & n2074;
assign n4798 = n766 | n9267;
assign n3559 = ~n1214;
assign n1451 = n13359 & n2286;
assign n7390 = n4447 | n5023;
assign n11814 = ~n13038;
assign n9843 = n12047 | n4548;
assign n3499 = n8213 & n13635;
assign n3689 = n10523 | n9938;
assign n12673 = ~n7814;
assign n3226 = ~(n478 | n453);
assign n12510 = n10394 | n4271;
assign n13611 = n2025 | n11102;
assign n5486 = ~n3776;
assign n334 = ~(n6085 | n5916);
assign n4884 = n11313 & n11659;
assign n10529 = ~n3344;
assign n11463 = n13364 & n3217;
assign n14233 = n12130 | n276;
assign n4642 = n9564 & n10213;
assign n5165 = n12101 & n11247;
assign n12000 = n6130 & n9753;
assign n1872 = n1662 & n5615;
assign n6919 = n865 & n2342;
assign n10682 = n6744 & n7897;
assign n3695 = n13860 & n8562;
assign n1039 = n234 | n10148;
assign n7891 = n501 & n6533;
assign n3307 = n5570 | n3339;
assign n352 = ~(n5132 | n10709);
assign n651 = ~(n1028 | n6715);
assign n14178 = ~n11404;
assign n4323 = n6857 | n7645;
assign n13496 = n5628 & n3072;
assign n9638 = n6596 | n6665;
assign n9944 = ~n12930;
assign n1753 = n6854 & n8924;
assign n12645 = n9285 | n5245;
assign n12860 = ~(n10323 | n1865);
assign n7863 = n5335 & n13936;
assign n399 = ~(n573 | n12492);
assign n4902 = n13342 & n12479;
assign n1643 = n11724 | n3451;
assign n11541 = n7676 & n8341;
assign n5604 = n7203 & n9358;
assign n5447 = n7211 & n6950;
assign n4507 = ~(n8527 | n8420);
assign n5905 = n3222 & n13968;
assign n204 = n1775 & n8570;
assign n12324 = ~n4550;
assign n9162 = n10191 | n635;
assign n7029 = n9716 | n3140;
assign n6730 = ~n81;
assign n629 = n504 | n11416;
assign n9381 = n8213 & n9048;
assign n4328 = n11336 & n4936;
assign n1512 = n839 | n11995;
assign n11152 = n3976 & n8220;
assign n1444 = n9230 | n6954;
assign n874 = n13227 & n594;
assign n5123 = n6288 | n5519;
assign n6303 = n457 & n6547;
assign n4004 = n9191 & n548;
assign n3372 = ~(n5065 | n8180);
assign n12017 = n9620 | n4893;
assign n5683 = n11392 | n11854;
assign n68 = ~(n11232 | n8762);
assign n11746 = n4052 | n13876;
assign n11381 = n13656 & n7872;
assign n13756 = n3958 | n1265;
assign n6666 = n12832 & n10315;
assign n10973 = ~n637;
assign n10268 = n808 & n6156;
assign n1002 = n4614 & n11326;
assign n5281 = n333 & n7408;
assign n9309 = ~(n2086 | n7431);
assign n2846 = ~n5435;
assign n11064 = n10516 & n2977;
assign n14349 = n13516 | n4389;
assign n838 = ~n9169;
assign n3782 = n6519 | n8156;
assign n3599 = n4877 | n7414;
assign n12654 = ~(n10309 | n11732);
assign n2029 = n3222 | n8315;
assign n11427 = ~(n1378 | n2390);
assign n8337 = ~n3155;
assign n13976 = n9747 | n1886;
assign n9771 = n3886 | n2228;
assign n5817 = n5472 | n9965;
assign n10465 = ~n7660;
assign n10410 = n4932 & n4683;
assign n13581 = n2761 | n7751;
assign n711 = n8575 | n12720;
assign n9080 = ~n7662;
assign n4607 = ~(n11047 | n708);
assign n1433 = n9035 | n52;
assign n14150 = ~n2417;
assign n8055 = n6867 | n12386;
assign n8293 = n8692 & n11149;
assign n4934 = n8582 | n9460;
assign n6967 = n8517 | n879;
assign n4083 = n2877 | n11060;
assign n14355 = n13501 | n6538;
assign n3657 = n8490 | n4392;
assign n7905 = ~n8631;
assign n13860 = ~n3313;
assign n9018 = n13755 & n10729;
assign n12572 = n11362 | n5725;
assign n9591 = n12013 & n59;
assign n9746 = n10913 | n6540;
assign n9317 = n8376 & n3113;
assign n3299 = n11300 & n9341;
assign n5827 = ~(n5715 | n5289);
assign n336 = n13096 & n6334;
assign n10784 = ~n3070;
assign n6168 = n4898 | n8457;
assign n3621 = ~(n7365 | n6345);
assign n4652 = ~(n2932 | n665);
assign n7187 = ~n11861;
assign n4167 = n7026 & n1593;
assign n13637 = ~(n9657 | n12911);
assign n13002 = ~n4082;
assign n3608 = ~n13000;
assign n12019 = ~n12444;
assign n1565 = n1834 | n14427;
assign n8109 = n8605 & n12560;
assign n10942 = n3743 & n13845;
assign n2890 = n5647 | n11408;
assign n3790 = n1006 | n2294;
assign n2754 = n1147 | n8005;
assign n1227 = n5764 & n12164;
assign n9997 = n8043 & n7399;
assign n2533 = ~n8122;
assign n1655 = n6013 & n9973;
assign n12544 = n11183 | n8632;
assign n7249 = ~n10889;
assign n5676 = ~(n4491 | n792);
assign n7818 = ~n11590;
assign n7877 = n9944 & n1574;
assign n6012 = n5225 & n11987;
assign n10727 = n12998 & n10740;
assign n11722 = ~n12776;
assign n572 = n100 | n2975;
assign n942 = n9898 & n10491;
assign n9954 = n9078 | n10228;
assign n8299 = n7700 | n5790;
assign n7144 = n13464 & n6297;
assign n4712 = n1588 & n6543;
assign n2772 = n6498 | n5430;
assign n5735 = ~(n11047 | n5915);
assign n12704 = n4803 & n6535;
assign n13943 = n8969 | n8646;
assign n13939 = ~(n4988 | n1822);
assign n4586 = n4574 & n8285;
assign n3635 = ~n5675;
assign n305 = n5548 | n6361;
assign n669 = n5710 | n5308;
assign n11302 = ~n13981;
assign n14326 = n2091 | n11590;
assign n4464 = ~n1076;
assign n2938 = n8209 | n4613;
assign n9424 = n695 | n4440;
assign n5290 = n6157 & n8202;
assign n12841 = n13246 & n10677;
assign n7670 = ~n1495;
assign n14512 = ~n6765;
assign n9456 = ~n4324;
assign n7294 = n13518 | n9334;
assign n10175 = n9015 & n10451;
assign n4228 = n13078 & n13623;
assign n6281 = n706 & n8956;
assign n10495 = ~(n4105 | n857);
assign n6196 = ~n1771;
assign n9780 = ~n7875;
assign n5365 = ~n670;
assign n6645 = n7767 & n6789;
assign n4714 = n2686 | n2528;
assign n6530 = n5236 | n9016;
assign n12531 = ~n6559;
assign n13705 = n3394 | n13871;
assign n6686 = n2082 & n621;
assign n5561 = n889 & n8636;
assign n8340 = n4498 | n14207;
assign n13801 = n11315 | n8948;
assign n4134 = ~n7754;
assign n2147 = n4233 | n8591;
assign n4923 = ~n9596;
assign n5560 = n6531 & n12556;
assign n4155 = n10781 | n11160;
assign n11426 = n9941 & n459;
assign n836 = n5553 & n5189;
assign n13709 = ~(n4233 | n1627);
assign n6508 = n9269 | n1549;
assign n8620 = ~n5601;
assign n3788 = n11739 | n1353;
assign n354 = n12461 & n3102;
assign n8326 = n11495 & n6437;
assign n6111 = ~n2320;
assign n12848 = n4347 & n10286;
assign n2347 = n3097 & n7515;
assign n7229 = ~n628;
assign n2011 = n10025 & n2611;
assign n8562 = n6205 | n7923;
assign n7403 = ~(n9529 | n6075);
assign n11059 = n3273 | n13073;
assign n487 = n7912 | n1980;
assign n673 = ~n10255;
assign n5678 = n1447 | n10283;
assign n1746 = n8151 | n388;
assign n9802 = n2412 | n10759;
assign n1838 = ~n8735;
assign n5475 = ~n5951;
assign n199 = ~(n7448 | n8794);
assign n14351 = ~n11668;
assign n3027 = ~(n2009 | n3760);
assign n632 = n9226 | n1533;
assign n8243 = n4821 | n14218;
assign n13010 = n10061 & n489;
assign n9545 = n12445 & n3150;
assign n8551 = ~(n4092 | n6790);
assign n8699 = n6046 | n7583;
assign n13008 = n13597 & n7173;
assign n4199 = ~n13696;
assign n5280 = n9069 & n12424;
assign n12667 = n13781 & n3949;
assign n10413 = n4554 & n4041;
assign n12400 = ~n2934;
assign n11170 = n12759 | n12516;
assign n14322 = n11980 | n13778;
assign n7999 = ~(n7519 | n7458);
assign n1774 = n6205 | n14325;
assign n7628 = n10351 | n8229;
assign n14345 = n12820 | n14143;
assign n12369 = n4844 & n1116;
assign n11553 = n4880 & n13475;
assign n636 = ~n4000;
assign n2016 = ~n12746;
assign n9199 = n13083 | n13798;
assign n597 = n13433 & n10011;
assign n1821 = ~n10108;
assign n289 = n4546 & n4796;
assign n963 = n11223 | n13309;
assign n11804 = ~n5242;
assign n3628 = ~n498;
assign n5747 = ~(n1342 | n4917);
assign n2557 = n533 & n973;
assign n4932 = ~n1784;
assign n4616 = n2089 | n6006;
assign n1908 = n12779 | n977;
assign n6485 = n1875 | n12610;
assign n8225 = n9804 | n3514;
assign n10469 = ~n10965;
assign n2241 = ~n1311;
assign n3525 = n7250 | n6915;
assign n5835 = n1613 | n8167;
assign n12134 = n89 | n9455;
assign n1750 = n10449 | n13488;
assign n3736 = ~n12218;
assign n308 = n2531 | n13587;
assign n8662 = n3435 & n4723;
assign n13497 = n1354 & n5962;
assign n7893 = n6649 & n9788;
assign n8003 = n14074 & n11283;
assign n4308 = n2724 & n7271;
assign n14380 = n9323 & n9782;
assign n11209 = n2527 & n1163;
assign n3098 = n10784 | n5436;
assign n7725 = ~(n8701 | n9436);
assign n11166 = n8969 | n9904;
assign n3558 = n6090 | n5386;
assign n7434 = n5468 | n1952;
assign n9932 = n11329 & n3589;
assign n2319 = n4614 & n13388;
assign n4331 = n11440 | n4316;
assign n12623 = n3169 & n851;
assign n1211 = n6891 | n11741;
assign n9363 = n4508 | n8852;
assign n12401 = ~n628;
assign n11476 = n1610 & n2489;
assign n2574 = ~(n10342 | n4259);
assign n10366 = n1266 & n12406;
assign n5263 = n11315 | n8559;
assign n9530 = n10229 & n2253;
assign n3146 = ~(n5715 | n4610);
assign n9214 = n888 & n1401;
assign n6761 = n9898 & n434;
assign n9151 = ~n14154;
assign n444 = n2387 | n10807;
assign n8269 = ~(n12248 | n12348);
assign n10884 = n7862 | n4350;
assign n8469 = n6596 | n12841;
assign n395 = n3715 & n10863;
assign n4893 = n8007 & n5889;
assign n6060 = n10229 & n8037;
assign n2282 = n769 | n7454;
assign n10600 = n5335 & n6219;
assign n11763 = n494 & n12995;
assign n5354 = ~n9967;
assign n6101 = n13297 & n10467;
assign n1810 = n1582 | n12181;
assign n6239 = ~(n6679 | n6421);
assign n10596 = n14109 & n6518;
assign n9088 = ~(n13153 | n12347);
assign n7906 = n392 & n6142;
assign n11366 = n11036 | n1982;
assign n3110 = n9151 | n12383;
assign n3068 = n10929 | n12097;
assign n2086 = ~n12444;
assign n14328 = n10084 & n4017;
assign n9657 = ~n10617;
assign n6609 = ~n920;
assign n10432 = n1391 | n39;
assign n4991 = n7612 & n4704;
assign n8639 = n11420 | n1488;
assign n903 = ~(n9984 | n5718);
assign n6954 = n9617 & n7910;
assign n5707 = n2111 | n6913;
assign n9938 = n8923 & n4914;
assign n7701 = ~(n6905 | n3027);
assign n3696 = ~n5221;
assign n13915 = n10960 | n7312;
assign n6393 = n11569 & n811;
assign n12351 = ~n9878;
assign n7085 = n10024 | n1618;
assign n10358 = ~n4633;
assign n4705 = ~(n1028 | n6613);
assign n3504 = n14063 & n4707;
assign n6133 = ~(n6971 | n11578);
assign n1257 = ~(n194 | n7008);
assign n6003 = n13276 | n13878;
assign n8344 = n1613 | n10587;
assign n4954 = n2904 & n1039;
assign n1020 = n4602 | n6079;
assign n13543 = n4104 & n13449;
assign n11245 = n1254 & n13879;
assign n10528 = ~(n14238 | n3906);
assign n14231 = n5587 | n13674;
assign n1386 = n7803 | n14493;
assign n12157 = n12295 | n2832;
assign n10767 = ~n12522;
assign n2194 = ~n8631;
assign n7077 = n7484 & n7502;
assign n11884 = n4435 | n3499;
assign n10081 = n8480 | n1528;
assign n1749 = n9811 & n1102;
assign n1202 = ~n7289;
assign n8654 = n6373 | n10038;
assign n1368 = n6051 & n3184;
assign n8504 = ~(n5848 | n399);
assign n3115 = n5480 | n9251;
assign n800 = n1711 | n3983;
assign n3881 = n1728 | n12928;
assign n299 = ~(n5504 | n7340);
assign n2316 = n5188 | n2334;
assign n7096 = n8045 | n6273;
assign n12795 = n9321 & n6469;
assign n4999 = n4791 | n7831;
assign n10585 = n3047 | n13463;
assign n3492 = ~n2164;
assign n2995 = n6697 & n1975;
assign n5505 = ~n10099;
assign n12426 = n10857 | n1157;
assign n3975 = n11313 & n8075;
assign n13710 = n9345 & n1499;
assign n7888 = ~n11331;
assign n9250 = n7693 & n12302;
assign n1022 = n11584 | n9871;
assign n1789 = n10784 | n9813;
assign n4866 = n10808 | n10872;
assign n6647 = n3435 & n4961;
assign n9808 = n8964 | n5568;
assign n6145 = n12202 & n983;
assign n4874 = n13107 & n10316;
assign n4300 = ~n10372;
assign n4577 = n14313 & n10887;
assign n1498 = n11804 | n7895;
assign n7046 = n4562 | n5961;
assign n5915 = ~(n3428 | n8086);
assign n10665 = n3986 & n12157;
assign n5375 = n4790 & n8171;
assign n7083 = n13941 | n8709;
assign n6563 = n13227 & n7666;
assign n12672 = ~(n10289 | n5879);
assign n8174 = n13142 | n6174;
assign n834 = n12037 & n3879;
assign n7554 = n11542 | n1169;
assign n7753 = n13518 | n5399;
assign n13859 = n1247 & n8355;
assign n7682 = n11384 | n6147;
assign n15 = ~n9563;
assign n2214 = n13338 & n780;
assign n11431 = n49 | n6220;
assign n244 = ~(n9807 | n12330);
assign n3487 = ~(n9567 | n5005);
assign n13894 = ~(n5172 | n4651);
assign n13468 = n3527 | n9897;
assign n2492 = n12683 & n7099;
assign n4177 = n12015 & n12215;
assign n8218 = n10197 & n8501;
assign n2644 = ~n2723;
assign n12637 = ~(n9423 | n9506);
assign n3642 = ~(n7920 | n4477);
assign n9955 = n14157 & n7478;
assign n3024 = n8458 | n12689;
assign n2126 = n4895 & n3798;
assign n3442 = n1705 | n11529;
assign n5527 = ~(n3344 | n2769);
assign n1282 = n13575 & n1177;
assign n6477 = ~(n3871 | n2813);
assign n14221 = n7245 | n6282;
assign n10056 = n10781 | n4598;
assign n1620 = n8232 & n9551;
assign n1811 = n1697 | n5325;
assign n11712 = n13407 & n1144;
assign n8377 = n9321 & n5373;
assign n1677 = ~n8884;
assign n3641 = n6672 | n1017;
assign n2231 = n9285 | n8599;
assign n8623 = n648 | n6776;
assign n11946 = ~(n13941 | n14300);
assign n12332 = n11950 & n8757;
assign n9971 = n12768 & n8868;
assign n4196 = ~(n13675 | n5722);
assign n8919 = n5012 & n11082;
assign n12189 = ~n5288;
assign n2755 = n3877 | n12074;
assign n4385 = n12768 & n8537;
assign n449 = n5575 | n3468;
assign n10975 = ~n2202;
assign n11009 = n6128 & n12426;
assign n13119 = n2750 | n5405;
assign n14211 = n12764 | n7059;
assign n3344 = ~n5886;
assign n1245 = n14313 & n7494;
assign n4520 = n13404 & n2003;
assign n12613 = n89 | n14396;
assign n12411 = n13130 | n13391;
assign n13673 = n12998 & n14288;
assign n8863 = ~(n2780 | n7439);
assign n14397 = n3569 | n11278;
assign n13576 = n14404 | n3077;
assign n4849 = n4435 | n9619;
assign n12960 = ~n5852;
assign n7030 = ~(n3870 | n8190);
assign n1752 = n13226 | n626;
assign n3370 = ~n5460;
assign n5084 = ~n777;
assign n14476 = ~(n2790 | n13839);
assign n6843 = n12633 | n6542;
assign n3268 = ~n3402;
assign n11899 = n79 & n2704;
assign n12700 = ~(n11558 | n7557);
assign n4166 = n98 & n14027;
assign n11130 = n7389 | n8997;
assign n14318 = ~(n8189 | n2798);
assign n340 = n69 | n9180;
assign n14009 = ~n6147;
assign n6989 = n9154 | n3833;
assign n13092 = n11951 | n11539;
assign n7237 = n898 & n5508;
assign n6076 = n4803 & n13938;
assign n13125 = n8983 | n14114;
assign n1632 = n974 | n5729;
assign n9789 = n13485 | n9625;
assign n4590 = n2783 & n1738;
assign n6568 = n6596 | n11317;
assign n12659 = n2236 | n14436;
assign n13594 = n13676 & n11821;
assign n12160 = n4690 & n2375;
assign n3476 = n6971 | n11723;
assign n8840 = ~(n7551 | n2163);
assign n4222 = n5823 & n252;
assign n6617 = n8432 & n10127;
assign n12750 = n1247 & n11138;
assign n4267 = ~n13992;
assign n3933 = n8986 | n11374;
assign n726 = n3401 & n6435;
assign n430 = ~(n10342 | n4086);
assign n8931 = n5823 & n14420;
assign n5821 = n5926 & n14491;
assign n12343 = n8242 | n8644;
assign n3989 = n2845 | n12142;
assign n11013 = n9315 & n11177;
assign n13786 = n10224 | n313;
assign n4270 = ~n12409;
assign n5540 = ~(n6426 | n2133);
assign n3258 = n14366 | n4884;
assign n6619 = n3569 | n2138;
assign n4197 = n7627 & n11970;
assign n14216 = ~n14365;
assign n1051 = ~n918;
assign n10066 = n13074 | n6043;
assign n1638 = ~n5333;
assign n5824 = ~(n13310 | n9732);
assign n1352 = n11838 & n13384;
assign n7117 = n12741 & n12382;
assign n9804 = ~n8813;
assign n11349 = n12542 & n6959;
assign n6141 = ~(n2212 | n4766);
assign n9725 = n12695 | n12071;
assign n7931 = n8721 & n2193;
assign n4383 = ~(n13522 | n2312);
assign n7959 = n9265 & n6230;
assign n641 = n5454 | n8859;
assign n7348 = n12250 & n3074;
assign n3543 = n7043 & n150;
assign n5047 = n222 & n12724;
assign n10756 = n9742 | n6065;
assign n5367 = n776 & n2231;
assign n14117 = ~(n4200 | n11910);
assign n5649 = ~(n8277 | n9841);
assign n13143 = n1494 | n7893;
assign n12951 = n14481 | n7958;
assign n5677 = n9226 | n14380;
assign n1939 = n2055 | n6993;
assign n2141 = n1772 & n4931;
assign n7517 = n1261 | n4845;
assign n1319 = ~(n8527 | n4836);
assign n6744 = ~n10828;
assign n8752 = ~n11617;
assign n2953 = ~n6067;
assign n7707 = n7060 & n9394;
assign n11056 = ~(n7418 | n4396);
assign n11940 = n9617 & n13250;
assign n7501 = n1356 | n5723;
assign n1250 = n13130 | n6071;
assign n13393 = n1669 | n6988;
assign n1418 = n8238 & n5797;
assign n12983 = n10229 & n14062;
assign n13638 = n13078 & n9789;
assign n7052 = ~n13135;
assign n12233 = n14088 | n12000;
assign n9727 = ~(n3107 | n8534);
assign n12844 = ~n4777;
assign n11271 = n6471 | n7566;
assign n9950 = ~n13725;
assign n2824 = n1254 & n12377;
assign n6749 = n8828 | n2156;
assign n6684 = n1071 & n10645;
assign n8098 = n10408 & n13589;
assign n7158 = n10506 & n2416;
assign n2676 = n5048 & n4537;
assign n3649 = n2686 | n1625;
assign n4930 = n808 & n10488;
assign n8157 = n11142 & n10777;
assign n1155 = n9972 & n14453;
assign n11227 = n6703 | n3893;
assign n8323 = n12023 | n8531;
assign n9871 = ~n13257;
assign n1459 = n10302 & n7735;
assign n12064 = n14188 | n9656;
assign n12791 = n9297 & n14256;
assign n7455 = ~n1378;
assign n7686 = n10516 & n9535;
assign n13633 = n787 | n462;
assign n10084 = ~n10376;
assign n14454 = n1452 & n7373;
assign n4382 = ~n8262;
assign n4968 = n8242 | n3713;
assign n1879 = n14446 & n5114;
assign n5031 = n3435 & n8862;
assign n7051 = n10294 | n11161;
assign n2730 = n9151 | n6166;
assign n14370 = ~n2472;
assign n2916 = n1582 | n5516;
assign n6253 = n7229 | n3666;
assign n9882 = n11379 | n14253;
assign n4826 = n4807 | n2157;
assign n4283 = ~(n5391 | n4523);
assign n11661 = n7212 | n11514;
assign n2703 = ~(n3019 | n11496);
assign n4183 = ~(n7130 | n2075);
assign n9020 = n695 | n13710;
assign n10838 = n11576 | n1289;
assign n1308 = n12013 & n13852;
assign n14093 = ~n442;
assign n3233 = n7590 | n7450;
assign n7526 = n1362 | n12961;
assign n3542 = n6600 | n14475;
assign n10289 = ~n14154;
assign n9523 = n2783 & n11366;
assign n2954 = n480 | n5539;
assign n3054 = ~n1462;
assign n7735 = n8242 | n5411;
assign n5738 = ~n12107;
assign n5727 = n3932 & n9043;
assign n12740 = ~(n2016 | n2344);
assign n13527 = n1775 & n3819;
assign n6230 = n10191 | n12791;
assign n1976 = ~(n11309 | n1091);
assign n13794 = n9507 | n9979;
assign n13759 = ~n7027;
assign n11323 = n2149 | n10813;
assign n600 = ~n10046;
assign n8131 = n2925 & n1946;
assign n5249 = n11183 | n12151;
assign n5904 = ~n5149;
assign n9213 = ~(n5197 | n13893);
assign n12107 = ~n11426;
assign n1066 = n10834 | n4291;
assign n11383 = n1189 | n11368;
assign n4130 = n5084 | n11487;
assign n14517 = ~(n3132 | n4287);
assign n6280 = n8007 & n762;
assign n11679 = ~n10376;
assign n10875 = n1834 | n6701;
assign n13122 = n11033 & n6767;
assign n6417 = n3212 & n994;
assign n6195 = ~(n13677 | n1263);
assign n9155 = n2064 & n7253;
assign n3377 = n6753 & n11921;
assign n10766 = n11157 & n3758;
assign n1651 = n6781 | n2736;
assign n19 = n12858 & n8773;
assign n6374 = ~(n13707 | n6407);
assign n8941 = n6242 | n7952;
assign n2003 = n11285 | n2426;
assign n13256 = n14404 | n11996;
assign n403 = n1431 & n12674;
assign n4482 = n5710 | n1573;
assign n1584 = n4261 & n1105;
assign n11010 = n9898 & n3259;
assign n4975 = n5414 & n7141;
assign n14230 = n6192 & n8042;
assign n1407 = n10015 & n6704;
assign n10029 = ~(n7920 | n12133);
assign n2350 = ~(n11988 | n6893);
assign n3016 = n3826 | n11826;
assign n10571 = ~n6536;
assign n949 = ~(n183 | n9744);
assign n7133 = n3076 | n8597;
assign n9370 = n12741 & n804;
assign n9371 = n12345 & n3946;
assign n13484 = ~n9994;
assign n6049 = n8801 & n7378;
assign n7569 = n14120 & n11458;
assign n8475 = n8378 | n1550;
assign n2186 = ~(n8301 | n12780);
assign n670 = ~n5118;
assign n12071 = n14157 & n14342;
assign n6740 = n2272 | n3950;
assign n9730 = n12500 | n7855;
assign n5841 = n1701 | n6881;
assign n6088 = ~n9971;
assign n937 = n10360 & n2080;
assign n7630 = n8300 & n12306;
assign n6492 = n12265 & n8781;
assign n2031 = n8034 | n8028;
assign n776 = ~n2744;
assign n5454 = ~n8695;
assign n8541 = n8476 | n9573;
assign n928 = ~(n10136 | n6949);
assign n6762 = n3401 & n8350;
assign n10030 = ~(n234 | n14126);
assign n14360 = ~n4895;
assign n14445 = n6730 | n12152;
assign n11409 = n7803 | n6306;
assign n7480 = n4359 & n8505;
assign n3477 = n904 & n13287;
assign n5410 = ~(n3876 | n8895);
assign n2331 = n2562 | n4734;
assign n3137 = n5084 | n3412;
assign n7607 = n1362 | n6385;
assign n8543 = ~n9172;
assign n3931 = n10197 & n1416;
assign n14300 = ~(n3395 | n4792);
assign n9313 = n2597 | n4094;
assign n7015 = ~n7146;
assign n4983 = n10556 & n5124;
assign n11915 = ~(n7334 | n2434);
assign n2382 = n533 & n13770;
assign n8641 = n10332 & n11340;
assign n740 = ~(n4534 | n4694);
assign n2665 = n13863 & n1634;
assign n9744 = n10458 & n7824;
assign n6306 = n12935 & n8804;
assign n5871 = ~n6451;
assign n2246 = ~n2484;
assign n11365 = n2367 & n8273;
assign n11871 = n2750 | n7699;
assign n9905 = n12990 & n947;
assign n7271 = n1198 | n202;
assign n7374 = n12092 & n10217;
assign n1720 = n4098 & n422;
assign n8868 = n11738 & n6861;
assign n1114 = n5625 | n1450;
assign n2561 = ~(n5986 | n7422);
assign n2875 = ~n11493;
assign n1481 = ~n11259;
assign n7732 = n13080 | n4837;
assign n11199 = n251 | n13891;
assign n5985 = n1876 & n1066;
assign n11784 = n2089 | n7712;
assign n22 = n12808 | n13890;
assign n4724 = n9716 | n9189;
assign n6752 = n3028 & n2172;
assign n4942 = n2857 | n2026;
assign n10522 = n6130 & n5995;
assign n11622 = n11142 & n4735;
assign n7887 = ~n9169;
assign n531 = n9650 & n2810;
assign n13138 = n7957 & n9839;
assign n7381 = n7810 & n3697;
assign n1950 = n412 | n2797;
assign n812 = n9944 & n11199;
assign n8831 = n1834 | n3082;
assign n13667 = n11748 & n4293;
assign n4743 = n10062 | n997;
assign n8660 = n904 & n4754;
assign n4066 = n10626 | n10601;
assign n1640 = ~n7972;
assign n3357 = n14219 & n4765;
assign n5908 = n10650 | n6074;
assign n10273 = n4806 & n11829;
assign n3670 = ~(n4913 | n9088);
assign n11279 = n11621 | n4846;
assign n10471 = n3332 & n2427;
assign n11934 = n12425 & n6169;
assign n8093 = n8638 | n3452;
assign n7494 = n11231 | n13582;
assign n5237 = ~n4146;
assign n10064 = n954 | n6929;
assign n3095 = n14029 | n2863;
assign n6866 = n13246 & n1485;
assign n5632 = n14366 | n1049;
assign n1608 = n2784 | n5264;
assign n4502 = ~n8002;
assign n12852 = ~n6791;
assign n7378 = n4045 | n13395;
assign n11587 = ~(n12136 | n3260);
assign n11225 = n6167 & n13808;
assign n12872 = ~n3918;
assign n4532 = n5647 | n2301;
assign n12770 = n100 | n2987;
assign n2970 = n6554 & n5595;
assign n3923 = ~n9416;
assign n14364 = n5450 | n12810;
assign n13233 = n7060 & n9602;
assign n8296 = n6690 | n5378;
assign n7826 = ~n6113;
assign n5062 = ~n2692;
assign n7389 = ~n3263;
assign n8261 = n12401 | n1043;
assign n9164 = n7527 | n11631;
assign n1896 = n1452 & n340;
assign n13037 = ~n11842;
assign n6979 = n8635 & n7999;
assign n4768 = n4581 & n891;
assign n12771 = n12935 & n139;
assign n13110 = n100 | n13398;
assign n13850 = ~n13181;
assign n10046 = ~n5429;
assign n10675 = n10457 & n9695;
assign n12936 = ~(n512 | n14336);
assign n10434 = n7673 & n14506;
assign n2414 = n7957 & n2478;
assign n9414 = ~n10341;
assign n1009 = n10367 & n12676;
assign n10982 = n12494 | n5421;
assign n10211 = n8513 | n11414;
assign n12708 = ~(n788 | n676);
assign n6661 = n5764 & n4226;
assign n11310 = n11313 & n3786;
assign n12785 = n8252 & n10998;
assign n14173 = n5012 & n2117;
assign n9497 = n10857 | n13296;
assign n10190 = n2158 & n5336;
assign n3566 = n12986 & n3085;
assign n1431 = ~n11668;
assign n10369 = n7156 | n13264;
assign n2034 = ~(n7179 | n9526);
assign n2431 = ~(n11285 | n818);
assign n8573 = ~(n8701 | n3991);
assign n735 = n1071 & n11708;
assign n9948 = ~(n10400 | n13238);
assign n12240 = n3914 | n97;
assign n5828 = n7697 | n10925;
assign n3936 = n5553 & n2921;
assign n2427 = n7530 | n3478;
assign n11421 = n10767 & n2567;
assign n8471 = n9544 & n7799;
assign n468 = n13863 & n605;
assign n2868 = ~n6053;
assign n10520 = n7914 | n958;
assign n9612 = ~(n11488 | n1910);
assign n10418 = n2322 & n6651;
assign n6347 = n573 | n204;
assign n5448 = n9015 & n5495;
assign n2793 = n13847 | n4566;
assign n10060 = n8232 & n1443;
assign n1479 = n930 | n11942;
assign n1394 = n12764 | n1949;
assign n11713 = ~n9721;
assign n6741 = n200 & n6911;
assign n9770 = n11710 | n8934;
assign n814 = n523 | n6808;
assign n12485 = n11551 | n2525;
assign n8155 = n9275 & n6238;
assign n9828 = n10019 | n10596;
assign n13090 = n1729 & n10928;
assign n9448 = n2412 | n7990;
assign n14438 = n2531 | n8152;
assign n10891 = n11183 | n9286;
assign n3167 = n5641 | n9895;
assign n3120 = ~n9354;
assign n8438 = n5007 | n1287;
assign n2176 = n8512 & n945;
assign n7253 = n14337 | n2539;
assign n5297 = n3826 | n8236;
assign n3069 = n8025 & n2053;
assign n11890 = n8490 | n3223;
assign n11760 = n8701 | n8455;
assign n3387 = n3672 & n7182;
assign n9520 = ~(n7683 | n13648);
assign n10001 = ~(n7588 | n12740);
assign n9878 = n9350 & n9640;
assign n3873 = ~n2409;
assign n8524 = ~n10787;
assign n6905 = ~n5151;
assign n14344 = n3332 & n875;
assign n11452 = n350 | n9977;
assign n11307 = n3888 | n8756;
assign n9452 = n4481 | n14061;
assign n4912 = n1772 & n3393;
assign n11518 = n11440 | n58;
assign n5967 = n2874 | n5437;
assign n10041 = ~(n3309 | n7013);
assign n11996 = n8047 & n696;
assign n951 = n4929 & n9014;
assign n6860 = n8638 | n5726;
assign n10734 = n9238 & n3243;
assign n7012 = n7779 & n10021;
assign n8096 = ~n1060;
assign n4933 = n3986 & n5286;
assign n4178 = n12351 | n8930;
assign n13585 = ~(n7971 | n3439);
assign n7791 = n3766 & n1412;
assign n7937 = n14446 & n14511;
assign n5336 = n11176 | n4862;
assign n9879 = ~(n13477 | n13586);
assign n9007 = n9232 & n2455;
assign n8276 = ~(n4296 | n8231);
assign n111 = n1391 | n10755;
assign n6257 = n12844 | n11417;
assign n8280 = n5553 & n4879;
assign n3583 = n12900 & n7476;
assign n3366 = ~n2048;
assign n7696 = ~n4047;
assign n13019 = n10234 | n1406;
assign n9929 = n4923 | n8082;
assign n8835 = n1741 | n5600;
assign n5347 = n2758 & n5998;
assign n12409 = n11837 & n7567;
assign n10707 = n9780 | n6200;
assign n7235 = n3710 & n11874;
assign n1574 = n2562 | n12702;
assign n2998 = ~n13383;
assign n12968 = ~n2383;
assign n7103 = n11406 & n8016;
assign n826 = n2643 & n13809;
assign n1929 = ~n6670;
assign n13671 = n9429 | n12326;
assign n12664 = ~(n14368 | n6686);
assign n7002 = n6316 & n9849;
assign n2193 = n3492 & n12572;
assign n376 = n14472 | n10894;
assign n12414 = ~n7441;
assign n7766 = n6206 | n1154;
assign n7243 = n11621 | n8563;
assign n542 = n1821 | n4336;
assign n6284 = ~(n13941 | n13353);
assign n7295 = n7443 & n11611;
assign n7614 = ~(n7334 | n613);
assign n13563 = n8701 | n8482;
assign n5276 = n12057 & n11860;
assign n11725 = n4908 | n7603;
assign n1382 = ~(n7940 | n12269);
assign n6727 = n2897 | n12941;
assign n14143 = n8025 & n5620;
assign n7038 = n185 | n2425;
assign n7663 = ~(n2790 | n5404);
assign n897 = n3952 & n8383;
assign n12522 = ~n6055;
assign n10809 = n511 | n9045;
assign n7087 = n10846 & n7390;
assign n8820 = n9856 | n7061;
assign n11254 = n446 & n3579;
assign n1440 = n1071 & n8740;
assign n3064 = n10516 & n5150;
assign n6640 = ~n12270;
assign n2802 = n4527 | n3652;
assign n5073 = n11839 | n10214;
assign n894 = n2587 & n8150;
assign n929 = n7934 | n1776;
assign n7568 = n9375 | n4489;
assign n10002 = n11837 & n7266;
assign n4751 = n14042 & n12093;
assign n5279 = ~n9456;
assign n9409 = n5823 & n12786;
assign n3185 = n4655 & n1355;
assign n9146 = n5815 | n7144;
assign n3078 = n2064 & n12558;
assign n8300 = ~n9416;
assign n1435 = n6128 & n306;
assign n2138 = n7826 & n9975;
assign n12897 = ~n1742;
assign n1626 = ~(n14419 | n10519);
assign n14366 = ~n4777;
assign n9434 = n783 & n1917;
assign n14186 = ~(n12705 | n12956);
assign n11488 = ~n8027;
assign n3452 = n4163 & n13026;
assign n11386 = n9780 | n9369;
assign n13605 = n3768 | n8080;
assign n12376 = n536 & n7568;
assign n2893 = n13806 | n2635;
assign n12505 = n13005 | n7388;
assign n13862 = n8252 | n203;
assign n8967 = n12620 & n13642;
assign n8087 = n1061 | n6008;
assign n4475 = n12092 & n11565;
assign n1581 = n10289 | n1304;
assign n3728 = n8828 | n11436;
assign n10782 = ~(n3768 | n1050);
assign n5869 = n12832 & n3136;
assign n10658 = n5570 | n3315;
assign n5930 = n2021 & n960;
assign n12752 = n6311 & n3376;
assign n9572 = n231 & n3866;
assign n11316 = ~n7681;
assign n13751 = n7627 & n60;
assign n9415 = n10825 | n14255;
assign n3038 = n7971 | n14122;
assign n14252 = ~n5033;
assign n3698 = n2888 | n1204;
assign n13805 = n390 | n7201;
assign n1281 = n12821 | n11532;
assign n9069 = ~n3967;
assign n5535 = n9952 & n5445;
assign n13340 = ~(n6039 | n13265);
assign n3217 = ~(n12179 | n8222);
assign n14033 = n8401 & n6493;
assign n4920 = n7443 & n7629;
assign n13515 = n11472 | n8318;
assign n10438 = n8452 | n11467;
assign n6501 = ~(n5840 | n10733);
assign n1792 = n3047 | n644;
assign n7070 = n7627 & n7830;
assign n8865 = n1876 & n2368;
assign n2448 = n13083 | n152;
assign n8674 = n5275 & n293;
assign n1001 = n6471 | n5727;
assign n7916 = n4525 & n5920;
assign n7993 = n12531 & n7559;
assign n2493 = n10936 | n6349;
assign n13983 = n3736 & n609;
assign n8000 = ~(n3400 | n4542);
assign n2117 = n9140 | n12586;
assign n5155 = n4498 | n11520;
assign n9211 = ~n409;
assign n2172 = n7116 | n9980;
assign n1197 = n14213 & n4306;
assign n428 = ~n11547;
assign n1441 = n5715 | n10679;
assign n12122 = n5800 | n9545;
assign n10968 = n7267 & n2206;
assign n10297 = n12169 | n7128;
assign n13103 = ~n8524;
assign n4911 = n4359 & n11956;
assign n3516 = n3219 | n12812;
assign n7723 = n7697 | n6974;
assign n966 = n13074 | n2774;
assign n11354 = n5139 | n6092;
assign n12728 = n12601 | n12822;
assign n393 = ~n7336;
assign n8988 = n1354 & n7656;
assign n1709 = n7043 & n691;
assign n8719 = n1772 & n11669;
assign n6782 = ~(n827 | n2235);
assign n13714 = n5786 | n8552;
assign n6589 = n14157 & n7571;
assign n8460 = n7862 | n3369;
assign n2961 = ~n6119;
assign n13065 = n501 & n5717;
assign n11736 = n11300 & n10455;
assign n5076 = ~(n8647 | n1395);
assign n9784 = n1125 & n11779;
assign n11395 = n12265 & n14209;
assign n11822 = n8746 & n1976;
assign n8425 = n4620 | n3465;
assign n14376 = ~n4907;
assign n5356 = n11093 & n10018;
assign n11367 = n8238 & n11653;
assign n5706 = n782 | n12216;
assign n13960 = n6090 | n2830;
assign n8265 = n12611 & n4866;
assign n5255 = ~(n3196 | n10924);
assign n2110 = n8581 | n3592;
assign n3718 = n8789 & n1916;
assign n3927 = ~(n7759 | n9022);
assign n13941 = ~n1010;
assign n11748 = ~n5871;
assign n2757 = ~(n12934 | n10460);
assign n9454 = n10523 | n1373;
assign n6273 = n1427 & n5693;
assign n509 = n3766 & n13004;
assign n5218 = n8528 | n2166;
assign n9059 = n12998 & n10989;
assign n12970 = ~n10423;
assign n11595 = n3268 & n11087;
assign n13481 = n8386 & n5867;
assign n11313 = ~n9865;
assign n8872 = n4657 & n14523;
assign n14066 = n8908 | n3987;
assign n8668 = n4973 & n2991;
assign n5032 = n6711 | n145;
assign n494 = ~n8997;
assign n13061 = ~n5702;
assign n109 = n6706 | n7891;
assign n11461 = n11411 & n3251;
assign n13169 = n5053 & n5202;
assign n7199 = n9265 & n14421;
assign n10964 = n5180 | n10599;
assign n5223 = n4840 | n62;
assign n859 = n11171 | n12565;
assign n970 = n5999 & n8703;
assign n11711 = ~(n4589 | n8257);
assign n5346 = n1844 | n4137;
assign n5338 = n5628 & n9962;
assign n6494 = n2901 | n13880;
assign n5825 = ~n2619;
assign n5990 = ~n12175;
assign n712 = n9856 | n10182;
assign n6594 = n9984 | n9470;
assign n2452 = n14327 & n6352;
assign n14038 = ~n5665;
assign n12246 = n5800 | n4661;
assign n8899 = ~n14075;
assign n5175 = n10331 | n11595;
assign n10284 = n48 | n9790;
assign n10042 = n14157 & n11276;
assign n6481 = n1137 | n4539;
assign n631 = n5348 & n4211;
assign n11701 = n6822 & n1690;
assign n14361 = n10300 | n14392;
assign n12565 = n678 & n1507;
assign n13547 = ~n4777;
assign n3152 = n9422 | n10743;
assign n5396 = ~(n4491 | n8861);
assign n11607 = ~n11861;
assign n13146 = n13780 & n6574;
assign n759 = n12620 & n11857;
assign n12457 = n6051 & n5837;
assign n1286 = n14282 | n9609;
assign n4423 = n2401 | n9468;
assign n4640 = n2949 | n10966;
assign n5515 = n9102 & n8864;
assign n11741 = n10357 & n10187;
assign n14077 = n1701 | n1895;
assign n10414 = n8304 | n991;
assign n5521 = ~(n7075 | n3874);
assign n6216 = n8768 & n6375;
assign n12725 = n103 & n8076;
assign n4157 = n11484 & n3891;
assign n2369 = ~n11771;
assign n1040 = ~(n4544 | n6137);
assign n12780 = ~(n12280 | n1375);
assign n7595 = n2645 | n9697;
assign n385 = n9885 & n11526;
assign n972 = n2158 & n5572;
assign n11506 = n9705 & n12463;
assign n4622 = n4102 & n12553;
assign n1958 = n4650 | n4615;
assign n1365 = n5512 | n4131;
assign n8415 = n12020 | n1151;
assign n421 = n394 | n1268;
assign n8971 = n13885 | n1449;
assign n8370 = ~(n2597 | n9968);
assign n9663 = n2224 & n3558;
assign n1112 = ~n2934;
assign n1201 = n6135 & n2457;
assign n13410 = n5603 | n6820;
assign n12415 = n251 | n13237;
assign n11484 = ~n7802;
assign n11731 = n6242 | n13624;
assign n4503 = ~(n10186 | n1626);
assign n12210 = n5139 | n732;
assign n4910 = n8897 | n335;
assign n4109 = ~(n9601 | n8467);
assign n8798 = ~n11343;
assign n10166 = ~n2958;
assign n8854 = n2724 & n3396;
assign n5952 = ~n4258;
assign n2384 = n13236 & n1303;
assign n12915 = n4627 & n12271;
assign n14494 = n1840 | n4159;
assign n12809 = n13745 & n1474;
assign n1242 = n13489 & n10510;
assign n6431 = n4468 | n9255;
assign n4295 = n6311 & n12104;
assign n2863 = n4657 & n13611;
assign n4901 = ~n9967;
assign n1902 = ~(n12569 | n10110);
assign n10479 = ~n2791;
assign n6165 = n7898 | n9646;
assign n12254 = ~n2069;
assign n7242 = n10855 & n8561;
assign n11780 = n9742 | n1282;
assign n640 = n12400 | n12072;
assign n14276 = n4422 & n8996;
assign n5477 = n7249 | n288;
assign n4045 = ~n14354;
assign n8017 = n8897 | n5311;
assign n4485 = n4239 | n6491;
assign n6401 = ~(n4091 | n5392);
assign n876 = n8476 | n4303;
assign n2885 = n77 | n642;
assign n11872 = n13096 & n5841;
assign n327 = ~n1458;
assign n10379 = n10820 & n11497;
assign n12828 = n4394 & n1264;
assign n12015 = ~n10372;
assign n2588 = n1231 & n250;
assign n3037 = ~n11151;
assign n9243 = n11980 | n3936;
assign n7558 = n1051 | n245;
assign n5141 = n12683 & n9249;
assign n3533 = n6606 & n2872;
assign n8084 = n10647 & n12753;
assign n7217 = n5450 | n7592;
assign n12706 = ~(n7052 | n9328);
assign n13575 = ~n12765;
assign n11828 = n1044 | n13311;
assign n1294 = n12042 & n14097;
assign n14523 = n2025 | n8728;
assign n1778 = n3777 | n5616;
assign n7683 = ~n9878;
assign n10264 = n14038 & n14503;
assign n8812 = ~n14464;
assign n3315 = n6343 & n13357;
assign n7650 = n11621 | n734;
assign n6312 = n4199 | n9466;
assign n9197 = ~n2778;
assign n13727 = n8386 & n4926;
assign n5511 = n405 & n9655;
assign n10101 = n1354 & n7510;
assign n5973 = n12226 & n4965;
assign n3930 = n5409 | n12813;
assign n1183 = n11033 & n12432;
assign n10807 = n13297 & n6176;
assign n2946 = n6436 | n11590;
assign n1996 = n4481 | n13176;
assign n13210 = n11097 | n12378;
assign n1729 = ~n4266;
assign n4156 = ~n13908;
assign n9029 = n7852 & n11413;
assign n3811 = n1006 | n11196;
assign n4519 = n5861 | n3105;
assign n9216 = ~n4716;
assign n3341 = n10383 | n2626;
assign n8768 = ~n12697;
assign n5617 = n12057 & n4593;
assign n553 = ~n4325;
assign n7593 = n5253 | n952;
assign n9688 = n12651 | n5794;
assign n12721 = ~n1911;
assign n165 = n10562 & n13739;
assign n14416 = ~(n13835 | n4547);
assign n6301 = n1047 & n4349;
assign n10785 = ~(n8825 | n5784);
assign n10956 = n8045 | n2978;
assign n13258 = n7912 | n12446;
assign n4887 = ~n13363;
assign n7856 = n69 | n5981;
assign n7639 = n1820 | n8900;
assign n12846 = ~n3309;
assign n6877 = n6822 & n3649;
assign n4410 = n1339 & n4234;
assign n783 = ~n8168;
assign n4101 = ~(n10824 | n4385);
assign n10203 = ~(n421 | n1062);
assign n11737 = ~n82;
assign n10709 = ~(n911 | n1341);
assign n8629 = ~n521;
assign n1303 = n12075 | n10734;
assign n5595 = n13466 & n7484;
assign n5886 = n13035 & n857;
assign n1876 = ~n8555;
assign n7548 = ~(n6122 | n1604);
assign n6878 = n2878 | n9858;
assign n5395 = n9429 | n9565;
assign n1172 = ~n6274;
assign n7168 = n13850 & n11222;
assign n11604 = n11123 | n6509;
assign n7290 = n10539 | n14258;
assign n4353 = n5825 & n6725;
assign n10096 = n10556 & n11615;
assign n1823 = n627 & n5639;
assign n2945 = n511 | n9817;
assign n11376 = ~(n742 | n4278);
assign n6045 = n4508 | n11978;
assign n11544 = n12998 & n4702;
assign n12639 = n6857 | n1935;
assign n7634 = ~(n1462 | n9021);
assign n7995 = n11495 & n38;
assign n11492 = ~n6196;
assign n14154 = n7376 & n1868;
assign n16 = n3710 & n7357;
assign n7081 = ~n6139;
assign n7884 = n9113 & n13044;
assign n13608 = n3277 & n10931;
assign n4592 = n7912 | n11009;
assign n5570 = ~n4891;
assign n11853 = n4619 & n12190;
assign n1141 = n1602 | n5187;
assign n12295 = ~n12106;
assign n733 = n4180 | n9288;
assign n7202 = n10815 & n6986;
assign n8259 = n10767 & n2252;
assign n12395 = n11315 | n6664;
assign n7516 = n9617 & n7867;
assign n13698 = ~n12489;
assign n6584 = ~(n6039 | n13740);
assign n2593 = n4239 | n153;
assign n9144 = n10731 | n8320;
assign n7587 = n3942 & n12352;
assign n12058 = n14093 & n7722;
assign n7420 = n6109 | n314;
assign n2920 = n14319 | n14002;
assign n4829 = ~n2996;
assign n201 = n5226 & n6600;
assign n11047 = ~n6123;
assign n7869 = n8983 | n12276;
assign n2146 = n10083 | n6182;
assign n2133 = ~(n329 | n11154);
assign n10207 = n1428 & n13873;
assign n216 = n8592 | n12172;
assign n12097 = n1268 | n4895;
assign n8732 = n13572 & n9486;
assign n4647 = n2367 & n4054;
assign n1149 = ~(n9291 | n7109);
assign n11068 = n12357 & n3008;
assign n1851 = ~(n13557 | n5805);
assign n5563 = n4156 & n2714;
assign n1455 = n11220 & n12083;
assign n5796 = n4300 & n13903;
assign n4545 = n10084 & n7535;
assign n2769 = ~(n619 | n12591);
assign n6050 = n3952 & n1160;
assign n12743 = ~(n5288 | n13208);
assign n10555 = n8372 & n3024;
assign n8482 = n4901 & n9479;
assign n12096 = ~n448;
assign n6778 = n10624 | n12422;
assign n11960 = n14093 & n4173;
assign n9107 = ~n8682;
assign n8970 = n1855 & n3531;
assign n5965 = n11710 | n5030;
assign n8777 = n11470 & n9398;
assign n7313 = n3366 & n7682;
assign n11743 = n14249 | n13636;
assign n13434 = n13017 & n1003;
assign n4924 = ~n14320;
assign n51 = n11420 | n12771;
assign n7949 = n4828 | n11610;
assign n10865 = n6754 & n3900;
assign n7715 = n10338 & n13761;
assign n5803 = n10678 & n1085;
assign n10753 = n12857 & n6454;
assign n9477 = n4239 | n3066;
assign n9101 = n8111 & n2495;
assign n3500 = n7810 & n11959;
assign n7840 = n7481 | n7140;
assign n13792 = n4239 | n11733;
assign n6198 = n3673 & n1194;
assign n9816 = n80 & n9763;
assign n4430 = ~(n8277 | n6117);
assign n6963 = ~(n9461 | n7087);
assign n5711 = n4574 & n2147;
assign n3035 = n9898 & n1118;
assign n9827 = n8747 | n12587;
assign n706 = ~n7507;
assign n11154 = ~(n5852 | n11587);
assign n11260 = ~(n9703 | n10006);
assign n2598 = n4929 & n11204;
assign n3772 = n965 & n961;
assign n5815 = ~n8695;
assign n3036 = n2877 | n750;
assign n10398 = n11510 | n3720;
assign n10601 = n12335 & n11728;
assign n7627 = ~n7023;
assign n1973 = n13885 | n5291;
assign n7834 = ~(n6466 | n6546);
assign n12252 = n5011 & n13506;
assign n11718 = n3161 | n6943;
assign n4552 = n11503 & n11545;
assign n4399 = n13074 | n9029;
assign n5760 = n4655 & n3683;
assign n1232 = n10294 | n10942;
assign n5514 = n8969 | n6656;
assign n7127 = ~(n506 | n6400);
assign n13868 = n2709 & n2102;
assign n7859 = n3320 | n12640;
assign n6924 = n13107 & n10130;
assign n5767 = n5012 & n13204;
assign n912 = n14404 | n2762;
assign n8325 = n7212 | n3613;
assign n7740 = ~(n8920 | n13816);
assign n1057 = n8747 | n6393;
assign n4672 = n12976 & n949;
assign n6191 = ~(n9176 | n11609);
assign n8088 = n14357 | n7748;
assign n4384 = n6354 & n6098;
assign n5935 = n12695 | n13301;
assign n77 = ~n4550;
assign n9678 = n251 | n9248;
assign n5533 = n11360 | n13402;
assign n2682 = ~n2744;
assign n9837 = n1225 | n6480;
assign n11868 = n10224 | n7782;
assign n7727 = n12934 | n10663;
assign n2471 = n6891 | n6441;
assign n3383 = n5764 & n11135;
assign n4518 = n9186 | n12336;
assign n3611 = n6525 & n9786;
assign n12363 = n5315 | n8305;
assign n6300 = ~(n12278 | n8365);
assign n7212 = ~n11308;
assign n13856 = n3011 | n11477;
assign n4600 = n6271 | n11506;
assign n1301 = n5940 & n7428;
assign n13376 = ~n11100;
assign n10077 = n11420 | n6960;
assign n6506 = n8748 | n13086;
assign n6209 = ~n13426;
assign n4708 = ~n9305;
assign n10969 = ~n7902;
assign n7588 = ~n9778;
assign n11948 = n11472 | n10448;
assign n1856 = n5064 | n8280;
assign n2323 = ~(n12823 | n13434);
assign n7939 = n7745 & n5395;
assign n12440 = ~(n13317 | n6521);
assign n12847 = n1117 & n10496;
assign n14078 = n2783 & n11468;
assign n11101 = ~(n12292 | n7788);
assign n12116 = ~(n4313 | n13442);
assign n5071 = ~n13360;
assign n5620 = n8490 | n5287;
assign n13446 = ~n9846;
assign n4333 = ~n9604;
assign n3568 = ~(n48 | n3940);
assign n11758 = n14091 & n7014;
assign n3750 = n13227 & n7840;
assign n3826 = ~n9169;
assign n649 = n8490 | n10920;
assign n7173 = n7249 | n14018;
assign n1968 = n6854 & n6982;
assign n6096 = n1210 | n9893;
assign n3852 = n3667 | n11577;
assign n2157 = n11816 & n7488;
assign n11908 = n4856 & n189;
assign n103 = ~n5951;
assign n10440 = n11679 & n4476;
assign n12939 = n5458 & n3058;
assign n14214 = n5092 & n6285;
assign n3222 = ~n5225;
assign n9712 = n9323 & n2178;
assign n7385 = n13755 & n3717;
assign n5644 = n533 & n11162;
assign n11533 = ~(n12046 | n5364);
assign n6673 = n2474 & n14326;
assign n8406 = n11176 | n923;
assign n11654 = n11824 | n3775;
assign n5660 = n4544 | n5142;
assign n14082 = n3886 | n9103;
assign n12697 = ~n12975;
assign n4180 = ~n7819;
assign n1572 = n3877 | n13419;
assign n7986 = n225 & n233;
assign n13035 = ~n9026;
assign n8013 = n4162 | n10498;
assign n4082 = n13109 | n9110;
assign n9015 = ~n9592;
assign n12388 = ~(n8458 | n12826);
assign n14503 = n7812 | n5476;
assign n7010 = n8372 & n10281;
assign n14169 = n1254 & n4124;
assign n1213 = n7693 & n2174;
assign n5885 = n7678 | n2349;
assign n8039 = n4162 | n10812;
assign n9471 = n9035 | n10525;
assign n9 = n9226 | n9062;
assign n5476 = n9745 & n7534;
assign n10989 = n2888 | n4412;
assign n8556 = n12461 & n2256;
assign n695 = ~n565;
assign n10909 = ~n7200;
assign n9374 = n7156 | n13565;
assign n1667 = n13074 | n9481;
assign n4587 = n3365 & n5382;
assign n10918 = n11336 & n4888;
assign n10654 = n6486 & n2986;
assign n2602 = n5732 | n8763;
assign n11803 = ~n10177;
assign n2380 = ~(n2098 | n7452);
assign n9005 = n2315 | n13339;
assign n8549 = n3047 | n6399;
assign n8637 = n12568 | n5082;
assign n11668 = ~n3324;
assign n6040 = n12802 & n6218;
assign n3089 = ~(n3871 | n5255);
assign n2979 = n7810 & n1996;
assign n12530 = ~(n13190 | n11165);
assign n6122 = ~n4634;
assign n6459 = n1006 | n11619;
assign n3369 = n9885 & n4055;
assign n2497 = ~n739;
assign n11752 = n9807 | n2700;
assign n12093 = n12020 | n11423;
assign n12312 = ~(n9924 | n2834);
assign n999 = n12858 & n7998;
assign n5435 = ~n744;
assign n3900 = n9864 | n8056;
assign n7571 = n2401 | n1110;
assign n14304 = n9285 | n7262;
assign n7405 = n7122 | n5283;
assign n12677 = ~(n228 | n9922);
assign n573 = ~n4847;
assign n9441 = n5236 | n12855;
assign n12353 = ~n6123;
assign n7021 = n1924 & n3653;
assign n14020 = n2180 & n11108;
assign n9615 = ~(n9078 | n11147);
assign n6188 = n12149 | n12160;
assign n11710 = ~n3021;
assign n12303 = ~n11875;
assign n14348 = n10089 | n8888;
assign n10295 = n12428 | n12208;
assign n4215 = n7909 & n4352;
assign n8388 = ~(n329 | n3325);
assign n6407 = ~(n14377 | n14208);
assign n8027 = ~n2919;
assign n14460 = n13342 & n2146;
assign n10713 = ~n12106;
assign n6166 = n6135 & n8261;
assign n202 = n7043 & n12613;
assign n6171 = n11406 & n12158;
assign n7798 = ~n10051;
assign n2829 = n5454 | n3245;
assign n2741 = n7745 & n6376;
assign n4804 = n1708 & n6862;
assign n3275 = n3777 | n5614;
assign n11882 = ~n1348;
assign n7035 = ~(n1685 | n4889);
assign n13263 = n9226 | n11025;
assign n3021 = n5029 & n7050;
assign n12671 = n9174 | n9484;
assign n11341 = n10294 | n567;
assign n4316 = n4486 & n8191;
assign n12358 = n12132 & n12933;
assign n2510 = ~n630;
assign n12153 = n11406 & n6773;
assign n13520 = ~n10828;
assign n465 = n13854 | n4517;
assign n10886 = n5641 | n11856;
assign n7852 = ~n5460;
assign n13058 = n13941 | n4;
assign n2537 = n4573 | n13511;
assign n865 = ~n12483;
assign n3176 = n3219 | n8454;
assign n4784 = n13379 & n9628;
assign n3905 = ~n10099;
assign n7950 = n227 | n10972;
assign n12148 = n1685 | n3456;
assign n466 = n12918 & n830;
assign n10499 = n12324 | n7573;
assign n3183 = n6654 | n13988;
assign n1787 = n7076 | n7006;
assign n5618 = ~n8809;
assign n9514 = n8401 & n5297;
assign n13074 = ~n4465;
assign n13578 = n12625 | n1718;
assign n14301 = n222 & n1965;
assign n9081 = n627 & n11827;
assign n9762 = n4973 & n5220;
assign n3178 = n10560 | n10806;
assign n3075 = n2310 & n8207;
assign n10128 = ~(n458 | n3633);
assign n5247 = ~(n4213 | n4430);
assign n12853 = ~(n7588 | n2948);
assign n6653 = n4657 & n342;
assign n4019 = n13226 | n5818;
assign n447 = n11679 & n14156;
assign n41 = n2246 | n1567;
assign n2236 = ~n1214;
assign n6430 = ~(n3497 | n7850);
assign n10935 = n3986 & n12774;
assign n2402 = n4128 | n13719;
assign n11206 = ~(n7188 | n1007);
assign n12553 = n13220 | n8977;
assign n6331 = n3559 | n1584;
assign n10337 = n55 & n11337;
assign n10253 = n7122 | n1709;
assign n14378 = n2820 & n11248;
assign n939 = n638 & n7703;
assign n11682 = n10855 & n2955;
assign n6745 = n10457 & n5768;
assign n9413 = n185 | n8474;
assign n3968 = n8045 | n13775;
assign n7018 = n5779 & n2549;
assign n10019 = ~n12776;
assign n5608 = n4525 & n2307;
assign n10922 = ~n4824;
assign n5919 = ~n8925;
assign n10454 = n11379 | n3648;
assign n7974 = n1362 | n2914;
assign n1491 = n11909 | n7506;
assign n4411 = n5132 | n2467;
assign n9057 = n647 | n7657;
assign n2495 = n5507 | n12963;
assign n57 = ~(n12630 | n9995);
assign n9501 = n9705 & n2506;
assign n8291 = ~n5197;
assign n5972 = n10154 | n9805;
assign n9303 = ~(n163 | n5521);
assign n6876 = n6428 | n9687;
assign n1236 = n1028 | n8850;
assign n6521 = n706 & n4743;
assign n12016 = n5483 | n5602;
assign n10996 = n13535 & n5212;
assign n10769 = n10969 & n8994;
assign n5739 = n10705 & n7930;
assign n9492 = n8172 | n11677;
assign n7228 = n7003 | n5167;
assign n7901 = n4407 | n6969;
assign n14255 = n12460 & n4799;
assign n5 = n12611 & n10335;
assign n9710 = n10209 & n12016;
assign n11588 = n4407 | n13822;
assign n9446 = n9726 & n1490;
assign n2139 = n11438 | n5408;
assign n14511 = n4498 | n12943;
assign n4318 = n7684 | n4088;
assign n6913 = n12226 & n525;
assign n7019 = n6711 | n11226;
assign n13455 = n11163 & n3881;
assign n12903 = n13338 & n2661;
assign n2171 = ~n3345;
assign n7149 = n251 | n10817;
assign n7124 = ~(n5952 | n1084);
assign n3746 = n80 & n12599;
assign n6363 = n6519 | n4933;
assign n1072 = n14227 & n5120;
assign n7408 = n2236 | n5125;
assign n3647 = n4806 & n12799;
assign n3237 = n5918 & n10722;
assign n6353 = n8821 | n11457;
assign n13811 = ~n11435;
assign n6322 = n9323 & n10120;
assign n1125 = ~n168;
assign n11992 = n8432 & n4915;
assign n7697 = ~n4847;
assign n954 = ~n11152;
assign n13843 = n10731 | n12704;
assign n11036 = ~n918;
assign n4119 = n1914 | n7363;
assign n9535 = n11722 | n759;
assign n12685 = n4244 & n9234;
assign n10506 = ~n10973;
assign n3980 = n7909 & n5492;
assign n4877 = ~n10889;
assign n7312 = n8768 & n1947;
assign n13114 = n10470 & n8269;
assign n14496 = n12295 | n9004;
assign n2874 = ~n10629;
assign n718 = ~n5525;
assign n9071 = n8692 & n9880;
assign n7143 = ~(n5665 | n1019);
assign n6637 = n7227 | n14301;
assign n11866 = n695 | n3534;
assign n10921 = ~(n2953 | n7202);
assign n5575 = ~n11308;
assign n8018 = n12265 & n443;
assign n8511 = ~n3946;
assign n9042 = n4394 & n7058;
assign n3769 = ~(n4913 | n7740);
assign n4566 = n9069 & n1001;
assign n9537 = n4267 & n6673;
assign n906 = ~n6053;
assign n4952 = n13525 & n7294;
assign n9739 = n3715 & n10208;
assign n1465 = n4657 & n2042;
assign n785 = n8786 & n11593;
assign n6138 = n12425 & n8694;
assign n13763 = n13484 & n11752;
assign n6532 = n4509 & n2271;
assign n6638 = ~n1548;
assign n2600 = n6316 & n13757;
assign n9595 = ~(n9266 | n3477);
assign n293 = n11572 | n4703;
assign n151 = ~n2354;
assign n3777 = ~n238;
assign n11198 = ~(n4741 | n8617);
assign n1848 = n7677 & n2329;
assign n4238 = n10332 & n2068;
assign n8867 = n9853 & n1498;
assign n11848 = n4445 & n14155;
assign n14115 = n12131 | n3941;
assign n4212 = ~(n14133 | n12380);
assign n13724 = n11510 | n784;
assign n11070 = n5266 | n5303;
assign n7817 = n4233 | n13445;
assign n13373 = n13484 & n11261;
assign n7619 = n3888 | n4265;
assign n5099 = n13220 | n8241;
assign n6226 = n14358 & n634;
assign n3534 = n9345 & n2402;
assign n6290 = ~(n6085 | n68);
assign n3105 = n8372 & n10068;
assign n9061 = n8825 | n2313;
assign n14336 = ~(n12934 | n13235);
assign n1802 = ~n4282;
assign n9329 = n263 | n4000;
assign n2263 = n11105 | n14339;
assign n7360 = n10626 | n1272;
assign n10262 = n9571 & n8826;
assign n10460 = ~(n7238 | n9177);
assign n12911 = ~(n4913 | n14170);
assign n2974 = n12149 | n6831;
assign n10893 = n5317 & n9296;
assign n2660 = ~(n6428 | n5527);
assign n8696 = n2465 & n9225;
assign n3304 = n12324 | n1142;
assign n11724 = ~n3357;
assign n1095 = n11484 & n6321;
assign n7033 = n3099 | n9591;
assign n13995 = n1854 & n14295;
assign n6056 = n13656 & n13068;
assign n12762 = n13656 & n11236;
assign n4090 = ~(n7245 | n2044);
assign n14208 = ~(n2218 | n11711);
assign n7356 = n13016 | n102;
assign n8452 = ~n2545;
assign n2666 = ~(n1383 | n9482);
assign n13418 = n7426 | n8933;
assign n11134 = n13707 | n3703;
assign n2628 = n7438 | n2242;
assign n13584 = ~(n2428 | n13999);
assign n1888 = n8517 | n2600;
assign n11664 = n13814 & n11332;
assign n7719 = n1047 & n1862;
assign n8802 = n13227 & n14197;
assign n6355 = n3715 & n5040;
assign n6593 = n11722 | n11499;
assign n10696 = n8250 & n4512;
assign n13466 = ~n9544;
assign n13259 = n12209 & n8233;
assign n10244 = ~(n12651 | n13596);
assign n6994 = n4255 | n962;
assign n6785 = n2461 & n6528;
assign n6832 = n2904 & n3824;
assign n6670 = ~n7662;
assign n12620 = ~n5268;
assign n5680 = n9218 | n2763;
assign n13255 = ~n8106;
assign n8499 = n5088 & n3660;
assign n6237 = n12772 & n7594;
assign n4570 = ~(n8023 | n4960);
assign n7642 = n5071 & n5972;
assign n12129 = n5695 | n7794;
assign n6297 = n1660 | n9644;
assign n8264 = n7673 & n2894;
assign n2884 = n11814 & n221;
assign n9293 = n2518 | n14490;
assign n4728 = n10331 | n4752;
assign n511 = ~n11331;
assign n7338 = n7208 & n12062;
assign n8428 = n8301 | n4582;
assign n7090 = n10820 & n6446;
assign n6847 = n11636 & n11625;
assign n8306 = n1093 & n3638;
assign n6856 = n4445 & n8624;
assign n849 = n865 & n3129;
assign n3851 = n14388 & n6292;
assign n12898 = n9230 | n1245;
assign n14513 = n9238 & n10580;
assign n9025 = n1172 | n680;
assign n9301 = n3120 | n1989;
assign n2219 = n14327 & n13486;
assign n4297 = n9188 & n8492;
assign n7280 = n9944 & n862;
assign n11806 = n12500 | n5922;
assign n10143 = n4199 | n10354;
assign n5038 = ~n9305;
assign n11361 = n1876 & n14167;
assign n11762 = ~(n5480 | n8000);
assign n6868 = n718 & n4695;
assign n9201 = n10822 & n8971;
assign n7952 = n10710 & n9770;
assign n6808 = n12620 & n6379;
assign n9004 = n12389 & n9808;
assign n4819 = n14088 | n2853;
assign n9848 = ~(n234 | n6325);
assign n4766 = ~(n11047 | n10723);
assign n13140 = ~(n4534 | n13168);
assign n8129 = n12324 | n5906;
assign n11729 = n10560 | n7031;
assign n5770 = n6596 | n4493;
assign n7069 = ~(n6085 | n14248);
assign n1288 = n11142 & n26;
assign n14469 = n14373 & n11007;
assign n4764 = n7852 & n6485;
assign n9646 = n55 & n1988;
assign n967 = n12455 & n364;
assign n6566 = n5406 | n902;
assign n13524 = n6109 | n9299;
assign n7797 = n7852 & n5924;
assign n12982 = ~(n13675 | n3560);
assign n11768 = n12460 & n3322;
assign n3134 = ~n1214;
assign n10546 = n2547 & n8107;
assign n12420 = n14449 | n8423;
assign n13045 = n12321 & n3410;
assign n13384 = n1362 | n8717;
assign n5199 = ~(n11558 | n8929);
assign n12467 = ~(n7889 | n6185);
assign n1336 = n4207 | n2045;
assign n1008 = n14110 | n5759;
assign n10311 = n3286 & n14059;
assign n13933 = n2843 | n5638;
assign n14118 = n2529 | n7988;
assign n8417 = ~(n12254 | n9879);
assign n7344 = n965 & n14144;
assign n12417 = n646 & n13117;
assign n12459 = n10015 & n7743;
assign n3079 = n7076 | n2580;
assign n14198 = ~n7322;
assign n9127 = n1614 | n3068;
assign n9571 = ~n11369;
assign n7164 = ~(n1713 | n9019);
assign n3932 = ~n7278;
assign n3747 = n619 | n6040;
assign n3853 = n4722 & n11014;
assign n11135 = n13477 | n877;
assign n10885 = ~(n8424 | n4575);
assign n9552 = ~(n7971 | n2584);
assign n10984 = n4407 | n897;
assign n8565 = n11738 & n9373;
assign n9126 = ~(n3309 | n809);
assign n10285 = ~n3191;
assign n2503 = ~n12904;
assign n886 = ~(n7192 | n3479);
assign n14027 = n5575 | n1095;
assign n3609 = n9127 | n9698;
assign n5428 = n12159 & n12713;
assign n605 = n3076 | n1518;
assign n9458 = ~(n2868 | n12677);
assign n12974 = n4394 & n11683;
assign n14473 = n6051 & n9887;
assign n12328 = n12576 | n8662;
assign n11217 = n116 | n13704;
assign n2659 = n8431 & n11849;
assign n8289 = n4486 & n4968;
assign n7079 = ~n871;
assign n7643 = ~(n3602 | n9704);
assign n6518 = n12112 | n6342;
assign n10327 = n8151 | n11255;
assign n14042 = ~n12450;
assign n8811 = n4840 | n4298;
assign n7400 = n7909 & n14516;
assign n5583 = n5359 | n2187;
assign n8075 = n4822 | n9923;
assign n8944 = n12802 & n5543;
assign n14337 = ~n12874;
assign n1028 = ~n630;
assign n1289 = n2682 & n11937;
assign n228 = ~n5901;
assign n3752 = n6854 & n5089;
assign n9604 = ~n12888;
assign n13542 = n9136 | n6422;
assign n9996 = n6625 & n9874;
assign n9785 = ~(n11180 | n7783);
assign n300 = ~n10787;
assign n7980 = ~n1377;
assign n12688 = n4407 | n13855;
assign n7620 = n12389 & n9991;
assign n5938 = ~(n3640 | n5966);
assign n6797 = ~n9740;
assign n11232 = ~n2257;
assign n10049 = n11121 | n3853;
assign n7014 = n13698 | n7106;
assign n2799 = ~n10046;
assign n13670 = ~(n5840 | n618);
assign n5926 = ~n11369;
assign n10899 = n1962 & n8211;
assign n5555 = n4359 & n5830;
assign n14365 = n8817 & n12785;
assign n7118 = n766 | n892;
assign n12424 = n2229 | n6031;
assign n2326 = n1044 | n7835;
assign n7185 = n776 & n11110;
assign n5920 = n9856 | n3780;
assign n3103 = n2461 & n7922;
assign n3041 = n10374 & n7483;
assign n3 = ~n14216;
assign n10892 = n8849 & n10184;
assign n5642 = n4468 | n4034;
assign n2145 = n13407 & n5302;
assign n9433 = n11620 | n10507;
assign n13905 = n9898 & n1957;
assign n10073 = n5234 | n7978;
assign n4358 = ~n1955;
assign n4915 = n11551 | n13607;
assign n3033 = n7391 & n1;
assign n3999 = n5088 & n13119;
assign n10032 = ~n12970;
assign n10714 = ~n6905;
assign n3009 = n11749 | n2073;
assign n13711 = n9529 | n2971;
assign n6039 = ~n12394;
assign n7206 = n4554 & n12840;
assign n9898 = ~n871;
assign n11113 = ~n8887;
assign n12375 = n5695 | n9357;
assign n6304 = n11621 | n12747;
assign n12801 = n6157 & n11168;
assign n9495 = n8768 & n6409;
assign n10178 = n9620 | n773;
assign n2498 = n9321 & n13960;
assign n10233 = ~n7704;
assign n5405 = n776 & n5865;
assign n7536 = ~(n5558 | n1959);
assign n5895 = n2846 & n419;
assign n13536 = n9375 | n1036;
assign n3164 = ~n2472;
assign n1687 = n4627 & n6620;
assign n9695 = n9804 | n4962;
assign n11288 = n48 | n7127;
assign n4813 = n9198 & n12242;
assign n1537 = n5253 | n4114;
assign n3552 = n8151 | n8433;
assign n9276 = ~(n703 | n9647);
assign n1264 = n11405 | n6432;
assign n13810 = ~(n4544 | n3351);
assign n12693 = ~n8500;
assign n10070 = n646 & n2493;
assign n10313 = n11153 & n11253;
assign n11979 = n5548 | n5541;
assign n2458 = n8605 & n10111;
assign n13287 = n11710 | n3279;
assign n3227 = n3204 & n5881;
assign n12127 = ~n10236;
assign n55 = ~n6787;
assign n10572 = n6271 | n8734;
assign n12371 = n283 | n3423;
assign n5792 = n10763 & n8911;
assign n2337 = n6957 & n10520;
assign n14086 = n3607 & n10104;
assign n12993 = n11702 & n12842;
assign n14324 = ~(n4207 | n14318);
assign n13152 = n8020 & n4075;
assign n10896 = n12018 & n10845;
assign n2162 = n553 | n4983;
assign n9299 = n8232 & n2400;
assign n4480 = n1613 | n8538;
assign n1102 = n11724 | n2333;
assign n14520 = ~(n584 | n13030);
assign n11749 = n12581 | n1022;
assign n12745 = n3672 & n6707;
assign n153 = n5062 & n6500;
assign n2619 = ~n3812;
assign n2832 = n12389 & n10997;
assign n13940 = n8986 | n1273;
assign n743 = n12013 & n4827;
assign n993 = n10234 | n7553;
assign n7803 = ~n10629;
assign n7382 = n844 & n2892;
assign n7177 = n12480 | n3655;
assign n363 = n9944 & n76;
assign n4562 = ~n7064;
assign n14060 = ~n12278;
assign n6478 = n4655 & n14108;
assign n5791 = n1775 & n13789;
assign n7224 = n5229 & n10414;
assign n11747 = ~(n2468 | n14112);
assign n8365 = n10059 & n7395;
assign n1922 = n11804 | n8906;
assign n13677 = ~n5294;
assign n9582 = n10154 | n3215;
assign n4931 = n8964 | n14020;
assign n9077 = n568 | n2192;
assign n8327 = n3800 | n279;
assign n960 = n13080 | n11021;
assign n9918 = n12620 & n9264;
assign n10789 = n13718 | n14160;
assign n10649 = ~n4708;
assign n5978 = ~(n4207 | n7496);
assign n10328 = n4807 | n3994;
assign n4703 = n8789 & n8160;
assign n13108 = ~n6264;
assign n13430 = n3025 | n7205;
assign n7653 = n10560 | n12754;
assign n12503 = ~n9193;
assign n12317 = n13698 | n7239;
assign n220 = n13035 & n6022;
assign n7319 = n10562 & n10398;
assign n1836 = n9174 | n8244;
assign n3004 = n706 & n12443;
assign n373 = n9890 & n10558;
assign n11998 = ~n11071;
assign n1853 = n11285 | n3631;
assign n4164 = ~(n9913 | n12848);
assign n757 = n1137 | n9129;
assign n1961 = n1391 | n10434;
assign n2642 = n1117 & n410;
assign n3898 = n5275 & n12285;
assign n102 = n6135 & n6420;
assign n7122 = ~n9686;
assign n6091 = n7421 & n2213;
assign n5357 = n6242 | n4236;
assign n13170 = n11950 & n9729;
assign n4194 = n5762 | n1666;
assign n3345 = ~n4589;
assign n10611 = n7530 | n8221;
assign n7449 = n5493 | n6240;
assign n4209 = n4806 & n9771;
assign n9839 = n13142 | n6856;
assign n12727 = ~n14016;
assign n11241 = n12169 | n9402;
assign n14458 = n85 | n5773;
assign n11449 = ~(n7229 | n4738);
assign n46 = n10080 & n7474;
assign n9220 = n3062 | n1502;
assign n12347 = ~(n8458 | n3651);
assign n3202 = n12351 | n7987;
assign n7982 = n2322 & n12363;
assign n1549 = n3276 & n4514;
assign n3630 = n11459 | n14;
assign n10804 = n14388 & n2207;
assign n8134 = n9245 & n416;
assign n8846 = n3062 | n10564;
assign n2866 = ~n6965;
assign n889 = ~n168;
assign n3582 = ~(n1243 | n14229);
assign n9086 = n9726 & n2139;
assign n14455 = ~n9172;
assign n9917 = n9015 & n11286;
assign n12407 = n5011 & n13949;
assign n8127 = ~(n13477 | n9521);
assign n13251 = n11157 & n14102;
assign n9569 = n13745 & n5552;
assign n593 = n850 | n6091;
assign n7023 = ~n8357;
assign n6186 = n536 & n13180;
assign n9550 = n3263 | n11345;
assign n5826 = n1481 & n10821;
assign n11694 = n6311 & n13092;
assign n10420 = n1711 | n11675;
assign n12237 = n1602 | n4873;
assign n11926 = ~(n151 | n10030);
assign n9664 = n14313 & n7194;
assign n11278 = n4627 & n10788;
assign n5421 = n5312 & n971;
assign n8422 = n2089 | n10171;
assign n12702 = n11406 & n9044;
assign n7466 = n74 | n13109;
assign n6223 = n5362 | n10039;
assign n10549 = n4045 | n2509;
assign n3335 = n5007 | n3913;
assign n12357 = ~n6810;
assign n58 = n13572 & n12395;
assign n8771 = n13531 | n8642;
assign n4955 = n4065 | n8503;
assign n3403 = n3777 | n7752;
assign n9473 = n9238 & n7022;
assign n2625 = n6263 | n12043;
assign n2196 = n11816 & n11540;
assign n12022 = n2181 | n9058;
assign n2878 = ~n622;
assign n4961 = n5266 | n4308;
assign n323 = n3512 | n14479;
assign n9761 = n12994 | n5439;
assign n7958 = n2082 & n6160;
assign n6713 = n13676 & n12399;
assign n2198 = n333 & n12240;
assign n13930 = n3914 | n8114;
assign n4687 = n7041 & n5856;
assign n13674 = n2445 & n9711;
assign n5472 = ~n12394;
assign n10456 = ~(n11580 | n9700);
assign n6068 = n4722 & n4026;
assign n1189 = ~n9580;
assign n12597 = n9804 | n8875;
assign n724 = n6085 | n12758;
assign n8496 = ~n4105;
assign n4431 = n12034 | n2941;
assign n7731 = n11839 | n3864;
assign n8097 = n9898 & n1536;
assign n2351 = n14042 & n13058;
assign n6591 = n6744 & n3115;
assign n11526 = n5861 | n6082;
assign n2941 = n3743 & n14355;
assign n14220 = n4908 | n10792;
assign n2524 = n4871 & n9587;
assign n8520 = n646 & n9832;
assign n880 = n7053 & n1475;
assign n4036 = n4443 | n1347;
assign n3363 = n10808 | n2270;
assign n5372 = n2843 | n13303;
assign n14320 = ~n7052;
assign n2030 = ~(n10929 | n12964);
assign n9428 = n9490 | n13514;
assign n10076 = n5807 | n14078;
assign n5325 = ~(n5897 | n4337);
assign n501 = ~n5108;
assign n11705 = n5861 | n10555;
assign n12584 = n13147 & n9235;
assign n4461 = n3815 | n13146;
assign n13160 = n1266 & n13178;
assign n12056 = n8980 | n1476;
assign n1157 = n5092 & n1621;
assign n9321 = ~n8798;
assign n14253 = n9972 & n11997;
assign n9382 = n1741 | n5290;
assign n5955 = n14088 | n10210;
assign n13538 = ~(n3602 | n11044);
assign n1760 = ~n2040;
assign n1604 = ~(n8701 | n9037);
assign n13804 = n10367 & n14043;
assign n13401 = n974 | n9219;
assign n1980 = n7427 & n415;
assign n12207 = n11171 | n12493;
assign n9659 = n4692 & n9452;
assign n9577 = ~n3345;
assign n1069 = n8431 & n11873;
assign n4272 = ~(n3768 | n10340);
assign n12048 = n1117 & n8174;
assign n26 = n2149 | n3303;
assign n6078 = n11405 | n3605;
assign n7690 = n5548 | n2007;
assign n581 = n4525 & n181;
assign n3634 = n8517 | n5003;
assign n3694 = ~(n4313 | n10739);
assign n290 = n2533 & n12529;
assign n10392 = n9069 & n11271;
assign n5778 = n8066 & n6886;
assign n5752 = n7887 | n3677;
assign n4162 = ~n6123;
assign n14288 = n7888 | n12789;
assign n7829 = n6867 | n7381;
assign n8859 = n13379 & n7732;
assign n3459 = n11028 & n7323;
assign n12670 = ~(n1383 | n4375);
assign n7618 = ~n702;
assign n13872 = n9238 & n323;
assign n11470 = ~n4296;
assign n9494 = ~n674;
assign n11704 = ~n8735;
assign n4055 = n5861 | n9281;
assign n3236 = n11542 | n4193;
assign n14422 = n9188 & n4473;
assign n4880 = ~n6990;
assign n7900 = ~n9236;
assign n13582 = n12542 & n8940;
assign n13947 = ~(n13707 | n6813);
assign n9470 = n2758 & n10982;
assign n1743 = n10084 & n8278;
assign n5355 = n10084 & n9861;
assign n62 = n5348 & n8834;
assign n13253 = n7443 & n12004;
assign n11063 = n7443 & n1077;
assign n2976 = n5139 | n1673;
assign n4658 = n808 & n11061;
assign n1794 = n10072 & n4431;
assign n13302 = n4509 & n11705;
assign n8608 = n782 | n325;
assign n4604 = n8302 & n12440;
assign n9023 = n8066 & n9670;
assign n10692 = n7427 & n13680;
assign n269 = n7249 | n10726;
assign n10363 = ~n3742;
assign n10627 = ~(n13675 | n7072);
assign n10488 = n185 | n5503;
assign n5187 = n5011 & n1386;
assign n2298 = n4382 & n10830;
assign n624 = n6343 & n10443;
assign n9880 = n8210 | n1298;
assign n1732 = n4614 & n2077;
assign n11234 = n7912 | n12314;
assign n2982 = n11909 | n9399;
assign n8132 = n14351 & n10427;
assign n13661 = ~(n5780 | n10106);
assign n6421 = ~(n6428 | n7955);
assign n1396 = n10024 | n11205;
assign n11040 = ~n5195;
assign n6074 = n8635 | n13814;
assign n7017 = n6242 | n12649;
assign n1881 = ~n6603;
assign n12165 = ~(n2597 | n11915);
assign n11727 = ~(n3287 | n3214);
assign n9721 = ~n10400;
assign n11448 = n6373 | n8546;
assign n5695 = ~n10204;
assign n8711 = n4546 & n14066;
assign n6454 = n3134 | n13777;
assign n3136 = n13130 | n14456;
assign n9320 = n8304 | n4214;
assign n13715 = n10247 & n13468;
assign n1207 = n12821 | n11167;
assign n9014 = n14337 | n12563;
assign n4665 = n10383 | n14314;
assign n11023 = ~(n12197 | n13474);
assign n12878 = ~(n14166 | n2125);
assign n13766 = n9111 | n1350;
assign n8923 = ~n2432;
assign n1510 = n12400 | n1969;
assign n186 = ~(n4210 | n2695);
assign n13641 = ~n5108;
assign n4504 = n11285 | n6932;
assign n10108 = n13230 & n398;
assign n7786 = n12741 & n8226;
assign n12408 = n965 & n6923;
assign n6833 = ~(n4439 | n14333);
assign n5149 = n14178 & n1850;
assign n7189 = n3164 | n401;
assign n9769 = n13420 | n10466;
assign n9265 = ~n7621;
assign n822 = n6730 | n2728;
assign n6467 = n5062 & n1579;
assign n3859 = ~(n13759 | n9615);
assign n8587 = n1414 & n6494;
assign n11435 = ~n12757;
assign n10014 = ~(n9577 | n7437);
assign n13762 = n3527 | n2143;
assign n10993 = n4562 | n12293;
assign n7402 = n6260 | n11930;
assign n6332 = n6844 & n937;
assign n14452 = n1520 & n1179;
assign n5369 = n11739 | n2689;
assign n7279 = n7419 & n5134;
assign n5720 = ~(n13677 | n6760);
assign n8796 = ~(n2057 | n12876);
assign n10966 = n6507 & n2625;
assign n13352 = ~(n7011 | n3719);
assign n4538 = n222 & n6834;
assign n3221 = n10245 | n10996;
assign n4614 = ~n7808;
assign n198 = n361 | n738;
assign n12073 = n8768 & n3933;
assign n9856 = ~n10985;
assign n12719 = n4722 & n4667;
assign n7876 = ~(n648 | n8603);
assign n5523 = n12130 | n9223;
assign n4851 = ~n14133;
assign n12100 = ~n1966;
assign n1933 = n4807 | n13241;
assign n7562 = n7011 | n2121;
assign n7559 = n11935 | n7777;
assign n4231 = ~(n5569 | n9475);
assign n1130 = n3273 | n455;
assign n12248 = ~n7521;
assign n11030 = n12425 & n6568;
assign n4800 = n13854 | n25;
assign n14315 = n9780 | n2568;
assign n4062 = n4508 | n1316;
assign n8759 = n6830 & n9988;
assign n3155 = n2012 & n10079;
assign n13480 = n8512 & n9068;
assign n14307 = n6480 & n7631;
assign n1819 = n8908 | n12715;
assign n10764 = n7426 | n5262;
assign n4289 = ~n2497;
assign n10125 = n2983 & n7565;
assign n14083 = n12622 | n14502;
assign n3722 = n11542 | n7786;
assign n7413 = n10302 & n10369;
assign n14199 = n14327 & n9488;
assign n12330 = ~(n11489 | n2623);
assign n7071 = n14408 & n12708;
assign n9609 = n4422 & n8437;
assign n152 = n7079 & n1014;
assign n6553 = n8432 & n4274;
assign n8035 = n4692 & n6252;
assign n13898 = n2645 | n3397;
assign n8442 = n7697 | n6203;
assign n4419 = n12037 & n5321;
assign n3574 = n9269 | n9405;
assign n979 = n4828 | n2935;
assign n13757 = n9429 | n13138;
assign n1816 = n523 | n11012;
assign n6246 = ~(n1028 | n6488);
assign n7770 = n12531 & n2546;
assign n11514 = n11484 & n8270;
assign n12050 = n4967 | n11215;
assign n3562 = n12130 | n7540;
assign n11935 = ~n11788;
assign n7181 = n3512 | n2459;
assign n13380 = n6288 | n9326;
assign n883 = n10019 | n5109;
assign n14488 = ~(n228 | n12891);
assign n9796 = n10374 & n10757;
assign n12302 = n5493 | n460;
assign n1559 = ~n5467;
assign n14470 = n6242 | n6823;
assign n1251 = ~(n10973 | n10431);
assign n8703 = n9211 | n3897;
assign n4268 = n11313 & n1438;
assign n1402 = n9724 & n8063;
assign n4540 = n13359 & n3751;
assign n5370 = n2904 & n10086;
assign n1605 = n6711 | n4364;
assign n6037 = n2897 | n4456;
assign n9671 = n2562 | n1641;
assign n10664 = n2064 & n4778;
assign n13494 = n5471 & n7828;
assign n8090 = ~(n8301 | n5599);
assign n7048 = n6205 | n3306;
assign n1815 = n13477 | n8953;
assign n1936 = n1640 | n3972;
assign n14274 = n8277 | n12520;
assign n9111 = ~n2472;
assign n3053 = n8825 | n3571;
assign n11745 = ~(n9340 | n6087);
assign n9724 = ~n3967;
assign n878 = ~(n7756 | n3817);
assign n1832 = n11636 & n3476;
assign n13439 = n13520 & n2606;
assign n11543 = ~(n4624 | n7372);
assign n4557 = n4313 | n3632;
assign n489 = ~(n7980 | n9059);
assign n8197 = ~n7710;
assign n10059 = ~n11605;
assign n1983 = n13112 | n12309;
assign n35 = n4407 | n6146;
assign n4021 = n6607 | n3384;
assign n11202 = n7736 | n13702;
assign n1594 = n9151 | n1201;
assign n10033 = n10930 & n5331;
assign n3546 = ~n3046;
assign n969 = n14188 | n13708;
assign n13398 = n638 & n14317;
assign n14440 = n10922 & n3554;
assign n1148 = n10084 & n5424;
assign n7376 = n2804 | n5009;
assign n521 = ~n14011;
assign n4541 = n5184 & n8051;
assign n3876 = ~n10864;
assign n10908 = n718 & n1207;
assign n12140 = n11748 & n10040;
assign n13628 = ~(n6000 | n3517);
assign n2775 = n80 & n6272;
assign n13830 = n12994 | n4457;
assign n14207 = n8025 & n1661;
assign n8203 = n9931 | n7279;
assign n3662 = n1701 | n14050;
assign n12769 = n5471 & n7342;
assign n14085 = n12455 & n14266;
assign n10925 = n1775 & n11632;
assign n4891 = n5788 & n8682;
assign n5200 = n4195 | n10570;
assign n3051 = n769 | n12887;
assign n6427 = n8897 | n11106;
assign n8861 = ~(n14198 | n3848);
assign n12636 = ~n13636;
assign n5310 = n4684 | n5696;
assign n9140 = ~n4203;
assign n250 = n361 | n11124;
assign n9056 = n231 & n11906;
assign n8106 = ~n9924;
assign n2632 = n8569 & n8316;
assign n9566 = ~(n4771 | n11762);
assign n2374 = n1924 & n10850;
assign n11017 = ~n13206;
assign n2072 = n4602 | n9947;
assign n8839 = n13700 & n3109;
assign n4347 = ~n6657;
assign n13212 = n7391 & n2870;
assign n653 = n3710 & n5910;
assign n1885 = n11090 | n6301;
assign n8031 = n573 | n3584;
assign n8614 = n7812 | n7285;
assign n1136 = ~n13295;
assign n13126 = n9885 & n9278;
assign n12458 = n12994 | n7939;
assign n3749 = ~(n8877 | n1411);
assign n7534 = n1582 | n5607;
assign n3381 = n6428 | n516;
assign n9510 = n11300 & n11288;
assign n4034 = n7691 & n13051;
assign n14181 = n14450 & n3996;
assign n2738 = ~n7904;
assign n402 = n8304 | n1779;
assign n2968 = n13446 | n5685;
assign n9941 = ~n12142;
assign n7214 = n6744 & n13125;
assign n10443 = n2562 | n1466;
assign n7207 = ~(n1685 | n13300);
assign n14505 = n11674 & n9055;
assign n1911 = ~n10341;
assign n7172 = n5475 & n7579;
assign n13863 = ~n3313;
assign n2264 = n2531 | n9104;
assign n525 = n7914 | n3189;
assign n4368 = ~(n10858 | n3996);
assign n1665 = n7392 & n2356;
assign n12402 = n6690 | n7951;
assign n2215 = n3401 & n6740;
assign n13154 = ~n2778;
assign n7781 = ~n650;
assign n2232 = n14472 | n9524;
assign n10623 = n14107 | n3121;
assign n1893 = n4358 & n3847;
assign n10582 = n10815 & n7297;
assign n13920 = n523 | n2084;
assign n10772 = n1006 | n13851;
assign n5854 = n329 | n10305;
assign n13207 = n5591 & n8088;
assign n9706 = n12475 & n7137;
assign n5120 = n8748 | n10260;
assign n8694 = n8490 | n2429;
assign n9183 = n12549 | n7306;
assign n7765 = n4354 & n13393;
assign n5624 = n5092 & n4056;
assign n7441 = n1076 & n1045;
assign n13272 = n286 & n1746;
assign n2717 = n8620 & n11473;
assign n8836 = n14150 & n4560;
assign n2464 = n986 & n969;
assign n2921 = n10731 | n7400;
assign n10442 = n12047 | n10085;
assign n10298 = n7887 | n5584;
assign n1627 = ~(n10368 | n4705);
assign n10079 = ~n666;
assign n13247 = n12494 | n10375;
assign n8790 = n12625 | n3992;
assign n3577 = ~n5631;
assign n2391 = n11470 & n9120;
assign n1214 = n7822 & n2609;
assign n14260 = ~n7902;
assign n9690 = ~(n355 | n3619);
assign n13006 = n12721 & n11746;
assign n7815 = n7419 & n9960;
assign n14109 = ~n5268;
assign n2208 = n2315 | n6845;
assign n13277 = n9864 | n13703;
assign n5302 = n5997 | n11912;
assign n8612 = ~(n12069 | n8090);
assign n3489 = n5695 | n6866;
assign n12535 = n2201 & n12718;
assign n11286 = n13432 | n505;
assign n12663 = n555 | n5355;
assign n12437 = n3193 | n3795;
assign n12138 = n5266 | n4921;
assign n14498 = n69 | n4642;
assign n11921 = n12543 | n417;
assign n1890 = n7697 | n5081;
assign n9636 = n7443 & n14519;
assign n13662 = n781 | n13763;
assign n13030 = ~(n7886 | n5192);
assign n8361 = ~n6714;
assign n11531 = ~(n4988 | n1902);
assign n210 = n11262 & n6087;
assign n12263 = n9218 | n1848;
assign n538 = n6629 | n3740;
assign n6629 = ~n3284;
assign n1755 = n9803 | n9830;
assign n4471 = ~(n30 | n4704);
assign n841 = n5007 | n10513;
assign n7632 = n6695 | n4060;
assign n7728 = n3877 | n4449;
assign n3593 = n9035 | n11772;
assign n3118 = n11090 | n13899;
assign n12062 = n12139 | n10359;
assign n5598 = n2058 & n7632;
assign n6998 = n89 | n2359;
assign n9872 = n5823 & n2499;
assign n8236 = n406 & n13346;
assign n6800 = n6343 & n11876;
assign n3077 = n8047 & n5020;
assign n6461 = n5053 & n367;
assign n1408 = n7043 & n2765;
assign n8981 = n14319 | n10057;
assign n13654 = n11315 | n11976;
assign n6942 = n10854 & n7671;
assign n8021 = ~n11244;
assign n3730 = ~(n4877 | n6712);
assign n9431 = n3526 & n2896;
assign n6471 = ~n4609;
assign n13213 = ~n9987;
assign n7730 = n9726 & n4942;
assign n9714 = ~(n13087 | n10483);
assign n4679 = n9297 & n3257;
assign n4288 = n4844 & n11561;
assign n6061 = n13252 & n5017;
assign n1822 = ~(n1617 | n13810);
assign n6308 = n6023 & n2475;
assign n7709 = ~(n10036 | n1042);
assign n13580 = n13501 | n10175;
assign n2813 = ~(n827 | n6906);
assign n4517 = n2583 & n3960;
assign n441 = n7551 | n9566;
assign n6982 = n12428 | n5241;
assign n3643 = n8702 & n5097;
assign n435 = n9111 | n4273;
assign n6116 = n1136 & n2802;
assign n14395 = n7438 | n9662;
assign n8618 = n3047 | n13174;
assign n5316 = n10626 | n12750;
assign n7657 = n5434 & n12862;
assign n2165 = n12091 | n13473;
assign n6057 = n3952 & n9536;
assign n7755 = ~n12658;
assign n10261 = n6706 | n13907;
assign n12244 = n11875 | n4117;
assign n3926 = ~n11001;
assign n860 = n428 & n13598;
assign n384 = n12034 | n12731;
assign n5696 = n14120 & n11450;
assign n12874 = n1936 & n13270;
assign n2584 = ~(n31 | n6502);
assign n10856 = ~(n11558 | n1064);
assign n14090 = n2318 | n5374;
assign n11766 = ~(n14466 | n9295);
assign n5781 = n7887 | n5593;
assign n9357 = n12461 & n2032;
assign n8508 = n3813 & n1647;
assign n13729 = n2942 & n5390;
assign n13216 = n12075 | n10906;
assign n7890 = ~(n1458 | n6963);
assign n3768 = ~n11308;
assign n4864 = n8242 | n14343;
assign n11046 = ~(n1628 | n9359);
assign n1472 = ~(n8404 | n12021);
assign n6587 = n7418 | n4283;
assign n1916 = n12353 | n14391;
assign n6939 = n3942 & n3469;
assign n990 = n7970 & n4194;
assign n12310 = n4502 & n9738;
assign n7308 = ~n8397;
assign n4351 = n4261 & n9293;
assign n8371 = n6754 & n14211;
assign n1110 = n5458 & n1654;
assign n7345 = ~n11218;
assign n1017 = ~(n3905 | n3321);
assign n6906 = ~(n2790 | n12678);
assign n957 = ~n6555;
assign n6084 = n4045 | n720;
assign n1619 = n3268 & n11877;
assign n1529 = n13433 & n13052;
assign n13049 = ~(n6041 | n14047);
assign n3992 = n7327 & n790;
assign n5773 = n12472 & n3288;
assign n8579 = n13860 & n13973;
assign n3337 = n12400 | n9073;
assign n4536 = ~(n13707 | n9948);
assign n5083 = n504 | n10242;
assign n9909 = ~(n11980 | n10347);
assign n12689 = n2998 & n4150;
assign n12455 = ~n11870;
assign n11473 = n5414 | n12270;
assign n5865 = n9285 | n14346;
assign n12087 = ~n10917;
assign n7860 = n7370 & n3188;
assign n14387 = n5647 | n735;
assign n3818 = n1729 & n8549;
assign n11267 = ~(n2017 | n6889);
assign n3866 = n7076 | n8258;
assign n3537 = n1602 | n12407;
assign n5045 = n1074 & n13015;
assign n7095 = n10394 | n13034;
assign n8380 = n2281 & n3192;
assign n11791 = ~(n12453 | n9239);
assign n2281 = ~n2752;
assign n11753 = n8358 & n3618;
assign n2396 = ~(n1480 | n13519);
assign n11519 = n7754 | n7889;
assign n9851 = n4508 | n258;
assign n3030 = n10396 | n3417;
assign n6604 = n7063 & n3363;
assign n12314 = n2064 & n7737;
assign n6970 = n4239 | n3482;
assign n2449 = n4880 & n9503;
assign n13021 = ~n12345;
assign n11033 = ~n9414;
assign n8477 = n11176 | n13701;
assign n4377 = n11748 & n2815;
assign n1646 = n4546 & n8263;
assign n9902 = n11316 & n9389;
assign n5408 = n3635 & n9343;
assign n9310 = n9853 & n423;
assign n13100 = n3126 | n826;
assign n12223 = n6271 | n8674;
assign n13909 = n12250 & n1826;
assign n8430 = n6724 & n12361;
assign n7227 = ~n6264;
assign n2195 = ~(n11481 | n1492);
assign n12747 = n8923 & n5328;
assign n9453 = n1421 & n298;
assign n13978 = ~n3681;
assign n12590 = n2149 | n11557;
assign n2519 = n14313 & n6580;
assign n12928 = n7026 & n11843;
assign n2585 = n11090 | n8484;
assign n5946 = n8147 & n13380;
assign n10591 = n3910 & n1546;
assign n9787 = ~(n8877 | n1859);
assign n10647 = ~n1378;
assign n5571 = n718 & n13027;
assign n6069 = n5062 & n5099;
assign n11598 = n5603 | n1948;
assign n2924 = ~n5046;
assign n10173 = n13547 | n607;
assign n8233 = n9245 | n9110;
assign n11614 = ~n6743;
assign n133 = n4207 | n9135;
assign n8987 = n2055 | n3103;
assign n4945 = n9035 | n7393;
assign n6753 = ~n7808;
assign n1488 = n10855 & n3515;
assign n12430 = n1011 & n4564;
assign n7605 = ~n9677;
assign n1515 = n103 & n12537;
assign n2624 = ~n1908;
assign n2203 = n4978 | n6151;
assign n25 = n10566 & n11103;
assign n1904 = ~n12697;
assign n8183 = ~n8122;
assign n12550 = n11411 & n1096;
assign n14048 = n9345 & n12411;
assign n12788 = n2694 | n10334;
assign n12746 = n56 & n201;
assign n11687 = ~n6114;
assign n13057 = n6316 & n12495;
assign n365 = n9745 & n50;
assign n13985 = n11953 | n10119;
assign n379 = n550 & n13539;
assign n10674 = n11951 | n3919;
assign n8308 = n6316 & n7848;
assign n6812 = n850 | n10388;
assign n7183 = n225 & n1692;
assign n9913 = ~n5683;
assign n4235 = n1193 & n6431;
assign n2387 = ~n8272;
assign n6863 = n11336 & n993;
assign n12172 = n13823 & n10971;
assign n3006 = n3743 & n4817;
assign n4558 = n4788 & n14092;
assign n8725 = n10083 | n12561;
assign n6164 = n13780 & n1088;
assign n5413 = n5480 | n3947;
assign n10286 = n6690 | n13497;
assign n5820 = n9275 & n13792;
assign n9703 = ~n8672;
assign n12950 = n3888 | n14353;
assign n11330 = n7909 & n7858;
assign n9200 = n1576 | n4731;
assign n14206 = n9824 & n4717;
assign n11172 = n4655 & n4140;
assign n12666 = ~(n5118 | n1767);
assign n2673 = n5936 | n2534;
assign n2545 = n12397 & n6928;
assign n725 = ~(n9806 | n14526);
assign n14128 = n2057 | n9155;
assign n2008 = n13641 & n6202;
assign n14391 = n14327 & n9756;
assign n1447 = ~n9921;
assign n8195 = n8386 & n5909;
assign n8953 = ~(n13394 | n3730);
assign n12447 = ~(n4953 | n11068);
assign n5426 = n4840 | n13065;
assign n7470 = n8769 & n3098;
assign n8362 = n8821 | n12123;
assign n1490 = n11438 | n12834;
assign n8718 = n1805 | n5592;
assign n10270 = n11816 & n8038;
assign n9541 = ~n4720;
assign n8689 = n1354 & n745;
assign n1007 = n7187 & n2481;
assign n11037 = n10539 | n6470;
assign n11156 = n6167 & n8951;
assign n8213 = ~n10377;
assign n11876 = n2562 | n6171;
assign n13921 = n492 | n608;
assign n12144 = n954 | n10708;
assign n9732 = ~(n11628 | n6405);
assign n8353 = ~n3572;
assign n1868 = n6640 & n1203;
assign n9888 = ~(n5977 | n3014);
assign n4897 = ~n749;
assign n13902 = n6867 | n3500;
assign n11977 = ~(n3922 | n12116);
assign n2013 = n11176 | n1150;
assign n13200 = n1247 & n2441;
assign n789 = ~(n906 | n8594);
assign n1454 = n6013 & n5589;
assign n1548 = n13882 | n6680;
assign n13530 = ~(n2415 | n4438);
assign n4253 = n3219 | n10631;
assign n9586 = ~(n8580 | n11778);
assign n11174 = n8786 & n1322;
assign n12099 = ~(n10323 | n9612);
assign n4237 = n9238 & n1034;
assign n14217 = n4562 | n1723;
assign n5984 = n5936 | n2295;
assign n1613 = ~n4606;
assign n488 = ~(n584 | n2999);
assign n13427 = n2099 & n6458;
assign n612 = n8620 | n2674;
assign n2375 = n6046 | n11525;
assign n998 = n8821 | n6612;
assign n8982 = ~(n10254 | n3890);
assign n12393 = n6596 | n2022;
assign n10991 = n10245 | n10968;
assign n9032 = n10857 | n13788;
assign n1405 = n11213 & n13198;
assign n925 = n12295 | n3746;
assign n5311 = n13676 & n4950;
assign n12779 = ~n10080;
assign n4184 = n7852 & n1446;
assign n7913 = ~(n7973 | n2303);
assign n12373 = n13626 & n13578;
assign n2050 = n14107 | n4081;
assign n11098 = n1480 | n11069;
assign n8366 = n5857 & n4814;
assign n5936 = ~n3007;
assign n13855 = n3952 & n6783;
assign n7423 = n12820 | n13769;
assign n2393 = n3826 | n8259;
assign n756 = n14091 & n4883;
assign n13968 = ~n13224;
assign n8810 = n13745 & n6236;
assign n6496 = n3277 & n452;
assign n11477 = n2310 & n7341;
assign n13861 = n3886 | n9651;
assign n8670 = ~(n2969 | n9493);
assign n14415 = n9726 & n10505;
assign n10198 = n7171 | n5046;
assign n1342 = ~n10603;
assign n6095 = n12101 & n7984;
assign n12003 = n2099 & n814;
assign n6221 = ~(n6768 | n903);
assign n10680 = n8432 & n13187;
assign n10323 = ~n2320;
assign n5170 = ~(n2781 | n9520);
assign n7370 = ~n12872;
assign n12577 = n12159 & n7082;
assign n4553 = n3169 & n13724;
assign n12610 = n687 & n3856;
assign n4311 = n320 | n12927;
assign n5422 = n1140 & n938;
assign n4922 = n12019 | n10769;
assign n14436 = n5582 & n13323;
assign n3800 = ~n10069;
assign n5596 = n13511 | n13364;
assign n1243 = n10147 | n14464;
assign n3812 = n12209 & n8134;
assign n10780 = n13464 & n143;
assign n3590 = n7438 | n7269;
assign n12806 = n4803 & n2265;
assign n6449 = ~(n7115 | n9031);
assign n13750 = n12057 & n10195;
assign n13190 = ~n739;
assign n8016 = n9442 | n12434;
assign n10622 = ~n10975;
assign n10599 = n4098 & n2915;
assign n5737 = n9811 & n1643;
assign n11095 = n100 | n939;
assign n9043 = n4602 | n2337;
assign n613 = ~(n5468 | n12312);
assign n5234 = ~n3455;
assign n8079 = n7053 & n1992;
assign n14247 = n10622 & n1581;
assign n11246 = ~(n10837 | n6418);
assign n9068 = n8726 | n5383;
assign n13311 = n10084 & n1698;
assign n9488 = n11360 | n5579;
assign n4702 = n7888 | n14081;
assign n9684 = n6531 & n8833;
assign n8099 = n1100 & n10073;
assign n4816 = n11438 | n10503;
assign n40 = n12549 | n2622;
assign n10179 = ~n7027;
assign n8351 = n4162 | n5811;
assign n14213 = ~n13219;
assign n5269 = n3204 & n7728;
assign n9987 = n12636 & n7811;
assign n2218 = ~n9959;
assign n6830 = ~n1771;
assign n13459 = n10678 & n209;
assign n10849 = n14038 & n6996;
assign n11910 = ~(n5715 | n6667);
assign n9956 = ~n10147;
assign n12156 = n8527 | n12128;
assign n578 = ~(n2766 | n3566);
assign n13658 = n7282 & n1277;
assign n7258 = n3628 & n8970;
assign n10390 = ~(n7900 | n6279);
assign n338 = n6695 | n4937;
assign n5787 = n3512 | n3915;
assign n1302 = n12622 | n4841;
assign n8595 = n2772 & n1334;
assign n2459 = n7026 & n5111;
assign n12428 = ~n8148;
assign n7582 = ~(n10402 | n3235);
assign n9208 = n14227 & n507;
assign n13722 = ~n4646;
assign n4811 = n10516 & n4402;
assign n9010 = n11576 | n12980;
assign n909 = n11411 & n12555;
assign n4653 = ~(n13675 | n12120);
assign n7907 = n2177 & n5557;
assign n5006 = ~(n9984 | n6124);
assign n11119 = n13718 | n10578;
assign n10971 = n8986 | n4758;
assign n1312 = ~n11305;
assign n11208 = n11036 | n182;
assign n10724 = n129 & n7774;
assign n3132 = ~n12776;
assign n8848 = n7429 & n11785;
assign n507 = n8748 | n9632;
assign n11282 = n5489 & n9430;
assign n7126 = n4806 & n13861;
assign n7851 = n10457 & n12329;
assign n4919 = n12475 & n3083;
assign n413 = ~(n2417 | n10329);
assign n5874 = n5458 & n12491;
assign n8866 = ~n5077;
assign n14121 = n1028 | n14172;
assign n7927 = ~(n3354 | n13089);
assign n5469 = ~(n1844 | n1527);
assign n2589 = n4844 & n5025;
assign n9246 = n12015 & n11734;
assign n8186 = ~(n13081 | n13352);
assign n12155 = ~(n7551 | n9630);
assign n11647 = ~n2130;
assign n3617 = n5234 | n14437;
assign n3868 = n405 & n4992;
assign n6293 = n12020 | n9661;
assign n5580 = n1804 & n10741;
assign n3338 = ~(n5118 | n878);
assign n12908 = n2246 | n3945;
assign n5997 = ~n751;
assign n2372 = n1431 & n9000;
assign n314 = n4546 & n9688;
assign n11792 = n9119 | n2895;
assign n1579 = n9780 | n11243;
assign n6444 = ~(n4978 | n4760);
assign n317 = ~n622;
assign n14210 = ~n7941;
assign n14003 = n5240 & n8050;
assign n7016 = n5940 & n12319;
assign n13301 = n12265 & n8175;
assign n9670 = n4052 | n3180;
assign n13982 = n1391 | n4332;
assign n10607 = ~(n9984 | n9701);
assign n13499 = n2224 & n2920;
assign n10492 = ~(n3132 | n8473);
assign n7509 = n2465 & n7901;
assign n4179 = n1535 | n3000;
assign n14026 = n11093 & n3221;
assign n2079 = n9931 | n12859;
assign n99 = n13509 | n2201;
assign n818 = ~(n1693 | n2631);
assign n11102 = n1427 & n9505;
assign n4883 = n3273 | n6433;
assign n4380 = n432 & n88;
assign n8102 = n7053 & n1644;
assign n11410 = ~(n4248 | n6268);
assign n6394 = n13641 & n12793;
assign n3301 = n387 | n2594;
assign n4242 = n2181 | n9872;
assign n3347 = n3134 | n12231;
assign n10254 = ~n4966;
assign n7741 = n8986 | n12684;
assign n5977 = ~n382;
assign n12539 = ~(n3873 | n705);
assign n4673 = ~(n10593 | n7695);
assign n9399 = n3607 & n1569;
assign n9982 = n13107 & n3124;
assign n9798 = n10969 & n7726;
assign n4497 = n2412 | n9930;
assign n2274 = n49 | n8275;
assign n5097 = n49 | n2641;
assign n3216 = n11047 | n6935;
assign n187 = n7358 | n9648;
assign n1804 = ~n10372;
assign n13731 = n4602 | n7049;
assign n1685 = ~n622;
assign n1166 = n7684 | n2578;
assign n3058 = n7359 | n14467;
assign n832 = n1582 | n13564;
assign n9226 = ~n5242;
assign n7216 = ~n2454;
assign n12722 = n6629 | n8414;
assign n2798 = ~(n8825 | n1385);
assign n9551 = n11171 | n4597;
assign n2036 = ~(n14135 | n11757);
assign n1520 = ~n10036;
assign n12482 = n781 | n8430;
assign n5903 = n3877 | n5244;
assign n275 = n14430 | n10162;
assign n5776 = n8828 | n9822;
assign n2390 = ~(n7227 | n8199);
assign n14305 = n3559 | n3872;
assign n14467 = n10338 & n12214;
assign n5374 = n6531 & n6896;
assign n1228 = n11220 & n832;
assign n13033 = n4502 | n2201;
assign n6630 = ~(n4049 | n13183);
assign n381 = n1225 & n11751;
assign n11145 = n7527 | n11896;
assign n1730 = n7677 & n7528;
assign n8883 = n2510 | n10652;
assign n11011 = ~n7404;
assign n10500 = n1602 | n14034;
assign n6004 = n1261 | n7994;
assign n10018 = n568 | n2581;
assign n3060 = n1494 | n2826;
assign n9361 = n11459 | n5731;
assign n7287 = n4289 & n3343;
assign n9266 = ~n12506;
assign n6241 = n11551 | n2119;
assign n4280 = ~(n2098 | n6443);
assign n6941 = ~n12322;
assign n3985 = n4899 | n4249;
assign n3687 = n11722 | n13144;
assign n11440 = ~n12746;
assign n14273 = ~n3893;
assign n3744 = n12730 & n10764;
assign n8232 = ~n8048;
assign n4429 = n3193 | n3957;
assign n4685 = n1137 | n5004;
assign n13587 = n533 & n9095;
assign n11043 = n12335 & n6587;
assign n13075 = n1431 & n5079;
assign n2765 = n49 | n11185;
assign n8676 = n8111 & n704;
assign n9450 = ~n6248;
assign n3713 = n6724 & n3688;
assign n7889 = n10765 | n4154;
assign n6769 = n13489 & n4665;
assign n14176 = n9747 | n13994;
assign n12481 = n2897 | n2936;
assign n2244 = n6891 | n3026;
assign n1924 = ~n3344;
assign n11962 = n8932 & n10916;
assign n4717 = n13432 | n2939;
assign n2017 = ~n13668;
assign n6774 = n12475 & n6035;
assign n6412 = n14029 | n6666;
assign n6505 = n333 & n4006;
assign n7246 = n13093 & n578;
assign n3177 = ~(n2677 | n12667);
assign n5529 = n12018 & n4823;
assign n10932 = n12772 & n2043;
assign n738 = n10589 & n6021;
assign n11917 = n98 & n8325;
assign n6784 = n8066 & n9791;
assign n6339 = n4276 & n10884;
assign n13483 = n5450 | n13170;
assign n10538 = n11953 | n4127;
assign n6949 = ~(n7739 | n8139);
assign n213 = n4289 & n1800;
assign n12961 = n10229 & n2263;
assign n131 = n766 | n1543;
assign n11320 = n12112 | n12327;
assign n4937 = n13359 & n11263;
assign n13243 = n12185 & n11133;
assign n12344 = n7076 | n2721;
assign n5114 = n4498 | n14129;
assign n1411 = ~(n7660 | n6583);
assign n14338 = n8575 | n4426;
assign n6743 = ~n13725;
assign n12865 = ~(n6953 | n10464);
assign n1445 = n6135 & n2803;
assign n828 = ~(n1820 | n3262);
assign n5420 = n10913 | n570;
assign n11958 = n4856 & n12662;
assign n2131 = n7156 | n6708;
assign n5144 = ~n426;
assign n3892 = n1914 | n8137;
assign n13508 = ~(n4233 | n13145);
assign n12887 = n6354 & n569;
assign n13648 = ~(n9818 | n13325);
assign n6476 = ~(n14419 | n13538);
assign n30 = n4659 | n12573;
assign n9296 = n11121 | n8074;
assign n14035 = n10678 & n4023;
assign n10362 = n5764 & n5594;
assign n12069 = ~n8927;
assign n14122 = n1662 & n12307;
assign n5855 = ~n13511;
assign n11795 = n11336 & n633;
assign n3684 = n361 | n4677;
assign n3787 = n2367 & n6796;
assign n9736 = n8213 & n1037;
assign n10606 = n14109 & n6173;
assign n1137 = ~n1041;
assign n2237 = n13074 | n2616;
assign n10543 = n6730 | n4139;
assign n13423 = n5779 & n13797;
assign n3142 = n5137 & n1005;
assign n520 = n13220 | n8676;
assign n3471 = n6838 & n12913;
assign n8547 = ~(n2251 | n9376);
assign n13701 = n9315 & n11049;
assign n13997 = ~(n6797 | n7876);
assign n10419 = n13700 & n10417;
assign n9139 = n9824 & n6549;
assign n13858 = n1278 & n1958;
assign n6826 = n5038 & n13366;
assign n10812 = n14327 & n5248;
assign n4646 = ~n4135;
assign n13395 = n11406 & n10614;
assign n7553 = n14063 & n14438;
assign n1903 = n5695 | n8556;
assign n13955 = n8714 | n10685;
assign n9676 = n172 | n7317;
assign n9073 = n3565 & n7892;
assign n12098 = n6016 & n5817;
assign n8507 = ~n12885;
assign n11378 = n10825 | n14422;
assign n3584 = n3 & n980;
assign n13081 = ~n12580;
assign n6046 = ~n4149;
assign n10976 = n12994 | n9409;
assign n987 = n6023 & n1054;
assign n6097 = n2784 | n8102;
assign n1496 = n1189 | n5054;
assign n10429 = n4840 | n6394;
assign n11980 = ~n6978;
assign n7250 = ~n3284;
assign n13465 = n13246 & n7243;
assign n6722 = n9232 & n1664;
assign n4579 = n9052 & n641;
assign n6052 = ~n6874;
assign n11347 = n12391 & n6368;
assign n13809 = n12211 | n4222;
assign n1775 = ~n3402;
assign n13226 = ~n1267;
assign n6267 = n10024 | n397;
assign n12033 = n2724 & n6503;
assign n9039 = ~(n7887 | n13414);
assign n4978 = ~n8695;
assign n6960 = n12935 & n13191;
assign n3613 = n11484 & n1599;
assign n12729 = n10913 | n9949;
assign n6759 = n11838 & n3842;
assign n12509 = n11702 & n11897;
assign n13888 = n2901 | n7235;
assign n1086 = ~n4595;
assign n2407 = n10147 & n4671;
assign n12229 = ~n1843;
assign n1562 = n2510 | n4029;
assign n11180 = ~n8704;
assign n12581 = n2946 | n5418;
assign n7145 = ~n7291;
assign n5863 = n6971 | n852;
assign n8267 = n5144 | n8294;
assign n6170 = n7116 | n13963;
assign n8560 = n4435 | n5560;
assign n13305 = n2518 | n13503;
assign n3430 = n5732 | n6069;
assign n736 = n13840 & n177;
assign n3491 = ~n9818;
assign n4713 = ~n2731;
assign n10199 = n11838 & n2031;
assign n10847 = n9230 | n4775;
assign n12082 = n12543 | n6226;
assign n7316 = n7081 & n2259;
assign n11083 = n12844 | n12598;
assign n10063 = n9375 | n14460;
assign n12587 = n6899 & n689;
assign n3541 = ~(n11111 | n165);
assign n13413 = ~n9596;
assign n9149 = n10247 & n14030;
assign n2505 = ~n1763;
assign n1328 = n7684 | n6995;
assign n1692 = n8821 | n12277;
assign n3550 = n4128 | n12735;
assign n12193 = ~n10465;
assign n8590 = ~(n7075 | n2844);
assign n11576 = ~n1041;
assign n1200 = n14058 | n6752;
assign n49 = ~n9306;
assign n10287 = ~(n10688 | n723);
assign n7291 = ~n10803;
assign n7925 = n6981 & n10672;
assign n1417 = ~n3324;
assign n10693 = n3424 & n14100;
assign n6907 = ~n12580;
assign n5858 = n7527 | n466;
assign n10156 = n12038 & n4987;
assign n5286 = n12295 | n7620;
assign n5176 = n13069 & n13827;
assign n7059 = n10763 & n1999;
assign n4113 = n1112 | n7457;
assign n11987 = ~(n14296 | n7791);
assign n10834 = ~n751;
assign n396 = n9705 & n7046;
assign n936 = n222 & n9075;
assign n3538 = n1202 | n1145;
assign n11027 = n8401 & n3016;
assign n7171 = ~n4039;
assign n6105 = n13877 & n675;
assign n11438 = ~n10346;
assign n3950 = n12265 & n12049;
assign n229 = n8304 | n9762;
assign n10158 = n3120 | n3039;
assign n3952 = ~n10828;
assign n10874 = n13525 & n8541;
assign n5054 = n1231 & n8367;
assign n3929 = n14521 | n7832;
assign n3821 = n14109 & n1921;
assign n11511 = n7781 | n9252;
assign n8667 = n2531 | n13066;
assign n6940 = n11329 & n10671;
assign n4814 = n283 | n4753;
assign n10920 = n12461 & n4310;
assign n4462 = n12101 & n5363;
assign n7510 = n976 | n11201;
assign n4533 = n14009 | n2048;
assign n3150 = n7898 | n3111;
assign n9046 = ~n2298;
assign n12608 = n10032 & n291;
assign n8814 = n9142 | n6460;
assign n5647 = ~n4939;
assign n4509 = ~n1178;
assign n5102 = n11403 & n10853;
assign n2973 = ~n9414;
assign n5662 = n11704 | n120;
assign n6725 = n6607 | n13812;
assign n10547 = n12202 & n12413;
assign n7645 = n1678 & n556;
assign n7093 = n8855 & n10023;
assign n9778 = ~n742;
assign n9786 = n5454 | n8405;
assign n12603 = n7736 | n8195;
assign n8700 = n12047 | n6415;
assign n2408 = n8821 | n7460;
assign n3837 = n12953 & n7564;
assign n7097 = n5493 | n12623;
assign n12132 = ~n8302;
assign n1610 = ~n2692;
assign n1366 = n10154 | n831;
assign n12559 = n13118 | n385;
assign n3503 = n12105 & n5259;
assign n2290 = n11360 | n4380;
assign n13453 = n10781 | n14414;
assign n7047 = n14198 | n9307;
assign n855 = n12034 | n597;
assign n5501 = n10209 & n8488;
assign n13853 = n3367 & n2768;
assign n4496 = n6428 | n2283;
assign n12748 = n2547 & n4940;
assign n10915 = n7667 & n12790;
assign n7465 = n10871 | n1832;
assign n4654 = ~(n6000 | n9552);
assign n7821 = n11157 & n4480;
assign n7328 = n9113 & n8610;
assign n13950 = ~(n1944 | n9303);
assign n13124 = ~(n12046 | n8312);
assign n12624 = n12101 & n7151;
assign n3251 = n14282 | n13744;
assign n3646 = n10449 | n10490;
assign n1583 = n8066 & n8477;
assign n7043 = ~n10269;
assign n13322 = n8702 & n1889;
assign n4544 = ~n7875;
assign n7373 = n69 | n1164;
assign n961 = n5266 | n5061;
assign n9179 = n11028 & n1845;
assign n2700 = n1255 & n3183;
assign n14190 = n3724 & n11690;
assign n3699 = n4791 | n1583;
assign n12839 = n3125 | n3513;
assign n6032 = n13005 | n7698;
assign n11315 = ~n7339;
assign n556 = n7971 | n3576;
assign n4092 = ~n565;
assign n6376 = n1576 | n11398;
assign n5864 = ~(n13394 | n8943);
assign n5437 = n14388 & n3604;
assign n2753 = n1678 & n12473;
assign n1078 = n12077 | n6917;
assign n748 = ~n2497;
assign n11398 = n1100 & n9320;
assign n1847 = n2378 & n12559;
assign n10731 = ~n9846;
assign n1140 = ~n11969;
assign n6772 = n4486 & n7626;
assign n2363 = n1821 | n5351;
assign n3683 = n6730 | n13369;
assign n4408 = n10909 & n1249;
assign n13149 = n387 | n4001;
assign n9964 = n7122 | n10174;
assign n8823 = n13860 & n11720;
assign n3849 = n5764 & n11658;
assign n9513 = n12101 & n3811;
assign n6829 = ~n4379;
assign n6266 = n8552 | n9589;
assign n2620 = n14446 & n13699;
assign n5763 = n5348 & n4592;
assign n5064 = ~n6978;
assign n10881 = n817 | n6771;
assign n8495 = n11379 | n6333;
assign n3707 = n965 & n4204;
assign n5027 = n3370 & n1562;
assign n48 = ~n777;
assign n8774 = n8358 & n9263;
assign n11263 = n1198 | n3643;
assign n2213 = n9151 | n8130;
assign n10160 = n13555 & n3575;
assign n2534 = n10822 & n13457;
assign n14047 = ~(n1028 | n5712);
assign n14525 = ~n11401;
assign n4143 = n2564 & n3404;
assign n9641 = n8401 & n5781;
assign n433 = n1147 | n5743;
assign n14232 = n15 & n10674;
assign n9153 = n10399 & n5464;
assign n1889 = n10396 | n3518;
assign n1735 = n11313 & n4327;
assign n1216 = n5641 | n2374;
assign n8468 = n5317 & n9411;
assign n11885 = n3449 | n650;
assign n3841 = n6754 & n13277;
assign n4602 = ~n7441;
assign n10786 = n10461 | n3601;
assign n5816 = n1610 & n5971;
assign n9715 = n13338 & n11354;
assign n10870 = n12449 & n4748;
assign n1948 = n12389 & n5928;
assign n12170 = ~(n11498 | n8551);
assign n10828 = ~n210;
assign n7442 = n5483 | n11030;
assign n10231 = ~n13093;
assign n1442 = n11572 | n3718;
assign n6824 = n3809 | n1835;
assign n13743 = n13484 & n9731;
assign n927 = n3888 | n1326;
assign n7011 = ~n7289;
assign n6129 = n12764 | n1435;
assign n11517 = n12620 & n11019;
assign n11927 = n3271 | n74;
assign n9467 = n3986 & n11598;
assign n1762 = ~(n6052 | n602);
assign n10435 = n4978 | n343;
assign n9058 = n5823 & n4825;
assign n6746 = n9885 & n2959;
assign n2266 = n1876 & n5377;
assign n1967 = n7803 | n7242;
assign n1474 = n8480 | n7344;
assign n10068 = n5625 | n8206;
assign n6227 = n7943 & n7310;
assign n6271 = ~n409;
assign n14508 = ~(n8458 | n1344);
assign n3651 = ~(n1929 | n6875);
assign n8585 = n12105 & n1275;
assign n4686 = n1711 | n2038;
assign n4599 = n2322 & n8140;
assign n11632 = n3871 | n11042;
assign n1897 = n10330 & n14158;
assign n8977 = n10166 & n1166;
assign n350 = ~n8315;
assign n4324 = n7934 & n1793;
assign n6615 = n11704 | n4930;
assign n12966 = ~(n8277 | n9606);
assign n12958 = n3710 & n10412;
assign n1357 = n10378 | n10080;
assign n2949 = ~n5901;
assign n13266 = ~(n5944 | n11862);
assign n971 = n8332 | n7172;
assign n11069 = ~(n11546 | n11812);
assign n4366 = ~(n3394 | n4252);
assign n3796 = n2006 & n3270;
assign n3390 = n13413 | n6153;
assign n12629 = n10624 | n12985;
assign n4481 = ~n9846;
assign n14147 = n13118 | n6250;
assign n1169 = n12741 & n1020;
assign n7398 = n390 | n11327;
assign n6894 = n6486 & n12696;
assign n9416 = ~n10115;
assign n1139 = n6867 | n9659;
assign n437 = n12475 & n6615;
assign n6988 = n2904 & n4367;
assign n14507 = n11153 & n1809;
assign n8260 = n4581 & n10131;
assign n10669 = n2149 | n4187;
assign n12527 = ~n6254;
assign n2512 = ~(n8656 | n9147);
assign n6588 = n3586 & n11208;
assign n5797 = n11360 | n11322;
assign n4881 = n2998 & n9854;
assign n1331 = n11737 & n10517;
assign n7028 = n3204 & n1367;
assign n13621 = n8304 | n4454;
assign n10377 = ~n8003;
assign n9388 = ~n2520;
assign n11950 = ~n12503;
assign n10903 = n4199 | n10602;
assign n2482 = n3672 & n8032;
assign n4465 = n11188 & n772;
assign n2324 = n783 & n953;
assign n11680 = ~n4786;
assign n2782 = n15 & n12804;
assign n1587 = n9745 & n5510;
assign n11175 = n4967 | n11925;
assign n7156 = ~n7339;
assign n7327 = ~n12904;
assign n12280 = ~n3587;
assign n3478 = n2521 & n3843;
assign n5699 = n11581 | n3209;
assign n10448 = n8147 & n3073;
assign n4783 = n783 & n3490;
assign n1150 = n8183 & n9425;
assign n10360 = ~n12782;
assign n1683 = n2878 | n10691;
assign n6255 = n9238 & n13563;
assign n4539 = n13240 & n3979;
assign n7054 = n6697 & n7034;
assign n13716 = n6109 | n6359;
assign n5151 = n6909 & n6185;
assign n21 = n11839 | n9208;
assign n11447 = n8213 & n503;
assign n10221 = n13531 | n11893;
assign n11999 = ~(n10289 | n1251);
assign n5512 = ~n4659;
assign n2794 = n5416 & n6705;
assign n69 = ~n11055;
assign n5862 = n428 & n4182;
assign n6731 = ~n4708;
assign n10525 = n8431 & n2216;
assign n2839 = n13477 | n5034;
assign n8011 = n7079 & n9758;
assign n9777 = n13005 | n2806;
assign n7984 = n5833 | n4903;
assign n9894 = n10913 | n10695;
assign n1401 = ~n10470;
assign n3724 = ~n5618;
assign n11769 = n14401 | n6759;
assign n10000 = n14065 | n13944;
assign n3502 = n1857 & n5749;
assign n7733 = n14465 & n13524;
assign n558 = ~(n7146 | n7281);
assign n3083 = n1838 | n8070;
assign n9493 = ~(n4195 | n5022);
assign n6838 = ~n7902;
assign n12863 = n3247 & n5369;
assign n6688 = n5891 | n8836;
assign n13900 = n7401 | n8873;
assign n12709 = n3394 | n11432;
assign n14414 = n10647 & n11448;
assign n3922 = ~n2816;
assign n12912 = ~(n3530 | n9707);
assign n1449 = n5279 & n6581;
assign n265 = n7673 & n6998;
assign n5756 = n7612 & n14283;
assign n189 = n5409 | n7214;
assign n10519 = ~(n6088 | n10774);
assign n14514 = n523 | n7680;
assign n13784 = ~n14133;
assign n1378 = ~n14071;
assign n5615 = n8592 | n13462;
assign n2864 = n12057 & n1922;
assign n6983 = n511 | n7311;
assign n2888 = ~n11331;
assign n1818 = ~(n12999 | n11198);
assign n14491 = n4357 | n502;
assign n3763 = n2318 | n9381;
assign n4448 = n5779 & n3699;
assign n9599 = n1051 | n3064;
assign n5331 = n5695 | n8426;
assign n10399 = ~n5182;
assign n14335 = n11909 | n7287;
assign n1029 = n13531 | n10576;
assign n6458 = n11722 | n7561;
assign n10177 = ~n14071;
assign n13783 = n12047 | n2365;
assign n5687 = n4803 & n9020;
assign n11941 = n13547 | n5933;
assign n9942 = n14093 & n8284;
assign n833 = n7426 | n11694;
assign n13878 = n6243 & n12663;
assign n1671 = n4092 | n1464;
assign n7868 = n3062 | n6902;
assign n4735 = n6629 | n10043;
assign n9439 = ~(n11581 | n1463);
assign n2705 = n533 & n13794;
assign n6420 = n2694 | n11968;
assign n8597 = n9890 & n10117;
assign n3133 = n13707 | n9476;
assign n3234 = ~n2788;
assign n4227 = n5553 & n7446;
assign n9469 = n1428 & n10957;
assign n11808 = n12039 & n2399;
assign n830 = n4807 | n10610;
assign n14031 = n3608 | n12025;
assign n6887 = ~(n2341 | n12099);
assign n4018 = ~n2432;
assign n3808 = n11171 | n3123;
assign n7661 = ~(n5569 | n12666);
assign n9876 = n12131 | n10101;
assign n11817 = n3212 & n3304;
assign n7749 = n6288 | n13025;
assign n12551 = n4156 & n9781;
assign n9889 = n6822 & n11380;
assign n11412 = ~n13213;
assign n1043 = n14042 & n13921;
assign n3208 = n747 | n9023;
assign n14191 = n1788 & n3023;
assign n60 = n10224 | n3647;
assign n1253 = n4162 | n13106;
assign n4976 = n7961 & n9868;
assign n4664 = ~(n9577 | n11796);
assign n2865 = n7079 & n10218;
assign n6990 = ~n4966;
assign n7922 = n4822 | n7236;
assign n3015 = ~n9810;
assign n13476 = ~n3870;
assign n11163 = ~n1955;
assign n3455 = n6903 & n10751;
assign n1339 = ~n9613;
assign n10721 = n8630 & n6353;
assign n13957 = n3320 | n11555;
assign n14061 = n8300 & n7492;
assign n5710 = ~n2794;
assign n9883 = n2583 & n12803;
assign n1414 = ~n6559;
assign n1469 = n7963 & n11981;
assign n8819 = n6428 | n5387;
assign n4563 = n6649 & n10118;
assign n9425 = n954 | n12145;
assign n12749 = ~(n478 | n11747);
assign n14148 = n7862 | n13054;
assign n12924 = n1640 & n7590;
assign n11852 = ~n3130;
assign n8760 = n5362 | n13459;
assign n12111 = n12852 & n9837;
assign n11969 = ~n1079;
assign n6295 = n14150 & n5804;
assign n11499 = n9113 & n8266;
assign n3067 = n820 | n9812;
assign n10475 = ~(n3546 | n4782);
assign n12258 = n432 & n1572;
assign n4516 = n2445 & n3144;
assign n8605 = ~n6829;
assign n2546 = n2686 | n9348;
assign n7474 = ~(n438 | n396);
assign n4848 = ~(n1023 | n4090);
assign n8978 = n7826 & n639;
assign n1670 = n646 & n1971;
assign n6185 = n9941 & n12126;
assign n7412 = n11303 | n6836;
assign n7163 = n6606 & n5689;
assign n13807 = ~(n8816 | n13526);
assign n8091 = n2099 & n13971;
assign n1475 = n10713 | n2775;
assign n5438 = n1278 & n14023;
assign n6513 = ~(n11628 | n6300);
assign n312 = ~(n1722 | n13993);
assign n4298 = n8247 & n10995;
assign n7032 = n3846 & n7805;
assign n4748 = n7697 | n9383;
assign n2217 = n3193 | n2364;
assign n14041 = n533 & n14409;
assign n5060 = n4806 & n5403;
assign n3672 = ~n13383;
assign n14291 = n9442 | n12660;
assign n13072 = ~n12897;
assign n3692 = n3134 | n9886;
assign n7088 = n6957 & n12545;
assign n9935 = n2510 | n10592;
assign n1143 = n9275 & n9319;
assign n892 = n8393 & n2507;
assign n11259 = ~n6364;
assign n8334 = ~(n9967 | n13842);
assign n239 = ~n5306;
assign n10604 = ~(n14466 | n8984);
assign n652 = n12968 | n5126;
assign n5278 = ~n7704;
assign n543 = n5185 & n4035;
assign n13554 = n4932 & n14008;
assign n492 = ~n1010;
assign n995 = n2006 & n10868;
assign n3215 = n10820 & n11863;
assign n6698 = n8183 & n12144;
assign n1553 = ~(n2822 | n6456);
assign n8461 = n12351 | n7251;
assign n11684 = n4018 & n1229;
assign n4214 = n6898 & n11692;
assign n6314 = n6999 & n10290;
assign n13449 = n4876 | n12110;
assign n6523 = n10083 | n11740;
assign n5966 = ~(n14466 | n3844);
assign n11165 = ~(n9423 | n360);
assign n3591 = n12611 & n13865;
assign n9631 = ~(n8353 | n3510);
assign n9773 = n9724 & n13431;
assign n3096 = n11551 | n2385;
assign n4623 = n3320 | n12465;
assign n10099 = ~n14524;
assign n2543 = ~(n4200 | n8671);
assign n13643 = n14107 | n7547;
assign n2617 = ~(n619 | n10481);
assign n12422 = n8697 & n12732;
assign n8483 = n10763 & n12429;
assign n10760 = ~n10573;
assign n11406 = ~n2497;
assign n8784 = ~(n13435 | n1234);
assign n1004 = ~(n1838 | n11280);
assign n1539 = ~n1342;
assign n13819 = n348 | n8439;
assign n6150 = n12015 & n7019;
assign n4246 = n317 | n365;
assign n7857 = n11422 & n12518;
assign n14402 = n1428 & n3430;
assign n11537 = n9726 & n1605;
assign n8120 = n1775 & n13288;
assign n8523 = n646 & n9415;
assign n3465 = n7609 | n4656;
assign n6500 = n11123 | n4084;
assign n1622 = n501 & n8478;
assign n12011 = n10032 & n5254;
assign n851 = n11510 | n13040;
assign n11334 = n227 | n8972;
assign n1839 = ~(n7809 | n7277);
assign n8272 = n8822 & n5412;
assign n1793 = n14521 & n659;
assign n6825 = n9265 & n8416;
assign n2613 = n11647 | n1799;
assign n6909 = ~n3388;
assign n12281 = n194 | n5565;
assign n9972 = ~n10469;
assign n9807 = ~n11813;
assign n1406 = n3861 & n8170;
assign n2990 = ~(n7662 | n7843);
assign n10542 = ~(n12112 | n1798);
assign n635 = n10854 & n9204;
assign n4971 = n1222 & n2034;
assign n1998 = n14366 | n9643;
assign n5890 = n13404 & n1787;
assign n5625 = ~n4550;
assign n2170 = ~(n12651 | n2360);
assign n11744 = n3164 | n14382;
assign n1809 = n13991 | n926;
assign n12843 = n8855 & n11334;
assign n313 = n4806 & n4048;
assign n13437 = ~n4535;
assign n6455 = n11008 & n7121;
assign n5390 = n9218 | n4315;
assign n10266 = n1834 | n4224;
assign n2104 = ~(n7365 | n8146);
assign n13436 = n10394 | n9842;
assign n13051 = n9289 | n3916;
assign n12730 = ~n1813;
assign n14223 = n2387 | n2273;
assign n10388 = n10229 & n1864;
assign n10783 = n9069 & n12618;
assign n11770 = ~(n9124 | n3735);
assign n11150 = n3025 | n12609;
assign n7307 = n1741 | n4666;
assign n1383 = ~n5242;
assign n9298 = n7462 | n11781;
assign n2123 = ~(n10977 | n11056);
assign n5543 = n2111 | n7716;
assign n11369 = ~n9971;
assign n5789 = n2784 | n3767;
assign n7599 = n4627 & n14138;
assign n12253 = ~(n5024 | n5381);
assign n3745 = n9211 | n9720;
assign n7049 = n7081 & n6611;
assign n12542 = ~n14501;
assign n8103 = n12353 | n6281;
assign n5525 = ~n1311;
assign n2175 = n13890 & n9047;
assign n1681 = ~n14512;
assign n5819 = n9811 & n9164;
assign n12552 = n4481 | n9666;
assign n7368 = n8431 & n3678;
assign n7687 = ~(n11713 | n9094);
assign n1283 = ~(n11094 | n7962);
assign n325 = n10302 & n5263;
assign n856 = n4045 | n12153;
assign n6872 = n5491 | n3151;
assign n9926 = n9230 | n6895;
assign n13833 = n251 | n213;
assign n7708 = ~n6270;
assign n2358 = n8517 | n2995;
assign n5133 = n7436 | n3540;
assign n7724 = n3126 | n7005;
assign n3342 = n4684 | n9801;
assign n9766 = ~n10050;
assign n8894 = n1428 & n12631;
assign n13063 = ~(n7660 | n5128);
assign n13865 = n10808 | n8993;
assign n7601 = ~(n12651 | n4212);
assign n13808 = n6085 | n9179;
assign n6408 = n8907 & n11660;
assign n9389 = n3134 | n2145;
assign n6734 = n13720 | n3673;
assign n11561 = n13220 | n3141;
assign n1784 = ~n12175;
assign n3124 = n1838 | n285;
assign n10473 = n4018 & n5661;
assign n8642 = n11020 & n3650;
assign n3458 = ~(n355 | n14476);
assign n12810 = n2177 & n14322;
assign n5160 = n14303 | n7667;
assign n7849 = n7438 | n11289;
assign n14111 = n2082 & n5067;
assign n1048 = n10539 | n2516;
assign n2235 = ~(n2790 | n3372);
assign n1586 = n3672 & n8069;
assign n6333 = n9972 & n208;
assign n13490 = n1071 & n10976;
assign n14238 = ~n4906;
assign n10205 = n1051 | n7866;
assign n11001 = n7798 & n12937;
assign n9248 = n748 & n12534;
assign n4139 = n13823 & n13424;
assign n12195 = n10332 & n13599;
assign n10210 = n1138 & n4386;
assign n6108 = n7862 | n3637;
assign n7379 = n9102 & n9775;
assign n4821 = ~n11415;
assign n2140 = n10234 | n8046;
assign n4904 = n4844 & n921;
assign n12055 = ~(n11713 | n13630);
assign n5669 = ~(n742 | n8058);
assign n10365 = n4261 & n5994;
assign n12435 = ~n8799;
assign n7971 = ~n2794;
assign n9067 = n541 & n5415;
assign n13359 = ~n13181;
assign n294 = n8300 & n10393;
assign n12307 = n9747 | n3116;
assign n809 = ~(n8419 | n12785);
assign n4359 = ~n4824;
assign n4170 = n3011 | n8333;
assign n1657 = n9423 | n10779;
assign n12442 = n4525 & n13149;
assign n8164 = n10969 & n8392;
assign n9302 = n6822 & n463;
assign n14453 = n2025 | n7461;
assign n13215 = n11576 | n3052;
assign n12345 = n12132 | n3166;
assign n3330 = n13108 | n12065;
assign n7148 = n7116 | n6317;
assign n3273 = ~n12489;
assign n1589 = n14400 | n13541;
assign n13834 = n10136 | n3912;
assign n12934 = ~n12588;
assign n14495 = n3527 | n7516;
assign n9125 = n12549 | n8775;
assign n8271 = n9069 & n9539;
assign n7503 = n5918 & n12239;
assign n14242 = n8964 | n1032;
assign n227 = ~n6274;
assign n12838 = ~(n3443 | n5941);
assign n8516 = n11674 & n5352;
assign n6677 = ~(n10285 | n10641);
assign n3806 = n7443 & n7526;
assign n1364 = n13367 & n3254;
assign n1518 = n10032 & n7976;
assign n1217 = n9230 | n11940;
assign n14202 = n8301 | n11696;
assign n5268 = ~n11375;
assign n13854 = ~n4891;
assign n12493 = n5240 & n9926;
assign n5951 = ~n2371;
assign n8314 = n3099 | n3481;
assign n14010 = n7693 & n13137;
assign n11444 = ~n5217;
assign n12464 = n2025 | n10899;
assign n7300 = n48 | n9869;
assign n13282 = n3800 | n13837;
assign n4070 = n12295 | n8853;
assign n6035 = n12149 | n7387;
assign n12710 = n9198 & n4800;
assign n13922 = n392 & n9212;
assign n2857 = ~n10346;
assign n14071 = n1011 & n9658;
assign n6789 = n6111 | n5862;
assign n126 = n4022 & n2664;
assign n1615 = ~(n228 | n14228);
assign n1154 = n392 & n216;
assign n6235 = n5053 & n13088;
assign n2806 = n11569 & n12839;
assign n2796 = n4422 & n9331;
assign n13877 = ~n7120;
assign n10557 = n2961 & n12017;
assign n11204 = n10857 | n8123;
assign n7783 = ~(n5833 | n10001);
assign n5030 = n9724 & n12337;
assign n13696 = n9829 & n5148;
assign n643 = n1193 & n13515;
assign n12475 = ~n1571;
assign n1920 = ~n9110;
assign n13588 = n6695 | n13179;
assign n3160 = n7462 | n290;
assign n12438 = n12259 & n11807;
assign n1593 = n13083 | n653;
assign n1124 = n271 & n9765;
assign n11831 = n387 | n11599;
assign n7611 = n185 | n2324;
assign n11636 = ~n13219;
assign n27 = n12421 & n4770;
assign n7674 = n1699 & n13032;
assign n6208 = n1028 | n106;
assign n8834 = n9864 | n5792;
assign n13424 = n3168 | n9028;
assign n12231 = n7057 & n14371;
assign n6628 = n8581 | n5080;
assign n2876 = n7779 & n7932;
assign n12291 = n4684 | n14381;
assign n13281 = n3120 | n12369;
assign n11437 = n4739 | n4938;
assign n7462 = ~n1060;
assign n9328 = ~(n4741 | n1012);
assign n3920 = ~(n10511 | n12283);
assign n4738 = ~(n7223 | n3909);
assign n10430 = n3715 & n8040;
assign n3454 = n12139 | n3828;
assign n539 = n7957 & n806;
assign n8772 = n11710 | n9049;
assign n1377 = n4320 | n11666;
assign n13070 = ~(n1722 | n3639);
assign n2261 = n4244 & n273;
assign n9369 = n3861 & n1596;
assign n862 = n4045 | n7451;
assign n13489 = ~n4490;
assign n13284 = n13142 | n11823;
assign n12833 = n7267 & n13136;
assign n2838 = n4255 | n9911;
assign n4633 = ~n1544;
assign n7349 = n8849 & n5514;
assign n12834 = n2322 & n3071;
assign n9521 = ~(n1769 | n86);
assign n1645 = n13432 | n2659;
assign n2361 = n3212 & n1817;
assign n574 = n10399 & n4526;
assign n3816 = ~(n11771 | n11275);
assign n3316 = n7250 | n5737;
assign n11674 = ~n6829;
assign n11690 = n10713 | n1558;
assign n5971 = n9780 | n2828;
assign n2182 = n10855 & n4834;
assign n7335 = n3405 & n3160;
assign n6857 = ~n4720;
assign n10439 = n11459 | n9510;
assign n9662 = n10854 & n529;
assign n835 = n9315 & n11806;
assign n5220 = n1261 | n4567;
assign n12787 = n12721 & n3827;
assign n3457 = ~n7546;
assign n10645 = n2181 | n13057;
assign n1452 = ~n1843;
assign n551 = n5240 & n5337;
assign n6342 = n7911 & n9258;
assign n5717 = n2057 | n13950;
assign n12480 = ~n13364;
assign n8783 = n1202 | n1736;
assign n4721 = n1804 & n2980;
assign n7665 = n695 | n1465;
assign n2633 = n12935 & n1068;
assign n8632 = n12592 & n5056;
assign n232 = n5252 & n2430;
assign n5305 = n7227 | n3999;
assign n2867 = n6971 | n4470;
assign n9782 = n11223 | n4952;
assign n6840 = ~(n11580 | n7625);
assign n10561 = n1258 | n2220;
assign n3328 = n14388 & n2469;
assign n10581 = n6316 & n3985;
assign n3666 = n8020 & n5896;
assign n13896 = n7430 | n7664;
assign n919 = ~n8814;
assign n2975 = n638 & n5699;
assign n5388 = n13572 & n12996;
assign n13361 = ~n7376;
assign n13144 = n9113 & n12997;
assign n5335 = ~n8963;
assign n2450 = n2412 | n6733;
assign n6311 = ~n5427;
assign n5942 = n10678 & n11549;
assign n3148 = ~(n10650 | n7567);
assign n1050 = ~(n11259 | n4344);
assign n12433 = ~(n4092 | n3971);
assign n2722 = n10562 & n1645;
assign n9527 = n5071 & n12849;
assign n2701 = n12259 & n13410;
assign n1543 = n986 & n12064;
assign n3276 = ~n11668;
assign n8821 = ~n622;
assign n3701 = n9747 | n11736;
assign n11382 = n1231 & n10009;
assign n7311 = n8432 & n4241;
assign n14127 = n5587 | n226;
assign n14447 = n7529 & n13665;
assign n1796 = n5997 | n13638;
assign n370 = n4840 | n8371;
assign n8246 = n904 & n6294;
assign n8355 = n172 | n9902;
assign n1248 = n1538 | n13289;
assign n5317 = ~n7346;
assign n2645 = ~n426;
assign n1170 = n8147 & n9367;
assign n13869 = ~n394;
assign n8531 = n12592 & n2203;
assign n1162 = n10209 & n7423;
assign n13374 = n3025 | n11115;
assign n13668 = n2967 & n12924;
assign n13596 = ~(n9557 | n1953);
assign n2028 = n6486 & n13801;
assign n5983 = n4359 & n13451;
assign n5224 = n5471 & n3330;
assign n13241 = n8047 & n12653;
assign n7625 = ~(n11988 | n4108);
assign n6621 = n3219 | n10833;
assign n6465 = n873 & n83;
assign n8056 = n10763 & n284;
assign n7640 = n103 & n11294;
assign n7615 = n10534 | n2500;
assign n6636 = n13863 & n7133;
assign n12615 = ~n6193;
assign n9756 = n10024 | n5578;
assign n5169 = n11008 & n14090;
assign n8250 = ~n230;
assign n6811 = n14449 | n4948;
assign n8754 = n6128 & n13482;
assign n3374 = n1772 & n4106;
assign n1156 = n6781 | n8823;
assign n2432 = ~n10861;
assign n1274 = ~(n4050 | n956);
assign n614 = n11647 | n7411;
assign n11601 = n10784 | n3289;
assign n5805 = ~(n12075 | n2209);
assign n686 = n12730 & n10551;
assign n4271 = n3536 & n10139;
assign n8519 = n7063 & n11346;
assign n10843 = ~(n1860 | n7204);
assign n14030 = n3527 | n1082;
assign n1024 = n12421 & n10170;
assign n2551 = n9315 & n11307;
assign n6041 = ~n13779;
assign n9232 = ~n10269;
assign n1531 = n1610 & n14315;
assign n12262 = n14435 | n4129;
assign n4799 = n7527 | n4979;
assign n6651 = n13847 | n14180;
assign n8305 = n12250 & n5671;
assign n13504 = n1125 & n1863;
assign n11538 = ~(n5159 | n11657);
assign n5327 = n11551 | n6592;
assign n775 = n5507 | n10696;
assign n12784 = n3813 & n190;
assign n4992 = n3088 | n10337;
assign n6269 = ~(n1681 | n6133);
assign n13283 = ~n1073;
assign n5440 = n12472 & n14053;
assign n7656 = n5986 | n10306;
assign n4605 = n7914 | n4736;
assign n14298 = n12034 | n14010;
assign n8658 = n8816 | n12313;
assign n11633 = n13186 | n8439;
assign n3468 = n10457 & n12085;
assign n10342 = ~n2607;
assign n774 = n11163 & n1470;
assign n11255 = n3586 & n1330;
assign n2880 = ~(n10289 | n6702);
assign n7425 = n10913 | n551;
assign n2731 = n3652 | n3799;
assign n6737 = n12998 & n13344;
assign n11681 = ~(n1685 | n10885);
assign n7647 = n8147 & n12814;
assign n3680 = n5948 & n8744;
assign n12732 = n11647 | n5028;
assign n7045 = n3062 | n64;
assign n12496 = n9174 | n6367;
assign n5784 = ~(n12191 | n4463);
assign n9001 = n85 | n5820;
assign n6895 = n9617 & n8760;
assign n678 = ~n11969;
assign n1458 = ~n14181;
assign n6871 = n13941 | n3966;
assign n8792 = n11472 | n3753;
assign n11103 = n251 | n12843;
assign n2817 = n11581 | n14117;
assign n1957 = n6350 | n8205;
assign n12136 = n4172 | n74;
assign n11534 = n6436 & n8298;
assign n8625 = n5948 & n5021;
assign n11772 = ~(n13979 | n7207);
assign n11638 = n4052 | n654;
assign n13746 = n7358 | n4027;
assign n10292 = n3286 & n1635;
assign n5171 = n8450 | n10378;
assign n307 = n4065 | n3732;
assign n5157 = n7678 | n12405;
assign n11692 = n4631 | n2586;
assign n11513 = n1937 & n5770;
assign n1477 = n4828 | n7986;
assign n13981 = ~n4500;
assign n4397 = n5071 & n3664;
assign n3043 = ~n5023;
assign n79 = ~n5795;
assign n8092 = n10229 & n3761;
assign n12646 = n2682 & n4097;
assign n12538 = n12019 | n5165;
assign n10864 = ~n2752;
assign n10632 = n14042 & n113;
assign n708 = ~(n7900 | n11267);
assign n14412 = n2951 & n10403;
assign n3424 = ~n6193;
assign n3356 = ~n5761;
assign n10411 = n9529 | n7100;
assign n4548 = n7284 & n440;
assign n11759 = n6654 | n4251;
assign n10773 = n13698 | n13006;
assign n4512 = n9507 | n5913;
assign n10644 = n9890 & n12951;
assign n7231 = n3986 & n4070;
assign n12963 = n8250 & n175;
assign n9350 = n7230 | n702;
assign n157 = n6318 & n9491;
assign n13073 = n3405 & n846;
assign n1942 = n6343 & n9678;
assign n5484 = n6848 | n12782;
assign n3576 = n7203 & n13550;
assign n9548 = n5317 & n2335;
assign n3475 = ~(n1357 | n7184);
assign n7574 = n8517 | n10581;
assign n13429 = n3673 | n5023;
assign n10403 = n10953 & n5226;
assign n7215 = n8581 | n5814;
assign n8830 = n974 | n1754;
assign n8182 = n7187 & n11323;
assign n1453 = n13626 & n13838;
assign n12979 = ~(n3107 | n7234);
assign n4680 = n6519 | n10665;
assign n11326 = n11047 | n3004;
assign n1480 = ~n5627;
assign n2310 = ~n8008;
assign n13699 = n5483 | n9064;
assign n434 = n9490 | n9914;
assign n6053 = ~n10254;
assign n12696 = n8242 | n7288;
assign n10106 = ~(n2236 | n13358);
assign n4906 = ~n11628;
assign n1142 = n13342 & n3998;
assign n3656 = n14481 | n6505;
assign n7326 = n4722 & n7688;
assign n9602 = n12625 | n6735;
assign n11581 = ~n11055;
assign n4551 = n8569 & n3593;
assign n4514 = n8748 | n3611;
assign n2904 = ~n1495;
assign n8307 = n11636 & n6190;
assign n1225 = ~n10283;
assign n8951 = n5362 | n2637;
assign n6324 = ~(n6397 | n1519);
assign n9526 = n11838 & n2114;
assign n7288 = n11153 & n14443;
assign n1863 = n11090 | n5534;
assign n121 = n6519 | n880;
assign n12228 = n10024 | n8098;
assign n9738 = n2760 | n13509;
assign n9803 = ~n7450;
assign n11169 = n2058 & n625;
assign n12226 = ~n6139;
assign n12705 = ~n12691;
assign n14125 = n3932 & n3241;
assign n9443 = n5053 & n7646;
assign n1569 = n1172 | n3567;
assign n13911 = n8786 & n12954;
assign n6013 = ~n9950;
assign n11777 = n12400 | n4451;
assign n3153 = n7284 & n4798;
assign n13949 = n7803 | n14294;
assign n2899 = ~(n13627 | n709);
assign n3578 = n14282 | n7750;
assign n9353 = ~n9169;
assign n5087 = n3273 | n12787;
assign n5063 = n8045 | n9548;
assign n9113 = ~n5268;
assign n4763 = n7708 & n1755;
assign n5069 = ~(n5132 | n8101);
assign n10498 = n706 & n10706;
assign n9174 = ~n6332;
assign n12322 = n10407 | n4659;
assign n8386 = ~n9197;
assign n7292 = n8581 | n3911;
assign n14166 = ~n12687;
assign n7302 = n706 & n10690;
assign n1390 = ~(n12112 | n7985);
assign n4939 = n9516 & n7336;
assign n1773 = n4757 & n8095;
assign n12563 = n6130 & n13100;
assign n7219 = ~n6357;
assign n1306 = n14419 | n12824;
assign n6916 = n8332 | n105;
assign n6225 = n7391 & n2708;
assign n5238 = n11036 | n12003;
assign n717 = ~n8291;
assign n14267 = n5475 & n2773;
assign n5323 = ~(n13072 | n9033);
assign n200 = ~n8048;
assign n10869 = n2521 & n6792;
assign n14407 = n3028 & n6042;
assign n5044 = n5800 | n13545;
assign n13391 = n1962 & n10476;
assign n1456 = n11803 & n12578;
assign n2438 = n7529 & n8173;
assign n8118 = n838 | n12921;
assign n11218 = n11479 | n8463;
assign n4417 = ~n93;
assign n6482 = n7934 & n3929;
assign n9251 = n646 & n5659;
assign n11351 = n8821 | n12006;
assign n6099 = ~n4656;
assign n12994 = ~n1220;
assign n12758 = ~(n10189 | n5299);
assign n10155 = n11980 | n2574;
assign n3731 = n6318 & n11955;
assign n1278 = ~n4785;
assign n7257 = n4722 & n2652;
assign n9347 = n8111 & n8807;
assign n3235 = ~(n1112 | n2579);
assign n12194 = ~(n946 | n12940);
assign n9842 = n3536 & n9935;
assign n847 = n7481 | n2997;
assign n12340 = n14107 | n5581;
assign n9202 = n10523 | n1580;
assign n1100 = ~n6326;
assign n14441 = n638 & n10297;
assign n11586 = n10622 & n6183;
assign n3997 = ~(n7720 | n11353);
assign n5675 = ~n13560;
assign n11616 = n7015 & n11846;
assign n5470 = n13547 | n6235;
assign n10200 = ~(n13350 | n1472);
assign n6336 = n8605 & n8560;
assign n8040 = n7219 | n351;
assign n14024 = n6989 | n30;
assign n13164 = n1937 & n6576;
assign n5459 = ~n10828;
assign n11418 = ~(n8607 | n1056);
assign n5115 = n10134 & n13217;
assign n11136 = n13535 & n1973;
assign n5103 = n6595 | n3796;
assign n1437 = n7691 & n5487;
assign n6199 = ~(n5480 | n2512);
assign n4121 = n5779 & n1130;
assign n3735 = ~(n48 | n11486);
assign n6739 = n14063 & n14439;
assign n12208 = n11093 & n5813;
assign n680 = n3846 & n4863;
assign n13038 = ~n6308;
assign n1906 = n13252 & n8394;
assign n9573 = n2527 & n14424;
assign n2822 = ~n481;
assign n12243 = ~n2009;
assign n5736 = n9102 & n5039;
assign n7820 = n85 | n12027;
assign n13441 = n10815 & n8192;
assign n5282 = n9890 & n2614;
assign n891 = n13706 | n8109;
assign n10575 = n3219 | n1454;
assign n7964 = n7421 & n7356;
assign n13095 = n769 | n4794;
assign n7895 = n12445 & n10037;
assign n2328 = n13240 & n12199;
assign n9619 = n2367 & n1188;
assign n9462 = n7249 | n3059;
assign n7130 = ~n8446;
assign n303 = n4365 | n7652;
assign n5849 = ~(n9529 | n5741);
assign n1129 = n12013 & n12419;
assign n12861 = n2645 | n9534;
assign n11026 = n11951 | n6366;
assign n10818 = n13525 & n11075;
assign n1391 = ~n9686;
assign n14018 = n8247 & n11895;
assign n700 = ~n201;
assign n13702 = n8427 & n1276;
assign n383 = n3826 | n7089;
assign n6181 = n1061 | n5292;
assign n6102 = n9211 | n3486;
assign n4186 = n541 & n12246;
assign n2781 = ~n6670;
assign n12692 = n5569 | n11709;
assign n4734 = n4289 & n6628;
assign n11292 = n9052 & n332;
assign n12286 = ~(n2017 | n237);
assign n922 = n7700 | n12583;
assign n7894 = ~(n4639 | n7355);
assign n6021 = n7116 | n14432;
assign n11773 = n10449 | n1016;
assign n13914 = n4445 & n4068;
assign n3239 = ~(n3255 | n7608);
assign n12361 = n12695 | n11395;
assign n11892 = n8332 | n8030;
assign n7275 = ~n13765;
assign n11079 = ~(n14058 | n322);
assign n1758 = ~(n12334 | n9007);
assign n12211 = ~n1220;
assign n9533 = n11804 | n7025;
assign n10088 = n5475 & n7307;
assign n12959 = n12592 & n6530;
assign n9160 = n6690 | n33;
assign n5748 = ~(n9807 | n7136);
assign n4293 = n7076 | n148;
assign n8456 = n4822 | n8995;
assign n10237 = n10089 | n11005;
assign n2883 = n2521 & n11083;
assign n10332 = ~n168;
assign n13781 = ~n12970;
assign n9946 = n1452 & n9363;
assign n2004 = n12960 & n4378;
assign n786 = n1937 & n649;
assign n6470 = n7208 & n9797;
assign n7966 = n3273 | n13122;
assign n7193 = n6206 | n10206;
assign n6201 = n12185 & n12458;
assign n8070 = n2422 & n9518;
assign n4716 = n6388 | n1568;
assign n9447 = n12782 & n9276;
assign n2308 = n9315 & n10716;
assign n5130 = n9972 & n12464;
assign n2060 = n4655 & n10533;
assign n6580 = n11231 | n12877;
assign n4791 = ~n12489;
assign n9180 = n13421 & n4801;
assign n345 = n13501 | n3020;
assign n9642 = n3710 & n7033;
assign n867 = n5144 | n3006;
assign n13417 = n6672 | n7542;
assign n7750 = n4422 & n1184;
assign n8253 = n898 & n12783;
assign n14056 = n172 | n3200;
assign n2671 = n2021 & n14025;
assign n11943 = n7909 & n10454;
assign n1694 = ~(n5035 | n2028);
assign n8937 = n1904 & n13341;
assign n5838 = n12625 | n2458;
assign n2226 = n3043 | n4225;
assign n10998 = n1011 | n8800;
assign n50 = n7219 | n10547;
assign n12044 = n6606 & n29;
assign n11364 = n5489 & n4119;
assign n10245 = ~n3007;
assign n139 = n6519 | n7738;
assign n6228 = ~(n900 | n2314);
assign n3199 = n8866 & n5576;
assign n5304 = n5483 | n5161;
assign n10770 = n11223 | n14234;
assign n13570 = n7370 & n5309;
assign n14299 = n6135 & n9162;
assign n1367 = n838 | n2440;
assign n8363 = ~n5690;
assign n12889 = n13501 | n14272;
assign n14275 = n5582 & n6154;
assign n11964 = ~(n9078 | n12979);
assign n2694 = ~n628;
assign n8557 = ~n9214;
assign n8196 = n8701 | n4959;
assign n13278 = ~(n2575 | n1233);
assign n4340 = ~n918;
assign n5832 = n1278 | n730;
assign n6929 = n4358 & n2821;
assign n3967 = ~n5886;
assign n10511 = ~n7291;
assign n11865 = n6507 & n9964;
assign n7779 = ~n2619;
assign n9420 = n8592 | n11770;
assign n5944 = ~n1979;
assign n8146 = ~(n1623 | n1852);
assign n4132 = n12185 & n4285;
assign n7874 = n10154 | n12607;
assign n76 = n4045 | n14021;
assign n5928 = n8964 | n6095;
assign n10483 = n7308 & n10518;
assign n3196 = ~n4711;
assign n2570 = n11620 | n3810;
assign n11445 = ~n12189;
assign n168 = ~n3331;
assign n1290 = n5084 | n3580;
assign n10017 = n3273 | n6180;
assign n12507 = n7429 & n11372;
assign n3436 = ~(n2086 | n302);
assign n9594 = n3914 | n5657;
assign n3902 = n8638 | n2650;
assign n11925 = n5348 & n3187;
assign n1146 = n2961 & n2702;
assign n9540 = n8378 | n849;
assign n11138 = n14481 | n1081;
assign n2759 = n573 | n13448;
assign n137 = n3724 & n8616;
assign n12410 = n555 | n1148;
assign n1476 = n8801 & n545;
assign n14341 = ~(n5217 | n459);
assign n2389 = n8769 & n470;
assign n10307 = n1855 | n11404;
assign n11878 = n3193 | n7789;
assign n12491 = n7359 | n4376;
assign n7194 = n5007 | n14146;
assign n1224 = n3846 & n6143;
assign n1235 = n8932 & n1281;
assign n4223 = n4095 & n5868;
assign n10637 = ~n10775;
assign n2433 = n13226 | n4647;
assign n2859 = n8412 & n9175;
assign n1310 = n12531 & n13612;
assign n2553 = n12401 | n6303;
assign n3554 = n8210 | n6772;
assign n1344 = ~(n2781 | n3924);
assign n2853 = n5252 & n12290;
assign n7248 = n12226 & n3337;
assign n5189 = n4481 | n12806;
assign n10963 = ~(n619 | n6419);
assign n10844 = n14419 | n5821;
assign n13787 = n2686 | n5000;
assign n2504 = n10854 & n21;
assign n10813 = n9811 & n5451;
assign n6120 = n8034 | n14247;
assign n7824 = n3168 | n5517;
assign n1592 = n2709 & n4981;
assign n4671 = ~(n10712 | n3231);
assign n11123 = ~n7875;
assign n14161 = n4840 | n3841;
assign n2317 = ~(n3696 | n5645);
assign n3484 = n3777 | n14179;
assign n8137 = n4509 & n14398;
assign n10425 = ~(n13276 | n1103);
assign n12359 = n9890 & n2153;
assign n14251 = n6090 | n8169;
assign n1206 = n5997 | n2884;
assign n594 = n13112 | n10279;
assign n1423 = ~n12714;
assign n3869 = n12169 | n3921;
assign n10806 = n8932 & n3858;
assign n4048 = n3886 | n2108;
assign n7128 = n5137 & n9511;
assign n11312 = n6629 | n10386;
assign n10810 = n2330 & n13282;
assign n11338 = n4289 & n2937;
assign n4601 = ~n14408;
assign n9840 = ~(n3845 | n8648);
assign n3254 = n8378 | n4262;
assign n14443 = n12695 | n2639;
assign n12091 = n11519 | n10225;
assign n11460 = n6527 & n1387;
assign n4285 = n12211 | n9559;
assign n10626 = ~n13234;
assign n14333 = ~(n13477 | n5864);
assign n12203 = n5999 & n5066;
assign n3198 = n2846 & n308;
assign n13456 = n3743 & n12873;
assign n3126 = ~n4939;
assign n14228 = ~(n4270 | n11727);
assign n4946 = n7812 | n14378;
assign n7138 = n930 | n9932;
assign n2835 = n1006 | n7827;
assign n12913 = n2761 | n3143;
assign n12513 = ~(n8361 | n12005);
assign n9115 = ~(n10936 | n8057);
assign n6572 = ~(n6672 | n5243);
assign n576 = n9442 | n1224;
assign n14123 = n4690 & n8870;
assign n2309 = n13754 | n2165;
assign n8404 = ~n918;
assign n11308 = n1932 & n5265;
assign n11597 = ~n9465;
assign n5703 = ~(n5977 | n2739);
assign n10356 = n5807 | n9584;
assign n5892 = n3861 & n800;
assign n8176 = n6013 & n10992;
assign n8053 = n5977 | n2764;
assign n2825 = n9650 & n13747;
assign n13521 = n6271 | n13242;
assign n1398 = n10622 & n9660;
assign n3305 = ~(n13557 | n10373);
assign n7594 = n11724 | n4165;
assign n8301 = ~n4939;
assign n2333 = n14213 & n1542;
assign n10464 = ~(n1820 | n10793);
assign n2284 = n14358 & n7029;
assign n5002 = n13518 | n10471;
assign n13912 = ~n6517;
assign n3601 = n2378 & n3067;
assign n7361 = n3923 & n11866;
assign n7769 = n10763 & n14127;
assign n7165 = n11406 & n5096;
assign n1849 = n5454 | n6066;
assign n8744 = n5144 | n6207;
assign n9812 = n9102 & n3508;
assign n9407 = n286 & n12595;
assign n930 = ~n3455;
assign n3291 = n7779 & n13275;
assign n13919 = n7430 | n719;
assign n9790 = n1526 & n13094;
assign n2778 = n8620 & n4975;
assign n13775 = n3286 & n11769;
assign n5415 = n1383 | n12901;
assign n1918 = n12092 & n11077;
assign n4373 = n9792 | n13992;
assign n14046 = n3088 | n6826;
assign n794 = n5570 | n2479;
assign n8001 = n2643 & n1811;
assign n7495 = n4791 | n11089;
assign n10038 = n5088 & n9384;
assign n1443 = n8908 | n114;
assign n3406 = n11484 & n8718;
assign n1484 = n10534 | n5973;
assign n3082 = n13755 & n14152;
assign n8581 = ~n6274;
assign n6229 = n2564 & n3674;
assign n9524 = n12472 & n7301;
assign n10330 = ~n7802;
assign n5993 = n8638 | n6346;
assign n4700 = n6854 & n4100;
assign n8332 = ~n4317;
assign n660 = n2179 | n12287;
assign n5546 = n5471 & n6017;
assign n1220 = n10012 & n887;
assign n784 = n2983 & n4946;
assign n7767 = ~n7920;
assign n9148 = n11405 | n4329;
assign n3761 = n11105 | n274;
assign n10716 = n11048 | n7847;
assign n9326 = n12105 & n13374;
assign n8328 = n5071 & n14192;
assign n10339 = n476 | n13542;
assign n10560 = ~n12588;
assign n14014 = n5253 | n5501;
assign n9138 = n4365 & n9270;
assign n12372 = n13991 | n4989;
assign n8566 = n13404 & n7226;
assign n569 = n1044 | n6483;
assign n7848 = n1576 | n5653;
assign n8352 = ~(n14058 | n14434);
assign n4442 = n8950 & n1512;
assign n872 = n12500 | n6255;
assign n1348 = n2201 | n6147;
assign n616 = n4180 | n1688;
assign n2163 = ~(n4771 | n9838);
assign n14479 = n1414 & n7790;
assign n6582 = n10399 & n5123;
assign n9085 = n8458 | n2482;
assign n974 = ~n6978;
assign n8459 = ~(n7683 | n6195);
assign n13867 = ~n11666;
assign n11333 = n4289 & n4644;
assign n6667 = ~(n4417 | n4185);
assign n11243 = n14063 & n11850;
assign n11265 = n3569 | n7473;
assign n13573 = ~(n2684 | n9629);
assign n13595 = ~(n7624 | n6840);
assign n3062 = ~n4720;
assign n8606 = n11422 & n11006;
assign n1864 = n1494 | n5529;
assign n12164 = n791 | n10095;
assign n5517 = n7060 & n9825;
assign n6977 = n2518 | n12701;
assign n3842 = n14198 | n1413;
assign n11688 = ~n11529;
assign n9423 = ~n6274;
assign n8935 = n12990 & n1029;
assign n13261 = n1526 & n67;
assign n13735 = n8638 | n13995;
assign n1298 = n10302 & n1846;
assign n7125 = n6111 | n603;
assign n8194 = n2401 | n6868;
assign n14177 = n7076 | n5927;
assign n13885 = ~n12249;
assign n13928 = n1875 | n1585;
assign n9294 = n7693 & n12652;
assign n8185 = n13978 | n11563;
assign n13948 = n950 | n2662;
assign n11035 = n13118 | n5490;
assign n1355 = n10960 | n5882;
assign n4030 = n10763 & n14231;
assign n11665 = n7961 & n8351;
assign n4190 = n8151 | n2267;
assign n7756 = ~n8220;
assign n10889 = n7871 & n3015;
assign n3047 = ~n10108;
assign n9341 = n48 | n7707;
assign n7584 = n6517 | n6999;
assign n10551 = n14188 | n13496;
assign n2280 = n6167 & n870;
assign n6995 = n8786 & n8713;
assign n5559 = n12100 | n4384;
assign n5866 = n1840 | n12646;
assign n11881 = n7249 | n8188;
assign n2033 = n8849 & n2254;
assign n7139 = n6971 | n2120;
assign n12034 = ~n426;
assign n6691 = n6109 | n3334;
assign n12257 = n820 | n5736;
assign n14184 = n7227 | n3441;
assign n13632 = ~(n6428 | n13844);
assign n6549 = n4828 | n10849;
assign n12036 = n8386 & n11729;
assign n7920 = ~n5178;
assign n1820 = ~n6804;
assign n2225 = n3715 & n14316;
assign n9170 = ~(n3546 | n9090);
assign n13066 = n8250 & n1153;
assign n2144 = n5312 & n4820;
assign n8657 = n11117 | n3833;
assign n3644 = n10922 & n13512;
assign n10616 = n11329 & n10532;
assign n4203 = n4744 & n8049;
assign n13137 = n13501 | n7602;
assign n13328 = n14063 & n11293;
assign n4989 = n8427 & n7727;
assign n7872 = n8513 | n12725;
assign n6131 = n9102 & n2066;
assign n1462 = ~n7533;
assign n6351 = n9564 & n12496;
assign n1831 = n1223 | n7674;
assign n6527 = ~n11548;
assign n6232 = n13555 & n4461;
assign n4437 = n8044 & n11641;
assign n4617 = n6838 & n2835;
assign n13824 = n9620 | n5617;
assign n5986 = ~n238;
assign n5148 = ~n6266;
assign n1309 = ~(n6313 | n10785);
assign n10641 = ~(n5468 | n3928);
assign n1063 = ~(n13061 | n115);
assign n2696 = n2218 | n6227;
assign n12035 = ~(n10179 | n13438);
assign n2760 = ~n10426;
assign n3759 = n9620 | n6980;
assign n12473 = n6206 | n5760;
assign n14420 = n4899 | n7107;
assign n10821 = n5180 | n13319;
assign n3104 = ~(n2624 | n8564);
assign n12151 = n9052 & n5461;
assign n6383 = ~n10407;
assign n5414 = ~n5009;
assign n9455 = n5948 & n14298;
assign n5022 = ~(n2212 | n5735);
assign n13099 = n12425 & n8584;
assign n12859 = n3212 & n10063;
assign n14029 = ~n565;
assign n8074 = n4722 & n118;
assign n848 = ~n1093;
assign n4696 = ~(n2332 | n13371);
assign n1722 = ~n11493;
assign n7903 = n12353 | n2284;
assign n1862 = n13806 | n7101;
assign n12042 = ~n3309;
assign n13320 = n5458 & n12379;
assign n4730 = ~(n648 | n12315);
assign n3244 = n5857 & n5754;
assign n9273 = n11816 & n5666;
assign n1503 = n8980 | n9451;
assign n9218 = ~n4149;
assign n2905 = n7961 & n8013;
assign n1295 = n13446 | n13934;
assign n6558 = n7436 | n9784;
assign n819 = n12820 | n3573;
assign n4192 = n12764 | n11602;
assign n8584 = n390 | n10075;
assign n958 = n3755 & n3885;
assign n3756 = n2843 | n13562;
assign n4583 = n3099 | n4434;
assign n1995 = n1061 | n3503;
assign n10226 = n5603 | n3731;
assign n14472 = ~n1894;
assign n7448 = ~n53;
assign n9334 = n10197 & n6749;
assign n9788 = n7229 | n8346;
assign n7301 = n1258 | n180;
assign n12690 = n317 | n7167;
assign n4372 = n7914 | n9997;
assign n5643 = n457 & n6508;
assign n7716 = n10134 & n4113;
assign n9817 = n7911 & n10840;
assign n4621 = n9509 & n5103;
assign n12523 = n9853 & n10415;
assign n11967 = ~n2644;
assign n12143 = ~(n8511 | n1307);
assign n10165 = n1074 & n10838;
assign n6515 = ~(n12280 | n6358);
assign n5650 = n13520 & n1631;
assign n7897 = n14107 | n178;
assign n932 = n1699 & n11321;
assign n9616 = n4573 & n5127;
assign n5582 = ~n9046;
assign n690 = n12712 | n13667;
assign n8502 = n10936 | n1749;
assign n3717 = n12100 | n12203;
assign n4501 = n4359 & n12835;
assign n1032 = n2180 & n10772;
assign n6372 = n10458 & n10284;
assign n14137 = n10191 | n2504;
assign n11002 = n12353 | n8791;
assign n6742 = n1447 & n14039;
assign n95 = n11495 & n7098;
assign n3322 = n11724 | n1349;
assign n10428 = ~n12121;
assign n696 = n10394 | n11451;
assign n9588 = n8452 | n4206;
assign n7802 = ~n6364;
assign n11363 = n11411 & n9412;
assign n6200 = n10166 & n4472;
assign n13407 = ~n8555;
assign n6657 = ~n5872;
assign n8240 = n13706 | n14505;
assign n211 = n6838 & n347;
assign n2604 = n9953 & n2248;
assign n9491 = n2086 | n10185;
assign n12570 = n2709 & n9448;
assign n3570 = n8172 | n14149;
assign n9141 = n3169 & n5083;
assign n5330 = n8452 | n188;
assign n9048 = n3093 | n12762;
assign n2360 = ~(n14133 | n4142);
assign n8663 = ~n3587;
assign n13377 = ~(n12483 | n13337);
assign n5962 = n5986 | n6774;
assign n12301 = n5815 | n6689;
assign n10094 = n85 | n1143;
assign n10187 = n10933 | n9579;
assign n795 = ~(n5977 | n6887);
assign n4788 = ~n10269;
assign n7065 = ~n1357;
assign n8166 = n11607 & n11887;
assign n9584 = n3586 & n2787;
assign n12856 = n10815 & n2340;
assign n7788 = ~(n4046 | n3899);
assign n1404 = n3093 | n254;
assign n10091 = ~n8572;
assign n5008 = n4095 & n7525;
assign n3705 = n12494 | n3314;
assign n12392 = n9285 | n4675;
assign n3368 = n7429 & n10325;
assign n12724 = n1840 | n8060;
assign n1158 = n12018 & n2628;
assign n10132 = n12918 & n12760;
assign n5377 = n8575 | n4228;
assign n10613 = n6128 & n1525;
assign n450 = ~n14510;
assign n13785 = n11953 | n557;
assign n6915 = n12460 & n13655;
assign n13840 = ~n5185;
assign n1834 = ~n3070;
assign n9156 = n3561 | n14163;
assign n3140 = n8401 & n10298;
assign n1959 = n348 & n4949;
assign n1991 = n13535 & n4626;
assign n11891 = n2016 | n7469;
assign n3197 = n6822 & n12831;
assign n11029 = n4128 | n6793;
assign n7795 = n8111 & n1328;
assign n8294 = n13433 & n13580;
assign n13267 = n457 & n1097;
assign n12145 = n7768 & n236;
assign n12488 = n2272 | n10042;
assign n9763 = n12870 | n3471;
assign n13015 = n2750 | n1751;
assign n8133 = n12389 & n11182;
assign n1985 = n7230 & n7401;
assign n2109 = n10713 | n7273;
assign n4224 = n5926 & n6732;
assign n12683 = ~n7575;
assign n14054 = n9218 | n2033;
assign n10913 = ~n2970;
assign n11797 = n4276 & n11655;
assign n9053 = n718 & n1882;
assign n9011 = n839 | n2060;
assign n6177 = n12449 & n4728;
assign n5645 = n14357 & n5484;
assign n1534 = ~(n4207 | n4652);
assign n8343 = n5335 & n5835;
assign n13403 = n11620 | n3509;
assign n8311 = n2091 & n13990;
assign n2704 = n553 | n10096;
assign n5914 = ~(n6428 | n6622);
assign n1905 = n1662 & n11193;
assign n3770 = n10534 | n8228;
assign n6439 = n7284 & n11892;
assign n2265 = n14029 | n14048;
assign n10927 = n776 & n10472;
assign n1727 = n9188 & n3206;
assign n6248 = n2091 & n11485;
assign n12698 = n10781 | n13308;
assign n780 = n4822 | n12974;
assign n10556 = ~n9613;
assign n9398 = n11036 | n13849;
assign n10691 = n2820 & n2916;
assign n13993 = ~(n478 | n1899);
assign n9617 = ~n1436;
assign n6361 = n2177 & n9243;
assign n4710 = n7250 | n195;
assign n4582 = ~(n8663 | n9847);
assign n8942 = ~n1780;
assign n6155 = n1494 | n10898;
assign n6245 = n5454 | n4784;
assign n14466 = ~n10204;
assign n9655 = n4199 | n3266;
assign n11252 = n536 & n6652;
assign n8580 = ~n5549;
assign n13600 = n8923 & n722;
assign n14501 = ~n2257;
assign n13776 = ~(n11445 | n14324);
assign n474 = ~n5029;
assign n9528 = n7481 | n11387;
assign n2457 = n2694 | n14193;
assign n6867 = ~n6978;
assign n728 = n12295 | n1710;
assign n1252 = n7249 | n10865;
assign n3351 = ~(n2194 | n9888);
assign n607 = n5053 & n8230;
assign n455 = n12721 & n10249;
assign n5949 = n13432 | n391;
assign n9629 = ~(n1383 | n3621);
assign n7447 = n2897 | n14372;
assign n9358 = n9747 | n6624;
assign n8829 = ~(n6011 | n6116);
assign n5319 = n12018 & n9752;
assign n6086 = n333 & n12942;
assign n3690 = n11405 | n9728;
assign n5568 = n6838 & n4043;
assign n2444 = n2486 & n2673;
assign n2647 = n12101 & n11571;
assign n5363 = n2761 | n10265;
assign n1514 = n12990 & n1156;
assign n6495 = n2016 | n13595;
assign n7343 = n6690 | n7293;
assign n7080 = n4156 & n13211;
assign n10040 = n13112 | n14454;
assign n10236 = n1850 & n11852;
assign n5712 = ~(n2000 | n9909);
assign n7371 = ~(n9404 | n10811);
assign n8594 = ~(n228 | n10391);
assign n7457 = n2961 & n5156;
assign n13650 = ~n14293;
assign n12060 = ~(n4233 | n14080);
assign n2052 = ~(n1838 | n12035);
assign n8645 = ~(n11428 | n13986);
assign n10441 = ~(n3959 | n8874);
assign n9116 = n8301 | n378;
assign n10919 = n6271 | n12001;
assign n3107 = ~n1997;
assign n14405 = n12576 | n7543;
assign n7102 = n10556 & n2681;
assign n7281 = ~(n5160 | n7811);
assign n5812 = n2111 | n13500;
assign n3520 = n11093 & n7593;
assign n6089 = ~(n14198 | n1280);
assign n7698 = n12404 & n8348;
assign n13307 = n541 & n4556;
assign n12661 = n8453 & n912;
assign n1803 = n4195 | n10859;
assign n3480 = n4880 & n1191;
assign n4651 = ~(n6085 | n4944);
assign n540 = n4468 | n1170;
assign n3872 = n1876 & n8904;
assign n6516 = n3419 & n11;
assign n13024 = n3715 & n7435;
assign n1769 = ~n10380;
assign n13589 = n3826 | n13272;
assign n5959 = ~n6387;
assign n2159 = n10032 & n12325;
assign n5404 = ~(n14106 | n14271);
assign n10341 = n11362 & n1056;
assign n6529 = ~(n9529 | n7701);
assign n6655 = n10197 & n6843;
assign n3813 = ~n1473;
assign n10408 = ~n7275;
assign n955 = ~n9272;
assign n11329 = ~n13003;
assign n14240 = n8213 & n4479;
assign n6275 = n666 & n12627;
assign n12955 = ~(n4313 | n14186);
assign n6654 = ~n12588;
assign n5034 = n13597 & n11175;
assign n2898 = n5710 | n2827;
assign n14521 = ~n11961;
assign n10225 = n9107 | n2332;
assign n2484 = n3623 & n235;
assign n6335 = ~(n6030 | n7524);
assign n1661 = n8490 | n6726;
assign n804 = n4602 | n6479;
assign n9188 = ~n6819;
assign n2679 = n930 | n643;
assign n12675 = n13507 & n4831;
assign n6764 = n11472 | n574;
assign n8634 = n7443 & n13955;
assign n7996 = n1741 | n7968;
assign n4824 = ~n241;
assign n2059 = n11316 & n2288;
assign n7692 = ~(n3577 | n12978);
assign n9142 = ~n12025;
assign n355 = ~n7915;
assign n4241 = n10539 | n6850;
assign n3928 = ~(n13255 | n4280);
assign n2340 = n13978 | n12509;
assign n12596 = n3485 & n5745;
assign n6945 = n7961 & n7654;
assign n9277 = ~(n1914 | n3823);
assign n8599 = n5459 & n13643;
assign n2461 = ~n9865;
assign n136 = n8453 & n4750;
assign n1707 = ~(n5018 | n11562);
assign n2301 = n2643 & n73;
assign n4456 = n12857 & n6930;
assign n10191 = ~n628;
assign n10065 = ~(n8424 | n14254);
assign n13244 = ~(n5715 | n2245);
assign n9021 = ~(n13429 | n8901);
assign n10897 = ~n11325;
assign n14112 = ~(n12244 | n10830);
assign n12907 = n6531 & n1404;
assign n7034 = n4899 | n7224;
assign n4248 = n12927 | n10050;
assign n517 = n4358 & n12114;
assign n2910 = ~n7584;
assign n8742 = n3709 | n1763;
assign n1843 = ~n13425;
assign n2680 = n930 | n10067;
assign n9479 = n2901 | n13905;
assign n12857 = ~n11771;
assign n4820 = n11953 | n242;
assign n11125 = ~(n234 | n3252);
assign n6854 = ~n6807;
assign n12327 = n12449 & n7225;
assign n11179 = n11472 | n1437;
assign n9158 = n1962 & n14274;
assign n11697 = ~n1868;
assign n10846 = ~n4225;
assign n209 = n13978 | n2735;
assign n3399 = n2111 | n272;
assign n6402 = n11379 | n4425;
assign n550 = ~n5502;
assign n3627 = n12428 | n13866;
assign n7831 = n3405 & n13974;
assign n4838 = n11867 & n12628;
assign n1275 = n5491 | n12769;
assign n11336 = ~n2692;
assign n6795 = n3169 & n1400;
assign n13765 = n12528 & n1388;
assign n13851 = n129 & n8593;
assign n13599 = n2874 | n12217;
assign n2636 = n2486 & n1457;
assign n11283 = n3628 & n10307;
assign n12273 = ~(n3394 | n8466);
assign n545 = n11909 | n249;
assign n10216 = n4899 | n3757;
assign n4460 = n2531 | n14041;
assign n1964 = n6288 | n8413;
assign n1686 = ~n5195;
assign n5387 = n1924 & n3236;
assign n5685 = n4803 & n1671;
assign n12682 = n12820 | n4161;
assign n13394 = ~n10314;
assign n2862 = n10408 & n3620;
assign n12657 = n9742 | n13567;
assign n13167 = n10523 | n11296;
assign n582 = ~n4172;
assign n2515 = ~(n11990 | n14101);
assign n2572 = n3263 & n13334;
assign n490 = n10615 & n10843;
assign n12977 = n5582 & n1578;
assign n1513 = ~(n6085 | n7024);
assign n2271 = n5861 | n1318;
assign n12755 = n9745 & n5133;
assign n11521 = n11951 | n12733;
assign n7570 = n13547 | n1735;
assign n9820 = ~(n3395 | n11924);
assign n9539 = n11542 | n14125;
assign n9027 = n3161 | n7823;
assign n11433 = n7691 & n8898;
assign n8145 = n6243 & n3346;
assign n10705 = ~n10400;
assign n13118 = ~n13901;
assign n7262 = n13520 & n11918;
assign n11551 = ~n4847;
assign n3801 = n619 | n9866;
assign n4493 = n4932 & n9454;
assign n9754 = ~n461;
assign n12020 = ~n1010;
assign n2655 = n4631 | n12716;
assign n12605 = ~(n5278 | n5849);
assign n13 = n2908 | n6329;
assign n6525 = ~n1724;
assign n7285 = n2820 & n1141;
assign n4869 = n9111 | n1636;
assign n1448 = n9403 | n8336;
assign n1795 = n6531 & n4474;
assign n13288 = n5570 | n11003;
assign n14130 = ~(n11581 | n2543);
assign n8569 = ~n9592;
assign n14051 = n6157 & n11026;
assign n12274 = ~(n2415 | n6572);
assign n454 = ~(n3871 | n526);
assign n7274 = n3877 | n6922;
assign n59 = n8897 | n3754;
assign n10424 = n12039 & n5637;
assign n7540 = n13297 & n3495;
assign n989 = ~(n8065 | n10425);
assign n14302 = n12633 | n13622;
assign n8671 = ~(n5715 | n5989);
assign n11493 = ~n6326;
assign n7970 = ~n7278;
assign n5314 = n11313 & n9036;
assign n13332 = n5471 & n895;
assign n6137 = ~(n5435 | n6816);
assign n4963 = ~n4953;
assign n65 = n3485 & n5752;
assign n11813 = n4786 & n4859;
assign n438 = ~n12850;
assign n8576 = n9977 | n13890;
assign n12094 = n227 | n12863;
assign n5332 = n6318 & n4416;
assign n14237 = n9620 | n6280;
assign n5273 = n13276 | n5227;
assign n4760 = ~(n13722 | n2276);
assign n14004 = n8881 | n7326;
assign n2258 = n4525 & n11644;
assign n12418 = n13103 & n1890;
assign n8741 = n817 | n14085;
assign n9758 = n9490 | n2004;
assign n9747 = ~n81;
assign n3277 = ~n11765;
assign n1089 = n446 & n6663;
assign n11275 = ~(n6544 | n5663);
assign n401 = n9617 & n4746;
assign n8946 = n14110 | n8516;
assign n5026 = ~n11130;
assign n11877 = n12139 | n7280;
assign n9239 = ~(n1112 | n14390);
assign n8528 = ~n2201;
assign n423 = n9226 | n544;
assign n4695 = n7359 | n7129;
assign n14053 = n5732 | n11504;
assign n6974 = n3 & n2858;
assign n6287 = n13952 & n9368;
assign n4500 = n3675 & n4763;
assign n10576 = n11403 & n5316;
assign n3462 = ~(n6422 | n7313);
assign n12452 = n8747 | n11917;
assign n7579 = n7426 | n107;
assign n11634 = ~(n9388 | n1040);
assign n10832 = n2246 | n9499;
assign n11261 = n13991 | n6589;
assign n12130 = ~n8272;
assign n13134 = n8015 | n5440;
assign n11396 = n14166 | n13018;
assign n11630 = ~(n1112 | n7634);
assign n5861 = ~n13165;
assign n6947 = n11121 | n14073;
assign n7511 = n3268 & n10658;
assign n9869 = n13626 & n5838;
assign n4873 = n5011 & n8639;
assign n12483 = ~n746;
assign n10013 = n8786 & n1057;
assign n13350 = ~n11809;
assign n12562 = n2874 | n2182;
assign n4889 = ~(n7407 | n6327);
assign n3606 = n781 | n11922;
assign n10587 = n200 & n5420;
assign n11942 = n11329 & n10990;
assign n4221 = n80 & n6524;
assign n3493 = n7308 & n14229;
assign n2918 = n14118 & n736;
assign n7908 = n7717 & n6412;
assign n8142 = n7914 | n8761;
assign n14446 = ~n10322;
assign n4670 = n5569 | n5648;
assign n6043 = n3370 & n6208;
assign n4097 = n9285 | n7039;
assign n5806 = n7652 & n11206;
assign n6699 = n392 & n3701;
assign n8278 = n9403 | n5174;
assign n8882 = ~(n1152 | n1388);
assign n9687 = n9724 & n12031;
assign n11481 = ~n11967;
assign n4530 = n8096 | n7541;
assign n4996 = n6013 & n3420;
assign n777 = n11743 & n6794;
assign n2359 = n10072 & n2406;
assign n8644 = n6724 & n8653;
assign n1580 = n5012 & n12054;
assign n6413 = ~n10403;
assign n5694 = n7156 | n6719;
assign n8052 = n5779 & n7966;
assign n9364 = n77 | n7784;
assign n7556 = n4162 | n4998;
assign n11195 = n4365 & n6948;
assign n10368 = ~n834;
assign n902 = n3932 & n1484;
assign n4525 = ~n304;
assign n3092 = n7943 & n13453;
assign n739 = n5574 & n3214;
assign n4251 = n12039 & n7261;
assign n5228 = n636 | n3506;
assign n9801 = n14120 & n2131;
assign n3332 = ~n5288;
assign n9066 = ~(n7375 | n3170);
assign n3839 = n12764 | n3078;
assign n1875 = ~n630;
assign n534 = n904 & n3371;
assign n12786 = n4899 | n11058;
assign n2638 = n10933 | n5619;
assign n6899 = ~n2919;
assign n4024 = n2949 | n4042;
assign n1742 = ~n10115;
assign n13831 = n2017 | n7028;
assign n135 = n8045 | n10893;
assign n7679 = n5252 & n7724;
assign n6382 = n11739 | n13499;
assign n11096 = ~(n7245 | n13498);
assign n7833 = n4821 | n11388;
assign n2409 = ~n2566;
assign n4189 = n478 | n11695;
assign n12232 = n13102 & n2690;
assign n14398 = n9931 | n7815;
assign n5848 = ~n11515;
assign n1783 = n11153 & n9336;
assign n3340 = n6824 | n3835;
assign n499 = n3193 | n3792;
assign n9713 = n13005 | n860;
assign n7084 = n14370 | n11156;
assign n5857 = ~n1724;
assign n11522 = n13413 | n4186;
assign n13886 = n2518 | n14393;
assign n9737 = n13240 & n2565;
assign n13189 = n4346 & n12585;
assign n14189 = n69 | n6674;
assign n5522 = n1805 | n3849;
assign n11038 = n12986 & n7501;
assign n5518 = ~(n6413 | n13989);
assign n14059 = n11121 | n3806;
assign n2842 = n5253 | n5701;
assign n2405 = ~n5117;
assign n191 = n4359 & n5742;
assign n813 = n7284 & n2142;
assign n1266 = ~n13139;
assign n4107 = n10089 | n10635;
assign n1972 = n13016 | n13409;
assign n3740 = n12772 & n7465;
assign n12591 = ~(n2644 | n9714);
assign n11580 = ~n7339;
assign n8282 = n12250 & n10343;
assign n4641 = n13342 & n3202;
assign n12851 = n3 & n7549;
assign n9028 = n13626 & n11396;
assign n5418 = ~n12279;
assign n11764 = n12185 & n1888;
assign n2068 = n2874 | n10904;
assign n12739 = ~(n500 | n7725);
assign n11413 = n1875 | n10444;
assign n5401 = n8427 & n4423;
assign n9560 = ~(n3870 | n4793);
assign n9673 = ~n1702;
assign n8369 = n1699 & n6799;
assign n9797 = n13854 | n2275;
assign n3725 = n13745 & n8243;
assign n3017 = n12421 & n13521;
assign n1277 = ~(n2571 | n7953);
assign n1079 = n550 & n1307;
assign n10999 = n10245 | n2620;
assign n7142 = n11710 | n13460;
assign n6504 = n6891 | n13771;
assign n8665 = n2181 | n328;
assign n281 = n7057 & n1796;
assign n12498 = n6724 & n9725;
assign n5628 = ~n5427;
assign n6816 = ~(n13714 | n2524);
assign n3991 = ~(n7352 | n488);
assign n3700 = n11950 & n5691;
assign n6509 = n2846 & n11214;
assign n12917 = n13407 & n13834;
assign n6712 = ~(n9703 | n8796);
assign n11480 = n3607 & n11691;
assign n13129 = n8476 | n445;
assign n1857 = ~n8008;
assign n9209 = n2387 | n7599;
assign n6206 = ~n2794;
assign n6398 = n9403 | n3880;
assign n7597 = n5710 | n1905;
assign n1106 = ~(n2969 | n13681);
assign n8607 = ~n1334;
assign n10552 = n3867 | n700;
assign n6309 = n4445 & n5642;
assign n8789 = ~n7808;
assign n5061 = n2724 & n6779;
assign n5630 = n3861 & n5049;
assign n14212 = n12202 & n12818;
assign n10855 = ~n11474;
assign n1546 = ~(n162 | n7761);
assign n12089 = n14373 & n2653;
assign n7796 = n7527 | n1389;
assign n1045 = n8812 & n2012;
assign n5371 = n7745 & n7576;
assign n2672 = n9977 & n3970;
assign n14457 = n1147 | n11254;
assign n14119 = n5317 & n366;
assign n4962 = n4098 & n8820;
assign n9506 = ~(n12107 | n11928);
assign n14001 = n9080 & n1977;
assign n12825 = n11011 | n7685;
assign n11657 = n13860 & n4066;
assign n13192 = n9285 | n13439;
assign n4957 = n4346 & n5380;
assign n4005 = n8372 & n7178;
assign n4522 = n1223 | n12948;
assign n13942 = n7677 & n10381;
assign n1567 = n1414 & n5145;
assign n6484 = n2874 | n7719;
assign n2611 = n1059 & n8742;
assign n4003 = n5833 | n8369;
assign n2997 = n9920 & n240;
assign n9903 = n9953 & n214;
assign n10154 = ~n13901;
assign n416 = n679 | n13109;
assign n9854 = n7683 | n122;
assign n2555 = n541 & n4260;
assign n4446 = n5240 & n2;
assign n5722 = ~(n9618 | n8578);
assign n3247 = ~n12107;
assign n9344 = n12712 | n8802;
assign n5341 = n9232 & n4253;
assign n12370 = n13103 & n8442;
assign n1064 = ~(n1760 | n6997);
assign n6735 = n7327 & n8992;
assign n13450 = n1711 | n6839;
assign n9100 = n4657 & n1250;
assign n2966 = n8304 | n4405;
assign n3843 = n2055 | n6785;
assign n8060 = n2465 & n14386;
assign n1928 = n1520 & n4648;
assign n11801 = n6046 | n8848;
assign n11944 = n568 | n9201;
assign n7552 = n13433 & n2801;
assign n3245 = n13379 & n2162;
assign n13306 = ~(n4988 | n11634);
assign n1163 = n8828 | n9105;
assign n1561 = n7448 | n2923;
assign n10656 = n7596 & n3782;
assign n2098 = ~n12249;
assign n6323 = ~n4465;
assign n13534 = n14157 & n5698;
assign n549 = n2874 | n3010;
assign n12798 = n10857 | n2485;
assign n1413 = n4757 & n2730;
assign n13172 = n13863 & n13461;
assign n2477 = n7427 & n368;
assign n634 = n9716 | n2135;
assign n8390 = n5458 & n3562;
assign n4845 = n627 & n2685;
assign n8902 = ~(n11040 | n2530);
assign n14356 = n13096 & n311;
assign n335 = n12412 & n5758;
assign n13478 = n3710 & n12154;
assign n8822 = n9766 | n4039;
assign n7968 = n8769 & n10266;
assign n9177 = ~(n7359 | n6072);
assign n10098 = n12601 | n6417;
assign n9668 = ~(n1820 | n3920);
assign n2726 = ~(n8023 | n8360);
assign n12202 = ~n14524;
assign n13464 = ~n5795;
assign n4828 = ~n8595;
assign n13622 = n3424 & n11864;
assign n113 = n9269 | n10540;
assign n9306 = n12714 & n11444;
assign n2483 = ~(n11285 | n9553);
assign n4422 = ~n4618;
assign n3417 = n12147 & n867;
assign n5239 = n3635 & n3381;
assign n4049 = ~n11016;
assign n6948 = n6849 & n13857;
assign n11567 = n5603 | n10681;
assign n11177 = n12075 | n7548;
assign n2453 = n3126 | n5251;
assign n11498 = ~n12897;
assign n5348 = ~n5108;
assign n6202 = n7003 | n10692;
assign n1919 = n5876 & n12944;
assign n5637 = n3569 | n8619;
assign n13634 = n11048 | n517;
assign n9708 = n6695 | n6106;
assign n9981 = n6242 | n4089;
assign n4994 = n4803 & n6678;
assign n7772 = n14401 | n9796;
assign n801 = n5815 | n9290;
assign n12877 = n10678 & n8299;
assign n1249 = n2246 | n9889;
assign n9075 = n9529 | n8696;
assign n7830 = n2412 | n13502;
assign n13917 = n6595 | n6687;
assign n6777 = n7670 & n10277;
assign n2401 = ~n12588;
assign n5267 = n646 & n8502;
assign n14295 = n4898 | n13385;
assign n5131 = ~n5596;
assign n2230 = n6857 | n2403;
assign n9995 = n8358 & n6462;
assign n2368 = n8575 | n11491;
assign n7720 = ~n8672;
assign n13443 = ~(n10289 | n8368);
assign n7515 = n3088 | n10502;
assign n13916 = ~(n2132 | n7837);
assign n12456 = ~(n1820 | n5181);
assign n2623 = ~(n12934 | n3380);
assign n2154 = ~n2451;
assign n7787 = n8582 | n3624;
assign n9476 = n627 & n6181;
assign n13365 = ~n12014;
assign n13969 = n6838 & n6459;
assign n3794 = n234 | n5778;
assign n12354 = ~(n1423 | n5402);
assign n12180 = n6111 | n9152;
assign n8717 = n10622 & n1972;
assign n2767 = n9931 | n12439;
assign n2206 = n4498 | n5672;
assign n12824 = n7391 & n5559;
assign n6143 = n11739 | n12098;
assign n1026 = ~(n8217 | n4231);
assign n7006 = n12953 & n4429;
assign n8283 = n1414 & n6842;
assign n6592 = n1775 & n4596;
assign n8304 = ~n3455;
assign n3780 = n5940 & n1371;
assign n2348 = n1261 | n7785;
assign n11637 = n8034 | n1773;
assign n13899 = n14388 & n6097;
assign n4076 = n10062 | n9514;
assign n13852 = n3320 | n14132;
assign n10453 = n3011 | n8329;
assign n4472 = n2531 | n3714;
assign n2039 = n8404 | n6247;
assign n11984 = n4851 & n10847;
assign n2346 = n12695 | n8018;
assign n4876 = ~n12776;
assign n3262 = ~(n10511 | n7066);
assign n12084 = ~n4830;
assign n4773 = ~(n12483 | n9282);
assign n8135 = ~(n8629 | n334);
assign n13296 = n5092 & n2491;
assign n7792 = n3886 | n10183;
assign n8324 = ~(n239 | n12982);
assign n3708 = n12611 & n9313;
assign n1915 = n13226 | n12907;
assign n2256 = n10523 | n13472;
assign n944 = n6607 | n4215;
assign n13845 = n5493 | n282;
assign n7702 = ~(n6883 | n5827);
assign n633 = n9780 | n5895;
assign n3127 = n2747 | n9387;
assign n2494 = n11422 & n8533;
assign n7472 = n12404 & n10536;
assign n13147 = ~n6787;
assign n13790 = n783 & n13134;
assign n9643 = n11313 & n4179;
assign n7230 = ~n8439;
assign n5110 = n9509 & n3529;
assign n13880 = n3710 & n5106;
assign n9354 = n3776 & n10276;
assign n9019 = ~(n14466 | n3467);
assign n14384 = ~(n9305 | n9634);
assign n11859 = n11803 & n4120;
assign n8589 = n2272 | n10105;
assign n5334 = n329 | n4343;
assign n12049 = n14430 | n1335;
assign n12021 = ~(n10638 | n14517);
assign n12469 = n6373 | n4538;
assign n7608 = ~(n5833 | n12525);
assign n6392 = n231 & n13110;
assign n11490 = n7938 & n7838;
assign n504 = ~n8595;
assign n3917 = n7245 | n8867;
assign n10489 = n9507 | n1606;
assign n5743 = n3565 & n2740;
assign n3667 = ~n5974;
assign n9914 = n7063 & n6077;
assign n4371 = n7551 | n6050;
assign n4808 = ~(n9388 | n9685);
assign n8678 = n12615 & n2560;
assign n9256 = n6606 & n5122;
assign n13385 = n13597 & n5684;
assign n11949 = n12960 & n10295;
assign n14383 = n2181 | n4900;
assign n2601 = n8877 | n9672;
assign n2479 = n2583 & n2982;
assign n4631 = ~n3616;
assign n8470 = n8210 | n4160;
assign n12175 = n3366 & n2871;
assign n7871 = n7484 | n6251;
assign n1623 = ~n13696;
assign n14256 = n492 | n7880;
assign n8336 = n8789 & n8036;
assign n4010 = n1701 | n4668;
assign n2841 = n1031 | n3501;
assign n8875 = n4163 & n9912;
assign n5837 = n2111 | n11616;
assign n6180 = n8066 & n3739;
assign n7789 = n10595 & n8296;
assign n14193 = n14042 & n583;
assign n8833 = n4925 | n623;
assign n10055 = n7938 & n1062;
assign n802 = n14388 & n5260;
assign n1384 = n8238 & n8985;
assign n10530 = n8151 | n12053;
assign n5389 = n116 | n3041;
assign n9051 = n3097 & n8251;
assign n12525 = ~(n3907 | n9969);
assign n14062 = n11105 | n9006;
assign n1385 = ~(n7575 | n9637);
assign n13184 = n5472 | n6832;
assign n9417 = n14446 & n819;
assign n6622 = ~(n3344 | n5894);
assign n4344 = ~(n7609 | n9373);
assign n2315 = ~n2918;
assign n4135 = ~n6534;
assign n11615 = n10933 | n4957;
assign n6082 = n536 & n1114;
assign n8433 = n3586 & n10453;
assign n1196 = ~(n2103 | n6439);
assign n212 = n6157 & n1648;
assign n4204 = n3815 | n4540;
assign n6321 = n1805 | n2911;
assign n5494 = n4508 | n6351;
assign n3771 = ~(n12112 | n10122);
assign n8895 = ~(n10309 | n13640);
assign n3232 = n638 & n7856;
assign n4718 = ~(n10363 | n10814);
assign n10007 = n4788 & n12499;
assign n11897 = n10626 | n10644;
assign n659 = n4433 | n1222;
assign n1825 = n5229 & n1479;
assign n7978 = n11329 & n8912;
assign n5492 = n8172 | n6653;
assign n13857 = n8721 | n6680;
assign n13325 = ~(n9806 | n2036);
assign n5296 = n8096 | n2384;
assign n1506 = n14273 | n8926;
assign n5086 = n504 | n9891;
assign n13381 = n9015 & n270;
assign n10808 = ~n8148;
assign n11589 = n11803 & n3935;
assign n5324 = ~(n4741 | n1274);
assign n5406 = ~n4609;
assign n14389 = n9890 & n2205;
assign n11228 = n14435 | n8321;
assign n4047 = n14178 | n498;
assign n4125 = n427 & n3104;
assign n3592 = n1729 & n2211;
assign n9275 = ~n5153;
assign n13175 = n283 | n2671;
assign n1409 = ~n5960;
assign n63 = n5975 | n4022;
assign n1949 = n7427 & n8690;
assign n1931 = n7970 & n9633;
assign n7009 = n748 & n7292;
assign n14381 = n14120 & n12482;
assign n4275 = n5575 | n12512;
assign n8349 = n848 & n12992;
assign n2520 = n3608 & n12932;
assign n10774 = ~(n13276 | n9907);
assign n6714 = n12357 & n4687;
assign n446 = ~n6119;
assign n6724 = ~n9994;
assign n5153 = ~n8224;
assign n257 = n14400 | n8164;
assign n6852 = n10083 | n959;
assign n10825 = ~n3284;
assign n2988 = ~(n2919 | n537);
assign n14474 = n4932 & n915;
assign n11304 = n1074 & n11356;
assign n11233 = ~(n10936 | n14250);
assign n4393 = n12130 | n8978;
assign n3783 = n12023 | n2336;
assign n7933 = n3120 | n12619;
assign n5934 = n7267 & n9487;
assign n7518 = ~n6397;
assign n13870 = n7972 & n8374;
assign n12714 = n12435 | n411;
assign n2446 = ~(n473 | n2186);
assign n6254 = ~n11259;
assign n4352 = n11379 | n8227;
assign n3632 = n5104 & n9011;
assign n1375 = ~(n1697 | n1652);
assign n10004 = n8964 | n8198;
assign n3760 = n11262 & n11885;
assign n11155 = ~(n12084 | n10203);
assign n14104 = ~(n8223 | n13584);
assign n3496 = n4655 & n6992;
assign n2847 = n10834 | n10102;
assign n14185 = n6323 | n7853;
assign n11667 = ~n3623;
assign n12737 = n573 | n12879;
assign n12377 = n1480 | n8084;
assign n197 = n12425 & n12247;
assign n8986 = ~n777;
assign n8993 = n1788 & n1380;
assign n12975 = n7041 & n10483;
assign n12594 = n13484 & n661;
assign n6142 = n11459 | n10272;
assign n6660 = ~n7889;
assign n8925 = ~n11232;
assign n8318 = n7691 & n7651;
assign n12589 = n4856 & n10984;
assign n9108 = n9953 & n4832;
assign n7524 = ~(n3445 | n13104);
assign n684 = n4481 | n1240;
assign n2809 = n6130 & n14202;
assign n2057 = ~n9371;
assign n10281 = n5625 | n12745;
assign n12794 = n8210 | n1766;
assign n14524 = ~n3331;
assign n526 = ~(n3196 | n7663);
assign n6159 = ~n6088;
assign n14363 = n13516 | n3868;
assign n249 = n3607 & n7215;
assign n2756 = n7026 & n6809;
assign n5840 = ~n10465;
assign n3156 = ~(n10363 | n4693);
assign n4042 = n6507 & n6276;
assign n8298 = ~(n7605 | n11407);
assign n6839 = n8250 & n4688;
assign n2915 = n4898 | n5842;
assign n13219 = ~n1984;
assign n10662 = n8513 | n8979;
assign n10541 = n13252 & n11301;
assign n6498 = ~n8746;
assign n5870 = n11438 | n10418;
assign n6425 = n8476 | n1866;
assign n6276 = n6263 | n10608;
assign n1244 = n7003 | n6541;
assign n2713 = n4828 | n7183;
assign n4426 = n13078 & n12328;
assign n8927 = n815 & n9022;
assign n6259 = n3132 | n4927;
assign n1173 = n9315 & n8736;
assign n1446 = n5450 | n6105;
assign n8010 = n8786 & n5465;
assign n4688 = n13005 | n901;
assign n913 = n9174 | n7860;
assign n9375 = ~n4550;
assign n9735 = n9811 & n7463;
assign n7746 = ~(n12999 | n11678);
assign n3840 = n11647 | n13405;
assign n1487 = n406 & n11159;
assign n8034 = ~n7322;
assign n8724 = n13413 | n9108;
assign n11717 = n10825 | n11768;
assign n20 = n11739 | n260;
assign n5937 = ~(n3907 | n2352);
assign n6018 = ~n5001;
assign n174 = n9529 | n2328;
assign n391 = n2983 & n10320;
assign n11781 = n2533 & n4980;
assign n1639 = ~n10172;
assign n14011 = ~n10485;
assign n4208 = n6111 | n2152;
assign n14063 = ~n2958;
assign n13445 = n7852 & n8613;
assign n12072 = n3565 & n11216;
assign n2580 = n1452 & n1786;
assign n3206 = n412 | n5105;
assign n3618 = n13108 | n8499;
assign n2185 = ~(n12075 | n12739);
assign n5463 = n228 | n6164;
assign n6305 = n10512 & n9611;
assign n3298 = n9229 | n11684;
assign n3359 = ~(n4913 | n4629);
assign n14504 = n7961 & n10142;
assign n13367 = ~n3361;
assign n3243 = n3512 | n7770;
assign n2367 = ~n10377;
assign n2652 = n8714 | n10521;
assign n5215 = n2533 & n12186;
assign n12774 = n12295 | n8022;
assign n8910 = n2177 & n1139;
assign n4330 = ~(n11498 | n14485);
assign n12041 = n14227 & n11429;
assign n853 = n100 | n1333;
assign n6926 = n10668 & n12182;
assign n9933 = n3932 & n2072;
assign n13230 = n10231 | n11902;
assign n11714 = n5033 | n4172;
assign n8506 = n820 | n10005;
assign n13268 = n5977 | n8952;
assign n1121 = ~(n13213 | n13097);
assign n11850 = n7684 | n13911;
assign n11830 = n12131 | n6187;
assign n10729 = n12100 | n3829;
assign n10275 = n10624 | n5939;
assign n1812 = ~n6058;
assign n13104 = ~(n4624 | n8352);
assign n207 = n10134 & n6100;
assign n1292 = n5570 | n9118;
assign n3440 = ~n10380;
assign n6836 = n333 & n8384;
assign n1887 = n6649 & n3310;
assign n13618 = n6857 | n8497;
assign n6835 = n9015 & n8159;
assign n8928 = n1356 | n9141;
assign n2285 = n3932 & n4972;
assign n9945 = n8582 | n7154;
assign n6804 = n7929 & n11113;
assign n13495 = n8789 & n4107;
assign n8494 = n7677 & n11166;
assign n7585 = n1741 | n11039;
assign n13358 = ~(n3003 | n6404);
assign n7942 = n5104 & n11249;
assign n14227 = ~n11668;
assign n8357 = n10310 & n6546;
assign n7654 = n12543 | n1418;
assign n9700 = ~(n4633 | n5748);
assign n11097 = ~n13234;
assign n5652 = n4340 | n5147;
assign n10497 = n4267 | n10407;
assign n3321 = ~(n13310 | n1552);
assign n146 = n5899 & n5854;
assign n14290 = ~(n6387 | n4831);
assign n6813 = ~(n10400 | n11439);
assign n13663 = n1669 | n5704;
assign n14392 = n9726 & n10579;
assign n5610 = n8427 & n4559;
assign n4806 = ~n13447;
assign n14444 = n1255 & n3729;
assign n12086 = ~n4270;
assign n8896 = n11231 | n5942;
assign n3238 = n478 | n11848;
assign n14091 = ~n1495;
assign n3719 = ~(n3876 | n9365);
assign n3912 = ~(n7739 | n10848);
assign n11612 = n2949 | n12033;
assign n3887 = n10330 & n530;
assign n13551 = ~(n8701 | n8334);
assign n1075 = n12990 & n1192;
assign n10394 = ~n4465;
assign n4309 = ~(n1686 | n8733);
assign n6612 = n11220 & n3641;
assign n3072 = n2877 | n12113;
assign n311 = n10624 | n6920;
assign n226 = n5252 & n8428;
assign n7151 = n1223 | n2381;
assign n5939 = n8697 & n3748;
assign n1427 = ~n7346;
assign n3884 = n9931 | n11817;
assign n10232 = n8907 | n4895;
assign n4416 = n2086 | n12612;
assign n1159 = ~(n4924 | n8860);
assign n10315 = n13130 | n9158;
assign n4128 = ~n3046;
assign n3059 = n13641 & n8871;
assign n13078 = ~n13038;
assign n6371 = n1427 & n7044;
assign n6024 = n10808 | n9009;
assign n9349 = n13016 | n5319;
assign n3734 = ~(n6209 | n6755);
assign n10907 = ~(n5977 | n3642);
assign n9518 = n6046 | n10892;
assign n163 = ~n12874;
assign n13874 = ~n6903;
assign n3453 = n12404 & n130;
assign n14175 = n8043 & n10274;
assign n6583 = ~(n3394 | n10597);
assign n8930 = n12015 & n12266;
assign n13545 = n12445 & n963;
assign n9270 = n6849 | n3804;
assign n13194 = ~n3367;
assign n8616 = n10713 | n8719;
assign n7109 = ~(n4313 | n6751);
assign n7606 = ~(n4897 | n12955);
assign n13105 = n1138 & n9669;
assign n11266 = n11020 & n10026;
assign n11827 = n9289 | n3131;
assign n14262 = n390 | n9431;
assign n13771 = n10556 & n4323;
assign n6030 = ~n10406;
assign n9576 = n2820 & n11203;
assign n1246 = ~(n3333 | n10257);
assign n5127 = n12357 | n666;
assign n8317 = n5012 & n2015;
assign n5496 = n10825 | n4297;
assign n5788 = n7216 | n14293;
assign n10536 = n7212 | n4157;
assign n5989 = ~(n4417 | n2561);
assign n3501 = n10330 & n9622;
assign n100 = ~n9453;
assign n10776 = ~(n12644 | n9963);
assign n8274 = n11722 | n10212;
assign n6418 = n8817 & n13862;
assign n5017 = n13130 | n14098;
assign n1852 = ~(n6731 | n3355);
assign n9095 = n6111 | n767;
assign n4484 = ~n760;
assign n10513 = n12542 & n10221;
assign n9752 = n12401 | n6942;
assign n7738 = n7053 & n11567;
assign n8316 = n13432 | n1069;
assign n4531 = n14319 | n6496;
assign n10009 = n11405 | n10901;
assign n5616 = n2709 & n11868;
assign n5809 = n5491 | n7917;
assign n14403 = n2016 | n8732;
assign n13887 = n7212 | n2536;
assign n9119 = ~n5184;
assign n3523 = ~n11227;
assign n2156 = n2521 & n6257;
assign n10888 = n9571 & n3756;
assign n12316 = ~(n4549 | n11751);
assign n13388 = n12353 | n2913;
assign n13879 = n3025 | n3551;
assign n7743 = n11105 | n6858;
assign n4749 = n4988 | n8885;
assign n9829 = n560 | n8486;
assign n5005 = ~(n163 | n2446);
assign n6773 = n1172 | n3830;
assign n9295 = ~(n5990 | n14168);
assign n5345 = n9191 & n7217;
assign n8178 = ~(n5042 | n9639);
assign n13414 = ~(n12522 | n2199);
assign n10114 = ~(n13937 | n5810);
assign n506 = ~n11412;
assign n7714 = ~(n4342 | n987);
assign n4974 = ~(n7362 | n2380);
assign n6570 = n11576 | n10927;
assign n3241 = n10534 | n3084;
assign n12125 = n12730 & n13454;
assign n3048 = n12039 & n8666;
assign n8756 = n11163 & n12146;
assign n10501 = n5053 & n9623;
assign n11240 = ~n8424;
assign n9121 = n4739 | n8009;
assign n2042 = n8045 | n6371;
assign n8862 = n5266 | n3256;
assign n7717 = ~n1742;
assign n6987 = n7429 & n2232;
assign n13569 = ~(n1623 | n6841);
assign n12656 = n4856 & n12645;
assign n13041 = ~n7920;
assign n4610 = ~(n12872 | n10495);
assign n14144 = n3815 | n7168;
assign n11200 = n6606 & n3119;
assign n9402 = n10595 & n8403;
assign n11100 = n14039 | n6791;
assign n13155 = ~n6264;
assign n10401 = ~(n1458 | n10746);
assign n7878 = n6471 | n12457;
assign n7870 = n678 & n14495;
assign n8419 = n203 | n5184;
assign n9150 = ~(n7418 | n9396);
assign n12474 = n6531 & n559;
assign n8258 = n1452 & n10666;
assign n5261 = n6744 & n10438;
assign n2511 = n1538 | n13444;
assign n8962 = n1582 | n12195;
assign n11809 = ~n4296;
assign n11142 = ~n11861;
assign n933 = ~(n8301 | n6515);
assign n9832 = n6629 | n10419;
assign n1871 = n10930 & n9992;
assign n5774 = n4840 | n7598;
assign n5322 = n14401 | n8508;
assign n4797 = ~(n1685 | n13530);
assign n6682 = n3506 & n1758;
assign n13150 = n13854 | n9547;
assign n12723 = n3062 | n5633;
assign n4844 = ~n2692;
assign n12306 = n4092 | n8872;
assign n1181 = n13130 | n5688;
assign n6624 = n10458 & n4130;
assign n10137 = n13359 & n246;
assign n723 = n6909 & n7816;
assign n13331 = n4722 & n2049;
assign n9729 = n974 | n11883;
assign n4391 = n1414 & n11904;
assign n13077 = n6596 | n13554;
assign n908 = n8789 & n13372;
assign n6390 = n8581 | n9989;
assign n4339 = n11459 | n8083;
assign n4098 = ~n304;
assign n4029 = n11950 & n13818;
assign n523 = ~n12776;
assign n3080 = n3164 | n10835;
assign n129 = ~n742;
assign n9896 = n7527 | n13906;
assign n10788 = n12712 | n431;
assign n10994 = n5226 | n13625;
assign n4547 = ~(n1623 | n10133);
assign n9036 = n1535 | n8434;
assign n12952 = n3785 & n305;
assign n8816 = ~n7600;
assign n1060 = n4341 & n6319;
assign n4900 = n6316 & n3049;
assign n9805 = n6527 & n7479;
assign n12519 = n6706 | n631;
assign n4903 = n129 & n9815;
assign n10120 = n4199 | n336;
assign n1965 = n1840 | n4958;
assign n9585 = n9078 | n9727;
assign n7691 = ~n5182;
assign n3163 = n10457 & n8225;
assign n7940 = ~n11401;
assign n1533 = n3097 & n2629;
assign n7537 = n647 | n3244;
assign n14016 = n2012 | n6810;
assign n2383 = n4373 & n6941;
assign n13007 = n14109 & n13919;
assign n12529 = n954 | n11141;
assign n8650 = ~n5257;
assign n8069 = n12351 | n4699;
assign n144 = n6350 | n8519;
assign n14180 = n9069 & n2992;
assign n292 = n3672 & n12163;
assign n8180 = ~(n9423 | n2726);
assign n138 = n10457 & n3902;
assign n3248 = ~n6806;
assign n3394 = ~n13234;
assign n3375 = n14472 | n8155;
assign n14239 = ~n14510;
assign n12593 = ~n9550;
assign n13540 = n11495 & n13976;
assign n13903 = n11438 | n6370;
assign n13864 = n14110 | n1300;
assign n13708 = n5628 & n9884;
assign n13260 = ~(n12934 | n681);
assign n5306 = ~n14367;
assign n10985 = n1908 & n8750;
assign n1296 = n2318 | n12474;
assign n13031 = n10015 & n9349;
assign n194 = ~n3357;
assign n6486 = ~n1120;
assign n8804 = n7364 | n4781;
assign n2925 = ~n13944;
assign n10805 = n7003 | n10613;
assign n7298 = n2055 | n9443;
assign n6603 = n11776 | n6873;
assign n13444 = n7060 & n13864;
assign n5041 = ~(n163 | n1126);
assign n2188 = ~n9186;
assign n13345 = n10595 & n11830;
assign n5664 = n13035 | n9186;
assign n13844 = ~(n6434 | n5400);
assign n13700 = ~n6819;
assign n10087 = n5475 & n12811;
assign n3353 = n13147 & n5002;
assign n5499 = n2486 & n8071;
assign n10652 = n2564 & n1761;
assign n3325 = ~(n1686 | n3658);
assign n5089 = n10808 | n2636;
assign n5846 = n12633 | n10693;
assign n13004 = n13537 | n5730;
assign n3742 = ~n12522;
assign n288 = n501 & n14128;
assign n11516 = n10035 | n4911;
assign n14209 = n6654 | n5191;
assign n426 = n5668 & n7546;
assign n12101 = ~n7902;
assign n5222 = n2758 & n13247;
assign n252 = n9429 | n5744;
assign n5075 = ~(n1028 | n1553);
assign n7867 = n5007 | n5803;
assign n13185 = n10300 | n14225;
assign n845 = n12414 | n9939;
assign n10183 = n327 & n14458;
assign n1 = n2843 | n12864;
assign n8845 = n5062 & n262;
assign n10361 = n6130 & n9121;
assign n4401 = n1247 & n11339;
assign n7135 = n13547 | n6461;
assign n5613 = ~n7258;
assign n8441 = ~(n2919 | n10782);
assign n4050 = ~n7931;
assign n10811 = ~(n7551 | n1338);
assign n66 = ~(n8887 | n9317);
assign n10182 = n5940 & n5774;
assign n11855 = n8213 & n7639;
assign n676 = n9275 & n9575;
assign n1419 = n1628 | n8099;
assign n2026 = n5876 & n13113;
assign n2027 = n4615 & n13980;
assign n3969 = n13240 & n5721;
assign n10409 = n5084 | n6014;
assign n13825 = n387 | n8409;
assign n7351 = n523 | n7747;
assign n9772 = n2998 & n10301;
assign n6135 = ~n7621;
assign n6249 = n5891 | n9741;
assign n2311 = n3804 & n7757;
assign n6577 = n5348 & n8364;
assign n13734 = ~n11347;
assign n9078 = ~n4149;
assign n6387 = n3833 | n6436;
assign n2605 = n5144 | n12007;
assign n11300 = ~n12697;
assign n8739 = n7717 & n7665;
assign n2882 = n10035 | n7480;
assign n12217 = n10855 & n10348;
assign n1178 = ~n11324;
assign n4017 = n4562 | n2319;
assign n5094 = n820 | n7379;
assign n2249 = n11223 | n3712;
assign n8911 = n14337 | n6805;
assign n7531 = n4844 & n10978;
assign n13039 = n12844 | n10501;
assign n3228 = n930 | n13914;
assign n9269 = ~n1010;
assign n11104 = n7156 | n2071;
assign n3569 = ~n8272;
assign n10249 = n8096 | n1381;
assign n4754 = n5641 | n8554;
assign n6136 = n3667 | n1753;
assign n6388 = ~n8635;
assign n7747 = n6830 & n408;
assign n8914 = n13516 | n5511;
assign n9065 = ~(n9871 | n13566);
assign n7635 = n4908 | n3548;
assign n9653 = ~(n3905 | n1733);
assign n6316 = ~n3926;
assign n11213 = ~n6426;
assign n12772 = ~n5944;
assign n5231 = n12615 & n6178;
assign n12095 = n648 | n6401;
assign n12117 = n7282 | n13944;
assign n938 = n9230 | n10150;
assign n11089 = n12721 & n6140;
assign n9963 = n13236 & n11573;
assign n461 = n1203 | n10426;
assign n2521 = ~n6193;
assign n9980 = n678 & n13285;
assign n12973 = n12449 & n8031;
assign n11429 = n647 | n8683;
assign n9292 = n13362 & n12540;
assign n2727 = ~n9041;
assign n195 = n9188 & n7304;
assign n4023 = n7700 | n8136;
assign n6556 = ~n9555;
assign n13286 = n8431 & n12148;
assign n6466 = n13364 | n2061;
assign n2305 = n3276 & n1901;
assign n13285 = n9111 | n13678;
assign n173 = n5861 | n4709;
assign n3913 = n10678 & n14329;
assign n2592 = n3193 | n9500;
assign n12866 = ~n8822;
assign n2160 = n3672 & n6669;
assign n2790 = ~n14354;
assign n11244 = n13194 | n9543;
assign n5058 = ~(n11285 | n1403);
assign n5519 = n12105 & n10981;
assign n13475 = n5266 | n3691;
assign n10533 = n6730 | n9627;
assign n3084 = n7081 & n1891;
assign n6156 = n185 | n4783;
assign n10636 = n14351 & n9057;
assign n12234 = n11737 & n12984;
assign n13686 = n387 | n7587;
assign n12811 = n7426 | n12752;
assign n13270 = ~n4561;
assign n8989 = n8386 & n3791;
assign n7259 = n11020 & n9974;
assign n8126 = ~(n12765 | n12388);
assign n7424 = n2310 & n11358;
assign n3623 = n13132 | n5960;
assign n5211 = n4828 | n4779;
assign n64 = n1678 & n12971;
assign n10389 = n49 | n8176;
assign n4827 = n8897 | n14191;
assign n570 = n10247 & n3080;
assign n3349 = n13362 & n9327;
assign n6514 = n11440 | n6910;
assign n11091 = n4407 | n5261;
assign n9626 = n839 | n10947;
assign n9016 = n2021 & n10493;
assign n1293 = ~(n13154 | n3716);
assign n9900 = n12404 & n1483;
assign n13040 = n225 & n2599;
assign n13713 = n8575 | n10468;
assign n1324 = n9323 & n10161;
assign n8611 = n8950 & n1285;
assign n42 = n3268 & n1873;
assign n5808 = n3871 | n6782;
assign n6806 = n11824 & n1447;
assign n10129 = n6606 & n6648;
assign n2099 = ~n8008;
assign n11618 = n12475 & n9802;
assign n13987 = n9726 & n8542;
assign n13557 = ~n670;
assign n8202 = n2877 | n13212;
assign n10902 = n14109 & n2945;
assign n4726 = n1711 | n2382;
assign n11700 = n14400 | n14261;
assign n14075 = ~n4324;
assign n8447 = n200 & n5775;
assign n11188 = n3364 | n6007;
assign n1223 = ~n1676;
assign n4207 = ~n2130;
assign n4210 = ~n8809;
assign n5096 = n9442 | n5765;
assign n11845 = n3320 | n13529;
assign n12576 = ~n11415;
assign n472 = n13379 & n7240;
assign n9661 = n3276 & n8623;
assign n8277 = ~n14412;
assign n13974 = n7462 | n914;
assign n8755 = n12185 & n7591;
assign n3019 = ~n6196;
assign n2259 = n1147 | n10557;
assign n360 = ~(n12107 | n11745);
assign n2766 = ~n5668;
assign n11377 = n9890 & n14056;
assign n11556 = n8692 & n11629;
assign n14013 = n14088 | n9241;
assign n8722 = n13485 | n5598;
assign n1585 = n11950 & n9449;
assign n12220 = ~(n14106 | n11050);
assign n9809 = n9705 & n1448;
assign n1080 = n6690 | n5538;
assign n6173 = n7888 | n5423;
assign n73 = n1697 | n5371;
assign n5158 = n4162 | n9254;
assign n9385 = n10566 & n11880;
assign n7392 = ~n300;
assign n23 = n3826 | n10851;
assign n2135 = n432 & n4020;
assign n1736 = n2281 & n10786;
assign n10028 = n7691 & n5996;
assign n374 = ~(n7229 | n9380);
assign n12823 = ~n736;
assign n10715 = ~n13779;
assign n9597 = n10731 | n11943;
assign n5308 = n1662 & n14176;
assign n2960 = n4255 | n11099;
assign n1317 = n10534 | n662;
assign n6112 = n2761 | n12938;
assign n3871 = ~n4891;
assign n13617 = n2645 | n7147;
assign n10384 = n1920 | n7104;
assign n11888 = n3097 & n3318;
assign n11787 = n13130 | n253;
assign n1049 = n13338 & n6328;
assign n11662 = ~(n8404 | n75);
assign n3324 = n11688 & n6268;
assign n24 = n9705 & n1442;
assign n895 = n7227 | n12605;
assign n2569 = n1428 & n12981;
assign n369 = n2179 | n2725;
assign n7961 = ~n7808;
assign n840 = n10461 | n6310;
assign n657 = n1820 | n10020;
assign n3625 = n9541 | n90;
assign n8279 = n1266 & n7118;
assign n14141 = n8386 & n11478;
assign n11270 = n8232 & n6681;
assign n10246 = n11223 | n14356;
assign n11989 = n11303 | n13749;
assign n4259 = ~(n12568 | n1524);
assign n11599 = n6192 & n12050;
assign n8226 = n12414 | n319;
assign n10515 = n4154 & n1180;
assign n6620 = n7358 | n1018;
assign n4035 = ~(n11761 | n1297);
assign n10436 = n4347 & n12671;
assign n12419 = n12428 | n5356;
assign n3914 = ~n1214;
assign n2473 = ~n10803;
assign n910 = n1875 | n11092;
assign n14285 = ~(n13350 | n8729);
assign n7178 = n8458 | n7233;
assign n6957 = ~n6139;
assign n10078 = n5628 & n8831;
assign n12997 = n2888 | n2855;
assign n9400 = ~(n8277 | n5396);
assign n4040 = n8238 & n2290;
assign n1272 = n13781 & n7447;
assign n11373 = n13108 | n2859;
assign n6886 = n11176 | n6698;
assign n13123 = n9429 | n539;
assign n3703 = n10399 & n4370;
assign n9610 = n1914 | n2950;
assign n10635 = n14145 & n5258;
assign n14055 = n14446 & n12777;
assign n1940 = n11576 | n6445;
assign n5498 = n6039 | n3733;
assign n3331 = n10619 & n4419;
assign n14136 = ~(n5418 | n6643);
assign n12078 = n6323 | n10397;
assign n5196 = n13867 & n4515;
assign n13556 = n6525 & n716;
assign n175 = n9507 | n11931;
assign n13964 = ~(n1838 | n4363);
assign n8525 = n4481 | n3980;
assign n13156 = n8881 | n13253;
assign n12567 = n11105 | n2243;
assign n10894 = n873 & n10561;
assign n6883 = ~n3094;
assign n6581 = n14466 | n13221;
assign n3414 = ~(n7551 | n299);
assign n10457 = ~n7802;
assign n5057 = ~(n882 | n12198);
assign n12514 = n7673 & n10798;
assign n6635 = n361 | n289;
assign n9683 = ~(n10121 | n12755);
assign n8855 = ~n13190;
assign n10743 = n9275 & n12068;
assign n5591 = ~n10278;
assign n10827 = n9507 | n2100;
assign n3396 = n1198 | n2190;
assign n6993 = n13338 & n9054;
assign n12867 = n3405 & n4530;
assign n2894 = n89 | n5162;
assign n5326 = n10705 & n3138;
assign n8245 = n9078 | n12507;
assign n3863 = ~(n12568 | n3779);
assign n9045 = n7911 & n3096;
assign n10282 = n7502 | n6758;
assign n14330 = n5725 & n2856;
assign n2134 = n7691 & n13517;
assign n11118 = n1044 | n604;
assign n6243 = ~n2566;
assign n7210 = ~(n11633 | n13207);
assign n5397 = n9218 | n7134;
assign n685 = ~(n8959 | n7865);
assign n3535 = n9745 & n5072;
assign n10752 = n10710 & n10886;
assign n6807 = ~n11441;
assign n14236 = ~(n5569 | n3338);
assign n9574 = n12994 | n2831;
assign n11235 = n3565 & n1279;
assign n3308 = ~(n1023 | n13471);
assign n9052 = ~n1086;
assign n13816 = ~(n8458 | n5170);
assign n3891 = n5180 | n8402;
assign n13991 = ~n11813;
assign n10640 = n1613 | n714;
assign n4060 = n13850 & n12156;
assign n3112 = n1112 | n7928;
assign n13001 = n11142 & n11717;
assign n11458 = n11315 | n14507;
assign n7350 = n3888 | n6511;
assign n13546 = n11403 & n2630;
assign n9410 = n7826 & n13746;
assign n2751 = n4422 & n6291;
assign n1061 = ~n9959;
assign n1530 = ~(n8209 | n9631);
assign n6792 = n12844 | n3862;
assign n9114 = n8404 | n3502;
assign n839 = ~n2794;
assign n13528 = ~(n7227 | n4636);
assign n9147 = ~(n1548 | n2193);
assign n10901 = n200 & n4360;
assign n12793 = n12764 | n14306;
assign n7252 = ~(n3418 | n3033);
assign n11441 = n9245 & n356;
assign n1082 = n2330 & n724;
assign n12564 = n2587 & n10639;
assign n1859 = ~(n12193 | n4366);
assign n1416 = n4207 | n1309;
assign n5600 = n8769 & n12478;
assign n185 = ~n4149;
assign n14049 = n7862 | n4400;
assign n2989 = n5641 | n5280;
assign n485 = n14446 & n6692;
assign n7528 = n14472 | n3362;
assign n6953 = ~n1312;
assign n4564 = n13650 | n8044;
assign n6964 = ~(n14166 | n6221);
assign n12595 = n12549 | n7896;
assign n1421 = n3820 | n674;
assign n3834 = n9650 & n13430;
assign n3063 = n11093 & n1537;
assign n10861 = n2760 & n2717;
assign n3230 = n6680 | n3804;
assign n11898 = ~(n5468 | n3774);
assign n14519 = n850 | n8092;
assign n13876 = n8183 & n12950;
assign n9625 = n13555 & n13229;
assign n10302 = ~n1120;
assign n2168 = n14319 | n8770;
assign n5391 = ~n2369;
assign n13603 = ~(n10620 | n8443);
assign n1524 = ~(n13072 | n12433);
assign n4104 = ~n6397;
assign n1097 = n492 | n6955;
assign n4240 = n904 & n8819;
assign n3266 = n55 & n1555;
assign n4150 = n10300 | n1601;
assign n8853 = n12389 & n10004;
assign n3294 = n9265 & n6299;
assign n13176 = n3923 & n4319;
assign n4338 = n3768 | n1897;
assign n1068 = n7364 | n4611;
assign n7042 = n2820 & n10500;
assign n3391 = n1857 & n2621;
assign n6370 = n2322 & n3825;
assign n13141 = n4147 & n14096;
assign n8876 = ~(n393 | n10880);
assign n13747 = n3025 | n5101;
assign n372 = n13446 | n8708;
assign n7676 = n8655 | n11143;
assign n7367 = n13885 | n786;
assign n4526 = n1061 | n2907;
assign n11767 = ~(n5172 | n6290);
assign n3449 = ~n11902;
assign n3748 = n8828 | n7394;
assign n6767 = n11176 | n10193;
assign n11602 = n7427 & n12798;
assign n3128 = n8242 | n6762;
assign n1688 = n9824 & n1477;
assign n12617 = n1140 & n435;
assign n7775 = ~(n2171 | n2396);
assign n5581 = n11607 & n218;
assign n301 = n480 | n7906;
assign n9274 = n550 | n9544;
assign n5745 = n3877 | n1009;
assign n13101 = n11153 & n5935;
assign n4122 = n7284 & n12227;
assign n2715 = n11816 & n2933;
assign n3739 = n8096 | n2184;
assign n12580 = ~n5990;
assign n3820 = ~n3910;
assign n5490 = n6527 & n2079;
assign n4770 = n6271 | n17;
assign n10792 = n6753 & n13491;
assign n6908 = n568 | n11991;
assign n2103 = ~n7929;
assign n10157 = n5574 & n5228;
assign n6602 = n3743 & n7097;
assign n11289 = n10854 & n8990;
assign n3639 = ~(n478 | n2707);
assign n5015 = ~(n14332 | n13826);
assign n2293 = n13413 | n12282;
assign n9967 = ~n11264;
assign n6578 = n13780 & n13982;
assign n10586 = n8983 | n5750;
assign n7742 = ~(n2875 | n3226);
assign n7660 = ~n4991;
assign n7364 = ~n7086;
assign n4100 = n10808 | n2444;
assign n4142 = ~(n14370 | n13945);
assign n6992 = n11459 | n9495;
assign n13432 = ~n8595;
assign n9985 = n2760 & n612;
assign n1988 = n10637 | n8218;
assign n1467 = n718 & n14397;
assign n2070 = n8232 & n4202;
assign n12598 = n2461 & n3805;
assign n7422 = ~(n7023 | n1004);
assign n11821 = n5253 | n10484;
assign n6882 = n11313 & n8456;
assign n918 = n9677 & n2269;
assign n3253 = n2562 | n1726;
assign n3172 = n2857 | n11501;
assign n5289 = ~(n12872 | n10263);
assign n7407 = ~n14461;
assign n13389 = ~(n2799 | n12431);
assign n2277 = n11316 & n8536;
assign n13518 = ~n10775;
assign n4523 = ~(n2236 | n7580);
assign n6022 = n10310 | n2061;
assign n3671 = n14319 | n4312;
assign n6093 = n14400 | n11536;
assign n864 = n13107 & n11238;
assign n4279 = n10736 & n10921;
assign n12275 = ~(n1342 | n858);
assign n4258 = n2925 | n7941;
assign n11296 = n5012 & n4787;
assign n2251 = ~n9829;
assign n13454 = n1741 | n6851;
assign n13956 = n11422 & n8460;
assign n12146 = n2747 | n6658;
assign n2451 = ~n7223;
assign n7106 = n12721 & n11638;
assign n6424 = ~n11654;
assign n11640 = n13991 | n6492;
assign n10653 = ~(n4195 | n3676);
assign n7943 = ~n4589;
assign n7105 = ~(n2405 | n9779);
assign n1575 = ~n5690;
assign n10510 = n14110 | n155;
assign n2582 = n14260 & n8234;
assign n2971 = n4856 & n134;
assign n10269 = ~n10219;
assign n6349 = ~(n7809 | n10353);
assign n7948 = n2747 | n7993;
assign n29 = n8404 | n10097;
assign n3661 = n12023 | n11144;
assign n4780 = n227 | n14447;
assign n8257 = ~(n1480 | n8249);
assign n11721 = n12421 & n561;
assign n2596 = n4261 & n711;
assign n2707 = ~(n3521 | n6374);
assign n2365 = n1266 & n6961;
assign n9247 = n5144 | n3896;
assign n13688 = ~(n8353 | n6584);
assign n5457 = n4276 & n8506;
assign n10 = n9423 | n7263;
assign n8952 = n13952 & n12505;
assign n12299 = n6243 & n4600;
assign n13336 = n3076 | n10937;
assign n10371 = n12018 & n5836;
assign n9228 = ~n8552;
assign n11055 = n5683 & n1985;
assign n6174 = n1193 & n540;
assign n6472 = n1193 & n11179;
assign n14421 = n10191 | n8303;
assign n10995 = n2057 | n2598;
assign n1420 = n11647 | n5623;
assign n8493 = n2021 & n9821;
assign n10016 = n12324 | n4603;
assign n9989 = n11411 & n8957;
assign n3117 = n1074 & n14182;
assign n11422 = ~n13360;
assign n8889 = n4340 | n8444;
assign n5439 = n7745 & n11057;
assign n8231 = ~(n2946 | n11485);
assign n10279 = n1452 & n14498;
assign n13276 = ~n1966;
assign n3791 = n12934 | n1235;
assign n9648 = n11748 & n1609;
assign n4550 = n12102 & n12533;
assign n13366 = n1701 | n9418;
assign n8633 = ~(n8015 | n13387);
assign n7330 = n1669 | n5485;
assign n2423 = n9807 | n9834;
assign n3057 = n3815 | n2912;
assign n9279 = n12250 & n3722;
assign n11132 = n79 & n6504;
assign n3039 = n11336 & n12632;
assign n4346 = ~n13908;
assign n2064 = ~n261;
assign n9366 = n1582 | n9332;
assign n8153 = ~(n4207 | n5343);
assign n10006 = ~(n2057 | n344);
assign n6345 = ~(n1623 | n2733);
assign n6853 = n11345 & n4580;
assign n1374 = n3743 & n779;
assign n248 = n2878 | n9739;
assign n3469 = n4967 | n2008;
assign n2158 = ~n1911;
assign n8908 = ~n2970;
assign n10583 = n3914 | n11712;
assign n4313 = ~n4720;
assign n10472 = n5409 | n4681;
assign n7092 = n5999 & n12066;
assign n4831 = n11117 & n13390;
assign n8828 = ~n2130;
assign n12391 = ~n5430;
assign n4812 = n11838 & n6120;
assign n378 = n2643 & n13830;
assign n286 = ~n82;
assign n2071 = n6724 & n2346;
assign n4858 = n3652 & n9683;
assign n6087 = n3449 & n6162;
assign n4612 = n986 & n6605;
assign n8903 = n1059 & n1765;
assign n13187 = n10331 | n1619;
assign n10318 = ~n3442;
assign n12880 = n4821 | n10124;
assign n3087 = n14435 | n12174;
assign n10393 = n8172 | n10642;
assign n10152 = n13342 & n11189;
assign n11201 = n3365 & n4497;
assign n11454 = n11011 | n2227;
assign n11387 = n12229 & n2217;
assign n5554 = n11621 | n6118;
assign n12536 = n8821 | n13024;
assign n10859 = ~(n11508 | n4607);
assign n6597 = n446 & n2293;
assign n810 = n11008 & n4171;
assign n33 = n2985 & n3484;
assign n11970 = n2412 | n10268;
assign n9136 = ~n8049;
assign n6858 = n10506 & n11402;
assign n12583 = n11020 & n13210;
assign n8368 = ~(n10730 | n374);
assign n625 = n6695 | n9474;
assign n8864 = n12601 | n4321;
assign n12348 = n11737 & n8347;
assign n7502 = ~n4147;
assign n3727 = n6205 | n14389;
assign n5544 = n2461 & n8255;
assign n12753 = n13155 | n5394;
assign n3003 = ~n11582;
assign n6639 = n11803 & n11373;
assign n11229 = n11935 | n146;
assign n1912 = n14370 | n8135;
assign n2418 = n8232 & n9746;
assign n1105 = n8575 | n12809;
assign n5182 = ~n12925;
assign n8558 = n11420 | n710;
assign n5444 = n12100 | n10008;
assign n9367 = n3161 | n11507;
assign n4276 = ~n13360;
assign n2488 = ~(n11832 | n9100);
assign n6219 = n361 | n3274;
assign n5399 = n2527 & n133;
assign n11107 = n1576 | n8515;
assign n6771 = n5088 & n8526;
assign n9559 = n7745 & n14187;
assign n10139 = n1875 | n9242;
assign n11903 = ~(n5986 | n1101);
assign n6386 = ~(n1577 | n10627);
assign n9534 = n12986 & n13742;
assign n1145 = n2281 & n7113;
assign n4220 = n3011 | n4811;
assign n3636 = n2025 | n10311;
assign n1921 = n2888 | n11992;
assign n8610 = n7888 | n12973;
assign n4252 = ~(n7919 | n3158);
assign n8235 = n3755 & n3759;
assign n2000 = ~n481;
assign n5918 = ~n2405;
assign n6072 = ~(n14239 | n13807);
assign n8849 = ~n8168;
assign n3964 = ~(n6018 | n8880);
assign n7549 = n8980 | n5203;
assign n8254 = n14319 | n13203;
assign n5929 = n1669 | n8052;
assign n5509 = ~n1780;
assign n10747 = n10245 | n5934;
assign n1611 = ~(n1112 | n5057);
assign n6406 = n116 | n10199;
assign n4061 = n817 | n8067;
assign n5981 = n5137 & n1080;
assign n5104 = ~n1812;
assign n7492 = n695 | n8322;
assign n11230 = n8923 & n917;
assign n1269 = n14091 & n10017;
assign n8188 = n8247 & n2063;
assign n1563 = n1427 & n13156;
assign n13666 = n4199 | n326;
assign n463 = n11935 | n8097;
assign n7416 = n1576 | n12847;
assign n9723 = n7211 & n2508;
assign n868 = n13359 & n13312;
assign n2911 = n4525 & n712;
assign n11080 = n986 & n7996;
assign n9372 = n9494 & n2357;
assign n11985 = n4435 | n6926;
assign n9633 = n4602 | n9355;
assign n4211 = n7912 | n6038;
assign n10917 = ~n10036;
assign n9931 = ~n13165;
assign n13866 = n1788 & n7434;
assign n8985 = n10024 | n4277;
assign n7454 = n6354 & n8891;
assign n5668 = n400 | n8073;
assign n12518 = n820 | n7090;
assign n12311 = ~n11515;
assign n2066 = n5861 | n6380;
assign n642 = n2998 & n11045;
assign n3285 = ~(n7418 | n3816);
assign n5193 = n783 & n3213;
assign n34 = ~n7466;
assign n4624 = ~n8291;
assign n14399 = n10765 & n13916;
assign n1779 = n4973 & n11134;
assign n1059 = ~n12009;
assign n13730 = n11674 & n7935;
assign n12932 = n14074 & n11726;
assign n5487 = n9289 | n5947;
assign n6002 = n13575 & n5093;
assign n8776 = n5038 & n13129;
assign n9485 = n12625 | n1461;
assign n2395 = ~(n14419 | n10459);
assign n7169 = n4923 | n7983;
assign n11088 = ~(n10318 | n13075);
assign n1018 = n11748 & n1983;
assign n9315 = ~n8122;
assign n4591 = n2310 & n7491;
assign n9503 = n228 | n47;
assign n6047 = ~(n7023 | n12447);
assign n591 = n8630 & n2408;
assign n7086 = n9182 & n14060;
assign n9307 = ~(n4299 | n7475);
assign n1101 = ~(n6052 | n5361);
assign n7819 = n1053 & n13298;
assign n5036 = n3888 | n3173;
assign n10416 = n1138 & n7522;
assign n3334 = n3028 & n9894;
assign n5142 = ~(n2194 | n795);
assign n8050 = n9230 | n1215;
assign n6391 = n5986 | n4080;
assign n3193 = ~n11055;
assign n10905 = n13147 & n14077;
assign n4195 = ~n7064;
assign n10458 = ~n12697;
assign n14509 = n8908 | n5277;
assign n3364 = ~n271;
assign n4274 = n10539 | n6234;
assign n11277 = ~(n228 | n5536);
assign n3460 = n511 | n6025;
assign n14187 = n1628 | n5375;
assign n8338 = n4313 | n8611;
assign n1578 = n10834 | n1797;
assign n7535 = n9403 | n6945;
assign n5116 = n13700 & n10974;
assign n7255 = ~n7354;
assign n13362 = ~n7802;
assign n4379 = n4447 & n8901;
assign n10679 = n2985 & n8651;
assign n7484 = ~n14072;
assign n5504 = ~n210;
assign n3446 = ~(n9567 | n12396);
assign n9316 = n10562 & n1359;
assign n11311 = n6507 & n10253;
assign n7304 = n412 | n12836;
assign n8071 = n568 | n9417;
assign n4376 = n7826 & n8998;
assign n2942 = ~n13447;
assign n14155 = n11472 | n11433;
assign n7879 = n815 & n1013;
assign n3171 = ~(n7359 | n7946);
assign n13022 = n8881 | n7967;
assign n7293 = n2985 & n5888;
assign n3846 = ~n4266;
assign n13945 = ~(n14011 | n8882);
assign n3447 = n13379 & n7337;
assign n9451 = n8801 & n1768;
assign n12205 = n11739 | n4737;
assign n13005 = ~n2320;
assign n1104 = n9174 | n7464;
assign n3300 = n7438 | n4751;
assign n7053 = ~n5618;
assign n9924 = ~n6516;
assign n6302 = ~(n8920 | n14508);
assign n1962 = ~n7346;
assign n1960 = n13421 & n13023;
assign n4325 = n14164 & n8540;
assign n6352 = n2017 | n4795;
assign n8408 = n2218 | n11018;
assign n8901 = n13720 & n14031;
assign n13761 = n5562 | n1168;
assign n3149 = n6242 | n4599;
assign n2100 = n11569 & n12471;
assign n8479 = n9151 | n1445;
assign n13254 = n976 | n4874;
assign n6457 = ~(n3457 | n14204);
assign n12986 = ~n11425;
assign n12290 = n4739 | n3237;
assign n5303 = n2724 & n5716;
assign n5726 = n1854 & n4529;
assign n10817 = n748 & n1657;
assign n6695 = ~n5901;
assign n14284 = ~(n1638 | n2917);
assign n14325 = n10032 & n1128;
assign n2706 = n638 & n12241;
assign n14124 = n13108 | n10165;
assign n0 = n8605 & n11884;
assign n12397 = n4404 | n10112;
assign n5055 = n13531 | n5143;
assign n2289 = n13978 | n12176;
assign n8116 = n5007 | n5622;
assign n5109 = n12998 & n11320;
assign n8838 = n6854 & n11914;
assign n12081 = n172 | n11707;
assign n4775 = n9617 & n2093;
assign n5666 = n6323 | n13846;
assign n12868 = n1708 & n12889;
assign n2496 = n678 & n6750;
assign n8476 = ~n10775;
assign n12742 = n8527 | n8324;
assign n3428 = ~n13544;
assign n13690 = n12844 | n12903;
assign n1899 = ~(n2468 | n13947);
assign n5048 = ~n6088;
assign n9212 = n8592 | n2618;
assign n11655 = n13118 | n13126;
assign n7777 = n5899 & n10852;
assign n5098 = ~(n234 | n4818);
assign n11971 = ~(n4633 | n159);
assign n11644 = n9856 | n13591;
assign n12582 = n4967 | n9070;
assign n1913 = n5569 | n11076;
assign n1065 = ~(n7345 | n1167);
assign n83 = n5732 | n2589;
assign n12964 = n14065 & n6134;
assign n3676 = ~(n11508 | n12681);
assign n13796 = n8786 & n14079;
assign n7347 = n2158 & n4670;
assign n8398 = ~n10688;
assign n771 = n10191 | n4078;
assign n5118 = ~n2250;
assign n12760 = n2315 | n9273;
assign n6697 = ~n7091;
assign n4580 = ~(n5026 | n10088);
assign n5485 = n5779 & n1909;
assign n8033 = n12802 & n9300;
assign n5759 = n2669 & n5270;
assign n3911 = n7529 & n20;
assign n13656 = ~n13139;
assign n8286 = ~(n13941 | n9352);
assign n11008 = ~n6829;
assign n2631 = ~(n11581 | n8330);
assign n8555 = ~n2298;
assign n720 = n748 & n5655;
assign n6272 = n12019 | n13800;
assign n14073 = n4722 & n13059;
assign n3224 = n286 & n10584;
assign n7500 = ~(n12322 | n12937);
assign n1989 = n1610 & n12566;
assign n14430 = ~n12588;
assign n7892 = n13413 | n14162;
assign n12957 = ~n14433;
assign n1115 = n7911 & n3348;
assign n5462 = n1699 & n6495;
assign n4479 = n4925 | n1898;
assign n7241 = n6981 | n427;
assign n8312 = ~(n9984 | n6);
assign n2800 = n5472 | n7018;
assign n8014 = n13016 | n7959;
assign n10300 = ~n9878;
assign n347 = n10035 | n191;
assign n9124 = ~n5921;
assign n13131 = n10969 & n2173;
assign n11627 = n9186 & n12423;
assign n13354 = ~n203;
assign n13988 = n1489 & n5523;
assign n9332 = n1125 & n3118;
assign n5719 = n8964 | n4617;
assign n9356 = n7812 | n7721;
assign n7223 = ~n10055;
assign n13522 = ~n13784;
assign n6014 = n13489 & n4676;
assign n10987 = n4973 & n6870;
assign n7935 = n10351 | n5222;
assign n1900 = n730 & n9444;
assign n5353 = n13850 & n10873;
assign n9846 = n513 & n34;
assign n3835 = n611 | n2309;
assign n9362 = n11804 | n9051;
assign n12030 = ~(n8825 | n6335);
assign n11257 = n7693 & n9976;
assign n2957 = n5312 & n10544;
assign n11003 = n2583 & n13833;
assign n13274 = ~(n6672 | n9653);
assign n8787 = n6016 & n13177;
assign n11779 = n11420 | n8680;
assign n564 = n7673 & n3176;
assign n6042 = n11171 | n12919;
assign n7596 = ~n11628;
assign n13665 = n3047 | n8377;
assign n3470 = n225 & n998;
assign n386 = ~(n10637 | n14174);
assign n4335 = n3126 | n8382;
assign n12206 = n5815 | n8493;
assign n7626 = n11315 | n5709;
assign n9172 = ~n2417;
assign n296 = n7529 & n8574;
assign n6930 = n3134 | n13615;
assign n3280 = n11117 & n12298;
assign n8453 = ~n13219;
assign n14160 = n13520 & n10586;
assign n1176 = n4347 & n13604;
assign n13951 = n13706 | n6455;
assign n11880 = n11909 | n7009;
assign n13182 = n10506 & n5107;
assign n14170 = ~(n13153 | n3990);
assign n8922 = n11157 & n13716;
assign n14100 = n12844 | n11310;
assign n12674 = n11183 | n11292;
assign n8727 = ~(n12127 | n11283);
assign n8158 = ~(n4572 | n6278);
assign n3925 = n2874 | n1025;
assign n1837 = n1535 | n10600;
assign n7220 = n4244 & n3347;
assign n337 = n1140 & n1360;
assign n179 = n7963 & n5654;
assign n14106 = ~n9863;
assign n12085 = n9804 | n581;
assign n7027 = ~n8361;
assign n5686 = n3546 | n1563;
assign n4527 = ~n10630;
assign n10317 = ~(n8767 | n5214);
assign n6845 = n11816 & n7817;
assign n1330 = n11036 | n7424;
assign n9667 = n2158 & n9480;
assign n11608 = n3815 | n6578;
assign n6531 = ~n10377;
assign n2634 = n7267 & n13330;
assign n3589 = n4631 | n9153;
assign n9862 = ~(n6933 | n7459);
assign n3011 = ~n918;
assign n11353 = ~(n2057 | n3446);
assign n14244 = n1701 | n2442;
assign n2801 = n1356 | n9917;
assign n7613 = n13464 & n2244;
assign n10035 = ~n1676;
assign n8350 = n13991 | n8989;
assign n12342 = n8490 | n14474;
assign n14250 = ~(n5944 | n10355);
assign n11210 = n7267 & n6179;
assign n11629 = n8210 | n1689;
assign n9860 = n12250 & n6566;
assign n13299 = n11090 | n10382;
assign n4794 = n6354 & n4571;
assign n788 = ~n2226;
assign n5163 = n10330 & n9210;
assign n10720 = n4357 | n970;
assign n7157 = n11153 & n2423;
assign n13062 = ~(n14198 | n11512);
assign n5092 = ~n5606;
assign n7254 = n10566 & n7149;
assign n5731 = n13823 & n1430;
assign n1700 = n11011 | n2782;
assign n9561 = n13885 | n1397;
assign n8063 = n619 | n1368;
assign n9620 = ~n9596;
assign n12804 = n2877 | n2676;
assign n4254 = n12292 | n14452;
assign n2834 = ~(n2098 | n6315);
assign n11635 = n2564 & n11527;
assign n2739 = ~(n2651 | n11535);
assign n13166 = n12039 & n4776;
assign n3426 = n8147 & n1964;
assign n7056 = n6147 | n11842;
assign n1231 = ~n5197;
assign n5360 = n1857 & n7351;
assign n12985 = n14321 & n5567;
assign n2657 = n2229 | n10164;
assign n1741 = ~n7404;
assign n1270 = n6128 & n7945;
assign n4921 = n6507 & n7405;
assign n3565 = ~n1462;
assign n14477 = n954 | n2861;
assign n8457 = n13597 & n1252;
assign n10451 = n13432 | n10721;
assign n1229 = n9140 | n14309;
assign n513 = n582 | n4774;
assign n11593 = n13005 | n3453;
assign n1680 = n6323 | n4764;
assign n1652 = ~(n7091 | n11469);
assign n8020 = ~n7223;
assign n5139 = ~n9580;
assign n1240 = n4803 & n7578;
assign n2937 = n1172 | n909;
assign n6798 = ~(n7364 | n14385);
assign n54 = n11814 & n9184;
assign n5287 = n12461 & n6304;
assign n7438 = ~n628;
assign n4936 = n10234 | n6728;
assign n10537 = n317 | n11524;
assign n9384 = n1840 | n7509;
assign n13682 = ~n10061;
assign n11355 = n974 | n4725;
assign n11894 = n3559 | n12977;
assign n901 = n98 & n4275;
assign n13769 = n1937 & n7398;
assign n11965 = n11620 | n4004;
assign n10941 = n2758 & n2338;
assign n6920 = n14321 & n10611;
assign n6010 = n3743 & n11509;
assign n2006 = ~n10177;
assign n9475 = ~(n5365 | n2185);
assign n3278 = n12226 & n10288;
assign n11446 = ~(n8527 | n6386);
assign n11851 = n9853 & n11735;
assign n8047 = ~n920;
assign n4741 = ~n7819;
assign n12355 = n14464 & n12766;
assign n6162 = n1361 | n13093;
assign n14484 = n5575 | n10675;
assign n924 = n10461 | n3326;
assign n4998 = n14145 & n484;
assign n6411 = n2527 & n614;
assign n3675 = ~n3166;
assign n3549 = n14210 | n8649;
assign n4089 = n2322 & n992;
assign n6658 = n7026 & n2088;
assign n4435 = ~n1267;
assign n4842 = n13252 & n8421;
assign n14350 = n2531 | n2557;
assign n8659 = n492 | n10636;
assign n12294 = ~n3704;
assign n4427 = n7957 & n12178;
assign n12212 = n7436 | n9224;
assign n13744 = n4354 & n3086;
assign n5081 = n9198 & n2051;
assign n816 = n1074 & n223;
assign n12840 = n553 | n3738;
assign n1041 = n7814 & n8398;
assign n9091 = n13850 & n10220;
assign n2508 = n9140 | n9093;
assign n4929 = ~n13981;
assign n7443 = ~n8451;
assign n5633 = n5104 & n1415;
assign n9013 = n12412 & n10747;
assign n13482 = n14088 | n10522;
assign n6968 = n1820 | n7409;
assign n9875 = ~(n1612 | n11051);
assign n12987 = n783 & n9117;
assign n10550 = n5997 | n497;
assign n1088 = n6263 | n13821;
assign n6215 = n8096 | n835;
assign n12139 = ~n4891;
assign n13203 = n14091 & n9459;
assign n10798 = n10396 | n10742;
assign n10602 = n13096 & n7123;
assign n4120 = n13155 | n4868;
assign n11771 = ~n3280;
assign n3622 = n4199 | n10905;
assign n14465 = ~n8963;
assign n1714 = ~(n9754 | n2233);
assign n3174 = n5048 & n1986;
assign n2058 = ~n10254;
assign n14296 = ~n9182;
assign n6802 = n1728 | n3022;
assign n10646 = ~n10378;
assign n6348 = n2583 & n11065;
assign n3962 = n11157 & n2779;
assign n6001 = n13641 & n149;
assign n10890 = n6595 | n6865;
assign n12854 = n1189 | n7863;
assign n1109 = n5873 | n10255;
assign n11874 = n3667 | n10577;
assign n8808 = n3904 & n2237;
assign n12604 = n10815 & n8185;
assign n3191 = ~n12403;
assign n12735 = n3286 & n7772;
assign n5159 = ~n1365;
assign n1895 = n10197 & n3728;
assign n516 = ~(n6434 | n10963);
assign n3879 = n1409 & n2316;
assign n10375 = n2473 & n8743;
assign n12478 = n1834 | n3174;
assign n8954 = n9944 & n14428;
assign n2558 = n1494 | n10718;
assign n12219 = n14358 & n12228;
assign n12765 = ~n10047;
assign n12942 = n3134 | n5753;
assign n13721 = n14366 | n5314;
assign n586 = n1391 | n9308;
assign n4185 = ~(n5986 | n12508);
assign n5214 = n3861 & n4318;
assign n4747 = ~(n3768 | n9395);
assign n1715 = n11163 & n5925;
assign n7521 = n888 | n12829;
assign n12630 = ~n7846;
assign n2881 = ~(n7584 | n609);
assign n11966 = n13354 | n737;
assign n4715 = n13017 & n3817;
assign n5478 = n553 | n2460;
assign n6925 = n4313 | n13628;
assign n11034 = n5335 & n7420;
assign n10970 = n4347 & n9876;
assign n6809 = n2686 | n6659;
assign n14429 = n1254 & n13836;
assign n14358 = ~n7507;
assign n9190 = ~n1417;
assign n637 = n5414 & n310;
assign n10717 = n12159 & n2249;
assign n12450 = ~n10055;
assign n11663 = n3886 | n13942;
assign n5385 = ~(n12548 | n13672);
assign n9427 = n5480 | n11023;
assign n4226 = n791 | n9961;
assign n8809 = n10059 & n13259;
assign n5011 = ~n168;
assign n1759 = n4276 & n6108;
assign n9222 = n6609 & n9433;
assign n6559 = ~n11264;
assign n1971 = n7250 | n5819;
assign n10294 = ~n426;
assign n8094 = n9952 & n8327;
assign n7226 = n7481 | n13171;
assign n5219 = n3025 | n5546;
assign n10174 = n7043 & n4855;
assign n10455 = n5084 | n8765;
assign n2746 = n2784 | n137;
assign n5795 = ~n6534;
assign n898 = ~n442;
assign n11018 = n12105 & n5809;
assign n9464 = n12472 & n9301;
assign n10685 = n10015 & n4578;
assign n7883 = n3914 | n2266;
assign n13793 = n7421 & n2287;
assign n3040 = ~(n5288 | n1534);
assign n12261 = n10913 | n9149;
assign n14287 = n9297 & n7731;
assign n7234 = ~(n8015 | n4110);
assign n1854 = ~n304;
assign n4487 = n10871 | n8307;
assign n9022 = n12528 & n1557;
assign n11368 = n5335 & n6635;
assign n3249 = n782 | n9873;
assign n1353 = n6016 & n5697;
assign n9281 = n8372 & n13832;
assign n2877 = ~n3070;
assign n3025 = ~n5627;
assign n9857 = n3800 | n13441;
assign n10335 = n2597 | n3063;
assign n9681 = n11183 | n854;
assign n5988 = n12169 | n6381;
assign n4683 = n9229 | n9723;
assign n9768 = ~(n1769 | n10349);
assign n6329 = n8965 & n1493;
assign n12996 = n8242 | n14489;
assign n4320 = ~n4117;
assign n13269 = n10710 & n10702;
assign n2831 = n7068 & n1313;
assign n5853 = n13781 & n9970;
assign n10657 = n3401 & n9435;
assign n13067 = n14373 & n6967;
assign n10121 = ~n7979;
assign n11120 = n8507 & n5196;
assign n8189 = ~n496;
assign n12463 = n11572 | n14032;
assign n8281 = n11748 & n3207;
assign n14246 = ~(n1623 | n14384);
assign n10036 = ~n1938;
assign n2656 = n9853 & n9533;
assign n9800 = n361 | n3814;
assign n4529 = n13477 | n3954;
assign n13064 = n13246 & n3298;
assign n6385 = n7421 & n8479;
assign n7020 = n873 & n11173;
assign n11515 = ~n300;
assign n4051 = n13404 & n14177;
assign n11585 = n4065 | n8235;
assign n11324 = n4698 & n1395;
assign n2721 = n1452 & n5494;
assign n10725 = n5064 | n4374;
assign n3192 = n10461 | n2494;
assign n12154 = n3099 | n1308;
assign n7369 = n12101 & n1831;
assign n14413 = n12543 | n7800;
assign n12568 = ~n9846;
assign n782 = ~n12746;
assign n11087 = n12139 | n7877;
assign n6787 = ~n885;
assign n829 = n4525 & n9168;
assign n415 = n14337 | n2435;
assign n5758 = n568 | n11210;
assign n12002 = ~(n5569 | n1851);
assign n5003 = n7068 & n1419;
assign n3111 = n55 & n5526;
assign n4084 = n3861 & n3411;
assign n3434 = ~n2029;
assign n11402 = n7438 | n5091;
assign n2082 = ~n7681;
assign n1648 = n11951 | n9324;
assign n858 = ~(n11047 | n3645);
assign n7693 = ~n11425;
assign n3175 = n6753 & n1187;
assign n12922 = ~n7077;
assign n7315 = n3485 & n11840;
assign n10814 = ~(n12968 | n10200);
assign n154 = n4435 | n2710;
assign n2142 = n11953 | n3744;
assign n10793 = ~(n7145 | n8818);
assign n120 = n4806 & n7611;
assign n8726 = ~n2545;
assign n10427 = n12023 | n8177;
assign n12024 = ~(n8363 | n6477);
assign n8136 = n11020 & n13758;
assign n10852 = n6350 | n907;
assign n8288 = ~n1086;
assign n12837 = n8825 | n5141;
assign n280 = n10784 | n13913;
assign n5713 = n8209 | n13470;
assign n9547 = n8801 & n2687;
assign n3594 = n12034 | n9250;
assign n8101 = ~(n1813 | n12316);
assign n914 = n2533 & n5417;
assign n11189 = n10083 | n10336;
assign n4846 = n7211 & n14442;
assign n6318 = ~n13723;
assign n2639 = n8427 & n11759;
assign n8220 = n2529 & n13840;
assign n7007 = ~n4210;
assign n2879 = ~(n4544 | n10980);
assign n6903 = n13682 | n12885;
assign n9990 = ~(n717 | n4201);
assign n5398 = n1225 & n11062;
assign n890 = n5762 | n5441;
assign n14482 = n11803 & n14124;
assign n6134 = n8866 | n7282;
assign n3419 = ~n2573;
assign n12938 = n1699 & n3249;
assign n1770 = n12986 & n7353;
assign n13440 = n10015 & n12567;
assign n3343 = n1172 | n7032;
assign n181 = n387 | n380;
assign n14499 = n3099 | n8838;
assign n7658 = ~(n8544 | n2666);
assign n12660 = n3247 & n8685;
assign n13755 = ~n11369;
assign n12413 = n2874 | n2327;
assign n182 = n2099 & n5528;
assign n7372 = ~(n14058 | n5902);
assign n7388 = n98 & n449;
assign n2456 = n2747 | n4167;
assign n3147 = n904 & n2989;
assign n3090 = n650 & n14222;
assign n322 = ~(n5509 | n2170);
assign n2474 = ~n5014;
assign n11394 = n3512 | n11701;
assign n3691 = n6507 & n3002;
assign n3918 = n6848 & n9031;
assign n6562 = n2908 | n3533;
assign n11983 = n5997 | n4257;
assign n11126 = n12034 | n6010;
assign n10683 = n412 | n13795;
assign n12209 = ~n7104;
assign n7451 = n3607 & n14425;
assign n1781 = n11440 | n5388;
assign n10614 = n227 | n7813;
assign n12106 = n5734 & n13002;
assign n3461 = ~n9563;
assign n13798 = n5899 & n6115;
assign n2239 = n14157 & n7653;
assign n11988 = ~n10358;
assign n11122 = n8649 & n7124;
assign n7973 = ~n7177;
assign n12338 = n8697 & n10768;
assign n8450 = ~n6758;
assign n7309 = n13728 | n13102;
assign n950 = n3287 | n8419;
assign n8381 = n12531 & n9083;
assign n3219 = ~n9306;
assign n11256 = n10624 | n1716;
assign n9516 = n1401 | n6693;
assign n7806 = ~(n4299 | n12672);
assign n3106 = n8404 | n7894;
assign n2490 = n6744 & n9427;
assign n12548 = ~n11435;
assign n7082 = n7898 | n7324;
assign n12537 = n14188 | n10078;
assign n3329 = n11647 | n5679;
assign n6106 = n6507 & n111;
assign n5402 = n6013 & n7595;
assign n3402 = ~n14365;
assign n589 = n3952 & n2050;
assign n13162 = n2820 & n3537;
assign n8212 = ~n7007;
assign n13368 = n12576 | n2449;
assign n6066 = n13379 & n3350;
assign n3395 = ~n9740;
assign n6286 = n3527 | n5535;
assign n493 = n10136 | n12773;
assign n5607 = n889 & n10940;
assign n14319 = ~n12394;
assign n8681 = n12169 | n7881;
assign n4727 = n647 | n7659;
assign n1641 = n4289 & n6803;
assign n13457 = n12820 | n11513;
assign n2043 = n7527 | n5545;
assign n10748 = n10323 | n7472;
assign n622 = n7979 & n4713;
assign n8375 = n428 & n11550;
assign n10359 = n9944 & n856;
assign n12870 = ~n12444;
assign n13651 = n55 & n7111;
assign n8832 = n5275 & n11197;
assign n4068 = n13707 | n7687;
assign n3279 = n2587 & n3801;
assign n12756 = n10035 | n4099;
assign n4693 = ~(n12968 | n6551);
assign n13655 = n7527 | n3614;
assign n12176 = n11702 & n6356;
assign n6415 = n7284 & n10538;
assign n8023 = ~n5738;
assign n9242 = n2564 & n414;
assign n12601 = ~n13165;
assign n6599 = n11231 | n1075;
assign n9233 = n405 & n10829;
assign n10043 = n13700 & n3711;
assign n2480 = n1031 | n3349;
assign n7467 = n13147 & n7384;
assign n10516 = ~n8008;
assign n9103 = n7429 & n362;
assign n10062 = ~n13668;
assign n2137 = ~n12136;
assign n98 = ~n11547;
assign n7464 = n14093 & n896;
assign n2065 = n8425 | n6938;
assign n5658 = n1031 | n668;
assign n7547 = n11607 & n5496;
assign n1412 = n10713 | n157;
assign n7513 = n10024 | n7734;
assign n9622 = n9804 | n11290;
assign n8440 = n3846 & n2268;
assign n10116 = n3942 & n14161;
assign n5941 = ~(n7466 | n7397);
assign n4988 = ~n9354;
assign n10142 = n10089 | n13712;
assign n12807 = ~n9769;
assign n12187 = n8480 | n13828;
assign n8036 = n11047 | n5425;
assign n6182 = n1804 & n3172;
assign n6965 = n9562 | n6586;
assign n9511 = n5715 | n10192;
assign n61 = n5603 | n6377;
assign n8248 = n647 | n7329;
assign n2204 = n2583 & n3398;
assign n13815 = n3485 & n2393;
assign n9308 = n9232 & n295;
assign n6217 = ~(n11980 | n430);
assign n5082 = n7717 & n9882;
assign n477 = n898 & n3403;
assign n2035 = n3164 | n10810;
assign n5138 = n2218 | n11245;
assign n2994 = n9716 | n65;
assign n3994 = n3904 & n2563;
assign n3786 = n1535 | n3220;
assign n8434 = n14465 & n6078;
assign n10111 = n10351 | n5347;
assign n2257 = n6556 & n10880;
assign n10699 = n10820 & n173;
assign n12684 = n13489 & n3341;
assign n7334 = ~n3191;
assign n1359 = n13432 | n7368;
assign n2514 = n4923 | n2864;
assign n5090 = n7596 & n7325;
assign n13304 = n4300 & n5357;
assign n9272 = n13869 | n8892;
assign n797 = n523 | n13799;
assign n2594 = n6192 & n12582;
assign n14196 = ~n752;
assign n6447 = n8372 & n6161;
assign n662 = n7015 & n6685;
assign n5921 = ~n4928;
assign n6669 = n7683 | n9446;
assign n4343 = n7063 & n6024;
assign n8061 = n5876 & n7142;
assign n3885 = n9620 | n11851;
assign n13892 = ~(n8816 | n12238);
assign n2525 = n1775 & n794;
assign n5113 = n9856 | n7016;
assign n7176 = n5236 | n4729;
assign n11919 = n2179 | n11618;
assign n4181 = n7810 & n6341;
assign n3903 = n6046 | n7131;
assign n11911 = ~(n6989 | n12298);
assign n2442 = n14321 & n14302;
assign n12534 = n9442 | n296;
assign n12814 = n3161 | n4015;
assign n13055 = ~n937;
assign n5154 = n2149 | n10167;
assign n10218 = n9490 | n1129;
assign n9850 = n4574 & n256;
assign n8138 = ~(n1706 | n14057);
assign n2691 = n2218 | n7775;
assign n5383 = n1588 & n11312;
assign n5684 = n6706 | n10259;
assign n13323 = n8575 | n10797;
assign n10678 = ~n14501;
assign n5657 = n7057 & n9554;
assign n13153 = ~n4007;
assign n6726 = n4932 & n9163;
assign n6649 = ~n7621;
assign n8721 = ~n5943;
assign n12545 = n1147 | n1089;
assign n11457 = n9745 & n5875;
assign n13165 = n11052 & n9751;
assign n6793 = n3286 & n9194;
assign n12047 = ~n6804;
assign n4854 = n8007 & n12122;
assign n956 = ~(n9035 | n2302);
assign n10965 = n3709 & n8794;
assign n172 = ~n11456;
assign n3517 = ~(n7971 | n8643);
assign n4973 = ~n13003;
assign n13531 = ~n3681;
assign n8364 = n7003 | n2477;
assign n4114 = n10822 & n5304;
assign n3376 = n2877 | n10888;
assign n2224 = ~n4618;
assign n6605 = n7426 | n12711;
assign n11574 = ~n4050;
assign n11358 = n4876 | n9918;
assign n38 = n10960 | n8937;
assign n7523 = ~n13102;
assign n8817 = ~n737;
assign n12121 = n13912 | n12218;
assign n9286 = n6525 & n12301;
assign n4264 = n12549 | n4590;
assign n11182 = n12870 | n9798;
assign n7710 = n2188 | n6114;
assign n10655 = ~(n7359 | n4455);
assign n8372 = ~n1478;
assign n9099 = n14388 & n5789;
assign n7003 = ~n9371;
assign n6819 = ~n1979;
assign n4985 = n7081 & n14457;
assign n2563 = n13074 | n12952;
assign n13248 = ~n9231;
assign n8991 = ~(n13874 | n12224);
assign n409 = n12850 & n13257;
assign n10740 = n511 | n1115;
assign n10803 = ~n3544;
assign n10943 = n3435 & n14292;
assign n6885 = n7043 & n3030;
assign n6837 = n7208 & n12056;
assign n13470 = n2224 & n2127;
assign n9260 = n5625 | n4881;
assign n10071 = n13069 & n6947;
assign n6139 = ~n3493;
assign n124 = n10589 & n6170;
assign n13492 = n10506 & n9734;
assign n3272 = ~(n10091 | n9400);
assign n3031 = n2229 | n6564;
assign n8992 = n10351 | n3539;
assign n9868 = n12543 | n13382;
assign n3941 = n1354 & n5885;
assign n8518 = ~(n3211 | n13121);
assign n4668 = n10197 & n6720;
assign n1219 = ~(n2171 | n14116);
assign n7191 = n8111 & n8667;
assign n1258 = ~n9354;
assign n7636 = n5132 | n5313;
assign n8465 = n5434 & n1212;
assign n2467 = ~(n11017 | n1432);
assign n11525 = n7429 & n508;
assign n11658 = n387 | n6939;
assign n6814 = n555 | n10440;
assign n5378 = n2985 & n6391;
assign n1625 = n5899 & n5334;
assign n7929 = n9228 | n1637;
assign n5291 = n10930 & n13805;
assign n12691 = ~n1812;
assign n11972 = n7426 | n212;
assign n7621 = ~n637;
assign n1713 = ~n8899;
assign n398 = n7781 & n12435;
assign n3100 = n2315 | n1517;
assign n4112 = n12615 & n1939;
assign n8206 = n9080 & n4178;
assign n14168 = ~(n99 | n9985);
assign n6801 = n6596 | n13064;
assign n7602 = n9015 & n11642;
assign n4245 = n12400 | n12905;
assign n7213 = n12034 | n13456;
assign n13826 = ~(n13055 | n12272);
assign n5705 = n3491 & n1500;
assign n2197 = n85 | n7321;
assign n11196 = n1699 & n10258;
assign n5480 = ~n2545;
assign n9130 = n13718 | n552;
assign n10779 = n1729 & n8618;
assign n12812 = n12147 & n610;
assign n10386 = n13700 & n12281;
assign n9092 = ~(n4535 | n3285);
assign n4389 = n405 & n14046;
assign n13181 = ~n12409;
assign n5456 = n12568 | n6197;
assign n2143 = n14313 & n8896;
assign n283 = ~n8695;
assign n3144 = n14435 | n1440;
assign n7365 = ~n12096;
assign n4956 = n1356 | n14206;
assign n3915 = n4901 & n13738;
assign n11536 = n10969 & n2882;
assign n13196 = n329 | n3807;
assign n3998 = n12351 | n7499;
assign n5691 = n4205 | n2876;
assign n5177 = ~(n11597 | n12103);
assign n14087 = n4276 & n10842;
assign n11730 = ~(n3400 | n7209);
assign n1552 = ~(n2005 | n6798);
assign n13523 = n28 | n6560;
assign n8080 = ~(n12527 | n13279);
assign n11215 = n5348 & n12204;
assign n2067 = ~n6693;
assign n6760 = ~(n9806 | n1226);
assign n10493 = n13080 | n3706;
assign n5366 = ~(n14239 | n13892);
assign n13555 = ~n6990;
assign n2341 = ~n13041;
assign n7411 = n7221 & n7298;
assign n12150 = n3904 & n1680;
assign n150 = n89 | n6579;
assign n8400 = n1074 & n6570;
assign n603 = n6899 & n2480;
assign n2415 = ~n14461;
assign n13837 = n10678 & n1651;
assign n11290 = n4163 & n4013;
assign n11205 = n10408 & n23;
assign n11114 = ~(n7624 | n9519);
assign n14156 = n11572 | n3175;
assign n12390 = ~(n14419 | n7965);
assign n2587 = ~n3967;
assign n371 = n5548 | n8310;
assign n3572 = ~n8798;
assign n13512 = n11440 | n196;
assign n9224 = n889 & n8391;
assign n2020 = n5807 | n7163;
assign n7525 = n11094 | n13881;
assign n13442 = ~(n1812 | n7834);
assign n2932 = ~n5438;
assign n11578 = ~(n4333 | n12060);
assign n5564 = n1660 | n982;
assign n11223 = ~n13696;
assign n8538 = n3028 & n11719;
assign n5122 = n3011 | n5785;
assign n1426 = ~(n7146 | n11630);
assign n817 = ~n6264;
assign n11623 = n4346 & n9626;
assign n10316 = n11704 | n14374;
assign n1805 = ~n8813;
assign n4362 = n4788 & n3516;
assign n13360 = ~n4830;
assign n8736 = n12075 | n13455;
assign n985 = n13220 | n3386;
assign n10775 = n11100 & n12593;
assign n7721 = n11220 & n6558;
assign n12141 = n3586 & n5238;
assign n5917 = n10784 | n6127;
assign n3207 = n13112 | n4565;
assign n8765 = n7060 & n10031;
assign n3858 = n12130 | n6921;
assign n1327 = ~(n7589 | n9848);
assign n1828 = n11558 | n14410;
assign n7560 = n1685 | n12274;
assign n86 = ~(n4877 | n554);
assign n6718 = n10394 | n9123;
assign n1460 = ~(n11148 | n2851);
assign n4054 = n12494 | n13160;
assign n585 = n4615 | n730;
assign n3162 = n14157 & n10140;
assign n10372 = ~n13047;
assign n11628 = ~n6212;
assign n4015 = n9650 & n3317;
assign n2688 = ~(n234 | n1026);
assign n3393 = n12019 | n3473;
assign n11922 = n2547 & n7586;
assign n6644 = ~(n8942 | n5626);
assign n8959 = ~n5218;
assign n7529 = ~n4266;
assign n3303 = n9811 & n11072;
assign n3151 = n5471 & n13962;
assign n2675 = n11422 & n9582;
assign n13908 = ~n6058;
assign n5814 = n7529 & n3578;
assign n6008 = n9509 & n10890;
assign n6034 = n12250 & n10509;
assign n13507 = ~n2699;
assign n8004 = n8897 | n8851;
assign n3045 = n7530 | n6103;
assign n6938 = n9134 | n2041;
assign n13034 = n9191 & n7690;
assign n8624 = n11472 | n9081;
assign n12526 = n4631 | n11221;
assign n8474 = n783 & n13318;
assign n11291 = n4447 & n6734;
assign n11981 = n9673 | n14072;
assign n7814 = n9280 | n3388;
assign n2381 = n1699 & n8608;
assign n1046 = n7267 & n71;
assign n6683 = n11220 & n6463;
assign n5068 = n13142 | n8583;
assign n2626 = n8605 & n4849;
assign n5250 = ~(n4233 | n13049);
assign n2032 = n10523 | n14173;
assign n75 = ~(n4639 | n10492);
assign n8973 = n9780 | n4188;
assign n13180 = n8458 | n13924;
assign n10206 = n11495 & n10034;
assign n5682 = n5548 | n10944;
assign n1668 = n14430 | n11808;
assign n7880 = n3276 & n10010;
assign n12989 = n3893 & n12253;
assign n988 = n748 & n11319;
assign n11530 = n11551 | n12710;
assign n3432 = n10854 & n13197;
assign n6893 = ~(n9807 | n1293);
assign n9508 = n13535 & n13579;
assign n12953 = ~n1843;
assign n530 = n1805 | n10362;
assign n10732 = n10834 | n8810;
assign n6298 = n4527 & n12738;
assign n943 = n10357 & n9143;
assign n8110 = n8569 & n5949;
assign n13952 = ~n230;
assign n7380 = n6854 & n4623;
assign n1256 = n8020 & n8415;
assign n8729 = ~(n8404 | n10480);
assign n3939 = n8697 & n2613;
assign n7078 = n7426 | n1674;
assign n9654 = ~n8044;
assign n3397 = n3743 & n12668;
assign n6733 = n4690 & n11801;
assign n6607 = ~n9846;
assign n13369 = n10458 & n1290;
assign n11728 = n7418 | n2198;
assign n12969 = n14351 & n4727;
assign n4729 = n79 & n11067;
assign n9639 = ~(n14419 | n989);
assign n10095 = n6625 & n370;
assign n12077 = n11086 | n10552;
assign n2697 = n9269 | n2305;
assign n9231 = ~n5944;
assign n11939 = n2942 & n1990;
assign n14002 = n3277 & n6149;
assign n11790 = n776 & n11588;
assign n6274 = n3989 & n6660;
assign n11540 = n11620 | n981;
assign n8879 = n12531 & n5453;
assign n3603 = n3130 & n6081;
assign n10509 = n5406 | n4850;
assign n14116 = ~(n1480 | n3685);
assign n2485 = n2445 & n2805;
assign n3494 = n7211 & n840;
assign n12222 = n4876 | n3821;
assign n3302 = ~(n11581 | n7702);
assign n2928 = ~(n3546 | n5247);
assign n1468 = ~(n4897 | n3694);
assign n8773 = n5891 | n4520;
assign n8918 = n8250 & n4208;
assign n8825 = ~n4777;
assign n4677 = n200 & n1819;
assign n9205 = ~(n6971 | n10588);
assign n3580 = n7060 & n12416;
assign n2370 = ~n5504;
assign n1901 = n647 | n8465;
assign n7266 = n14286 | n3893;
assign n554 = ~(n11975 | n12143);
assign n2819 = n11183 | n10643;
assign n5689 = n4340 | n4591;
assign n12427 = n13359 & n4432;
assign n12267 = n9890 & n12767;
assign n13089 = n5279 & n4176;
assign n12163 = n12759 | n13931;
assign n10181 = n4631 | n1259;
assign n5980 = n13466 | n1702;
assign n4701 = n3088 | n10874;
assign n4958 = n2682 & n12688;
assign n5105 = n12918 & n4934;
assign n408 = n511 | n1987;
assign n8778 = n3672 & n11170;
assign n6613 = ~(n7120 | n4348);
assign n8458 = ~n4550;
assign n4031 = n14166 | n11533;
assign n6026 = n3088 | n11872;
assign n2933 = n6323 | n11187;
assign n10997 = n8964 | n13131;
assign n10553 = n4261 & n10550;
assign n11287 = n12401 | n13267;
assign n11197 = n9403 | n13841;
assign n5382 = n10224 | n10273;
assign n2814 = n2445 & n10385;
assign n8007 = ~n11428;
assign n3757 = n5229 & n2679;
assign n1830 = n13240 & n2595;
assign n1717 = n11213 & n14257;
assign n14008 = n9229 | n10473;
assign n9564 = ~n6657;
assign n5798 = n13407 & n2745;
assign n12182 = n4925 | n9916;
assign n4777 = n12658 & n482;
assign n231 = ~n5871;
assign n10858 = n7667 | n10147;
assign n14379 = n14373 & n7574;
assign n3451 = n8453 & n7787;
assign n4765 = ~n8487;
assign n2820 = ~n3356;
assign n4486 = ~n1120;
assign n14079 = n13005 | n9900;
assign n10648 = ~n1109;
assign n583 = n12020 | n403;
assign n5674 = n3332 & n12300;
assign n10476 = n14401 | n9722;
assign n7858 = n8172 | n5843;
assign n11007 = n2181 | n10800;
assign n10331 = ~n4847;
assign n481 = ~n7120;
assign n10162 = n718 & n11265;
assign n11856 = n9069 & n1058;
assign n4152 = ~(n1348 | n12310);
assign n3187 = n9864 | n10749;
assign n9507 = ~n2320;
assign n765 = n7768 & n9593;
assign n12039 = ~n5525;
assign n8431 = ~n13734;
assign n7333 = n12494 | n3723;
assign n13220 = ~n7875;
assign n1332 = ~n6703;
assign n6820 = n1772 & n1589;
assign n3113 = n5634 | n8552;
assign n7603 = n7961 & n11672;
assign n1511 = n8412 & n5866;
assign n11226 = n3635 & n4496;
assign n9986 = n13080 | n4838;
assign n978 = n10294 | n14279;
assign n7182 = n10300 | n1108;
assign n11802 = ~(n7418 | n13661);
assign n2352 = ~(n2016 | n11114);
assign n5556 = n7697 | n11689;
assign n5300 = n4433 & n7313;
assign n13620 = n9650 & n12698;
assign n4133 = ~(n7362 | n7197);
assign n14294 = n1047 & n6363;
assign n2648 = n5948 & n4886;
assign n11832 = ~n12949;
assign n9207 = ~(n12757 | n8138);
assign n7629 = n850 | n6450;
assign n5590 = n2224 & n5929;
assign n9855 = n8897 | n9578;
assign n8843 = n2272 | n3162;
assign n12346 = n7697 | n6598;
assign n1659 = n4357 | n11721;
assign n1508 = n10619 | n11776;
assign n1664 = n89 | n339;
assign n8900 = ~(n7145 | n352);
assign n11793 = n12900 | n2164;
assign n9922 = ~(n4608 | n11446);
assign n4392 = n4932 & n13167;
assign n3809 = n7744 | n2065;
assign n8095 = n1494 | n13182;
assign n11153 = ~n9994;
assign n8239 = n5312 & n9844;
assign n11501 = n3635 & n11834;
assign n10584 = n12549 | n13592;
assign n8851 = n1788 & n9227;
assign n10569 = n10330 & n12235;
assign n3706 = n10357 & n7045;
assign n5128 = ~(n2808 | n6673);
assign n1047 = ~n11474;
assign n14297 = ~(n4829 | n2660);
assign n1740 = n718 & n1970;
assign n1160 = n8452 | n11622;
assign n1660 = ~n4325;
assign n8609 = n1261 | n10028;
assign n12726 = n6111 | n8375;
assign n12555 = n1821 | n6927;
assign n4444 = n6519 | n6489;
assign n3875 = ~n5160;
assign n13566 = n1802 & n5171;
assign n14135 = ~n13560;
assign n7267 = ~n10322;
assign n306 = n5587 | n2809;
assign n13679 = n839 | n13540;
assign n7577 = ~(n5509 | n10244);
assign n6721 = ~(n7696 | n1719);
assign n2559 = n7832 & n1694;
assign n8292 = n11551 | n12851;
assign n8385 = n1576 | n9079;
assign n3870 = ~n9608;
assign n5183 = n350 & n12308;
assign n4892 = n12935 & n2746;
assign n2528 = n7079 & n2711;
assign n3317 = n6595 | n6639;
assign n11214 = n7684 | n11174;
assign n2689 = n6016 & n13965;
assign n5655 = n9423 | n5037;
assign n12037 = ~n6007;
assign n14411 = n11163 & n11760;
assign n12965 = ~(n11492 | n6189);
assign n13420 = ~n6680;
assign n12171 = n6909 | n4154;
assign n1127 = ~n5294;
assign n3889 = ~(n6030 | n13060);
assign n9536 = n8726 | n5267;
assign n8980 = ~n4891;
assign n12259 = ~n4210;
assign n6443 = ~(n14075 | n11766);
assign n12341 = n9853 & n4441;
assign n6896 = n3093 | n11799;
assign n1052 = n1202 | n3494;
assign n5040 = n7219 | n4369;
assign n4006 = n3559 | n14275;
assign n13726 = n13108 | n4281;
assign n9206 = ~n13814;
assign n3482 = n11336 & n5660;
assign n3798 = ~(n6700 | n8390);
assign n13168 = ~(n13875 | n11977);
assign n11491 = n13078 & n12557;
assign n12236 = n11867 & n4557;
assign n8356 = n3526 & n7650;
assign n7843 = ~(n7683 | n8857);
assign n7475 = ~(n10289 | n7094);
assign n11566 = ~(n12323 | n4419);
assign n7225 = n7697 | n6837;
assign n7684 = ~n382;
assign n11475 = n7057 & n493;
assign n1656 = n11262 | n8799;
assign n3200 = n11316 & n11773;
assign n9368 = n10323 | n4002;
assign n14271 = ~(n9423 | n9694);
assign n5473 = n10245 | n9710;
assign n12571 = n8453 & n10328;
assign n8601 = n12460 & n9896;
assign n8767 = ~n3765;
assign n5446 = n3164 | n3437;
assign n6507 = ~n13181;
assign n7273 = n1772 & n6175;
assign n639 = n5891 | n2981;
assign n8421 = n2025 | n5176;
assign n1945 = ~(n4424 | n13013);
assign n3805 = n3445 | n9990;
assign n11085 = n6891 | n9322;
assign n3595 = n12019 | n4462;
assign n4611 = n3766 & n4745;
assign n5394 = n8412 & n13111;
assign n13505 = ~(n1628 | n312);
assign n3265 = n8332 | n6244;
assign n13772 = n10556 & n968;
assign n2297 = n12139 | n363;
assign n11707 = n4244 & n8878;
assign n2996 = ~n14135;
assign n4588 = n9353 | n4326;
assign n9558 = n7419 & n9260;
assign n11895 = n2057 | n4030;
assign n1691 = n7430 | n12370;
assign n13646 = n1431 & n11424;
assign n4350 = n9885 & n8567;
assign n1483 = n7212 | n10569;
assign n8860 = ~(n4741 | n7512);
assign n8856 = ~n10617;
assign n3250 = n3526 & n5078;
assign n6634 = ~(n9529 | n9185);
assign n5998 = n4925 | n8279;
assign n7965 = ~(n6088 | n10554);
assign n3766 = ~n5618;
assign n10910 = n13240 & n11119;
assign n1363 = n11008 & n2433;
assign n7409 = n7284 & n13985;
assign n3180 = n309 & n8686;
assign n13341 = n1538 | n14347;
assign n698 = n4898 | n14230;
assign n6092 = n14465 & n198;
assign n6183 = n11105 | n7158;
assign n5807 = ~n2383;
assign n13848 = n11020 & n8193;
assign n2439 = n12549 | n10048;
assign n4629 = ~(n12765 | n6828);
assign n436 = n12020 | n10433;
assign n7437 = ~(n1480 | n11427);
assign n12881 = n1428 & n11786;
assign n1044 = ~n409;
assign n12251 = n13806 | n14190;
assign n8426 = n3526 & n11279;
assign n14103 = n4574 & n3838;
assign n13334 = ~(n13376 | n11209);
assign n7987 = n4300 & n7017;
assign n11117 = ~n11933;
assign n13422 = ~(n8825 | n424);
assign n12495 = n4899 | n1825;
assign n12805 = n6135 & n771;
assign n2943 = n13367 & n3745;
assign n10265 = n129 & n5232;
assign n380 = n6192 & n11004;
assign n2153 = n11303 | n2277;
assign n8734 = n5275 & n2404;
assign n11820 = n13850 & n13883;
assign n7394 = n12521 & n10168;
assign n6075 = ~(n4174 | n3528);
assign n831 = n10820 & n3884;
assign n127 = n2064 & n11794;
assign n12381 = n13525 & n12629;
assign n1800 = n227 | n3818;
assign n266 = ~(n2086 | n3239);
assign n13630 = ~(n2218 | n10014);
assign n1081 = n2082 & n13927;
assign n11564 = n6271 | n3898;
assign n5465 = n10323 | n9908;
assign n14373 = ~n11715;
assign n3260 = n10025 & n456;
assign n9484 = n7370 & n369;
assign n10722 = n12211 | n7320;
assign n8478 = n7003 | n94;
assign n1092 = ~(n8656 | n11233);
assign n12827 = ~n5980;
assign n4398 = n3886 | n1603;
assign n5262 = n8769 & n1789;
assign n13579 = n5483 | n3069;
assign n5020 = n10394 | n5345;
assign n2745 = n2518 | n54;
assign n9958 = n10338 & n1021;
assign n9006 = n9265 & n14395;
assign n7546 = n10231 & n7781;
assign n11990 = ~n5354;
assign n1316 = n13421 & n10911;
assign n7799 = ~(n12800 | n9097);
assign n8563 = n7211 & n11643;
assign n7557 = ~(n4439 | n8127);
assign n14357 = ~n7272;
assign n10422 = n6167 & n8827;
assign n8210 = ~n12746;
assign n5194 = n3247 & n542;
assign n7947 = n5071 & n1734;
assign n13023 = n12131 | n9942;
assign n2339 = n10351 | n8268;
assign n9542 = n12960 & n9261;
assign n4980 = n12500 | n1893;
assign n14334 = n8828 | n5119;
assign n8211 = n8277 | n4740;
assign n6118 = n4018 & n1560;
assign n7445 = n2006 & n9794;
assign n12278 = n5225 | n9977;
assign n10598 = n6531 & n8700;
assign n2091 = ~n11143;
assign n533 = ~n230;
assign n562 = n12100 | n8145;
assign n1323 = ~(n48 | n13009);
assign n4176 = n390 | n4867;
assign n9395 = ~(n6788 | n13669);
assign n9337 = n12986 & n12115;
assign n2621 = n3132 | n13673;
assign n9253 = ~(n8592 | n3524);
assign n12541 = n5833 | n12853;
assign n595 = n11142 & n5154;
assign n3844 = ~(n5990 | n11299);
assign n5351 = n2224 & n13184;
assign n4146 = n10079 | n11756;
assign n2951 = n13037 | n1027;
assign n2481 = n6629 | n5010;
assign n8454 = n11614 & n13617;
assign n1676 = n13426 & n9793;
assign n8347 = n2908 | n12044;
assign n519 = n6090 | n8165;
assign n467 = ~(n7004 | n8841);
assign n14022 = n13367 & n1351;
assign n7550 = n2473 & n3265;
assign n11380 = n584 | n2865;
assign n9440 = ~(n12084 | n9277);
assign n3261 = n2510 | n4143;
assign n6285 = n3126 | n6684;
assign n13411 = n1538 | n12135;
assign n5333 = ~n12084;
assign n3441 = n12455 & n1940;
assign n9679 = n2002 | n11933;
assign n5867 = n10560 | n1824;
assign n13300 = ~(n7407 | n13274);
assign n78 = n13700 & n12972;
assign n2887 = n13706 | n1363;
assign n7713 = n8427 & n1668;
assign n13818 = n4205 | n7622;
assign n389 = n2061 & n7913;
assign n4736 = n8043 & n7169;
assign n316 = ~n6426;
assign n11751 = n6537 & n5832;
assign n9003 = n13700 & n12364;
assign n9505 = n8277 | n3857;
assign n11994 = ~(n2752 | n10700);
assign n14007 = n504 | n7440;
assign n770 = n8213 & n44;
assign n8472 = n6937 | n10470;
assign n10624 = ~n10775;
assign n13703 = n4929 & n14013;
assign n5906 = n13342 & n8461;
assign n8966 = n4788 & n13998;
assign n12557 = n12576 | n1238;
assign n254 = n13656 & n131;
assign n4772 = n1125 & n13299;
assign n7141 = n11676 | n8780;
assign n5368 = ~(n11325 | n9318);
assign n5888 = n3777 | n315;
assign n5634 = ~n8486;
assign n9607 = n6730 | n9040;
assign n6687 = n2006 & n6710;
assign n13704 = n10374 & n11637;
assign n14280 = n3164 | n10422;
assign n5260 = n2784 | n8947;
assign n5265 = ~n585;
assign n13324 = ~n5333;
assign n746 = n1802 & n7184;
assign n2797 = n11503 & n6107;
assign n6158 = ~(n2218 | n1219);
assign n7265 = n1776 & n7927;
assign n12256 = n11028 & n3422;
assign n5802 = n11336 & n10052;
assign n13893 = ~(n14058 | n5513);
assign n458 = ~n4373;
assign n1865 = ~(n4284 | n4272);
assign n7493 = n9353 | n1487;
assign n4077 = n11008 & n1752;
assign n6127 = n9571 & n3051;
assign n3214 = n636 & n12171;
assign n10876 = ~(n10637 | n1945);
assign n7960 = n5475 & n12825;
assign n3010 = n1047 & n2893;
assign n6914 = ~(n48 | n1121);
assign n2531 = ~n382;
assign n709 = ~(n8592 | n1707);
assign n13211 = n839 | n11172;
assign n6123 = n12909 & n12358;
assign n5562 = ~n7600;
assign n4247 = ~(n10648 | n6582);
assign n10593 = ~n2370;
assign n6176 = n5562 | n7471;
assign n3710 = ~n871;
assign n3561 = ~n8550;
assign n515 = n8828 | n2883;
assign n14353 = n4358 & n1808;
assign n8429 = n2901 | n6761;
assign n13846 = n3370 & n910;
assign n13027 = n7359 | n5366;
assign n8544 = ~n4216;
assign n7842 = ~n8576;
assign n1748 = n11837 | n2454;
assign n1907 = n12421 & n12410;
assign n11839 = ~n1010;
assign n4890 = n4422 & n5230;
assign n12585 = n480 | n10819;
assign n7956 = n492 | n8132;
assign n10577 = n12013 & n11703;
assign n3575 = n228 | n5353;
assign n9393 = n6857 | n12606;
assign n14126 = ~(n8217 | n7661);
assign n11651 = n10309 | n2603;
assign n2081 = n4359 & n6514;
assign n2108 = n8849 & n9925;
assign n1473 = ~n5300;
assign n14131 = n1857 & n1816;
assign n7793 = n28 | n6339;
assign n13642 = n7430 | n7180;
assign n10444 = n687 & n13401;
assign n3659 = n3088 | n13651;
assign n7794 = n12461 & n13079;
assign n3293 = n6838 & n13581;
assign n7912 = ~n9371;
assign n2733 = ~(n6731 | n4059);
assign n9405 = n14227 & n8248;
assign n1495 = ~n407;
assign n13069 = ~n13458;
assign n5947 = n9650 & n5219;
assign n976 = ~n238;
assign n5417 = n12500 | n1715;
assign n5933 = n2461 & n10563;
assign n10304 = n1875 | n3700;
assign n9859 = n10871 | n6847;
assign n14448 = n687 & n10155;
assign n5516 = n5011 & n11409;
assign n2435 = n5092 & n3087;
assign n9841 = ~(n1473 | n4152);
assign n5844 = n8965 & n8012;
assign n5431 = n8238 & n7513;
assign n1315 = n12449 & n5556;
assign n11397 = n10234 | n9347;
assign n4656 = n6480 | n3263;
assign n7734 = n432 & n4588;
assign n5907 = n6697 & n14083;
assign n9911 = n7053 & n12967;
assign n13347 = n14109 & n7637;
assign n11031 = n8768 & n10202;
assign n6210 = ~(n2866 | n12736);
assign n13297 = ~n6113;
assign n4281 = n222 & n3282;
assign n2076 = n8151 | n1221;
assign n2993 = n11647 | n14089;
assign n13664 = n10449 | n4506;
assign n609 = n7997 & n7241;
assign n1372 = ~(n151 | n2688);
assign n14417 = n9297 & n436;
assign n1494 = ~n14154;
assign n1171 = n80 & n257;
assign n9969 = ~(n2016 | n7030);
assign n2540 = ~(n3445 | n9213);
assign n12920 = ~(n11489 | n13260);
assign n7921 = ~(n3882 | n13508);
assign n11671 = ~(n7245 | n8645);
assign n10141 = n4358 & n2456;
assign n7153 = ~(n13399 | n13644);
assign n13157 = n3125 | n12490;
assign n14346 = n13520 & n9588;
assign n6369 = n10309 | n14284;
assign n3354 = ~n10994;
assign n13629 = n5458 & n13653;
assign n1696 = n14351 & n12544;
assign n2101 = n12802 & n1317;
assign n13400 = ~(n11094 | n789);
assign n12118 = n1354 & n14486;
assign n284 = n163 | n707;
assign n8160 = n12543 | n5431;
assign n11203 = n7436 | n7764;
assign n10558 = n11303 | n12685;
assign n10690 = n2017 | n11027;
assign n3311 = n14373 & n2900;
assign n6663 = n9620 | n13307;
assign n610 = n10294 | n6602;
assign n1190 = n7187 & n3316;
assign n1346 = n28 | n5457;
assign n5974 = n8163 & n10801;
assign n6538 = n3169 & n14007;
assign n11274 = n12455 & n4685;
assign n2288 = n3559 | n5798;
assign n10417 = n412 | n6931;
assign n6357 = n11244 & n1881;
assign n14418 = n3888 | n774;
assign n12515 = n12449 & n6241;
assign n12931 = n8923 & n377;
assign n14264 = n1854 & n2837;
assign n10609 = ~n2967;
assign n4534 = ~n4646;
assign n12204 = n7912 | n10664;
assign n13042 = n8569 & n2713;
assign n11603 = n9620 | n14270;
assign n8487 = n8746 | n8550;
assign n9927 = ~(n12968 | n1460);
assign n5902 = ~(n8942 | n8121);
assign n1669 = ~n12394;
assign n1555 = n1701 | n6655;
assign n9161 = n10857 | n2814;
assign n7132 = n11590 & n6430;
assign n10224 = ~n8735;
assign n13977 = ~n2973;
assign n3527 = ~n2472;
assign n11673 = n3942 & n11881;
assign n805 = n3846 & n6382;
assign n2747 = ~n2484;
assign n7232 = n12018 & n4941;
assign n1254 = ~n2906;
assign n10733 = ~(n3394 | n2123);
assign n13026 = n791 | n9996;
assign n3857 = ~(n4637 | n13062);
assign n10370 = n2082 & n2683;
assign n5636 = n10089 | n2219;
assign n3883 = n4346 & n13679;
assign n11006 = n10154 | n10699;
assign n10689 = n9745 & n13417;
assign n4836 = ~(n239 | n10387);
assign n8423 = n5489 & n11035;
assign n3581 = ~(n12568 | n12010);
assign n1168 = n14150 & n572;
assign n12528 = ~n10945;
assign n13344 = n7888 | n1665;
assign n3560 = ~(n12957 | n13657);
assign n12566 = n10234 | n13328;
assign n2047 = n7212 | n3887;
assign n3450 = ~(n8021 | n8679);
assign n7060 = ~n4490;
assign n1554 = n9804 | n1720;
assign n10274 = n4033 | n2656;
assign n1138 = ~n12069;
assign n5970 = ~(n2000 | n2541);
assign n10074 = n2961 & n11295;
assign n2429 = n12461 & n3689;
assign n11579 = n2518 | n9569;
assign n12264 = n5317 & n14004;
assign n1909 = n3273 | n524;
assign n6326 = ~n6248;
assign n9118 = n8801 & n2698;
assign n4938 = n2643 & n5898;
assign n11659 = n4822 | n8029;
assign n1761 = n6867 | n3498;
assign n7641 = n2983 & n6878;
assign n7377 = ~(n8798 | n13340);
assign n5963 = n9747 | n11031;
assign n4056 = n5647 | n13343;
assign n1845 = n7700 | n7259;
assign n850 = ~n7322;
assign n3445 = ~n9580;
assign n12006 = n11240 & n4008;
assign n10346 = n12506 & n5221;
assign n1099 = n1198 | n12946;
assign n6534 = n13209 & n10697;
assign n11957 = n13537 | n8133;
assign n11670 = n10922 & n1781;
assign n8141 = n5625 | n10738;
assign n7160 = ~(n8798 | n6121);
assign n13777 = n7057 & n7545;
assign n6996 = n317 | n10689;
assign n5050 = n3923 & n6402;
assign n13652 = n5762 | n4011;
assign n10305 = ~(n11040 | n12165);
assign n1011 = ~n8204;
assign n11062 = n6537 | n9921;
assign n537 = ~(n585 | n14023);
assign n12300 = n8828 | n13205;
assign n10257 = ~(n6971 | n5573);
assign n5208 = ~(n8216 | n7925);
assign n2714 = n839 | n8208;
assign n2037 = n5641 | n1402;
assign n11708 = n12211 | n3336;
assign n2397 = n12620 & n13896;
assign n3864 = n14351 & n9681;
assign n3472 = n4821 | n3772;
assign n2189 = ~(n4135 | n7210);
assign n13083 = ~n11788;
assign n6205 = ~n13234;
assign n8975 = ~n10736;
assign n10395 = n4601 & n14249;
assign n5134 = n12324 | n4475;
assign n13343 = n12185 & n11819;
assign n4137 = n6311 & n11601;
assign n7664 = n13103 & n11037;
assign n11115 = n10647 & n7718;
assign n13310 = ~n10629;
assign n8169 = n7670 & n7495;
assign n1808 = n2747 | n8879;
assign n5274 = n781 | n726;
assign n140 = n8821 | n13895;
assign n12906 = n8183 & n7350;
assign n6573 = n3861 & n13803;
assign n11343 = n3449 & n14204;
assign n4299 = ~n10897;
assign n7726 = n1223 | n2081;
assign n6356 = n3076 | n5282;
assign n11451 = n9191 & n8883;
assign n6937 = ~n12829;
assign n7847 = n9238 & n6936;
assign n12517 = n7673 & n11952;
assign n1381 = n13236 & n927;
assign n1946 = ~n8649;
assign n8869 = n3011 | n9881;
assign n8647 = n5046 | n394;
assign n4745 = n13537 | n11032;
assign n12076 = n405 & n7490;
assign n8208 = n11495 & n5963;
assign n9968 = ~(n12403 | n199);
assign n8207 = n4876 | n7328;
assign n3418 = ~n8521;
assign n1536 = n6350 | n3591;
assign n8672 = ~n11975;
assign n4584 = n898 & n8331;
assign n4511 = n13555 & n11923;
assign n2491 = n14435 | n13490;
assign n9185 = ~(n6905 | n3414);
assign n442 = ~n3918;
assign n514 = n4018 & n10877;
assign n9437 = n12614 & n12354;
assign n13678 = n2330 & n4009;
assign n11294 = n11011 | n2389;
assign n10540 = n14227 & n4390;
assign n3073 = n3161 | n2824;
assign n7101 = n3724 & n14496;
assign n10951 = n2645 | n1770;
assign n9109 = n11503 & n2208;
assign n5641 = ~n3021;
assign n31 = ~n14134;
assign n7785 = n8147 & n3865;
assign n8057 = ~(n13248 | n1257);
assign n4549 = ~n6742;
assign n11331 = n12168 & n12192;
assign n10480 = ~(n10638 | n592);
assign n6842 = n2686 | n8011;
assign n10277 = n13698 | n10758;
assign n7954 = ~(n4682 | n8311);
assign n8062 = n10825 | n1727;
assign n6596 = ~n10204;
assign n10069 = n6067 & n4769;
assign n2136 = n3846 & n1792;
assign n13583 = n4445 & n12526;
assign n43 = n13338 & n119;
assign n6973 = n12351 | n9086;
assign n2421 = n817 | n936;
assign n9241 = n6130 & n4058;
assign n4719 = n8047 & n4158;
assign n331 = n13755 & n9978;
assign n1658 = n12149 | n166;
assign n5164 = ~(n2932 | n9408);
assign n9289 = ~n9959;
assign n10842 = n13118 | n881;
assign n3607 = ~n2497;
assign n7479 = n9931 | n2922;
assign n5953 = n10134 & n3553;
assign n12374 = n9190 & n2649;
assign n14219 = n3895 | n760;
assign n6161 = n77 | n2160;
assign n2468 = ~n11120;
assign n8749 = n8714 | n14480;
assign n11653 = n11360 | n8745;
assign n6569 = n7618 | n844;
assign n1350 = n6167 & n3229;
assign n1070 = n8768 & n7741;
assign n9598 = n10394 | n8936;
assign n5407 = n14435 | n13067;
assign n4981 = n11704 | n12477;
assign n12054 = n10461 | n11282;
assign n3061 = n889 & n3925;
assign n8480 = ~n11415;
assign n12356 = ~(n11445 | n5978);
assign n677 = n12149 | n3186;
assign n12643 = ~(n5505 | n5824);
assign n6818 = n231 & n8738;
assign n377 = n28 | n11797;
assign n12929 = n9650 & n10923;
assign n4458 = ~(n4978 | n13140);
assign n11524 = n9745 & n1810;
assign n11019 = n2888 | n1315;
assign n3310 = n12401 | n14487;
assign n2412 = ~n8735;
assign n13616 = ~(n5977 | n10029);
assign n12919 = n10247 & n2035;
assign n1704 = n11316 & n14305;
assign n5507 = ~n382;
assign n12640 = n2486 & n8411;
assign n8513 = ~n4317;
assign n4508 = ~n11055;
assign n5614 = n3365 & n12090;
assign n7150 = n1701 | n184;
assign n8805 = n4690 & n4398;
assign n1564 = n2158 & n13767;
assign n5277 = n5240 & n5446;
assign n11547 = ~n381;
assign n9753 = n4739 | n8001;
assign n984 = n10224 | n4209;
assign n9923 = n4394 & n147;
assign n4810 = n5710 | n6478;
assign n7284 = ~n13139;
assign n11699 = n8431 & n4246;
assign n4213 = ~n8572;
assign n10916 = n12130 | n2930;
assign n13986 = ~(n1383 | n7981);
assign n14076 = n14074 | n3130;
assign n2509 = n8855 & n2110;
assign n7655 = n13882 & n8214;
assign n10507 = n7852 & n14121;
assign n2749 = n12425 & n1903;
assign n10796 = n12772 & n10790;
assign n273 = n3914 | n8865;
assign n7812 = ~n622;
assign n141 = n8043 & n6766;
assign n8827 = n11231 | n9106;
assign n1340 = n309 & n14477;
assign n2019 = n2908 | n6222;
assign n13056 = n8881 | n9181;
assign n6511 = n4358 & n7948;
assign n3205 = n7812 | n1228;
assign n12754 = n12039 & n13553;
assign n5771 = n446 & n3917;
assign n414 = n6867 | n9852;
assign n1855 = ~n10750;
assign n10700 = ~(n10309 | n11155);
assign n4825 = n12622 | n2642;
assign n12502 = n11316 & n6331;
assign n4882 = n12295 | n4221;
assign n6625 = ~n3440;
assign n9002 = n4357 | n3663;
assign n952 = n10209 & n5155;
assign n1334 = n3561 & n12900;
assign n12949 = n4887 | n6054;
assign n1485 = n9229 | n13294;
assign n8448 = n1051 | n8626;
assign n2437 = n6898 & n6764;
assign n7286 = n6867 | n2718;
assign n2436 = n3125 | n7851;
assign n7396 = n5861 | n7010;
assign n11508 = ~n11453;
assign n2084 = n9113 & n1343;
assign n7100 = ~(n4174 | n12155);
assign n4543 = n12741 & n845;
assign n6475 = ~(n2236 | n3963);
assign n2227 = n6157 & n13602;
assign n907 = n12611 & n4910;
assign n11959 = n13446 | n294;
assign n7397 = n3271 & n2262;
assign n10336 = n4300 & n5870;
assign n7453 = n13016 | n12188;
assign n6373 = ~n6264;
assign n4360 = n10913 | n13028;
assign n7541 = n13236 & n9730;
assign n7355 = ~(n3132 | n12965);
assign n6641 = n5986 | n13751;
assign n8852 = n13421 & n10574;
assign n3619 = ~(n11227 | n10157);
assign n14497 = n10857 | n11219;
assign n9436 = ~(n9967 | n13249);
assign n3385 = n80 & n10149;
assign n1772 = ~n13723;
assign n510 = ~n11714;
assign n2278 = n4690 & n9954;
assign n10491 = n9490 | n3708;
assign n6189 = ~(n12112 | n12626);
assign n8858 = n769 | n1024;
assign n14084 = n12038 & n11841;
assign n8972 = n1729 & n2938;
assign n1860 = ~n1936;
assign n13096 = ~n6787;
assign n2243 = n6135 & n1358;
assign n9312 = n12592 & n13175;
assign n2445 = ~n5606;
assign n14114 = n11607 & n11774;
assign n13214 = ~(n4928 | n6914);
assign n1984 = n4484 & n6116;
assign n13684 = n103 & n11454;
assign n11424 = n11183 | n5186;
assign n11231 = ~n10069;
assign n3947 = n7187 & n12590;
assign n7530 = ~n2130;
assign n9959 = n11792 & n8115;
assign n8631 = ~n5435;
assign n13657 = ~(n900 | n1818);
assign n5181 = ~(n10803 | n5069);
assign n9325 = n976 | n11390;
assign n1602 = ~n6357;
assign n12888 = ~n4715;
assign n6448 = ~(n3182 | n5293);
assign n6124 = ~(n3290 | n828);
assign n12284 = n6706 | n3737;
assign n5126 = n8965 & n10205;
assign n12849 = n13118 | n11194;
assign n9962 = n1834 | n13820;
assign n6073 = n1481 & n14241;
assign n11075 = n10624 | n3939;
assign n13080 = ~n4325;
assign n5299 = ~(n8877 | n6501);
assign n3119 = n3011 | n7686;
assign n13644 = ~(n8378 | n803);
assign n3259 = n9490 | n12296;
assign n6524 = n12870 | n9157;
assign n2869 = n10936 | n10932;
assign n4990 = n12324 | n8917;
assign n565 = n12949 & n10239;
assign n7310 = n6595 | n12650;
assign n3938 = n8825 | n3889;
assign n11238 = n1838 | n14000;
assign n12862 = n5236 | n472;
assign n12850 = n10646 | n4282;
assign n2854 = n5634 & n13791;
assign n5004 = n13240 & n4371;
assign n14489 = n13484 & n11936;
assign n7041 = ~n12012;
assign n9490 = ~n5974;
assign n10126 = n1582 | n13946;
assign n147 = n11405 | n8447;
assign n4255 = ~n7086;
assign n8335 = n4162 | n7302;
assign n12831 = n11935 | n1405;
assign n10097 = n10516 & n11462;
assign n12618 = n2229 | n8640;
assign n6541 = n6128 & n4819;
assign n13626 = ~n4490;
assign n343 = ~(n13722 | n2610);
assign n11004 = n4967 | n8290;
assign n3287 = n3506 | n6703;
assign n7989 = n5335 & n1200;
assign n13151 = n2064 & n9497;
assign n1177 = n77 | n14001;
assign n2478 = n930 | n2437;
assign n8687 = n4468 | n5946;
assign n3916 = n9509 & n8571;
assign n1313 = n12622 | n6063;
assign n9994 = ~n1544;
assign n6263 = ~n9686;
assign n3604 = n2784 | n6320;
assign n4438 = ~(n6672 | n12643);
assign n12687 = n6965 & n359;
assign n9079 = n5229 & n9287;
assign n1598 = n11580 | n13373;
assign n11611 = n1362 | n13793;
assign n10695 = n10247 & n7084;
assign n9223 = n13297 & n6249;
assign n1616 = ~(n12866 | n842);
assign n1153 = n13005 | n6763;
assign n6539 = n6744 & n1926;
assign n11221 = n10399 & n11718;
assign n9734 = n10191 | n14417;
assign n9187 = n11722 | n13601;
assign n176 = n5491 | n5224;
assign n3371 = n5315 | n894;
assign n10005 = n10820 & n11780;
assign n10478 = n10166 & n4686;
assign n14266 = n2750 | n3969;
assign n5842 = n5940 & n6904;
assign n745 = n3777 | n4197;
assign n1870 = n11036 | n3075;
assign n106 = n687 & n11355;
assign n3996 = n12636 & n5059;
assign n6027 = n9190 & n8323;
assign n4699 = n9726 & n11731;
assign n2873 = n12202 & n8558;
assign n3957 = n13421 & n7343;
assign n5534 = n1047 & n8793;
assign n12744 = n8714 | n1407;
assign n3052 = n2682 & n10789;
assign n4102 = ~n9388;
assign n9831 = n2181 | n6545;
assign n1801 = ~n11776;
assign n5528 = n523 | n13347;
assign n14500 = ~(n14367 | n14341);
assign n8904 = n10834 | n7675;
assign n12349 = n8630 & n10537;
assign n5257 = n13720 & n13999;
assign n7436 = ~n6357;
assign n7881 = n9564 & n12402;
assign n351 = n10332 & n160;
assign n10481 = ~(n2644 | n9390);
assign n10259 = n8247 & n3995;
assign n3944 = ~n6874;
assign n6891 = ~n4325;
assign n7022 = n8701 | n9302;
assign n4852 = n7745 & n1302;
assign n713 = n4300 & n9981;
assign n2907 = n12105 & n12462;
assign n8818 = ~(n5132 | n6944);
assign n82 = ~n6055;
assign n13500 = n12226 & n4245;
assign n5964 = n6354 & n11828;
assign n12339 = n4205 | n4353;
assign n11301 = n4128 | n8468;
assign n14286 = ~n11269;
assign n12468 = n6857 | n7942;
assign n12403 = ~n2011;
assign n3795 = n4347 & n1441;
assign n10090 = n11804 | n12076;
assign n12158 = n1172 | n2136;
assign n1721 = n13240 & n11810;
assign n7572 = n14188 | n12801;
assign n9238 = ~n1955;
assign n10754 = n12990 & n2289;
assign n8085 = n8800 & n57;
assign n799 = ~n7871;
assign n13132 = ~n2334;
assign n5976 = n6690 | n8689;
assign n12648 = n3932 & n3770;
assign n6497 = n11551 | n13527;
assign n1238 = n4880 & n975;
assign n8815 = n1202 | n514;
assign n10122 = ~(n300 | n6277);
assign n10883 = ~n4744;
assign n3751 = n1391 | n5341;
assign n14044 = ~(n8856 | n32);
assign n9892 = n769 | n5964;
assign n7209 = ~(n10936 | n13266);
assign n12956 = ~(n7971 | n1382);
assign n5210 = n12935 & n2838;
assign n4739 = ~n4939;
assign n1703 = ~(n11017 | n10934);
assign n8806 = n10294 | n1374;
assign n9376 = n13147 & n9674;
assign n9483 = n4092 | n1434;
assign n620 = n4340 | n11258;
assign n699 = ~(n13811 | n2928);
assign n7855 = n11163 & n8196;
assign n11482 = ~(n2566 | n6070);
assign n2787 = n11036 | n8091;
assign n5557 = n974 | n321;
assign n14224 = n5641 | n12564;
assign n11975 = ~n179;
assign n5236 = ~n8695;
assign n6341 = n10731 | n7908;
assign n13339 = n8047 & n104;
assign n13645 = n8476 | n4678;
assign n14367 = ~n10219;
assign n5301 = n501 & n13258;
assign n3789 = ~(n8378 | n8670);
assign n8025 = ~n9456;
assign n9666 = n3923 & n8495;
assign n10397 = n9191 & n14364;
assign n362 = n8015 | n483;
assign n7218 = n14029 | n12641;
assign n11485 = n13507 & n8657;
assign n7186 = n7970 & n13954;
assign n5434 = ~n1724;
assign n9779 = ~(n1697 | n1111);
assign n431 = n13227 & n9217;
assign n10239 = n2505 & n14252;
assign n3825 = n13847 | n8271;
assign n5931 = n13537 | n3374;
assign n67 = n14110 | n8161;
assign n4823 = n2694 | n7539;
assign n13086 = n5434 & n1849;
assign n7099 = n1189 | n3267;
assign n4451 = n446 & n9339;
assign n7778 = n317 | n3535;
assign n5441 = n7015 & n763;
assign n11847 = n203 & n1065;
assign n9288 = n10562 & n645;
assign n5868 = n13485 | n6232;
assign n1599 = n5180 | n11212;
assign n13111 = n1137 | n4951;
assign n1780 = ~n13365;
assign n4635 = n2179 | n6499;
assign n773 = n9953 & n4290;
assign n9235 = n13518 | n3931;
assign n9699 = n2904 & n3794;
assign n5072 = n7219 | n5561;
assign n12817 = n6625 & n12284;
assign n2275 = n9944 & n2331;
assign n11167 = n4627 & n4217;
assign n8175 = n6654 | n6601;
assign n12010 = ~(n1742 | n2420);
assign n12776 = n1377 & n9406;
assign n10948 = n9015 & n5086;
assign n4095 = ~n13038;
assign n10940 = n11420 | n4970;
assign n10904 = n10855 & n4444;
assign n2830 = n14091 & n3208;
assign n8878 = n3914 | n2129;
assign n11955 = n14400 | n2523;
assign n6966 = ~(n8015 | n8784);
assign n8885 = ~(n12569 | n9378);
assign n7352 = ~n5354;
assign n946 = ~n1506;
assign n710 = n7596 & n6994;
assign n14522 = n3861 & n10420;
assign n14327 = ~n7507;
assign n6218 = n10534 | n4985;
assign n4188 = n2846 & n3382;
assign n12864 = n5999 & n8475;
assign n10220 = n7122 | n84;
assign n12905 = n2961 & n14221;
assign n9951 = n6167 & n3269;
assign n2599 = n1685 | n4809;
assign n13183 = n446 & n11656;
assign n4969 = n747 | n3190;
assign n5474 = n13404 & n1853;
assign n1891 = n4065 | n13559;
assign n2318 = ~n1267;
assign n8462 = ~n11188;
assign n11573 = n11048 | n14411;
assign n7358 = ~n7600;
assign n304 = ~n2040;
assign n962 = n3766 & n12647;
assign n5646 = n6343 & n9671;
assign n5811 = n14327 & n12436;
assign n1036 = n13342 & n6852;
assign n11577 = n7063 & n7859;
assign n171 = n11572 | n486;
assign n2603 = n5489 & n7874;
assign n8156 = n3766 & n61;
assign n11765 = ~n407;
assign n11092 = n687 & n12339;
assign n4761 = n13362 & n1554;
assign n8907 = ~n1265;
assign n11455 = ~n11743;
assign n8354 = n1821 | n4890;
assign n10247 = ~n11969;
assign n5156 = n13413 | n2604;
assign n2776 = n5137 & n12051;
assign n4567 = n10705 & n9983;
assign n3094 = ~n14332;
assign n11816 = ~n920;
assign n12574 = n4614 & n11002;
assign n11542 = ~n4609;
assign n424 = ~(n12191 | n2540);
assign n5573 = ~(n12888 | n8751);
assign n14149 = n13252 & n2678;
assign n2388 = n13147 & n4010;
assign n905 = n3527 | n9024;
assign n10688 = n4154 | n3506;
assign n13461 = n6205 | n11377;
assign n12871 = n10072 & n855;
assign n3336 = n7068 & n11107;
assign n6103 = n12521 & n7570;
assign n1786 = n4508 | n2291;
assign n2167 = n7810 & n8712;
assign n524 = n8066 & n12692;
assign n1894 = n2226 & n10395;
assign n722 = n14449 | n9527;
assign n2463 = n11484 & n4356;
assign n10003 = n9541 | n4442;
assign n7705 = n428 & n13737;
assign n11151 = n4895 | n8780;
assign n2434 = ~(n5468 | n4133);
assign n893 = n7912 | n8754;
assign n11148 = ~n11809;
assign n11870 = ~n10172;
assign n8983 = ~n2545;
assign n3141 = n10166 & n14350;
assign n13097 = ~(n6044 | n11291);
assign n4205 = ~n6978;
assign n7240 = n1660 | n12236;
assign n1767 = ~(n12075 | n14310);
assign n10381 = n85 | n429;
assign n11041 = ~(n7223 | n8286);
assign n9336 = n7736 | n12036;
assign n12185 = ~n11715;
assign n778 = n13310 | n11500;
assign n9821 = n13875 | n11109;
assign n6148 = n10822 & n7367;
assign n11947 = n7187 & n11359;
assign n7432 = ~(n7011 | n11000);
assign n13623 = n4821 | n12408;
assign n7325 = n4255 | n12438;
assign n1883 = n14188 | n5338;
assign n6463 = n7219 | n2873;
assign n4657 = ~n10469;
assign n8704 = ~n9546;
assign n7917 = n11803 & n1422;
assign n3204 = ~n5429;
assign n12425 = ~n9456;
assign n6710 = n817 | n5045;
assign n1188 = n3093 | n3433;
assign n6616 = n8726 | n10633;
assign n10749 = n2064 & n14492;
assign n1867 = n11814 & n13368;
assign n12282 = n541 & n2161;
assign n9940 = n7551 | n10682;
assign n1094 = n6555 & n3296;
assign n13252 = ~n10469;
assign n460 = n8569 & n10590;
assign n4365 = ~n10112;
assign n9538 = n8816 | n6295;
assign n11015 = n6318 & n3595;
assign n6675 = n4908 | n4976;
assign n4648 = n12019 | n224;
assign n8712 = n12568 | n5687;
assign n11648 = n10302 & n11104;
assign n5852 = ~n11441;
assign n12943 = n8025 & n3657;
assign n10240 = n5548 | n8910;
assign n10579 = n6711 | n8660;
assign n12283 = ~(n5132 | n1703);
assign n13313 = ~(n6971 | n8154);
assign n4315 = n8849 & n8149;
assign n233 = n1685 | n1587;
assign n10396 = ~n9306;
assign n9825 = n14166 | n5799;
assign n7598 = n501 & n7845;
assign n10020 = n2473 & n10662;
assign n13970 = n4484 | n8746;
assign n4193 = n3932 & n7406;
assign n9618 = ~n14433;
assign n806 = n478 | n8668;
assign n12946 = n8702 & n1205;
assign n10539 = ~n4847;
assign n11683 = n1613 | n6741;
assign n11478 = n14430 | n1740;
assign n5746 = n6128 & n358;
assign n208 = n2025 | n6083;
assign n7885 = n14110 | n10243;
assign n10357 = ~n9613;
assign n827 = ~n4711;
assign n7247 = n9742 | n6186;
assign n14158 = n1805 | n5608;
assign n2908 = ~n2383;
assign n5593 = n11737 & n4264;
assign n13201 = ~n11606;
assign n5024 = ~n13012;
assign n7804 = ~(n3873 | n3789);
assign n1635 = n14401 | n7295;
assign n9291 = ~n749;
assign n5079 = n12023 | n14036;
assign n12446 = n4929 & n5955;
assign n854 = n5857 & n37;
assign n13953 = n11158 & n3177;
assign n8571 = n5491 | n11859;
assign n10229 = ~n10975;
assign n7366 = n4739 | n12089;
assign n10819 = n1662 & n9361;
assign n9234 = n10449 | n2596;
assign n6763 = n98 & n11483;
assign n8996 = n5472 | n9076;
assign n456 = n1059 | n5033;
assign n14139 = ~n9516;
assign n7456 = n12015 & n3965;
assign n13202 = n4199 | n9063;
assign n13615 = n5582 & n6977;
assign n6473 = n1805 | n6661;
assign n3674 = n5064 | n12161;
assign n13148 = ~(n13941 | n13997);
assign n12935 = ~n11474;
assign n2567 = n5807 | n5844;
assign n11978 = n9564 & n5976;
assign n2306 = n6695 | n868;
assign n14282 = ~n10108;
assign n6803 = n8581 | n11363;
assign n13501 = ~n7819;
assign n6277 = ~(n573 | n3951);
assign n4528 = n7745 & n13370;
assign n14492 = n5587 | n13105;
assign n6716 = n9490 | n9542;
assign n4535 = ~n10423;
assign n4494 = n4468 | n9504;
assign n8653 = n2272 | n9955;
assign n3792 = n4347 & n14205;
assign n9430 = n7862 | n6532;
assign n10953 = ~n1222;
assign n12644 = ~n4341;
assign n5550 = n5046 & n1616;
assign n8151 = ~n2383;
assign n11672 = n10089 | n11367;
assign n2552 = n974 | n2413;
assign n12235 = n5180 | n2258;
assign n10322 = ~n6516;
assign n4847 = n11966 & n5839;
assign n14277 = n5315 | n3373;
assign n11436 = n12615 & n5470;
assign n5233 = n2747 | n8108;
assign n11264 = n1409 & n12103;
assign n8697 = ~n9583;
assign n11788 = n2029 & n7842;
assign n10296 = n5936 | n14055;
assign n6085 = ~n10069;
assign n13174 = n4354 & n1379;
assign n12333 = n6744 & n6442;
assign n3181 = n3526 & n9556;
assign n205 = n10556 & n2638;
assign n12768 = ~n656;
assign n11073 = ~(n5762 | n330);
assign n7270 = n14401 | n7257;
assign n14200 = ~n2061;
assign n13873 = n5732 | n6467;
assign n4266 = ~n11426;
assign n3778 = n13518 | n10153;
assign n13107 = ~n1571;
assign n11086 = n13356 | n8647;
assign n1221 = n2783 & n7558;
assign n4524 = ~(n6971 | n7921);
assign n9783 = n12265 & n6438;
assign n694 = n1875 | n7907;
assign n1304 = ~(n10730 | n13910);
assign n5125 = n13407 & n2847;
assign n6585 = n13338 & n7497;
assign n2737 = n9229 | n9502;
assign n10309 = ~n4203;
assign n1937 = ~n9456;
assign n2398 = ~(n7905 | n5703);
assign n14279 = n13433 & n6490;
assign n101 = ~(n10571 | n9513);
assign n14374 = n2422 & n9585;
assign n2296 = n3952 & n9268;
assign n13349 = n1362 | n11886;
assign n7198 = n5362 | n1514;
assign n7850 = n7957 & n13621;
assign n8890 = n3485 & n14068;
assign n11190 = n11362 & n4894;
assign n5887 = n4195 | n908;
assign n295 = n13675 | n1655;
assign n4342 = n13814 | n4022;
assign n2187 = n7584 | n3248;
assign n10744 = n11679 & n14220;
assign n8032 = n12351 | n13304;
assign n4163 = ~n1760;
assign n3386 = n10166 & n13450;
assign n4644 = n1172 | n8440;
assign n5810 = ~(n9035 | n3139);
assign n406 = ~n82;
assign n10564 = n4156 & n6827;
assign n4314 = n6471 | n7117;
assign n10353 = ~(n194 | n14362);
assign n5777 = n7888 | n11342;
assign n5899 = ~n871;
assign n10320 = n2878 | n395;
assign n3114 = n13885 | n7762;
assign n8295 = n2510 | n7992;
assign n11112 = ~(n7905 | n10907);
assign n1886 = n1904 & n5482;
assign n4925 = ~n6804;
assign n13932 = n976 | n9982;
assign n3732 = n3755 & n2514;
assign n6969 = n8512 & n6616;
assign n9696 = n2367 & n7333;
assign n8963 = ~n1861;
assign n7476 = ~n13882;
assign n5782 = ~n8419;
assign n14095 = n12500 | n7159;
assign n5751 = n8581 | n2438;
assign n3427 = ~n9640;
assign n9677 = n12167 | n2699;
assign n2902 = n7011 | n5447;
assign n10628 = n4581 & n11272;
assign n2848 = ~n6422;
assign n2183 = ~(n3234 | n5755);
assign n5912 = ~(n1178 | n3359);
assign n10092 = n4877 | n12177;
assign n3685 = ~(n6020 | n13528);
assign n11807 = n10713 | n4136;
assign n3762 = ~n2895;
assign n7485 = n6090 | n1269;
assign n2965 = n6471 | n990;
assign n4758 = n13489 & n8710;
assign n5411 = n6724 & n8843;
assign n13197 = n9269 | n12041;
assign n2985 = ~n442;
assign n9070 = n5348 & n487;
assign n10351 = ~n1267;
assign n6132 = ~(n5480 | n8628);
assign n6766 = n4923 | n5276;
assign n5957 = ~(n3290 | n9668);
assign n89 = ~n9306;
assign n7264 = n7116 | n3203;
assign n3653 = n2229 | n2550;
assign n6821 = n4562 | n1002;
assign n9865 = ~n8565;
assign n8140 = n5315 | n10392;
assign n4354 = ~n4618;
assign n7108 = n8748 | n7729;
assign n4689 = n2111 | n7088;
assign n1073 = n14006 | n4785;
assign n14410 = n4163 & n5113;
assign n1370 = n4244 & n7883;
assign n2267 = n2783 & n6694;
assign n3908 = n7596 & n12251;
assign n9904 = n12038 & n4485;
assign n8636 = n13310 | n10528;
assign n2303 = n13107 & n12470;
assign n2670 = n11033 & n5296;
assign n333 = ~n7681;
assign n134 = n5409 | n9760;
assign n7512 = ~(n13937 | n14028);
assign n11248 = n1602 | n9749;
assign n1884 = n1258 | n11795;
assign n3598 = n5489 & n9610;
assign n682 = n5033 & n101;
assign n4361 = n14063 & n13268;
assign n13624 = n2322 & n6756;
assign n8028 = n4757 & n7453;
assign n4660 = n9102 & n7247;
assign n5136 = n13755 & n5444;
assign n863 = n12130 | n9410;
assign n6313 = ~n496;
assign n7700 = ~n3681;
assign n12224 = n4973 & n2655;
assign n14310 = ~(n7200 | n4759);
assign n2614 = n172 | n2261;
assign n10871 = ~n3357;
assign n14339 = n6649 & n6253;
assign n1987 = n12449 & n10659;
assign n7426 = ~n7404;
assign n6231 = n13575 & n10499;
assign n2321 = n8025 & n9082;
assign n5065 = ~n9863;
assign n7997 = ~n9893;
assign n5285 = n3512 | n7175;
assign n2222 = n7419 & n8141;
assign n12873 = n13501 | n4553;
assign n6360 = n7249 | n7383;
assign n368 = n14337 | n2668;
assign n8078 = n3276 & n3661;
assign n7506 = n4289 & n9025;
assign n14343 = n11153 & n8600;
assign n6551 = ~(n4296 | n6365);
assign n7564 = n11581 | n2776;
assign n8104 = ~(n11151 | n6408);
assign n3737 = n501 & n6561;
assign n13529 = n2486 & n11944;
assign n10837 = n5184 | n8635;
assign n12802 = ~n7278;
assign n5070 = n5562 | n8566;
assign n10668 = ~n11305;
assign n12884 = n89 | n13333;
assign n7200 = ~n6305;
assign n11453 = ~n1342;
assign n14317 = n12169 | n13345;
assign n555 = ~n409;
assign n6606 = ~n10303;
assign n10735 = n480 | n1872;
assign n11798 = n1610 & n13321;
assign n9601 = ~n11574;
assign n11093 = ~n6975;
assign n11723 = n11816 & n11965;
assign n8602 = n7421 & n1594;
assign n6153 = n9953 & n5044;
assign n2114 = n8714 | n1398;
assign n10580 = n1728 | n4391;
assign n10660 = ~n14483;
assign n14359 = n4790 & n2680;
assign n495 = n8358 & n4061;
assign n13965 = n6039 | n4121;
assign n10565 = ~(n2355 | n13116);
assign n7477 = n7250 | n5140;
assign n2967 = n8975 | n10945;
assign n7091 = ~n11001;
assign n9304 = n10019 | n10606;
assign n2804 = ~n8780;
assign n8443 = ~(n12292 | n11078);
assign n6426 = ~n9757;
assign n2935 = n2983 & n7778;
assign n7121 = n13226 | n3787;
assign n1522 = ~n4415;
assign n11362 = ~n14163;
assign n10082 = ~(n8543 | n2431);
assign n9637 = ~(n3445 | n10447);
assign n3018 = n3161 | n5110;
assign n4127 = n8393 & n8921;
assign n7066 = ~(n5132 | n247);
assign n7561 = n12620 & n3460;
assign n14449 = ~n4203;
assign n1434 = n12832 & n10634;
assign n6240 = n8569 & n979;
assign n11420 = ~n10629;
assign n13712 = n706 & n13831;
assign n1502 = n8950 & n9937;
assign n2500 = n7015 & n433;
assign n8857 = ~(n9818 | n2317);
assign n12472 = ~n8223;
assign n9531 = n8950 & n3038;
assign n12173 = n11804 | n5428;
assign n2121 = n2281 & n1346;
assign n968 = n6857 | n12551;
assign n12007 = n12986 & n3781;
assign n5053 = ~n9865;
assign n5822 = n2180 & n11516;
assign n8512 = ~n5504;
assign n4855 = n10396 | n935;
assign n12901 = n3097 & n10903;
assign n5878 = n10300 | n5705;
assign n13718 = ~n1833;
assign n4395 = n4631 | n5739;
assign n5192 = ~(n329 | n4309);
assign n2116 = n10457 & n3463;
assign n1393 = ~(n5621 | n11681);
assign n1678 = ~n13908;
assign n4470 = n3904 & n7095;
assign n13502 = n4690 & n10816;
assign n11706 = ~n9406;
assign n14480 = n7421 & n2558;
assign n217 = n317 | n6683;
assign n8740 = n12994 | n7002;
assign n9522 = n7245 | n4243;
assign n13627 = ~n14134;
assign n9650 = ~n2906;
assign n675 = n974 | n836;
assign n5329 = n10062 | n12258;
assign n5979 = n12576 | n11169;
assign n3495 = n8816 | n9572;
assign n12543 = ~n6123;
assign n7527 = ~n3357;
assign n4433 = ~n1027;
assign n13071 = n4481 | n5050;
assign n12560 = n4435 | n10967;
assign n2729 = ~n12168;
assign n626 = n6531 & n3389;
assign n9445 = n3435 & n13588;
assign n5609 = n1254 & n11150;
assign n1877 = n9323 & n6312;
assign n4837 = n1339 & n12468;
assign n13548 = n406 & n6623;
assign n14369 = n5628 & n3056;
assign n4573 = ~n11756;
assign n13098 = n13850 & n1099;
assign n9693 = n2445 & n11437;
assign n4046 = ~n10917;
assign n13060 = ~(n3445 | n11543);
assign n11212 = n4098 & n11835;
assign n1259 = n10399 & n9027;
assign n4723 = n2949 | n13613;
assign n3229 = n6085 | n10949;
assign n14107 = ~n2545;
assign n4744 = n14360 | n8598;
assign n10831 = n10626 | n3159;
assign n9711 = n5647 | n8755;
assign n6256 = ~n7282;
assign n6844 = n14245 | n4292;
assign n10570 = n1539 & n14413;
assign n5900 = n1582 | n4772;
assign n8877 = ~n3681;
assign n2586 = n10399 & n5138;
assign n6315 = ~(n14075 | n3462);
assign n5671 = n11542 | n9933;
assign n2212 = ~n11453;
assign n1807 = n9188 & n5858;
assign n6346 = n1854 & n2532;
assign n10706 = n11360 | n8890;
assign n7073 = n5023 & n6210;
assign n4926 = n10560 | n5571;
assign n2678 = n3546 | n287;
assign n13355 = n2897 | n1370;
assign n11715 = ~n5117;
assign n7314 = n7079 & n144;
assign n13467 = ~n3976;
assign n5761 = n4527 & n13434;
assign n13717 = n12858 & n12063;
assign n6328 = n5139 | n12828;
assign n665 = ~(n2462 | n8868);
assign n6918 = ~(n14011 | n7069);
assign n7353 = n4741 | n11844;
assign n7331 = n7211 & n11651;
assign n14099 = n4525 & n11831;
assign n3620 = n3877 | n1331;
assign n13158 = ~n10973;
assign n9928 = n1031 | n12026;
assign n11686 = n9898 & n4583;
assign n13631 = n4876 | n10902;
assign n348 = ~n11854;
assign n10256 = n10399 & n2696;
assign n470 = n14419 | n5612;
assign n8045 = ~n3046;
assign n7208 = ~n3402;
assign n518 = n11047 | n14199;
assign n579 = n1255 & n11570;
assign n2373 = n9323 & n13202;
assign n11642 = n504 | n12245;
assign n4287 = ~(n1771 | n1390);
assign n1806 = ~(n4313 | n4654);
assign n2349 = n3365 & n469;
assign n10952 = ~(n1697 | n8730);
assign n3715 = ~n3356;
assign n4597 = n1140 & n11744;
assign n11298 = n8908 | n12617;
assign n10618 = n1697 | n7054;
assign n4559 = n14430 | n10908;
assign n7566 = n12802 & n890;
assign n4767 = n9807 | n13481;
assign n11045 = n10300 | n13987;
assign n716 = n5815 | n9581;
assign n5162 = n5948 & n8806;
assign n14153 = n406 & n10327;
assign n1764 = n2461 & n12210;
assign n10119 = n103 & n12962;
assign n10590 = n504 | n7641;
assign n1768 = n4045 | n14086;
assign n6510 = n5180 | n14099;
assign n2040 = n9819 & n10900;
assign n5106 = n3099 | n3752;
assign n13018 = n2669 & n154;
assign n13121 = n3526 & n8287;
assign n11443 = n7693 & n6676;
assign n2299 = n10357 & n8913;
assign n2750 = ~n1041;
assign n9268 = n5480 | n13697;
assign n5698 = n2401 | n9053;
assign n13357 = n2562 | n7165;
assign n9553 = ~(n1693 | n14130);
assign n8801 = ~n12930;
assign n8393 = ~n5951;
assign n13552 = n4486 & n663;
assign n5956 = ~(n2727 | n1046);
assign n13477 = ~n10985;
assign n1982 = n2099 & n13920;
assign n887 = ~n30;
assign n2774 = n3370 & n10962;
assign n5275 = ~n10376;
assign n4454 = n4445 & n3133;
assign n8192 = n13531 | n5455;
assign n630 = n4036 & n5549;
assign n12133 = ~(n4656 | n5398);
assign n11956 = n782 | n10958;
assign n1195 = n3365 & n13786;
assign n2354 = ~n11765;
assign n11837 = ~n8926;
assign n10306 = ~(n3944 | n13964);
assign n4759 = ~(n11901 | n3879);
assign n983 = n11090 | n3851;
assign n6708 = n3401 & n219;
assign n5765 = n7529 & n10058;
assign n272 = n12226 & n3112;
assign n12797 = n4574 & n13436;
assign n688 = n12990 & n2601;
assign n4546 = ~n8048;
assign n4950 = n5936 | n1879;
assign n3002 = n6263 | n1941;
assign n2269 = ~n2946;
assign n13016 = ~n14154;
assign n8219 = n2089 | n7936;
assign n13827 = n116 | n7563;
assign n12984 = n12968 | n8777;
assign n547 = n6781 | n1482;
assign n12471 = n3125 | n2463;
assign n12701 = n11814 & n14263;
assign n1614 = n6466 | n11633;
assign n13485 = ~n11415;
assign n14248 = ~(n11232 | n4984);
assign n7452 = ~(n3640 | n2150);
assign n7583 = n7677 & n3375;
assign n407 = n6849 & n5166;
assign n10102 = n13745 & n4151;
assign n13173 = n10710 & n2037;
assign n8785 = n1481 & n6860;
assign n10340 = ~(n12527 | n12700);
assign n6705 = ~n6466;
assign n2295 = n10822 & n7442;
assign n261 = ~n4500;
assign n4071 = n5710 | n8326;
assign n3362 = n12038 & n4302;
assign n2330 = ~n1436;
assign n4032 = n6753 & n1253;
assign n11487 = n7060 & n2292;
assign n218 = n10825 | n1807;
assign n9463 = n9113 & n4168;
assign n13487 = n2058 & n11070;
assign n6264 = n13012 & n8345;
assign n3085 = n4180 | n6671;
assign n1379 = n1669 | n4448;
assign n941 = n4095 & n11430;
assign n8533 = n1914 | n12052;
assign n1179 = n12870 | n13969;
assign n5424 = n4908 | n9257;
assign n2663 = ~(n500 | n8573);
assign n10209 = ~n9924;
assign n1470 = n2246 | n2756;
assign n945 = n8983 | n12899;
assign n142 = ~(n9136 | n310);
assign n9397 = n2387 | n13717;
assign n11726 = n3628 | n4175;
assign n1969 = n3755 & n12896;
assign n843 = n8300 & n7882;
assign n7421 = ~n10975;
assign n5059 = n10660 | n14303;
assign n8405 = n79 & n8693;
assign n473 = ~n13408;
assign n12059 = n309 & n7619;
assign n2720 = n8043 & n8724;
assign n9885 = ~n11548;
assign n13068 = n8513 | n1515;
assign n12937 = n4267 & n8498;
assign n9340 = ~n398;
assign n6900 = n4844 & n985;
assign n7573 = n12092 & n9271;
assign n4632 = n6711 | n8061;
assign n7538 = ~(n12254 | n3610);
assign n2828 = n10166 & n14471;
assign n5688 = n5317 & n14067;
assign n4569 = n10822 & n3114;
assign n1361 = ~n8073;
assign n8600 = n2272 | n9783;
assign n3781 = n4741 | n12230;
assign n1297 = n11816 & n10066;
assign n934 = n3132 | n8759;
assign n5754 = n5815 | n13694;
assign n12126 = n5640 | n12614;
assign n2550 = n12802 & n13652;
assign n1273 = n13489 & n9485;
assign n14268 = n5562 | n4377;
assign n4914 = n14449 | n318;
assign n6244 = n5475 & n8399;
assign n4206 = n11607 & n3525;
assign n12894 = n100 | n3837;
assign n6944 = ~(n911 | n5469);
assign n6520 = n1776 | n13102;
assign n1634 = n6205 | n12267;
assign n8591 = ~(n10715 | n651);
assign n6423 = ~(n14198 | n5368);
assign n3814 = n10589 & n7264;
assign n5702 = n1946 & n1705;
assign n11272 = n10383 | n3988;
assign n2469 = n13806 | n9467;
assign n12362 = n2877 | n14331;
assign n3823 = ~(n1178 | n11410);
assign n11520 = n5279 & n3489;
assign n10193 = n13236 & n14418;
assign n8346 = n457 & n7956;
assign n3564 = n1610 & n11164;
assign n9583 = ~n13593;
assign n2870 = n12100 | n7092;
assign n1192 = n7700 | n6636;
assign n5007 = ~n10069;
assign n9858 = n2820 & n9366;
assign n546 = n10351 | n9736;
assign n1376 = n12611 & n8004;
assign n8144 = n8780 & n6897;
assign n10877 = n10309 | n1847;
assign n10957 = n1258 | n1531;
assign n4663 = ~(n6426 | n6567);
assign n10567 = n10015 & n11591;
assign n5259 = n6595 | n11589;
assign n1737 = n10936 | n78;
assign n11997 = n13130 | n9131;
assign n8640 = n7970 & n7615;
assign n14404 = ~n2918;
assign n803 = ~(n6018 | n10653);
assign n10867 = n8066 & n4630;
assign n6009 = n10302 & n3128;
assign n1956 = n5011 & n51;
assign n2779 = n14058 | n14426;
assign n4935 = n6527 & n8203;
assign n13847 = ~n3021;
assign n13084 = ~n8656;
assign n8515 = n4790 & n4189;
assign n2734 = n6703 & n11805;
assign n13553 = n3569 | n12915;
assign n8320 = n8300 & n9483;
assign n2371 = n494 & n12111;
assign n8107 = n12695 | n14141;
assign n522 = ~(n7011 | n11994);
assign n3965 = n2857 | n5239;
assign n2748 = n7156 | n12498;
assign n14265 = n10302 & n12343;
assign n1814 = n3204 & n2755;
assign n7204 = n6130 & n4532;
assign n13821 = n4788 & n2789;
assign n3600 = n718 & n14233;
assign n6554 = n12933 | n5502;
assign n13370 = n1628 | n8464;
assign n13676 = ~n6975;
assign n6881 = n14321 & n13926;
assign n5197 = ~n1861;
assign n14058 = ~n4606;
assign n3439 = ~(n7940 | n1501);
assign n12063 = n5562 | n4051;
assign n13139 = ~n3544;
assign n5681 = n5012 & n7793;
assign n11016 = n4601 | n14483;
assign n7930 = n6288 | n14429;
assign n10568 = ~n10239;
assign n3586 = ~n10303;
assign n4069 = n2709 & n2450;
assign n2024 = ~(n8629 | n1513);
assign n734 = n7211 & n12420;
assign n9587 = n494 | n11345;
assign n1591 = n1266 & n5466;
assign n10801 = n1920 & n13968;
assign n6747 = ~n13230;
assign n3410 = ~(n13021 | n8483);
assign n5482 = n1538 | n3803;
assign n4986 = n8453 & n9005;
assign n1970 = n12130 | n11646;
assign n3970 = ~(n3434 | n7314);
assign n4144 = ~n11412;
assign n5704 = n7670 & n5769;
assign n11931 = n11569 & n658;
assign n11696 = n5918 & n9831;
assign n12764 = ~n9371;
assign n4230 = n6192 & n10151;
assign n10710 = ~n5675;
assign n2926 = n13252 & n5686;
assign n7979 = n13840 | n10630;
assign n10745 = n11580 | n13101;
assign n12718 = ~(n1677 | n10567);
assign n6065 = n536 & n9364;
assign n1621 = n3126 | n667;
assign n13910 = ~(n7229 | n1712);
assign n11954 = n79 & n5478;
assign n242 = n8393 & n8835;
assign n6565 = ~(n8592 | n1392);
assign n6499 = n2709 & n5831;
assign n5925 = n2246 | n3197;
assign n7305 = n8250 & n10827;
assign n7722 = n7678 | n9600;
assign n12448 = n748 & n5751;
assign n12120 = ~(n6743 | n6457);
assign n4357 = ~n1966;
assign n3252 = ~(n9414 | n8829);
assign n7386 = ~(n5833 | n5937);
assign n9890 = ~n12970;
assign n10201 = n1548 | n2009;
assign n417 = n14358 & n4724;
assign n11162 = n8747 | n7705;
assign n6870 = n13707 | n5326;
assign n7807 = n954 | n765;
assign n6079 = n6957 & n4605;
assign n11403 = ~n7660;
assign n6489 = n7053 & n4882;
assign n11164 = n10234 | n3504;
assign n5940 = ~n3440;
assign n6805 = n5252 & n4335;
assign n646 = ~n11861;
assign n12650 = n2006 & n8654;
assign n7192 = ~n1421;
assign n6110 = n5940 & n6360;
assign n14372 = n12857 & n9594;
assign n13472 = n5012 & n6869;
assign n9097 = n10247 & n4869;
assign n6869 = n9140 | n2956;
assign n9976 = n4180 | n13381;
assign n8539 = n1820 | n1591;
assign n7813 = n1729 & n2363;
assign n13462 = n11300 & n3474;
assign n3774 = ~(n9924 | n4064);
assign n6456 = ~(n11980 | n3145);
assign n8955 = n309 & n12124;
assign n9799 = ~(n1628 | n7742);
assign n11317 = n6389 & n7;
assign n8435 = n7736 | n13727;
assign n8775 = n3586 & n13856;
assign n4375 = ~(n448 | n14246);
assign n10482 = n1623 | n6125;
assign n6400 = ~(n14166 | n1791);
assign n12820 = ~n12249;
assign n12238 = ~(n14455 | n10344);
assign n11550 = n3125 | n6073;
assign n5056 = n4978 | n7206;
assign n10860 = n14466 | n3181;
assign n8702 = ~n14367;
assign n8241 = n10166 & n4726;
assign n8022 = n80 & n11700;
assign n12930 = ~n7915;
assign n9517 = n6625 & n109;
assign n11066 = n7818 | n5014;
assign n8621 = ~(n12311 | n10180);
assign n11116 = ~(n6397 | n13193);
assign n4216 = ~n11428;
assign n1325 = n2908 | n1841;
assign n7633 = n6595 | n995;
assign n5594 = n9856 | n4230;
assign n2287 = n9151 | n12805;
assign n7810 = ~n2619;
assign n8709 = n3276 & n6506;
assign n7838 = n4698 | n394;
assign n5085 = n3755 & n9929;
assign n6776 = n6525 & n7176;
assign n13232 = n3923 & n8105;
assign n5471 = ~n10177;
assign n4406 = n14029 | n4842;
assign n3897 = n11679 & n1684;
assign n5491 = ~n5627;
assign n4402 = n4876 | n13007;
assign n11906 = n11285 | n6296;
assign n6704 = n10289 | n4563;
assign n7983 = n12057 & n9362;
assign n9794 = n13155 | n11304;
assign n10822 = ~n10322;
assign n10759 = n2942 & n9413;
assign n359 = n3043 & n4601;
assign n8244 = n898 & n9325;
assign n13549 = n13531 | n13172;
assign n2238 = n10933 | n11623;
assign n10762 = n5252 & n14387;
assign n2410 = n9174 | n8253;
assign n8263 = n7116 | n4446;
assign n7098 = n10960 | n11559;
assign n4420 = n7462 | n12906;
assign n13560 = n14357 & n12272;
assign n2191 = ~(n7364 | n186);
assign n6828 = ~(n12117 | n3199);
assign n3976 = n1801 | n10912;
assign n3420 = n12034 | n11257;
assign n11191 = n8372 & n13392;
assign n12759 = ~n9878;
assign n687 = ~n12503;
assign n4840 = ~n10889;
assign n10934 = ~(n1844 | n4503);
assign n2903 = n13854 | n6348;
assign n2087 = ~n8288;
assign n12161 = n5553 & n684;
assign n12926 = n5432 | n10858;
assign n267 = n5695 | n13465;
assign n9818 = ~n13047;
assign n8673 = n12169 | n1960;
assign n9132 = n2857 | n4240;
assign n13290 = n1602 | n14269;
assign n156 = n2058 & n5481;
assign n10291 = n11315 | n13743;
assign n1566 = n766 | n14394;
assign n1927 = n8737 & n7252;
assign n11571 = n2761 | n4501;
assign n12695 = ~n11813;
assign n4418 = n13572 & n13654;
assign n5392 = ~(n4978 | n740);
assign n10109 = ~(n2889 | n7536);
assign n13739 = n4828 | n13286;
assign n8066 = ~n1911;
assign n8333 = n2099 & n797;
assign n10382 = n14388 & n5052;
assign n11022 = n8969 | n10694;
assign n14043 = n8151 | n9523;
assign n3637 = n10820 & n4519;
assign n13832 = n9375 | n1586;
assign n12497 = n5562 | n9056;
assign n13592 = n8965 & n2039;
assign n11459 = ~n81;
assign n4560 = n7076 | n3232;
assign n10215 = n13407 & n11579;
assign n7875 = n3765 & n5149;
assign n11281 = n3546 | n13076;
assign n14204 = n1361 & n303;
assign n440 = n5132 | n14267;
assign n5042 = ~n3461;
assign n7362 = ~n8106;
assign n5458 = ~n5525;
assign n9178 = n3785 & n8295;
assign n6652 = n12324 | n10152;
assign n2684 = ~n4216;
assign n1175 = n12622 | n1030;
assign n4792 = ~(n648 | n1672);
assign n2327 = n12935 & n121;
assign n6343 = ~n12930;
assign n8920 = ~n4007;
assign n9645 = n1904 & n2511;
assign n13971 = n11722 | n9463;
assign n3012 = n14321 & n2096;
assign n2950 = ~(n9657 | n3670);
assign n2300 = n6046 | n13802;
assign n3802 = ~n9350;
assign n3966 = n9190 & n7537;
assign n9287 = n8304 | n11335;
assign n9359 = ~(n6326 | n12749);
assign n2090 = ~n74;
assign n4793 = ~(n7056 | n2871);
assign n10845 = n7229 | n10632;
assign n9338 = n1193 & n11948;
assign n12453 = ~n12088;
assign n3862 = n13338 & n11383;
assign n2097 = n11674 & n1915;
assign n787 = ~n3506;
assign n11924 = ~(n648 | n1509);
assign n10185 = n14260 & n9012;
assign n4260 = n9226 | n655;
assign n8193 = n10626 | n1629;
assign n8568 = n2709 & n9899;
assign n4674 = n4614 & n5198;
assign n8256 = n2098 | n1871;
assign n8130 = n9265 & n7849;
assign n7507 = ~n13544;
assign n1091 = n11636 & n1725;
assign n4818 = ~(n13977 | n9087);
assign n3188 = n976 | n7070;
assign n3505 = n11510 | n823;
assign n628 = n9272 & n12694;
assign n2344 = ~(n3959 | n10456);
assign n302 = ~(n9546 | n13996);
assign n1198 = ~n9686;
assign n12890 = n4481 | n6076;
assign n8844 = n1198 | n12517;
assign n4041 = n13080 | n11853;
assign n9685 = ~(n5904 | n8970);
assign n12533 = ~n12117;
assign n619 = ~n4609;
assign n9960 = n77 | n3387;
assign n12292 = ~n12106;
assign n10848 = ~(n11094 | n9458);
assign n6036 = n8007 & n11698;
assign n5352 = n9984 | n14240;
assign n247 = ~(n1813 | n10321);
assign n12352 = n6706 | n1622;
assign n7025 = n3097 & n10482;
assign n9567 = ~n11302;
assign n12494 = ~n6804;
assign n2517 = n3424 & n5632;
assign n10946 = n9541 | n108;
assign n11864 = n12844 | n5168;
assign n14510 = ~n3577;
assign n7520 = n6354 & n2535;
assign n9751 = ~n4248;
assign n2702 = n4923 | n9903;
assign n4620 = n4561 | n9810;
assign n9076 = n7670 & n12317;
assign n9290 = n13464 & n1424;
assign n5995 = n3126 | n3597;
assign n4666 = n6311 & n10844;
assign n10589 = ~n8048;
assign n3194 = n7436 | n8641;
assign n1144 = n8575 | n3725;
assign n3954 = n6625 & n5223;
assign n10737 = ~(n573 | n8006);
assign n1203 = ~n2674;
assign n2394 = n14260 & n12541;
assign n2304 = n9742 | n1133;
assign n13237 = n3607 & n10;
assign n2929 = ~(n9557 | n9215);
assign n2843 = ~n1966;
assign n12914 = n4898 | n11673;
assign n7463 = n10871 | n11314;
assign n9087 = ~(n5569 | n3305);
assign n8114 = n13407 & n5547;
assign n2470 = ~n1473;
assign n2542 = n8480 | n10943;
assign n10687 = n8183 & n10064;
assign n177 = ~n3652;
assign n9920 = ~n2889;
assign n6178 = n14366 | n2214;
assign n852 = ~(n3882 | n5250);
assign n2254 = n9422 | n14084;
assign n5749 = n523 | n7884;
assign n2270 = n1788 & n10296;
assign n5344 = n965 & n768;
assign n10933 = ~n4720;
assign n1733 = ~(n13310 | n11024);
assign n353 = n12576 | n6487;
assign n9391 = n12494 | n2957;
assign n11430 = n13485 | n9445;
assign n7236 = n14465 & n2466;
assign n4927 = n14109 & n4669;
assign n3614 = n12918 & n2046;
assign n8152 = n8250 & n10489;
assign n12308 = n10059 | n5225;
assign n926 = n1255 & n6233;
assign n193 = n3193 | n10436;
assign n11051 = ~(n6039 | n1185);
assign n3488 = ~(n9618 | n5577);
assign n11385 = n6023 | n13814;
assign n3886 = ~n4149;
assign n7718 = n6373 | n11274;
assign n7648 = n12759 | n9966;
assign n10977 = ~n13437;
assign n1107 = ~(n10479 | n14026);
assign n5240 = ~n11969;
assign n13680 = n14337 | n10345;
assign n2377 = n13083 | n3629;
assign n975 = n6695 | n13098;
assign n11973 = n6263 | n4362;
assign n11328 = ~n11345;
assign n2969 = ~n5001;
assign n4905 = n3877 | n13548;
assign n7482 = n11674 & n10612;
assign n9974 = n10626 | n6618;
assign n14347 = n4581 & n13951;
assign n13609 = n5764 & n6168;
assign n12443 = n9716 | n2862;
assign n14145 = ~n3428;
assign n6192 = ~n3440;
assign n8913 = n9541 | n741;
assign n13938 = n11379 | n4839;
assign n2664 = ~(n2729 | n12515);
assign n12694 = ~n12097;
assign n12104 = n2877 | n6225;
assign n6706 = ~n10889;
assign n8399 = n1844 | n10676;
assign n4556 = n1383 | n2104;
assign n4598 = n5471 & n5305;
assign n6113 = ~n5631;
assign n8111 = ~n2958;
assign n13333 = n10072 & n9050;
assign n3888 = ~n11152;
assign n8179 = n8812 | n12012;
assign n7 = n9229 | n8380;
assign n11923 = n3815 | n11211;
assign n1400 = n11510 | n11699;
assign n2173 = n1223 | n7581;
assign n7195 = n10668 & n2362;
assign n4301 = n1854 & n7776;
assign n9999 = n10589 & n10841;
assign n2833 = n1044 | n2221;
assign n11216 = n4033 | n6036;
assign n13980 = ~(n11251 | n9292);
assign n13539 = n3675 | n12321;
assign n11052 = n1946 | n5950;
assign n11503 = ~n6765;
assign n6955 = n3276 & n12095;
assign n10527 = n5764 & n3301;
assign n12103 = n5188 & n22;
assign n4263 = n12229 & n2592;
assign n263 = ~n4154;
assign n1016 = n4261 & n6414;
assign n9215 = ~(n14370 | n13894);
assign n6910 = n6486 & n4638;
assign n5364 = ~(n9984 | n12865);
assign n5312 = ~n13139;
assign n12635 = n6957 & n7861;
assign n9227 = n5468 | n4974;
assign n13672 = ~(n3546 | n3272);
assign n3585 = n2510 | n3195;
assign n10031 = n10383 | n4077;
assign n2901 = ~n11788;
assign n2499 = n4899 | n12048;
assign n4013 = n791 | n13008;
assign n3131 = n9509 & n10703;
assign n6149 = n747 | n2670;
assign n2818 = n2089 | n1878;
assign n6540 = n1140 & n8976;
assign n2392 = n2857 | n1919;
assign n3817 = n10512 & n1508;
assign n1633 = n9198 & n7505;
assign n4650 = ~n13561;
assign n11340 = n13310 | n4892;
assign n5653 = n5229 & n6330;
assign n2978 = n1962 & n13056;
assign n5049 = n1711 | n6287;
assign n4269 = n11621 | n8707;
assign n9549 = n8983 | n8157;
assign n5813 = n5468 | n9351;
assign n5948 = ~n9950;
assign n14192 = n13118 | n11460;
assign n2291 = n9564 & n13685;
assign n5753 = n7057 & n11983;
assign n10136 = ~n751;
assign n9000 = n8748 | n13556;
assign n6560 = n4276 & n259;
assign n8163 = n8112 | n13231;
assign n5067 = n3914 | n10215;
assign n9244 = n7803 | n10656;
assign n10423 = n2474 & n8311;
assign n9502 = n4018 & n3352;
assign n1261 = ~n3616;
assign n1874 = n13362 & n5522;
assign n321 = n7810 & n3836;
assign n7395 = n12209 | n13224;
assign n3733 = n3277 & n9998;
assign n10853 = n3076 | n10169;
assign n10873 = n1198 | n4558;
assign n357 = n13547 | n13169;
assign n6561 = n12764 | n13151;
assign n1963 = n2669 & n12781;
assign n12988 = ~(n14524 | n5177);
assign n14050 = n8697 & n3840;
assign n8252 = ~n8463;
assign n13289 = n1526 & n7885;
assign n10380 = n6981 & n13566;
assign n4111 = n14042 & n5073;
assign n6250 = n9885 & n10756;
assign n11512 = ~(n6062 | n13443);
assign n645 = n11510 | n10264;
assign n287 = ~(n10091 | n12119);
assign n10195 = n13516 | n2347;
assign n14329 = n7700 | n2665;
assign n4110 = ~(n1522 | n13306);
assign n747 = ~n12489;
assign n70 = n5823 & n11889;
assign n8249 = ~(n1378 | n3148);
assign n9084 = n4932 & n8815;
assign n7458 = n1254 & n10056;
assign n6689 = n13464 & n11502;
assign n8006 = ~(n1575 | n3089);
assign n793 = n3923 & n3327;
assign n11285 = ~n9453;
assign n419 = n7684 | n6645;
assign n13409 = n12018 & n14137;
assign n364 = n1137 | n1551;
assign n3158 = ~(n7418 | n297);
assign n2010 = ~(n10280 | n1530);
assign n12068 = n3120 | n7623;
assign n8015 = ~n1894;
assign n6690 = ~n6332;
assign n11735 = n1383 | n10717;
assign n12549 = ~n2383;
assign n2923 = ~n10801;
assign n14243 = ~(n2236 | n1595);
assign n8392 = n10035 | n4294;
assign n5584 = n10767 & n10530;
assign n439 = n10357 & n3693;
assign n9823 = n4346 & n2886;
assign n7631 = ~(n12200 | n1756);
assign n13473 = n11818 | n1561;
assign n8201 = ~(n7364 | n8691);
assign n13738 = n2686 | n1717;
assign n105 = n12730 & n11139;
assign n7763 = n13147 & n1000;
assign n2934 = n11016 & n3875;
assign n12184 = n12404 & n4338;
assign n5179 = n7026 & n8429;
assign n11560 = ~(n13627 | n6565);
assign n5107 = n12401 | n8485;
assign n9570 = n4172 & n1107;
assign n5039 = n12601 | n10524;
assign n11819 = n8517 | n4528;
assign n1209 = n4631 | n2134;
assign n3797 = ~(n3019 | n10542);
assign n11886 = n10622 & n6289;
assign n8679 = n10332 & n192;
assign n5565 = n11636 & n9702;
assign n3313 = ~n4991;
assign n1349 = n12918 & n4826;
assign n663 = n11315 | n12594;
assign n2260 = n7418 | n11442;
assign n5932 = ~(n2731 | n6298);
assign n12832 = ~n12757;
assign n4108 = ~(n9807 | n12936);
assign n9267 = n8393 & n833;
assign n14516 = n14029 | n4467;
assign n9159 = n8096 | n1173;
assign n13448 = n9198 & n10961;
assign n1747 = n10083 | n4721;
assign n2646 = ~(n7887 | n3156);
assign n11857 = n7430 | n10680;
assign n14174 = ~(n4424 | n8153);
assign n5768 = n9804 | n1227;
assign n5913 = n11569 & n14484;
assign n4126 = n2006 & n2421;
assign n14331 = n5926 & n3319;
assign n1829 = n5144 | n4804;
assign n8313 = n6085 | n2107;
assign n6213 = n2412 | n8805;
assign n7346 = ~n14406;
assign n11825 = n1431 & n2819;
assign n9198 = ~n3402;
assign n11379 = ~n565;
assign n11077 = n10083 | n5580;
assign n4984 = ~(n8557 | n5756);
assign n12655 = n9275 & n2593;
assign n13749 = n4244 & n7672;
assign n10103 = n8111 & n775;
assign n3658 = ~(n2597 | n6677);
assign n2245 = ~(n1262 | n2947);
assign n4638 = n11580 | n12748;
assign n6190 = n14404 | n9850;
assign n1285 = n5710 | n7995;
assign n10217 = n12759 | n3154;
assign n7542 = n10332 & n2112;
assign n1880 = n5088 & n13711;
assign n8409 = n3942 & n9462;
assign n12052 = n9102 & n12657;
assign n8958 = n6205 | n3855;
assign n8229 = n8213 & n8539;
assign n18 = ~(n13707 | n580);
assign n4684 = ~n12746;
assign n9781 = n5710 | n95;
assign n2413 = n7810 & n12890;
assign n1532 = n9269 | n8078;
assign n1003 = n10512 | n6873;
assign n1647 = n8714 | n2210;
assign n10597 = ~(n4535 | n14290);
assign n3050 = n1613 | n11270;
assign n12600 = n13096 & n3662;
assign n13133 = n5312 & n13785;
assign n12045 = n9724 & n3031;
assign n278 = n12025 & n123;
assign n4067 = n8817 | n5184;
assign n7666 = n13112 | n12367;
assign n2209 = ~(n6122 | n4093);
assign n9611 = n10619 & n2001;
assign n2803 = n2694 | n3432;
assign n8341 = n7818 & n9792;
assign n1021 = n7358 | n5890;
assign n13904 = n10332 & n9244;
assign n3755 = ~n6119;
assign n732 = n1231 & n6691;
assign n14486 = n2179 | n8960;
assign n796 = n12335 & n12360;
assign n754 = n13806 | n5358;
assign n8695 = n13900 & n931;
assign n11309 = ~n14219;
assign n5656 = n12229 & n8673;
assign n128 = n13103 & n11530;
assign n8884 = n9008 | n8002;
assign n1311 = n8907 & n11490;
assign n7277 = ~(n194 | n1246);
assign n14025 = n13875 | n1468;
assign n1790 = ~(n8527 | n14500);
assign n2356 = n10331 | n8120;
assign n5693 = n8881 | n3588;
assign n11352 = n7026 & n2023;
assign n10923 = n3025 | n7445;
assign n4681 = n5459 & n3974;
assign n11419 = n12615 & n7706;
assign n997 = n3485 & n8652;
assign n8664 = n2082 & n11894;
assign n13607 = n1775 & n2903;
assign n4020 = n9353 | n13804;
assign n3958 = ~n1268;
assign n14311 = ~(n8816 | n3557);
assign n3497 = ~n7676;
assign n7123 = n10624 | n12338;
assign n10851 = n10367 & n10356;
assign n9219 = n7810 & n1471;
assign n2812 = n200 & n10494;
assign n4249 = n1117 & n4044;
assign n13279 = ~(n11558 | n6833);
assign n1333 = n9920 & n12437;
assign n3764 = n13096 & n14244;
assign n443 = n6654 | n2538;
assign n4457 = n5823 & n10216;
assign n8994 = n1006 | n349;
assign n4052 = ~n1060;
assign n3327 = n11379 | n6224;
assign n14201 = n2318 | n11365;
assign n1873 = n12139 | n6410;
assign n5587 = ~n12874;
assign n8536 = n3559 | n11475;
assign n4594 = n5807 | n6588;
assign n2681 = n3062 | n12504;
assign n10402 = ~n12088;
assign n8407 = ~(n1299 | n379);
assign n11652 = n13847 | n10783;
assign n10642 = n12832 & n10956;
assign n4294 = n4359 & n5310;
assign n6422 = n11842 | n1222;
assign n12653 = n6323 | n14165;
assign n13438 = ~(n9078 | n10401);
assign n11327 = n13246 & n8783;
assign n703 = ~n6844;
assign n10045 = n11231 | n14035;
assign n1797 = n11814 & n12187;
assign n2202 = n4502 & n9985;
assign n1541 = n8172 | n5869;
assign n704 = n5507 | n5644;
assign n8330 = ~(n14332 | n3146);
assign n6897 = ~(n10883 | n7857);
assign n1014 = n3667 | n8824;
assign n6646 = ~(n11546 | n12008);
assign n5209 = ~n9236;
assign n2780 = ~n10864;
assign n3157 = n3212 & n10016;
assign n5283 = n4788 & n10575;
assign n7736 = ~n11813;
assign n12586 = n5489 & n5094;
assign n14401 = ~n14412;
assign n13318 = n14472 | n158;
assign n3943 = n5312 & n11181;
assign n7688 = n8034 | n6396;
assign n7179 = ~n2951;
assign n10431 = ~(n12097 | n11490);
assign n192 = n11420 | n11682;
assign n8758 = n7670 & n4999;
assign n7944 = n12633 | n4112;
assign n4390 = n647 | n8366;
assign n7827 = n10922 & n12794;
assign n4899 = ~n11541;
assign n8148 = n2791 & n2137;
assign n4278 = ~(n2016 | n9560);
assign n601 = n333 & n13664;
assign n3663 = n6354 & n2833;
assign n5762 = ~n7441;
assign n1326 = n11163 & n5393;
assign n12546 = n4791 | n7335;
assign n4096 = ~(n9078 | n8359);
assign n7387 = n2942 & n12263;
assign n10608 = n4788 & n7174;
assign n240 = n69 | n10970;
assign n4409 = ~(n7887 | n9614);
assign n12679 = n5088 & n3281;
assign n3296 = ~(n14139 | n4132);
assign n11058 = n5229 & n8661;
assign n9305 = ~n885;
assign n10057 = n5779 & n866;
assign n11504 = n5062 & n3682;
assign n5190 = n3942 & n10092;
assign n9498 = ~(n2868 | n14488);
assign n9512 = n9984 | n5957;
assign n3904 = ~n12888;
assign n8522 = n7068 & n8782;
assign n9722 = n10374 & n7047;
assign n4608 = ~n12086;
assign n14257 = n6350 | n5;
assign n12439 = n7419 & n12616;
assign n4202 = n12651 | n13715;
assign n9102 = ~n11548;
assign n10594 = n2682 & n9130;
assign n14461 = ~n8424;
assign n8076 = n11011 | n4295;
assign n2119 = n9198 & n761;
assign n6643 = n6937 & n5256;
assign n9037 = ~(n11990 | n14520);
assign n10290 = ~(n10428 | n2943);
assign n9323 = ~n5613;
assign n2242 = n10854 & n1199;
assign n5489 = ~n13360;
assign n2549 = n4791 | n6784;
assign n11916 = ~(n3768 | n11371);
assign n5775 = n8908 | n2240;
assign n5585 = ~(n2236 | n8158);
assign n11466 = n13641 & n6129;
assign n12102 = n1559 | n5077;
assign n4964 = n9864 | n2169;
assign n7580 = ~(n4572 | n928);
assign n4466 = n4346 & n7766;
assign n5847 = ~n11966;
assign n751 = n4716 & n11938;
assign n3464 = ~(n2241 | n5076);
assign n1037 = n12494 | n9038;
assign n3610 = ~(n13477 | n3466);
assign n10406 = ~n7575;
assign n11028 = ~n11232;
assign n14425 = n227 | n13090;
assign n10631 = n11614 & n384;
assign n12678 = ~(n5065 | n12637);
assign n9500 = n5137 & n913;
assign n387 = ~n10985;
assign n10524 = n536 & n11084;
assign n4405 = n1193 & n10181;
assign n2338 = n4925 | n10673;
assign n2322 = ~n5675;
assign n2272 = ~n11813;
assign n12575 = n11867 & n3679;
assign n7532 = n10815 & n5055;
assign n8284 = n7678 | n8568;
assign n4862 = n9315 & n13634;
assign n6197 = n8300 & n9492;
assign n11273 = n2310 & n9187;
assign n5204 = n1728 | n13695;
assign n12941 = n11316 & n3692;
assign n12271 = n12712 | n6563;
assign n13639 = n12927 & n1744;
assign n1084 = n13404 & n12894;
assign n2112 = n7803 | n10804;
assign n110 = n3132 | n3797;
assign n4997 = n11157 & n7773;
assign n2952 = ~(n2154 | n11946);
assign n8990 = n11839 | n9867;
assign n453 = ~(n6933 | n4536);
assign n5856 = n7308 | n14464;
assign n14162 = n9853 & n632;
assign n13773 = n11804 | n6322;
assign n6717 = n8517 | n5907;
assign n529 = n11839 | n12969;
assign n13379 = ~n5795;
assign n6350 = ~n5974;
assign n9709 = n6609 & n4399;
assign n13994 = n11300 & n11554;
assign n4322 = n1489 & n12680;
assign n6799 = n8210 | n7413;
assign n12110 = n12998 & n10809;
assign n6618 = n12335 & n6037;
assign n12225 = n9353 | n3224;
assign n10694 = n12038 & n92;
assign n7222 = n1117 & n13884;
assign n6154 = n2518 | n1294;
assign n80 = ~n13723;
assign n13460 = n9724 & n3747;
assign n3046 = n3542 & n2850;
assign n13681 = ~(n4195 | n6141);
assign n4129 = n14373 & n3741;
assign n8068 = n13363 & n5956;
assign n8065 = ~n6159;
assign n12319 = n7249 | n5301;
assign n11841 = n4239 | n11476;
assign n5147 = n4104 & n883;
assign n566 = n14481 | n7220;
assign n12773 = n12042 & n12880;
assign n9651 = n7677 & n13943;
assign n5859 = n11724 | n3850;
assign n11496 = ~(n12112 | n8504);
assign n4273 = n6167 & n6223;
assign n5362 = ~n10069;
assign n10133 = ~(n10649 | n10876);
assign n6590 = ~(n2742 | n9652);
assign n6608 = n13781 & n6727;
assign n6598 = n3268 & n5121;
assign n1547 = n12615 & n599;
assign n11389 = n4033 | n7486;
assign n8329 = n2310 & n8274;
assign n13741 = n4276 & n12257;
assign n821 = n8247 & n893;
assign n8019 = n5253 | n1991;
assign n2791 = n14252 | n4755;
assign n8290 = n5348 & n2712;
assign n1738 = n4340 | n13048;
assign n6780 = n7427 & n12233;
assign n8628 = ~(n12197 | n9115);
assign n11049 = n954 | n10141;
assign n11131 = ~(n3922 | n6449);
assign n5495 = n504 | n591;
assign n13425 = n9494 & n13116;
assign n258 = n13421 & n8219;
assign n13227 = ~n5871;
assign n9998 = n13698 | n9379;
assign n7393 = n225 & n12536;
assign n13740 = ~(n7589 | n5098);
assign n1184 = n6090 | n8758;
assign n5294 = ~n9818;
assign n13778 = n4692 & n2964;
assign n14194 = n116 | n9060;
assign n4959 = ~(n7352 | n6817);
assign n13486 = n10062 | n14033;
assign n9988 = n7430 | n128;
assign n10214 = n14227 & n7780;
assign n6193 = ~n5438;
assign n4645 = ~(n12075 | n2663);
assign n3466 = ~(n3210 | n3421);
assign n1523 = n8969 | n8894;
assign n8436 = n6157 & n5917;
assign n6943 = n7943 & n7604;
assign n12431 = ~(n7887 | n1033);
assign n1006 = ~n1676;
assign n4762 = n13446 | n3055;
assign n3448 = n10705 & n7749;
assign n7675 = n13745 & n3472;
assign n112 = n11157 & n12792;
assign n12886 = ~n7115;
assign n13225 = n13464 & n11085;
assign n12461 = ~n1784;
assign n5718 = ~(n11305 | n8999);
assign n13326 = n14465 & n9148;
assign n8517 = ~n1220;
assign n13568 = n7043 & n8669;
assign n7375 = ~n11967;
assign n502 = n12421 & n8797;
assign n2107 = n12990 & n13396;
assign n3877 = ~n9169;
assign n12606 = n8950 & n301;
assign n3339 = n2583 & n6610;
assign n4742 = ~n10529;
assign n7681 = ~n3280;
assign n11417 = n12683 & n1837;
assign n7957 = ~n9450;
assign n2073 = n13659 | n12926;
assign n12423 = ~(n474 | n12045);
assign n8871 = n9864 | n7769;
assign n5201 = n390 | n3773;
assign n11883 = n5825 & n944;
assign n11810 = n7551 | n2176;
assign n1335 = n1489 & n14223;
assign n755 = n12625 | n5169;
assign n8198 = n14260 & n598;
assign n4445 = ~n13003;
assign n3776 = n11852 | n13000;
assign n8537 = n11738 | n2615;
assign n11483 = n5575 | n6745;
assign n12835 = n782 | n6894;
assign n3901 = n12573 & n11538;
assign n7166 = n2318 | n11447;
assign n4386 = n5647 | n13243;
assign n6059 = n2055 | n5544;
assign n7909 = ~n9416;
assign n10723 = ~(n5209 | n12286);
assign n4105 = n2061 | n9186;
assign n598 = n1006 | n11670;
assign n5318 = n2236 | n6474;
assign n2886 = n6206 | n3179;
assign n2758 = ~n10377;
assign n11799 = n5312 & n10211;
assign n3865 = n9289 | n14518;
assign n13085 = ~(n717 | n11079);
assign n11535 = ~(n10323 | n2115);
assign n8984 = ~(n6907 | n522);
assign n4414 = n11163 & n5787;
assign n9750 = n13537 | n1171;
assign n824 = n5253 | n5384;
assign n1118 = n3099 | n6642;
assign n14342 = n10560 | n12939;
assign n2523 = n14260 & n12756;
assign n2041 = n4953 | n13055;
assign n2719 = n6607 | n11330;
assign n3874 = ~(n8301 | n3937);
assign n10326 = n9803 & n13091;
assign n341 = ~(n12904 | n11624);
assign n9319 = n4988 | n5816;
assign n9038 = n2473 & n6916;
assign n3389 = n4925 | n11381;
assign n4250 = n1660 | n4453;
assign n2579 = ~(n1462 | n11096);
assign n7175 = n12531 & n13888;
assign n4839 = n9345 & n6770;
assign n9050 = n10294 | n1529;
assign n310 = n11676 & n10232;
assign n762 = n9226 | n5992;
assign n3352 = n9140 | n3598;
assign n224 = n2180 & n3790;
assign n1015 = n4239 | n12895;
assign n5258 = n10062 | n5269;
assign n6399 = n2224 & n9689;
assign n8162 = ~n13154;
assign n13780 = ~n4270;
assign n8666 = n12821 | n999;
assign n8680 = n12935 & n1608;
assign n1233 = n6167 & n1925;
assign n2981 = n231 & n4504;
assign n3629 = n5899 & n3852;
assign n12174 = n14373 & n11284;
assign n6794 = ~n10858;
assign n1628 = ~n11541;
assign n12297 = n3088 | n7467;
assign n12399 = n10245 | n11136;
assign n8824 = n7063 & n4074;
assign n5742 = n11440 | n3948;
assign n10170 = n555 | n9167;
assign n12669 = n12414 | n207;
assign n9098 = n5891 | n874;
assign n3510 = ~(n6039 | n1327);
assign n478 = ~n3455;
assign n1165 = n11687 | n12336;
assign n10228 = n327 & n7067;
assign n1595 = ~(n9046 | n10548);
assign n4878 = n14435 | n14379;
assign n4218 = ~(n2098 | n5597);
assign n3753 = n627 & n1995;
assign n9660 = n10289 | n1158;
assign n9169 = n7521 & n12279;
assign n4404 = ~n3804;
assign n11489 = ~n8162;
assign n14101 = ~(n584 | n5540);
assign n8387 = n11909 | n11333;
assign n10514 = n6039 | n5370;
assign n6936 = n3512 | n13966;
assign n14235 = n1193 & n346;
assign n5909 = n12934 | n2640;
assign n6410 = n6343 & n14335;
assign n911 = ~n13206;
assign n1262 = ~n93;
assign n14423 = n392 & n3630;
assign n1723 = n1539 & n8335;
assign n12569 = ~n264;
assign n11889 = n12622 | n7222;
assign n8181 = n3536 & n10250;
assign n8976 = n14370 | n8117;
assign n13768 = n11814 & n14405;
assign n2129 = n4261 & n1206;
assign n8743 = n766 | n10087;
assign n2127 = n5472 | n2743;
assign n8545 = n4357 | n7969;
assign n6823 = n10710 & n3167;
assign n9263 = n817 | n7616;
assign n9167 = n11679 & n2849;
assign n8159 = n13432 | n10125;
assign n8793 = n6519 | n7231;
assign n11024 = ~(n2005 | n2191);
assign n4099 = n8692 & n11186;
assign n2044 = ~(n2684 | n12670);
assign n10192 = ~(n1262 | n11903);
assign n6952 = n13109 & n12761;
assign n12736 = n2669 & n7628;
assign n5245 = n5459 & n12109;
assign n7914 = ~n2934;
assign n792 = ~(n14198 | n7806);
assign n5783 = n333 & n10583;
assign n13416 = n1962 & n5389;
assign n7196 = n7076 | n5419;
assign n5379 = n14435 | n3311;
assign n5898 = n12211 | n2792;
assign n2735 = n13863 & n87;
assign n2216 = n7812 | n13162;
assign n14432 = n678 & n1217;
assign n5567 = n7530 | n12699;
assign n2200 = n3168 | n1453;
assign n9581 = n79 & n1119;
assign n7790 = n584 | n527;
assign n12135 = n1526 & n1556;
assign n14400 = ~n12444;
assign n13925 = n10062 | n13815;
assign n14142 = n2486 & n10333;
assign n9764 = n648 | n4579;
assign n8339 = n7250 | n9735;
assign n3292 = n12683 & n1496;
assign n2891 = n12147 & n11341;
assign n8646 = n1428 & n7933;
assign n705 = ~(n8378 | n4773);
assign n8707 = n8923 & n13523;
assign n10866 = n13531 | n13848;
assign n5135 = n14400 | n12624;
assign n779 = n13501 | n6835;
assign n7774 = n782 | n4418;
assign n5506 = n747 | n1564;
assign n14272 = n3169 & n7949;
assign n8451 = ~n5300;
assign n4606 = n10282 & n7065;
assign n10663 = ~(n11998 | n8548);
assign n6728 = n8111 & n2264;
assign n7514 = n457 & n6293;
assign n5037 = n3247 & n9877;
assign n2900 = n12211 | n2741;
assign n10123 = n4544 | n5892;
assign n12813 = n13520 & n5330;
assign n6875 = ~(n7683 | n5720);
assign n13426 = n7523 | n10573;
assign n10212 = n9113 & n5777;
assign n8583 = n4445 & n1209;
assign n2130 = n1073 & n6806;
assign n1693 = ~n2577;
assign n6958 = n4877 | n9192;
assign n432 = ~n7275;
assign n13246 = ~n1784;
assign n9284 = ~(n10323 | n8441);
assign n11160 = n8358 & n6637;
assign n4443 = ~n9977;
assign n4159 = n4856 & n441;
assign n8414 = n12460 & n9859;
assign n921 = n10234 | n13574;
assign n14283 = n7798 | n4659;
assign n6912 = n10309 | n13956;
assign n2486 = ~n6975;
assign n6662 = n5491 | n4126;
assign n9580 = n6096 & n2910;
assign n9255 = n8147 & n3018;
assign n14098 = n1962 & n9360;
assign n10836 = n8980 | n2204;
assign n4436 = n12159 & n3622;
assign n3896 = n7693 & n733;
assign n5493 = ~n7819;
assign n14023 = n4650 & n1260;
assign n14434 = ~(n13365 | n7601);
assign n6292 = n4255 | n8079;
assign n9128 = n1254 & n6872;
assign n13217 = n1147 | n14175;
assign n366 = n11121 | n12719;
assign n12389 = ~n13723;
assign n7975 = n4065 | n2720;
assign n3602 = ~n6159;
assign n8484 = n1047 & n754;
assign n7825 = n11404 & n10317;
assign n1345 = n7909 & n6632;
assign n2653 = n12211 | n4815;
assign n1134 = n5234 | n9171;
assign n4412 = n7911 & n2759;
assign n7357 = n6350 | n1376;
assign n11012 = n14109 & n2513;
assign n8437 = n5472 | n6777;
assign n13032 = n8210 | n9835;
assign n6997 = ~(n13477 | n9768);
assign n11528 = n6109 | n1620;
assign n5001 = ~n12483;
assign n11858 = n4627 & n12029;
assign n12216 = n4486 & n10745;
assign n8402 = n4098 & n698;
assign n4306 = n8582 | n45;
assign n4296 = ~n9537;
assign n8603 = ~(n2087 | n8586);
assign n5545 = n12918 & n3100;
assign n480 = ~n2794;
assign n13386 = n4162 | n11207;
assign n9460 = n8047 & n12078;
assign n11554 = n8986 | n13683;
assign n3319 = n13276 | n12318;
assign n9181 = n10374 & n8749;
assign n12633 = ~n2130;
assign n8238 = ~n7507;
assign n7969 = n5999 & n11564;
assign n8575 = ~n751;
assign n10044 = n12625 | n13730;
assign n8757 = n4205 | n3201;
assign n12947 = n3366 | n11842;
assign n6702 = ~(n10973 | n11449);
assign n5000 = n5899 & n6716;
assign n10887 = n3800 | n7532;
assign n8266 = n7888 | n4037;
assign n10661 = n12404 & n9928;
assign n2062 = ~(n10285 | n13273);
assign n1734 = n10154 | n6746;
assign n9864 = ~n9371;
assign n12641 = n4657 & n11281;
assign n6260 = ~n7667;
assign n7782 = n2942 & n8699;
assign n6442 = n8726 | n11947;
assign n6017 = n6373 | n5047;
assign n2518 = ~n751;
assign n9134 = n5904 | n9461;
assign n14451 = n13080 | n11400;
assign n9096 = n6680 & n3541;
assign n14028 = ~(n9035 | n1393);
assign n2693 = n6243 & n6102;
assign n3540 = n889 & n778;
assign n11014 = n8034 | n6060;
assign n3847 = n1728 | n11352;
assign n3431 = n10330 & n13428;
assign n3588 = n10374 & n593;
assign n10024 = ~n13668;
assign n13348 = n4739 | n2940;
assign n6493 = n3826 | n11421;
assign n12717 = n13885 | n13164;
assign n7651 = n9289 | n4691;
assign n8578 = ~(n900 | n13163);
assign n9145 = n5475 & n807;
assign n9694 = ~(n10280 | n5945);
assign n2411 = n3062 | n9531;
assign n6671 = n8569 & n9471;
assign n11314 = n14213 & n12991;
assign n6051 = ~n2644;
assign n9230 = ~n2472;
assign n9692 = n6111 | n1540;
assign n2207 = n4255 | n10728;
assign n2763 = n7677 & n2197;
assign n11646 = n4627 & n5070;
assign n6664 = n2547 & n12603;
assign n6167 = ~n1436;
assign n12511 = n8697 & n14334;
assign n12609 = n10647 & n13726;
assign n12625 = ~n12687;
assign n3401 = ~n9994;
assign n2764 = ~(n2651 | n12860);
assign n8881 = ~n14412;
assign n12061 = n13108 | n12679;
assign n10164 = n12741 & n5812;
assign n2789 = n49 | n3680;
assign n1993 = n9509 & n13239;
assign n691 = n10396 | n2891;
assign n11695 = ~(n3521 | n18);
assign n5271 = ~n3583;
assign n6378 = n3435 & n11612;
assign n8373 = n283 | n10413;
assign n7551 = ~n1833;
assign n10083 = ~n9878;
assign n10712 = ~n7402;
assign n13669 = ~(n11558 | n8417);
assign n11575 = n11008 & n13036;
assign n3435 = ~n6990;
assign n6038 = n10763 & n5298;
assign n10967 = n2758 & n657;
assign n12504 = n1678 & n669;
assign n7152 = n9830 & n13278;
assign n8184 = n930 | n10987;
assign n3474 = n5084 | n12255;
assign n13235 = ~(n7238 | n2544);
assign n13770 = n9507 | n11357;
assign n11826 = n286 & n4388;
assign n7990 = n2422 & n7792;
assign n8945 = n8569 & n3505;
assign n3008 = n7041 | n12976;
assign n5729 = n7779 & n9144;
assign n7233 = n9080 & n1747;
assign n10025 = ~n4755;
assign n9899 = n10224 | n7126;
assign n644 = n4354 & n14251;
assign n12741 = ~n7278;
assign n2378 = ~n12084;
assign n1827 = n394 & n6184;
assign n5241 = n11093 & n8019;
assign n753 = n986 & n13418;
assign n10085 = n1266 & n7636;
assign n2708 = n12100 | n12299;
assign n2002 = ~n9154;
assign n4073 = n11123 | n7795;
assign n12487 = n2082 & n12659;
assign n4861 = n4602 | n6631;
assign n4977 = n13297 & n3668;
assign n7801 = ~(n4742 | n2617);
assign n12040 = ~n9156;
assign n2049 = n8034 | n4918;
assign n9669 = n5647 | n7503;
assign n2577 = ~n2889;
assign n3882 = ~n9604;
assign n8485 = n457 & n12703;
assign n13958 = ~(n13276 | n11482);
assign n7076 = ~n9453;
assign n397 = n432 & n12225;
assign n10260 = n5857 & n12305;
assign n13488 = n1876 & n10732;
assign n8345 = n14273 & n7216;
assign n9702 = n4807 | n9709;
assign n8105 = n695 | n5130;
assign n6366 = n9571 & n1659;
assign n648 = ~n12331;
assign n4630 = n7462 | n10687;
assign n2424 = ~(n2057 | n5883);
assign n12460 = ~n6819;
assign n1672 = ~(n1086 | n5958);
assign n8190 = ~(n11580 | n11971);
assign n6488 = ~(n7120 | n7161);
assign n13571 = n13096 & n13645;
assign n10960 = ~n81;
assign n3512 = ~n2484;
assign n9466 = n13096 & n6778;
assign n6855 = n3762 & n6418;
assign n8082 = n9953 & n9;
assign n13614 = n11470 & n8869;
assign n2247 = n8358 & n12061;
assign n3553 = n1112 | n3308;
assign n3088 = ~n13696;
assign n238 = n7177 & n8496;
assign n3257 = n12020 | n4896;
assign n13562 = n13367 & n11118;
assign n13474 = ~(n10936 | n9675);
assign n5741 = ~(n9404 | n8840);
assign n13375 = n9898 & n13733;
assign n9387 = n7026 & n13412;
assign n3712 = n13525 & n5207;
assign n9593 = n2747 | n8381;
assign n3878 = n11950 & n1632;
assign n4987 = n1258 | n3564;
assign n12842 = n11097 | n13200;
assign n4009 = n5362 | n12256;
assign n13404 = ~n5871;
assign n4355 = n10330 & n4219;
assign n2912 = n2724 & n10432;
assign n2376 = n5434 & n2829;
assign n5785 = n2310 & n6593;
assign n2132 = ~n3989;
assign n297 = ~(n11771 | n6475);
assign n9478 = n10330 & n13735;
assign n1705 = ~n12927;
assign n8358 = ~n10177;
assign n12287 = n3365 & n984;
assign n4378 = n10808 | n6265;
assign n13223 = n7211 & n6369;
assign n6732 = n13276 | n7153;
assign n4473 = n10871 | n12571;
assign n871 = ~n9757;
assign n12162 = ~(n2752 | n142);
assign n9225 = n9285 | n5650;
assign n13959 = n2334 & n8577;
assign n11067 = n553 | n13772;
assign n14332 = ~n5872;
assign n13127 = n11748 & n3079;
assign n11656 = n4033 | n9067;
assign n879 = n7745 & n10350;
assign n14313 = ~n1436;
assign n1033 = ~(n12288 | n9927);
assign n4149 = n7402 & n5129;
assign n9838 = ~(n5480 | n11730);
assign n8209 = ~n10108;
assign n10189 = ~n8925;
assign n7190 = n4554 & n4103;
assign n7491 = n10019 | n11544;
assign n9472 = n11213 & n5700;
assign n3743 = ~n11425;
assign n2419 = n5603 | n10299;
assign n5503 = n327 & n10094;
assign n4153 = n13226 | n11583;
assign n1966 = n12121 & n11606;
assign n10324 = n2949 | n1451;
assign n4835 = n8866 & n9372;
assign n10878 = ~(n7229 | n11041);
assign n7299 = n1071 & n13764;
assign n11995 = n11495 & n13915;
assign n7136 = ~(n13154 | n8104);
assign n2927 = n11316 & n375;
assign n7363 = n10820 & n2984;
assign n11936 = n12695 | n5401;
assign n2262 = n10025 | n4172;
assign n3467 = ~(n6907 | n7432);
assign n8382 = n2643 & n4242;
assign n9499 = n4901 & n4714;
assign n6564 = n7970 & n4421;
assign n4321 = n536 & n8766;
assign n12647 = n12292 | n6650;
assign n11168 = n10784 | n9018;
assign n11698 = n13516 | n9233;
assign n9034 = n2949 | n215;
assign n2105 = n6695 | n11820;
assign n588 = ~n10384;
assign n9815 = n4684 | n7569;
assign n8540 = ~n11633;
assign n1606 = n98 & n11661;
assign n11161 = n13433 & n345;
assign n7918 = n2758 & n3705;
assign n1771 = ~n11375;
assign n3209 = n4347 & n1836;
assign n11025 = n9323 & n10770;
assign n1341 = ~(n1844 | n13011);
assign n8503 = n8043 & n4499;
assign n8147 = ~n5182;
assign n10980 = ~(n5435 | n13616);
assign n5579 = n432 & n8118;
assign n3721 = ~(n2154 | n1858);
assign n8688 = ~(n8363 | n13975);
assign n1371 = n4967 | n5763;
assign n3065 = n4898 | n2018;
assign n3738 = n10556 & n9220;
assign n5891 = ~n7600;
assign n11276 = n10560 | n4322;
assign n1731 = n10562 & n1433;
assign n2343 = ~n12244;
assign n552 = n5459 & n12340;
assign n8321 = n1071 & n12022;
assign n13013 = ~(n4207 | n5164);
assign n12242 = n12139 | n5646;
assign n2345 = ~(n13458 | n5518);
assign n5221 = n2080 & n11392;
assign n3286 = ~n7346;
assign n6354 = ~n3361;
assign n3109 = n412 | n6668;
assign n1977 = n12759 | n4177;
assign n3988 = n8605 & n4019;
assign n10634 = n4128 | n7112;
assign n14292 = n5266 | n8854;
assign n11596 = n7670 & n12546;
assign n9465 = n13132 & n3364;
assign n14222 = ~(n6747 | n8787);
assign n1711 = ~n382;
assign n9579 = n4346 & n7193;
assign n2871 = n11384 & n13033;
assign n6932 = ~(n1218 | n9439);
assign n10504 = n838 | n1132;
assign n11408 = n2643 & n2358;
assign n10415 = n1383 | n6709;
assign n12686 = n5253 | n7937;
assign n10034 = n9747 | n1070;
assign n6888 = ~n2607;
assign n916 = n865 & n6821;
assign n2302 = ~(n5665 | n5932);
assign n3070 = n8521 & n3977;
assign n13745 = ~n13038;
assign n6610 = n2562 | n11338;
assign n13800 = n12101 & n5969;
assign n749 = ~n3922;
assign n11800 = n10367 & n3552;
assign n4581 = ~n4490;
assign n12065 = n5088 & n12816;
assign n6233 = n2401 | n11962;
assign n10666 = n4508 | n9719;
assign n12775 = n13952 & n590;
assign n6650 = n1772 & n5719;
assign n13537 = ~n12106;
assign n8669 = n10396 | n13748;
assign n9863 = ~n13190;
assign n8715 = n11607 & n7477;
assign n12815 = n2533 & n9335;
assign n452 = n4791 | n10190;
assign n2840 = n2645 | n9337;
assign n4853 = n2021 & n169;
assign n10763 = ~n261;
assign n2607 = ~n3443;
assign n12088 = ~n7146;
assign n9030 = n6318 & n6093;
assign n6428 = ~n3021;
assign n12893 = n480 | n6699;
assign n12923 = ~(n9563 | n4101);
assign n5132 = ~n4317;
assign n7251 = n1804 & n9132;
assign n12250 = ~n3967;
assign n4182 = n3768 | n4761;
assign n4568 = n1854 & n13825;
assign n5833 = ~n1676;
assign n13419 = n11737 & n9183;
assign n13984 = ~(n12757 | n13159);
assign n7000 = n2533 & n3507;
assign n12521 = ~n6193;
assign n13378 = ~(n6788 | n10856);
assign n12763 = n13516 | n11888;
assign n13405 = n2521 & n12837;
assign n1392 = ~(n5018 | n3568);
assign n8677 = n2158 & n9159;
assign n9249 = n4822 | n9042;
assign n7953 = n2998 & n6340;
assign n10959 = ~(n7229 | n2952);
assign n10026 = n3076 | n2159;
assign n11137 = n2387 | n12183;
assign n11434 = ~(n1522 | n11531);
assign n8205 = n7063 & n9855;
assign n1103 = ~(n13399 | n164);
assign n973 = n8747 | n13660;
assign n3951 = ~(n14216 | n5112);
assign n5359 = n1152 | n1299;
assign n729 = n9931 | n2222;
assign n10863 = n7219 | n7162;
assign n4317 = n11130 & n2548;
assign n6985 = n7909 & n4406;
assign n253 = n1962 & n13022;
assign n6864 = n1678 & n10735;
assign n4807 = ~n2918;
assign n7644 = n5574 | n6703;
assign n2535 = n555 | n4545;
assign n12971 = n6206 | n8041;
assign n8748 = ~n12331;
assign n4455 = ~(n450 | n14311);
assign n3633 = n8965 & n620;
assign n8217 = ~n2973;
assign n4490 = ~n9987;
assign n1844 = ~n7404;
assign n9210 = n11558 | n10527;
assign n4731 = n1100 & n13284;
assign n1550 = n5275 & n171;
assign n159 = ~(n3867 | n2717);
assign n14081 = n7911 & n12737;
assign n2425 = n8849 & n7820;
assign n4636 = ~(n11870 | n6529);
assign n10391 = ~(n6211 | n117);
assign n14133 = ~n1079;
assign n4733 = n8480 | n9680;
assign n2178 = n11223 | n10818;
assign n268 = n12147 & n8267;
assign n14057 = n13728 & n929;
assign n5143 = n11702 & n12709;
assign n10872 = n1788 & n10999;
assign n12364 = n11724 | n4986;
assign n4008 = n7436 | n14212;
assign n10659 = n10331 | n1633;
assign n10367 = ~n82;
assign n4643 = n2985 & n6641;
assign n8270 = n5180 | n5173;
assign n13329 = n6781 | n12993;
assign n2936 = n333 & n5318;
assign n7278 = ~n2723;
assign n11862 = ~(n194 | n10271);
assign n11335 = n4973 & n8792;
assign n2630 = n10626 | n5853;
assign n13293 = n6596 | n354;
assign n13048 = n1857 & n13631;
assign n4138 = n7767 & n7125;
assign n13271 = n392 & n10439;
assign n5095 = n12092 & n13185;
assign n9515 = n4358 & n1934;
assign n8215 = n10407 & n10128;
assign n13342 = ~n13383;
assign n11401 = n14376 & n9616;
assign n12368 = n8513 | n13684;
assign n8627 = n12858 & n1892;
assign n764 = n4128 | n12264;
assign n6146 = n3952 & n5413;
assign n9759 = n3161 | n3092;
assign n6163 = n6266 | n13429;
assign n1695 = n85 | n6859;
assign n12320 = n8453 & n7139;
assign n90 = n1678 & n4482;
assign n14426 = n4546 & n12207;
assign n5654 = n9673 & n9274;
assign n12978 = ~(n8816 | n413);
assign n13128 = ~n421;
assign n8412 = ~n1639;
assign n10208 = n1602 | n12252;
assign n10348 = n4255 | n5206;
assign n4234 = n10933 | n5563;
assign n8733 = ~(n2597 | n7841);
assign n6696 = n6517 & n2054;
assign n2234 = ~(n4928 | n4368);
assign n3686 = ~(n14367 | n4653);
assign n7410 = n185 | n5193;
assign n6381 = n5137 & n9160;
assign n13029 = n13297 & n14268;
assign n11568 = n12870 | n14215;
assign n11619 = n1699 & n11518;
assign n5623 = n3424 & n10173;
assign n8395 = n5038 & n10275;
assign n4304 = n11980 | n2979;
assign n10548 = ~(n10136 | n9126);
assign n14354 = n13633 & n3523;
assign n4027 = n231 & n7196;
assign n3014 = ~(n2341 | n9284);
assign n5576 = n9494 | n5467;
assign n14040 = n5587 | n10416;
assign n6898 = ~n2468;
assign n1577 = ~n5306;
assign n9529 = ~n1041;
assign n4037 = n8432 & n5175;
assign n2823 = n10367 & n2076;
assign n8228 = n6957 & n13469;
assign n5080 = n3846 & n10585;
assign n12436 = n9716 | n1814;
assign n815 = ~n3972;
assign n1649 = n4354 & n2168;
assign n2406 = n10294 | n7552;
assign n1925 = n3800 | n9905;
assign n8122 = ~n2250;
assign n7068 = ~n3926;
assign n96 = n6830 & n12910;
assign n11425 = ~n13135;
assign n6083 = n1427 & n6406;
assign n13544 = n7708 & n10326;
assign n560 = ~n5786;
assign n3056 = n11951 | n6019;
assign n4236 = n10710 & n13218;
assign n1133 = n3212 & n13536;
assign n10186 = ~n3461;
assign n8965 = ~n10303;
assign n10534 = ~n7441;
assign n3479 = n638 & n5349;
assign n3306 = n13781 & n7412;
assign n7600 = n4258 & n5702;
assign n1322 = n10323 | n4521;
assign n1650 = n3424 & n10054;
assign n6984 = n3492 | n13882;
assign n13923 = n5406 | n8033;
assign n3987 = n4851 & n12869;
assign n4349 = n6519 | n5801;
assign n7998 = n5891 | n6392;
assign n11471 = n898 & n1778;
assign n4918 = n10622 & n6155;
assign n9480 = n4052 | n7000;
assign n12819 = n5908 | n14024;
assign n3831 = n3370 & n10304;
assign n7161 = ~(n11980 | n12838);
assign n13998 = n10396 | n268;
assign n7673 = ~n10269;
assign n3129 = n4908 | n11665;
assign n11305 = ~n8003;
assign n13728 = ~n14475;
assign n10223 = n5459 & n3264;
assign n5206 = n3986 & n2109;
assign n1305 = n11300 & n5757;
assign n4059 = ~(n10637 | n3040);
assign n4063 = ~(n13255 | n4218);
assign n1120 = ~n9608;
assign n3824 = n13698 | n6557;
assign n5207 = n8476 | n10144;
assign n8912 = n4631 | n5520;
assign n4863 = n3047 | n14276;
assign n6405 = ~(n7364 | n532);
assign n5217 = n12614 | n10765;
assign n5640 = ~n411;
assign n6627 = n3755 & n10178;
assign n13088 = n5139 | n10766;
assign n5108 = ~n179;
assign n10303 = ~n9537;
assign n7508 = n873 & n1035;
assign n8593 = n782 | n4585;
assign n5315 = ~n3021;
assign n9672 = ~(n12193 | n12273);
assign n5697 = n14319 | n4954;
assign n4833 = n3724 & n9750;
assign n6846 = n5434 & n14005;
assign n1226 = ~(n14135 | n5914);
assign n7911 = ~n8524;
assign n3437 = n14313 & n8438;
assign n12995 = n12852 | n3263;
assign n2526 = n1535 | n13326;
assign n6674 = n5137 & n11784;
assign n3123 = n5240 & n1444;
assign n4993 = n5454 | n2658;
assign n9704 = ~(n13276 | n7804);
assign n9806 = ~n10346;
assign n10235 = ~(n7971 | n2899);
assign n4305 = n2454 & n12194;
assign n11494 = n9265 & n3590;
assign n8932 = ~n2241;
assign n10535 = ~n6096;
assign n10021 = n13446 | n3483;
assign n14032 = n8789 & n5158;
assign n13841 = n1539 & n7556;
assign n7646 = n1535 | n8922;
assign n837 = n2315 | n10270;
assign n14419 = ~n3070;
assign n7668 = n4684 | n7415;
assign n5012 = ~n2432;
assign n5911 = n1223 | n932;
assign n14456 = n13069 & n14194;
assign n10176 = n8453 & n837;
assign n12105 = ~n2906;
assign n6462 = n6373 | n1880;
assign n1757 = n1840 | n12589;
assign n4400 = n4509 & n12728;
assign n8123 = n2445 & n2890;
assign n6203 = n7208 & n3454;
assign n7401 = ~n844;
assign n14068 = n9353 | n14153;
assign n9496 = ~(n6679 | n7444);
assign n14088 = ~n12874;
assign n12921 = n286 & n9125;
assign n13330 = n13885 | n10033;
assign n2152 = n428 & n8938;
assign n5945 = ~(n8209 | n7377);
assign n4757 = ~n11325;
assign n12013 = ~n6807;
assign n11486 = ~(n4144 | n10625);
assign n2001 = n12037 | n3367;
assign n6600 = ~n1776;
assign n10545 = n8480 | n6647;
assign n4085 = n2401 | n11306;
assign n9442 = ~n6274;
assign n13889 = n5548 | n13222;
assign n9623 = n3445 | n11382;
assign n6160 = n3559 | n12917;
assign n2547 = ~n4633;
assign n117 = ~(n8527 | n3686);
assign n2268 = n14282 | n1649;
assign n3429 = n9747 | n13314;
assign n13188 = n11724 | n1197;
assign n4886 = n900 | n11443;
assign n8691 = ~(n8212 | n3032);
assign n2792 = n7068 & n9200;
assign n14314 = n11008 & n14201;
assign n6144 = n10760 | n7354;
assign n1113 = n3401 & n12486;
assign n13675 = ~n9306;
assign n8619 = n4627 & n9344;
assign n9173 = n12531 & n13787;
assign n899 = n695 | n1906;
assign n1436 = ~n10485;
assign n965 = ~n6990;
assign n11372 = n9422 | n12881;
assign n4118 = ~(n11148 | n11662);
assign n4302 = n5732 | n14151;
assign n4348 = ~(n10651 | n13259);
assign n14113 = n4205 | n7012;
assign n14183 = ~(n14166 | n341);
assign n8530 = n5569 | n1340;
assign n9874 = n4877 | n821;
assign n1975 = n9429 | n11523;
assign n2292 = n14110 | n11575;
assign n9749 = n5011 & n11932;
assign n10681 = n6318 & n11568;
assign n13053 = ~(n10637 | n12743);
assign n8396 = n13948 | n5583;
assign n4868 = n8412 & n1757;
assign n9992 = n8490 | n10410;
assign n5690 = ~n14216;
assign n3615 = n4508 | n11833;
assign n3973 = ~(n2017 | n13389);
assign n2658 = n13379 & n4250;
assign n1182 = n14313 & n841;
assign n1997 = ~n1458;
assign n8117 = n2330 & n10045;
assign n12186 = n11048 | n4414;
assign n1617 = ~n264;
assign n14442 = n10461 | n4397;
assign n6067 = n957 | n9555;
assign n1126 = ~(n12069 | n8876);
assign n1725 = n2315 | n4586;
assign n4369 = n889 & n10077;
assign n9324 = n13755 & n9122;
assign n6364 = n4650 & n4385;
assign n4165 = n11636 & n5013;
assign n6815 = n13226 | n9684;
assign n13242 = n11679 & n6675;
assign n125 = n2401 | n13629;
assign n13694 = n2021 & n5564;
assign n823 = n14038 & n13590;
assign n8121 = ~(n12651 | n1174);
assign n10447 = ~(n5197 | n3475);
assign n9726 = ~n10372;
assign n7751 = n10922 & n14403;
assign n9811 = ~n6819;
assign n1119 = n13080 | n14478;
assign n4173 = n7678 | n13868;
assign n3921 = n9564 & n8422;
assign n1343 = n7430 | n1083;
assign n11350 = ~n5665;
assign n7297 = n8877 | n5102;
assign n2661 = n4822 | n4334;
assign n7590 = ~n10615;
assign n9640 = n7401 & n3820;
assign n1679 = n5575 | n2116;
assign n3415 = n12821 | n2095;
assign n4394 = ~n8963;
assign n2849 = n11572 | n3377;
assign n11133 = n1697 | n12751;
assign n13906 = n12918 & n1933;
assign n10741 = n2857 | n13269;
assign n7737 = n163 | n11945;
assign n14306 = n7427 & n9032;
assign n13112 = ~n9453;
assign n13849 = n2099 & n9304;
assign n245 = n2310 & n9836;
assign n3547 = n4880 & n11608;
assign n12298 = n8507 & n8847;
assign n10857 = ~n12874;
assign n459 = n5640 & n1656;
assign n6757 = n8726 | n1190;
assign n1034 = n2246 | n1505;
assign n9137 = ~(n10233 | n6634);
assign n6542 = n12615 & n13721;
assign n8051 = ~(n5847 | n5791);
assign n2022 = n3526 & n7562;
assign n5373 = n1669 | n13608;
assign n1788 = ~n6975;
assign n1990 = n6046 | n7349;
assign n1108 = n3491 & n4632;
assign n3255 = ~n8704;
assign n11111 = ~n1053;
assign n12214 = n12712 | n7256;
assign n14261 = n10969 & n2944;
assign n3283 = n976 | n4919;
assign n6282 = ~(n8544 | n1090);
assign n14478 = n11867 & n2230;
assign n13706 = ~n12687;
assign n5894 = ~(n5596 | n9616);
assign n8693 = n553 | n5524;
assign n81 = n8179 & n3155;
assign n12628 = n4313 | n2753;
assign n1054 = n3762 | n8635;
assign n5651 = n4790 & n229;
assign n9342 = n8439 & n4164;
assign n2591 = n7481 | n2706;
assign n664 = n6013 & n3594;
assign n14034 = n1125 & n549;
assign n857 = n10310 & n4072;
assign n4187 = n9188 & n11145;
assign n3529 = n5491 | n10486;
assign n2148 = n748 & n576;
assign n9691 = n8045 | n14119;
assign n9697 = n7693 & n7649;
assign n5605 = ~n13633;
assign n3509 = n3785 & n11979;
assign n11140 = n3800 | n12604;
assign n8449 = ~(n648 | n5216);
assign n2811 = ~(n1612 | n1486);
assign n11774 = n10825 | n4028;
assign n3940 = ~(n506 | n6964);
assign n9259 = n2422 & n8245;
assign n9300 = n12414 | n5115;
assign n8683 = n5857 & n6245;
assign n7427 = ~n261;
assign n10352 = n4052 | n2308;
assign n2233 = n4018 & n10159;
assign n11591 = n1494 | n10896;
assign n4732 = n13489 & n10044;
assign n2151 = n4973 & n6004;
assign n5016 = n8183 & n4875;
assign n167 = n4619 & n3625;
assign n5648 = n13236 & n8916;
assign n11339 = n11303 | n14111;
assign n3773 = n3526 & n3538;
assign n10496 = n13142 | n14235;
assign n4488 = n9804 | n4885;
assign n11896 = n14213 & n10698;
assign n14097 = n13485 | n10160;
assign n3425 = n6263 | n8966;
assign n1056 = n12391 & n13970;
assign n12445 = ~n5613;
assign n14052 = ~(n8212 | n11101);
assign n1542 = n8582 | n7711;
assign n9870 = n6625 & n5426;
assign n4967 = ~n10889;
assign n3269 = n11231 | n10754;
assign n12651 = ~n2970;
assign n9682 = n9289 | n12929;
assign n4574 = ~n920;
assign n3867 = ~n4859;
assign n12638 = n13078 & n4995;
assign n12845 = n11737 & n2020;
assign n1098 = n11569 & n2841;
assign n10022 = n3635 & n615;
assign n750 = n7391 & n8545;
assign n808 = ~n8361;
assign n6261 = n4988 | n4328;
assign n12323 = n3367 | n11776;
assign n14515 = n8151 | n12196;
assign n4002 = ~(n11488 | n4747);
assign n10958 = n4486 & n3606;
assign n8089 = n13246 & n4269;
assign n3049 = n1576 | n5651;
assign n658 = n3125 | n9478;
assign n1718 = n11674 & n9512;
assign n5566 = n12038 & n9477;
assign n12394 = n9769 & n4134;
assign n13758 = n11097 | n373;
assign n5923 = n11090 | n9099;
assign n10243 = n7327 & n2339;
assign n7703 = n69 | n11900;
assign n1271 = n2318 | n1795;
assign n4595 = n14065 & n3199;
assign n9435 = n7736 | n8893;
assign n13975 = ~(n3871 | n3458);
assign n9834 = ~(n512 | n2757);
assign n1076 = n9956 | n8397;
assign n5670 = n11011 | n14369;
assign n13316 = n5467 & n886;
assign n12241 = n11581 | n3312;
assign n940 = n10229 & n3110;
assign n5850 = n3846 & n1284;
assign n6435 = n7736 | n1745;
assign n10180 = ~(n573 | n12024);
assign n1882 = n2387 | n7715;
assign n6319 = ~n6011;
assign n1710 = n12389 & n13291;
assign n12255 = n4581 & n5954;
assign n2063 = n7912 | n951;
assign n1429 = n5507 | n7305;
assign n14036 = n6525 & n3982;
assign n9365 = ~(n10309 | n9440);
assign n536 = ~n1478;
assign n5757 = n3168 | n4057;
assign n3438 = n12057 & n10090;
endmodule
