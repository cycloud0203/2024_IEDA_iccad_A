// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Fri Jun 14 22:43:34 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604,
    n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112,
    n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288,
    n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558,
    n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738,
    n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088,
    n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272,
    n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479,
    n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816,
    n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136,
    n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349,
    n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618,
    n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952,
    n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319,
    n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722,
    n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031,
    n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213,
    n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443,
    n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822,
    n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379,
    n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590,
    n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790,
    n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305,
    n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566,
    n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731,
    n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963,
    n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305,
    n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614,
    n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827,
    n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251,
    n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493,
    n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926,
    n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117,
    n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514,
    n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763,
    n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220,
    n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479,
    n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667,
    n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121,
    n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398,
    n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650,
    n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900,
    n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263,
    n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494,
    n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783,
    n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230,
    n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603,
    n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899,
    n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271,
    n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546,
    n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918,
    n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247,
    n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524,
    n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968,
    n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095,
    n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954,
    n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227,
    n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496,
    n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880,
    n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107,
    n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327,
    n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531,
    n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770,
    n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040,
    n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259,
    n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478,
    n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946,
    n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287,
    n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674,
    n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898,
    n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068,
    n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309,
    n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492,
    n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764,
    n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068,
    n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333,
    n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657,
    n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912,
    n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129,
    n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485,
    n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023,
    n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240,
    n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435,
    n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643,
    n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926,
    n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191,
    n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512,
    n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752,
    n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089,
    n27104, n27120, n27134, n27188,
    n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194  );
  input  n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583,
    n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099,
    n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279,
    n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536,
    n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689,
    n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035,
    n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210,
    n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421,
    n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809,
    n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030,
    n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324,
    n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582,
    n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945,
    n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306,
    n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665,
    n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026,
    n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211,
    n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438,
    n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752,
    n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369,
    n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556,
    n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785,
    n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149,
    n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524,
    n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721,
    n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949,
    n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285,
    n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581,
    n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806,
    n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246,
    n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460,
    n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872,
    n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096,
    n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411,
    n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739,
    n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201,
    n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473,
    n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630,
    n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113,
    n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384,
    n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626,
    n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892,
    n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190,
    n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490,
    n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781,
    n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148,
    n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576,
    n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826,
    n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258,
    n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539,
    n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884,
    n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223,
    n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521,
    n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911,
    n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090,
    n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911,
    n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171,
    n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483,
    n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745,
    n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081,
    n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282,
    n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515,
    n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701,
    n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036,
    n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250,
    n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470,
    n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929,
    n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276,
    n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654,
    n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839,
    n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043,
    n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290,
    n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470,
    n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660,
    n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065,
    n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304,
    n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586,
    n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895,
    n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093,
    n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374,
    n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937,
    n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168,
    n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381,
    n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629,
    n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923,
    n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180,
    n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510,
    n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748,
    n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037,
    n27089, n27104, n27120, n27134, n27188;
  output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355_1, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361_1, new_n2362, new_n2363_1, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374_1, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387_1, new_n2388_1, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409_1, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416_1, new_n2417, new_n2418, new_n2419, new_n2420_1,
    new_n2421_1, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440_1, new_n2441, new_n2442, new_n2443, new_n2444_1,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479_1, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513_1, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533_1, new_n2534,
    new_n2535_1, new_n2536, new_n2537_1, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547_1, new_n2548, new_n2549, new_n2550, new_n2551, new_n2552,
    new_n2553_1, new_n2554, new_n2555_1, new_n2556, new_n2557, new_n2558,
    new_n2559, new_n2560_1, new_n2561_1, new_n2562, new_n2563, new_n2564,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570_1,
    new_n2571, new_n2572, new_n2573_1, new_n2574, new_n2575, new_n2576,
    new_n2577, new_n2578_1, new_n2579, new_n2580, new_n2581, new_n2582_1,
    new_n2583, new_n2584, new_n2585, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2593, new_n2594, new_n2595,
    new_n2596, new_n2597, new_n2598, new_n2599, new_n2601, new_n2602_1,
    new_n2603, new_n2604, new_n2605, new_n2606, new_n2607, new_n2608,
    new_n2609, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619_1, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646_1, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659_1, new_n2660, new_n2661_1, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680_1, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693_1,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703_1, new_n2704, new_n2705,
    new_n2706_1, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711_1,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731_1, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743_1, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761_1, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774_1, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779_1, new_n2780, new_n2781, new_n2782, new_n2783_1,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809_1, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816_1, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826_1, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2848, new_n2849,
    new_n2850, new_n2851, new_n2852, new_n2853_1, new_n2854, new_n2855,
    new_n2856, new_n2857, new_n2858_1, new_n2859, new_n2860_1, new_n2861,
    new_n2862, new_n2863, new_n2864, new_n2865, new_n2866, new_n2867,
    new_n2868, new_n2869, new_n2870, new_n2871, new_n2872, new_n2873,
    new_n2874, new_n2875, new_n2876, new_n2877, new_n2878, new_n2879,
    new_n2880, new_n2881, new_n2882, new_n2883, new_n2884, new_n2885,
    new_n2886_1, new_n2887_1, new_n2888, new_n2889, new_n2890, new_n2891,
    new_n2892, new_n2893, new_n2894, new_n2895, new_n2896, new_n2897,
    new_n2898, new_n2899, new_n2900, new_n2901, new_n2902, new_n2903,
    new_n2904, new_n2905, new_n2906, new_n2907, new_n2908, new_n2909,
    new_n2910, new_n2911, new_n2912, new_n2913, new_n2914, new_n2915,
    new_n2916, new_n2917, new_n2918, new_n2919, new_n2920, new_n2921,
    new_n2922, new_n2923, new_n2924, new_n2925, new_n2926, new_n2927,
    new_n2928, new_n2929_1, new_n2930, new_n2931, new_n2932, new_n2933,
    new_n2934, new_n2935, new_n2936, new_n2937, new_n2938, new_n2939,
    new_n2940, new_n2941, new_n2942, new_n2943, new_n2944_1, new_n2945,
    new_n2946, new_n2947, new_n2948_1, new_n2949, new_n2950, new_n2951,
    new_n2952, new_n2953, new_n2954, new_n2955, new_n2956, new_n2957,
    new_n2958, new_n2959, new_n2960, new_n2961_1, new_n2962, new_n2963,
    new_n2964, new_n2965, new_n2966, new_n2967, new_n2968, new_n2969,
    new_n2970, new_n2971_1, new_n2972, new_n2973, new_n2974, new_n2975,
    new_n2976, new_n2977, new_n2978_1, new_n2979_1, new_n2980, new_n2981,
    new_n2983, new_n2984, new_n2985_1, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999_1, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010_1, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017_1, new_n3018_1,
    new_n3019, new_n3020_1, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030_1,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067_1, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076_1, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3085, new_n3086, new_n3087, new_n3088, new_n3089_1, new_n3090,
    new_n3091, new_n3092, new_n3093, new_n3094, new_n3095, new_n3096,
    new_n3097, new_n3098, new_n3099, new_n3100, new_n3101, new_n3102,
    new_n3103, new_n3104, new_n3105, new_n3106, new_n3107, new_n3108,
    new_n3109, new_n3110, new_n3111, new_n3112, new_n3113, new_n3114,
    new_n3115, new_n3116, new_n3117, new_n3118, new_n3119, new_n3120,
    new_n3121, new_n3122, new_n3123, new_n3124, new_n3125_1, new_n3126_1,
    new_n3127, new_n3128, new_n3129, new_n3130, new_n3131, new_n3132,
    new_n3133, new_n3134, new_n3135, new_n3136_1, new_n3137, new_n3138,
    new_n3139, new_n3140, new_n3141, new_n3142, new_n3143, new_n3144,
    new_n3145, new_n3146, new_n3147, new_n3148, new_n3149, new_n3150,
    new_n3151, new_n3152, new_n3153, new_n3154, new_n3155, new_n3156,
    new_n3157, new_n3158, new_n3159, new_n3160, new_n3161_1, new_n3162,
    new_n3163, new_n3164_1, new_n3165, new_n3166, new_n3167, new_n3168,
    new_n3169, new_n3170, new_n3171, new_n3172, new_n3173, new_n3174,
    new_n3175, new_n3176, new_n3177, new_n3178, new_n3179, new_n3180,
    new_n3181, new_n3182, new_n3183, new_n3184, new_n3185, new_n3186,
    new_n3187, new_n3188, new_n3189, new_n3190, new_n3191, new_n3192,
    new_n3193, new_n3194, new_n3195, new_n3196, new_n3197, new_n3198,
    new_n3199, new_n3200, new_n3201, new_n3202, new_n3203, new_n3204,
    new_n3205, new_n3206, new_n3207, new_n3208_1, new_n3209, new_n3210,
    new_n3211, new_n3212, new_n3213, new_n3214, new_n3215, new_n3216,
    new_n3217, new_n3218, new_n3219_1, new_n3220, new_n3221, new_n3222,
    new_n3223, new_n3224, new_n3225, new_n3226, new_n3227, new_n3228_1,
    new_n3229, new_n3230, new_n3231, new_n3232, new_n3233, new_n3234,
    new_n3235_1, new_n3236, new_n3237, new_n3238, new_n3239, new_n3240,
    new_n3241, new_n3242, new_n3243, new_n3244_1, new_n3245, new_n3246,
    new_n3247, new_n3248, new_n3249, new_n3250, new_n3251, new_n3252,
    new_n3253_1, new_n3254, new_n3255, new_n3256, new_n3257, new_n3258,
    new_n3259, new_n3260_1, new_n3261, new_n3262, new_n3263_1, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279_1, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289_1,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301_1,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306_1, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316_1, new_n3317, new_n3318, new_n3319,
    new_n3320_1, new_n3321, new_n3322, new_n3323, new_n3324_1, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332_1, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343_1,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349_1,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366_1, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390_1, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3404, new_n3405, new_n3406, new_n3407, new_n3408, new_n3409,
    new_n3410, new_n3411, new_n3412, new_n3413, new_n3414, new_n3415,
    new_n3416, new_n3417, new_n3418, new_n3419, new_n3420, new_n3421,
    new_n3422, new_n3423, new_n3424, new_n3425_1, new_n3426_1, new_n3427,
    new_n3428, new_n3429, new_n3430, new_n3431, new_n3432, new_n3433,
    new_n3434, new_n3435, new_n3436, new_n3437, new_n3438, new_n3439,
    new_n3440, new_n3441, new_n3442, new_n3443, new_n3444, new_n3445,
    new_n3446, new_n3447, new_n3448, new_n3449, new_n3450, new_n3451_1,
    new_n3452, new_n3453, new_n3454, new_n3455, new_n3456, new_n3457,
    new_n3458, new_n3459_1, new_n3460_1, new_n3461, new_n3462, new_n3463,
    new_n3464, new_n3465, new_n3466, new_n3467, new_n3468_1, new_n3469,
    new_n3470, new_n3471, new_n3472, new_n3473, new_n3474, new_n3475,
    new_n3476, new_n3477, new_n3478, new_n3479, new_n3480_1, new_n3481,
    new_n3482, new_n3483, new_n3484, new_n3485, new_n3486, new_n3487,
    new_n3488, new_n3489, new_n3490, new_n3491, new_n3492, new_n3493,
    new_n3494, new_n3495, new_n3496, new_n3497, new_n3498, new_n3499,
    new_n3500, new_n3501, new_n3502_1, new_n3503, new_n3504, new_n3505,
    new_n3506_1, new_n3507, new_n3508, new_n3509, new_n3510, new_n3511,
    new_n3512, new_n3513, new_n3514, new_n3515, new_n3516_1, new_n3517,
    new_n3518, new_n3519, new_n3520, new_n3521, new_n3522, new_n3523,
    new_n3524, new_n3525, new_n3526, new_n3527, new_n3528_1, new_n3529,
    new_n3530, new_n3531, new_n3532, new_n3533, new_n3534, new_n3535,
    new_n3536, new_n3537, new_n3538, new_n3539, new_n3540, new_n3541_1,
    new_n3542, new_n3543, new_n3544, new_n3545, new_n3546, new_n3547,
    new_n3548, new_n3549, new_n3550, new_n3551, new_n3552, new_n3553,
    new_n3554, new_n3555_1, new_n3556, new_n3557, new_n3558, new_n3559,
    new_n3560, new_n3561_1, new_n3562, new_n3563_1, new_n3564, new_n3565,
    new_n3566, new_n3567, new_n3568, new_n3569, new_n3570_1, new_n3571,
    new_n3572, new_n3573, new_n3574, new_n3575, new_n3576, new_n3577,
    new_n3578, new_n3579, new_n3580, new_n3581, new_n3582_1, new_n3583,
    new_n3584, new_n3585, new_n3586, new_n3587, new_n3588, new_n3589,
    new_n3590, new_n3591, new_n3592, new_n3593, new_n3594, new_n3595,
    new_n3596, new_n3597, new_n3598, new_n3599, new_n3600, new_n3601,
    new_n3602, new_n3603, new_n3604, new_n3605, new_n3606, new_n3607,
    new_n3608, new_n3609, new_n3610, new_n3611, new_n3612, new_n3613,
    new_n3614, new_n3615, new_n3616, new_n3617_1, new_n3618_1, new_n3619,
    new_n3620, new_n3621, new_n3622, new_n3623, new_n3624, new_n3625,
    new_n3626, new_n3627, new_n3628, new_n3629, new_n3630, new_n3631,
    new_n3632, new_n3633, new_n3634, new_n3635, new_n3636, new_n3637,
    new_n3638, new_n3639, new_n3640, new_n3641, new_n3642_1, new_n3643,
    new_n3644, new_n3645, new_n3646, new_n3647, new_n3648, new_n3649_1,
    new_n3650, new_n3651, new_n3652, new_n3653, new_n3654, new_n3655,
    new_n3656, new_n3657, new_n3658, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665_1, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679_1, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710_1,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3724, new_n3725_1, new_n3726, new_n3727, new_n3728,
    new_n3729, new_n3730, new_n3731, new_n3732, new_n3733_1, new_n3734,
    new_n3735, new_n3736, new_n3737, new_n3738, new_n3739, new_n3740_1,
    new_n3741, new_n3742, new_n3743, new_n3744, new_n3745, new_n3746,
    new_n3747, new_n3748, new_n3749, new_n3750, new_n3751, new_n3752,
    new_n3753, new_n3754, new_n3755_1, new_n3756, new_n3757, new_n3758_1,
    new_n3759, new_n3760_1, new_n3761, new_n3762, new_n3763, new_n3764,
    new_n3765, new_n3766, new_n3767, new_n3768, new_n3769, new_n3770,
    new_n3771, new_n3772, new_n3773, new_n3774, new_n3775, new_n3776,
    new_n3777, new_n3778, new_n3779, new_n3780, new_n3781_1, new_n3782,
    new_n3783, new_n3784, new_n3785_1, new_n3786, new_n3787, new_n3788,
    new_n3789, new_n3790, new_n3791, new_n3792, new_n3793, new_n3794_1,
    new_n3795_1, new_n3796, new_n3797, new_n3798, new_n3799, new_n3800,
    new_n3801, new_n3802, new_n3803, new_n3804, new_n3805, new_n3806,
    new_n3807, new_n3808, new_n3809, new_n3810, new_n3811, new_n3812,
    new_n3813, new_n3814, new_n3815, new_n3816, new_n3817, new_n3818,
    new_n3819, new_n3820, new_n3821, new_n3822, new_n3823, new_n3824,
    new_n3825, new_n3826, new_n3827, new_n3828_1, new_n3829, new_n3830,
    new_n3831, new_n3832, new_n3833, new_n3834, new_n3835, new_n3836,
    new_n3837, new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1,
    new_n3843, new_n3844, new_n3845, new_n3846, new_n3847, new_n3848,
    new_n3849, new_n3850_1, new_n3851, new_n3852, new_n3853, new_n3854,
    new_n3855, new_n3856, new_n3857, new_n3858, new_n3859, new_n3860,
    new_n3861, new_n3862, new_n3863, new_n3864, new_n3865, new_n3866,
    new_n3867, new_n3868, new_n3869_1, new_n3870, new_n3871_1, new_n3872,
    new_n3873, new_n3874, new_n3875, new_n3876, new_n3877, new_n3878,
    new_n3879, new_n3880, new_n3881, new_n3882, new_n3883, new_n3884,
    new_n3885, new_n3886, new_n3887, new_n3888, new_n3889, new_n3890,
    new_n3891_1, new_n3892, new_n3893, new_n3894, new_n3895, new_n3896,
    new_n3897, new_n3898, new_n3899, new_n3900, new_n3901, new_n3902,
    new_n3903, new_n3904, new_n3905, new_n3906, new_n3907, new_n3908,
    new_n3909_1, new_n3910, new_n3911, new_n3912, new_n3913, new_n3914,
    new_n3915, new_n3916, new_n3917, new_n3918_1, new_n3919, new_n3920,
    new_n3921, new_n3922, new_n3923, new_n3924, new_n3925_1, new_n3926,
    new_n3927, new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1,
    new_n3933, new_n3934_1, new_n3935, new_n3936, new_n3937, new_n3938,
    new_n3939, new_n3940, new_n3941, new_n3942, new_n3943, new_n3944,
    new_n3945_1, new_n3946, new_n3947, new_n3948, new_n3949, new_n3950,
    new_n3951, new_n3952_1, new_n3953, new_n3954, new_n3955, new_n3956,
    new_n3957, new_n3958, new_n3959_1, new_n3960, new_n3961, new_n3962_1,
    new_n3963, new_n3964, new_n3965, new_n3966, new_n3967, new_n3968,
    new_n3969, new_n3970, new_n3971_1, new_n3972, new_n3973, new_n3974,
    new_n3975, new_n3976, new_n3977, new_n3978, new_n3979, new_n3980,
    new_n3981, new_n3982, new_n3983_1, new_n3984_1, new_n3985, new_n3986,
    new_n3987, new_n3988, new_n3989, new_n3990, new_n3991, new_n3992,
    new_n3993, new_n3994, new_n3995, new_n3996, new_n3997, new_n3998,
    new_n3999, new_n4000_1, new_n4001, new_n4002, new_n4003, new_n4004,
    new_n4005, new_n4006, new_n4007, new_n4008, new_n4009, new_n4010_1,
    new_n4011, new_n4012, new_n4013, new_n4014_1, new_n4015, new_n4016,
    new_n4017, new_n4018, new_n4019, new_n4020, new_n4021, new_n4022,
    new_n4023, new_n4024, new_n4025, new_n4026, new_n4027, new_n4028,
    new_n4029, new_n4030, new_n4031, new_n4032, new_n4033, new_n4034,
    new_n4035, new_n4036, new_n4037, new_n4038, new_n4039, new_n4040,
    new_n4041, new_n4042, new_n4043, new_n4044, new_n4045, new_n4046,
    new_n4047, new_n4048, new_n4049, new_n4050, new_n4051, new_n4052,
    new_n4053, new_n4054, new_n4055, new_n4056, new_n4057, new_n4058,
    new_n4059, new_n4060, new_n4061, new_n4062, new_n4063, new_n4064,
    new_n4065, new_n4066, new_n4067, new_n4068, new_n4069, new_n4070,
    new_n4071_1, new_n4072, new_n4074, new_n4075, new_n4076, new_n4077,
    new_n4078, new_n4079, new_n4080, new_n4081, new_n4082, new_n4083,
    new_n4084, new_n4085_1, new_n4086, new_n4087, new_n4088_1, new_n4089_1,
    new_n4090, new_n4091, new_n4092, new_n4093, new_n4094, new_n4095,
    new_n4096, new_n4097, new_n4098, new_n4099, new_n4100_1, new_n4101,
    new_n4102, new_n4103_1, new_n4104, new_n4105, new_n4106, new_n4107,
    new_n4108, new_n4109, new_n4110, new_n4111, new_n4112, new_n4113,
    new_n4114, new_n4115, new_n4116, new_n4117, new_n4118, new_n4119_1,
    new_n4120, new_n4121, new_n4122, new_n4123_1, new_n4124, new_n4125,
    new_n4126, new_n4127, new_n4128, new_n4129, new_n4130, new_n4131,
    new_n4132, new_n4133, new_n4134_1, new_n4135, new_n4136, new_n4137,
    new_n4138, new_n4139, new_n4140, new_n4141, new_n4142, new_n4143,
    new_n4144, new_n4145, new_n4146_1, new_n4147, new_n4148, new_n4149,
    new_n4150_1, new_n4151_1, new_n4152_1, new_n4153_1, new_n4154,
    new_n4155, new_n4156, new_n4157, new_n4158, new_n4159, new_n4160,
    new_n4161, new_n4162, new_n4163, new_n4164, new_n4165_1, new_n4166,
    new_n4167, new_n4168, new_n4169, new_n4170, new_n4171, new_n4172_1,
    new_n4173_1, new_n4174, new_n4175, new_n4176_1, new_n4177, new_n4178,
    new_n4179, new_n4180, new_n4181, new_n4182, new_n4183, new_n4184,
    new_n4185, new_n4186_1, new_n4187, new_n4188, new_n4189, new_n4190,
    new_n4191, new_n4192, new_n4193, new_n4194, new_n4195, new_n4196,
    new_n4197, new_n4198, new_n4199, new_n4200, new_n4201, new_n4202,
    new_n4203, new_n4204_1, new_n4205_1, new_n4206, new_n4207, new_n4208,
    new_n4209, new_n4210, new_n4211, new_n4212, new_n4213, new_n4214,
    new_n4215_1, new_n4216, new_n4217, new_n4218, new_n4219, new_n4220,
    new_n4221_1, new_n4222, new_n4223, new_n4224_1, new_n4225, new_n4226,
    new_n4227, new_n4228, new_n4229, new_n4230, new_n4231_1, new_n4232,
    new_n4233, new_n4234, new_n4235, new_n4236, new_n4237, new_n4238,
    new_n4239, new_n4240, new_n4241, new_n4242, new_n4243, new_n4244,
    new_n4245, new_n4246, new_n4247, new_n4248, new_n4249, new_n4250,
    new_n4251, new_n4252, new_n4253, new_n4254, new_n4255, new_n4256_1,
    new_n4257, new_n4258, new_n4259, new_n4260, new_n4261, new_n4262,
    new_n4263, new_n4264, new_n4265, new_n4266_1, new_n4267, new_n4268,
    new_n4269, new_n4270, new_n4271, new_n4272_1, new_n4273, new_n4274,
    new_n4275, new_n4276, new_n4277, new_n4278, new_n4279, new_n4280,
    new_n4281, new_n4282, new_n4283, new_n4284, new_n4285, new_n4286,
    new_n4287, new_n4288, new_n4289, new_n4290, new_n4291, new_n4292,
    new_n4293, new_n4294, new_n4295, new_n4296, new_n4297, new_n4298,
    new_n4299, new_n4300, new_n4301, new_n4302, new_n4303, new_n4304,
    new_n4305, new_n4306_1, new_n4307, new_n4308, new_n4309, new_n4310,
    new_n4311, new_n4312, new_n4313, new_n4314, new_n4315, new_n4316,
    new_n4317, new_n4318, new_n4319_1, new_n4320, new_n4321, new_n4322,
    new_n4323, new_n4324, new_n4325_1, new_n4326_1, new_n4327, new_n4328,
    new_n4329, new_n4330, new_n4331, new_n4332, new_n4334, new_n4335,
    new_n4336, new_n4337, new_n4338, new_n4339, new_n4340_1, new_n4341,
    new_n4342, new_n4343, new_n4344, new_n4345, new_n4346, new_n4347,
    new_n4348, new_n4349, new_n4350, new_n4351, new_n4352, new_n4353,
    new_n4354, new_n4355, new_n4356, new_n4357, new_n4358, new_n4359,
    new_n4360, new_n4361, new_n4362, new_n4363, new_n4364, new_n4365,
    new_n4366, new_n4367, new_n4368, new_n4369, new_n4370, new_n4371,
    new_n4372, new_n4373, new_n4374_1, new_n4375, new_n4376_1, new_n4377,
    new_n4378, new_n4379, new_n4380, new_n4381, new_n4382, new_n4383,
    new_n4384, new_n4385, new_n4386, new_n4387, new_n4388, new_n4389,
    new_n4390, new_n4391, new_n4392, new_n4393, new_n4394, new_n4395,
    new_n4396, new_n4397, new_n4398, new_n4399, new_n4400, new_n4401_1,
    new_n4402, new_n4403, new_n4404, new_n4405, new_n4406, new_n4407,
    new_n4408, new_n4409_1, new_n4410, new_n4411, new_n4412, new_n4413,
    new_n4414, new_n4415, new_n4416, new_n4417, new_n4418, new_n4419,
    new_n4420, new_n4421, new_n4422, new_n4423, new_n4424_1, new_n4425,
    new_n4426_1, new_n4427, new_n4428, new_n4429, new_n4430, new_n4431,
    new_n4432_1, new_n4433, new_n4434, new_n4435, new_n4436, new_n4437,
    new_n4438, new_n4439, new_n4440, new_n4441_1, new_n4442, new_n4443,
    new_n4444, new_n4445, new_n4446, new_n4447, new_n4448, new_n4449,
    new_n4450, new_n4451_1, new_n4452, new_n4453, new_n4454, new_n4455,
    new_n4456, new_n4457, new_n4458, new_n4459, new_n4460, new_n4461,
    new_n4462, new_n4463, new_n4464, new_n4465, new_n4466, new_n4467,
    new_n4468, new_n4469, new_n4470, new_n4471, new_n4472, new_n4473,
    new_n4474, new_n4475, new_n4476_1, new_n4477, new_n4478_1, new_n4479,
    new_n4480, new_n4481, new_n4482, new_n4483, new_n4484, new_n4485,
    new_n4486, new_n4487, new_n4488, new_n4489, new_n4490, new_n4491,
    new_n4492, new_n4493, new_n4494, new_n4495, new_n4496, new_n4497,
    new_n4498, new_n4499, new_n4500, new_n4501, new_n4502, new_n4503,
    new_n4504, new_n4505, new_n4506, new_n4507, new_n4508, new_n4509,
    new_n4510, new_n4511, new_n4512, new_n4513, new_n4514_1, new_n4515,
    new_n4516, new_n4517, new_n4518, new_n4519, new_n4520, new_n4521,
    new_n4522, new_n4523, new_n4524, new_n4525, new_n4526, new_n4527,
    new_n4528, new_n4529_1, new_n4530, new_n4531, new_n4532, new_n4533,
    new_n4534, new_n4535, new_n4536, new_n4537, new_n4538, new_n4539,
    new_n4540, new_n4541, new_n4542, new_n4543, new_n4544, new_n4545,
    new_n4546, new_n4547, new_n4548, new_n4549, new_n4550, new_n4551,
    new_n4552_1, new_n4553, new_n4554, new_n4555, new_n4556, new_n4557,
    new_n4558, new_n4559, new_n4560, new_n4561, new_n4562, new_n4563,
    new_n4564, new_n4565, new_n4566, new_n4567, new_n4568, new_n4569,
    new_n4570, new_n4571, new_n4572, new_n4573, new_n4574, new_n4575,
    new_n4576, new_n4577, new_n4578, new_n4579, new_n4580, new_n4581,
    new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587,
    new_n4588_1, new_n4589, new_n4591, new_n4592, new_n4593, new_n4594,
    new_n4595_1, new_n4596, new_n4597, new_n4598, new_n4599, new_n4600,
    new_n4601, new_n4602, new_n4603, new_n4604, new_n4605, new_n4606,
    new_n4607, new_n4608, new_n4609, new_n4610, new_n4611, new_n4612,
    new_n4613, new_n4614, new_n4615, new_n4616, new_n4617, new_n4618,
    new_n4619, new_n4620, new_n4621, new_n4622, new_n4623, new_n4624_1,
    new_n4625, new_n4626, new_n4627, new_n4628, new_n4629, new_n4630,
    new_n4631, new_n4632, new_n4633, new_n4634, new_n4635, new_n4636,
    new_n4637, new_n4638, new_n4639, new_n4640, new_n4641, new_n4642,
    new_n4643, new_n4644, new_n4645, new_n4646_1, new_n4647, new_n4648,
    new_n4649, new_n4650, new_n4651, new_n4652, new_n4653, new_n4654,
    new_n4655, new_n4656, new_n4657, new_n4658, new_n4659, new_n4660,
    new_n4661, new_n4662, new_n4663, new_n4664, new_n4665_1, new_n4666,
    new_n4668, new_n4669, new_n4670, new_n4671, new_n4672, new_n4673,
    new_n4674_1, new_n4675, new_n4676, new_n4677, new_n4678, new_n4679,
    new_n4680, new_n4681, new_n4682, new_n4683, new_n4684, new_n4685,
    new_n4686, new_n4687, new_n4688, new_n4689, new_n4690, new_n4691,
    new_n4692, new_n4693_1, new_n4694, new_n4695, new_n4696, new_n4697,
    new_n4698, new_n4699, new_n4700, new_n4701, new_n4702, new_n4703,
    new_n4704, new_n4705, new_n4706, new_n4707, new_n4708, new_n4709,
    new_n4710, new_n4711, new_n4712, new_n4713, new_n4714, new_n4715,
    new_n4716, new_n4717, new_n4718, new_n4719, new_n4720, new_n4721,
    new_n4722_1, new_n4723, new_n4724, new_n4725, new_n4726, new_n4727,
    new_n4728, new_n4729, new_n4730, new_n4731_1, new_n4732, new_n4733,
    new_n4734, new_n4735, new_n4736, new_n4737, new_n4738, new_n4739,
    new_n4740, new_n4741, new_n4742, new_n4743, new_n4744, new_n4745_1,
    new_n4746, new_n4747_1, new_n4748, new_n4749, new_n4750, new_n4751,
    new_n4752, new_n4753, new_n4754, new_n4755, new_n4756, new_n4757,
    new_n4758, new_n4759, new_n4760, new_n4761, new_n4762, new_n4763,
    new_n4764, new_n4765, new_n4766_1, new_n4767, new_n4768, new_n4769,
    new_n4770_1, new_n4771, new_n4772, new_n4773, new_n4774, new_n4775,
    new_n4776, new_n4777_1, new_n4778, new_n4779, new_n4780, new_n4781,
    new_n4782, new_n4783, new_n4784, new_n4785_1, new_n4786, new_n4787,
    new_n4788, new_n4789, new_n4790, new_n4791, new_n4792, new_n4793,
    new_n4794, new_n4795, new_n4796, new_n4797, new_n4798, new_n4799,
    new_n4800, new_n4801, new_n4802, new_n4803, new_n4804_1, new_n4805,
    new_n4806, new_n4807, new_n4808, new_n4809, new_n4810_1, new_n4811,
    new_n4812_1, new_n4813, new_n4814_1, new_n4815, new_n4816, new_n4817,
    new_n4818, new_n4819, new_n4820, new_n4821, new_n4822, new_n4823,
    new_n4824, new_n4825, new_n4826, new_n4827, new_n4828, new_n4829,
    new_n4830, new_n4831, new_n4832, new_n4833, new_n4834, new_n4835,
    new_n4836, new_n4837, new_n4838, new_n4839, new_n4840, new_n4841,
    new_n4842, new_n4843, new_n4844, new_n4845, new_n4846, new_n4847,
    new_n4848, new_n4849, new_n4850_1, new_n4851, new_n4853, new_n4854,
    new_n4855, new_n4856, new_n4857, new_n4858_1, new_n4859, new_n4860,
    new_n4861, new_n4862, new_n4863, new_n4864, new_n4865, new_n4866,
    new_n4867, new_n4868, new_n4869, new_n4870, new_n4871, new_n4872,
    new_n4873, new_n4874, new_n4875, new_n4876, new_n4877, new_n4878,
    new_n4879, new_n4880, new_n4881, new_n4882, new_n4883, new_n4884,
    new_n4885, new_n4886, new_n4887, new_n4888, new_n4889, new_n4890,
    new_n4891_1, new_n4892, new_n4893, new_n4894, new_n4895, new_n4896,
    new_n4897, new_n4898, new_n4899, new_n4900, new_n4901, new_n4902,
    new_n4903, new_n4904, new_n4905, new_n4906, new_n4907, new_n4908,
    new_n4909, new_n4910, new_n4911, new_n4912, new_n4913_1, new_n4914,
    new_n4915, new_n4916, new_n4917, new_n4918, new_n4919, new_n4920,
    new_n4921, new_n4922, new_n4923, new_n4924, new_n4925_1, new_n4926,
    new_n4927, new_n4928, new_n4929, new_n4930, new_n4931, new_n4932,
    new_n4933, new_n4934, new_n4935, new_n4936, new_n4937, new_n4938,
    new_n4939_1, new_n4940, new_n4941, new_n4942, new_n4943, new_n4944,
    new_n4945, new_n4946, new_n4947_1, new_n4948, new_n4949, new_n4950,
    new_n4951, new_n4952_1, new_n4953, new_n4954, new_n4955, new_n4956,
    new_n4957_1, new_n4958, new_n4959, new_n4960, new_n4961, new_n4962,
    new_n4963, new_n4964_1, new_n4965, new_n4966_1, new_n4967_1, new_n4968,
    new_n4969, new_n4970, new_n4971, new_n4972_1, new_n4973, new_n4974,
    new_n4975, new_n4976, new_n4977, new_n4978, new_n4979, new_n4980,
    new_n4981, new_n4982, new_n4983, new_n4984, new_n4985, new_n4986,
    new_n4987, new_n4988, new_n4989, new_n4990, new_n4991, new_n4992,
    new_n4993, new_n4994, new_n4995, new_n4996, new_n4997, new_n4998,
    new_n4999, new_n5000, new_n5001, new_n5002, new_n5003, new_n5004,
    new_n5005, new_n5006, new_n5007, new_n5008, new_n5009, new_n5010,
    new_n5011_1, new_n5012, new_n5013, new_n5014, new_n5015, new_n5016,
    new_n5017, new_n5018, new_n5019, new_n5020_1, new_n5021, new_n5022,
    new_n5023, new_n5024_1, new_n5025_1, new_n5026_1, new_n5027, new_n5028,
    new_n5029, new_n5030, new_n5031_1, new_n5032, new_n5033, new_n5034,
    new_n5035, new_n5036, new_n5037, new_n5038, new_n5039, new_n5040,
    new_n5041, new_n5042, new_n5043, new_n5044, new_n5045, new_n5046_1,
    new_n5047, new_n5048, new_n5049, new_n5050, new_n5051, new_n5052,
    new_n5053, new_n5054, new_n5055, new_n5056, new_n5057, new_n5058,
    new_n5059, new_n5060_1, new_n5061, new_n5062_1, new_n5063, new_n5064_1,
    new_n5065, new_n5066, new_n5067, new_n5068, new_n5069, new_n5070,
    new_n5071, new_n5072, new_n5073, new_n5074, new_n5075, new_n5076,
    new_n5077_1, new_n5078, new_n5079, new_n5080, new_n5081, new_n5082_1,
    new_n5083, new_n5084, new_n5085, new_n5086, new_n5087, new_n5088,
    new_n5089, new_n5090, new_n5091, new_n5092, new_n5093, new_n5094,
    new_n5095, new_n5096, new_n5097, new_n5098_1, new_n5099, new_n5100,
    new_n5101_1, new_n5102, new_n5103, new_n5104, new_n5105, new_n5106,
    new_n5107, new_n5108, new_n5109, new_n5110, new_n5111, new_n5112,
    new_n5113, new_n5114, new_n5115_1, new_n5116, new_n5117, new_n5118,
    new_n5119, new_n5120_1, new_n5121, new_n5122, new_n5123, new_n5124,
    new_n5125, new_n5126, new_n5127, new_n5128_1, new_n5129, new_n5130,
    new_n5131_1, new_n5132, new_n5133, new_n5134, new_n5135, new_n5136,
    new_n5137, new_n5138, new_n5139, new_n5140_1, new_n5141, new_n5142,
    new_n5143, new_n5144, new_n5145, new_n5146, new_n5147, new_n5148,
    new_n5149, new_n5150, new_n5151, new_n5152, new_n5153, new_n5154,
    new_n5155, new_n5156, new_n5157, new_n5158_1, new_n5159, new_n5160,
    new_n5161, new_n5162, new_n5163, new_n5164, new_n5165, new_n5166,
    new_n5167, new_n5168_1, new_n5169, new_n5170, new_n5171, new_n5172,
    new_n5173, new_n5174, new_n5175, new_n5176, new_n5177, new_n5178,
    new_n5179, new_n5180, new_n5181, new_n5182, new_n5183, new_n5184_1,
    new_n5185, new_n5186, new_n5187, new_n5188, new_n5189, new_n5190,
    new_n5191, new_n5192, new_n5193, new_n5194, new_n5195, new_n5196,
    new_n5197, new_n5198, new_n5199, new_n5200, new_n5201, new_n5202,
    new_n5203, new_n5204, new_n5205, new_n5206, new_n5207, new_n5208,
    new_n5209, new_n5210, new_n5211_1, new_n5212, new_n5213_1, new_n5214,
    new_n5215, new_n5216, new_n5217, new_n5218, new_n5219, new_n5220,
    new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226_1,
    new_n5227, new_n5229, new_n5230, new_n5231, new_n5232, new_n5233,
    new_n5234, new_n5235, new_n5236, new_n5237, new_n5238, new_n5239,
    new_n5240, new_n5241, new_n5242, new_n5243, new_n5244, new_n5245,
    new_n5246, new_n5247, new_n5248, new_n5249, new_n5250, new_n5251,
    new_n5252, new_n5253, new_n5254, new_n5255_1, new_n5256_1, new_n5257,
    new_n5258, new_n5259, new_n5260, new_n5261, new_n5262, new_n5263,
    new_n5264, new_n5265_1, new_n5266, new_n5267, new_n5268, new_n5269,
    new_n5270, new_n5271, new_n5272, new_n5273_1, new_n5274_1, new_n5275,
    new_n5276, new_n5277, new_n5278, new_n5279, new_n5280, new_n5281,
    new_n5282, new_n5283, new_n5284, new_n5285, new_n5286, new_n5287,
    new_n5288, new_n5289, new_n5290, new_n5291, new_n5292, new_n5293,
    new_n5294, new_n5295, new_n5296, new_n5297, new_n5298, new_n5299,
    new_n5300_1, new_n5301, new_n5302_1, new_n5303, new_n5304, new_n5305,
    new_n5306, new_n5307, new_n5308, new_n5309, new_n5310, new_n5311,
    new_n5312, new_n5313, new_n5314, new_n5315, new_n5316, new_n5317,
    new_n5318, new_n5319, new_n5320, new_n5321, new_n5322, new_n5323,
    new_n5324, new_n5325_1, new_n5326, new_n5327, new_n5328, new_n5329,
    new_n5330_1, new_n5331, new_n5332, new_n5333, new_n5334, new_n5335,
    new_n5336, new_n5337_1, new_n5338, new_n5339, new_n5340, new_n5341,
    new_n5342, new_n5343, new_n5344, new_n5345, new_n5346, new_n5347,
    new_n5348, new_n5349, new_n5350, new_n5351_1, new_n5352, new_n5353_1,
    new_n5354, new_n5355, new_n5356, new_n5357, new_n5358, new_n5359,
    new_n5360, new_n5361, new_n5362, new_n5363, new_n5364, new_n5365,
    new_n5366, new_n5367, new_n5368, new_n5369, new_n5370, new_n5371,
    new_n5372, new_n5373, new_n5374, new_n5375, new_n5376_1, new_n5377,
    new_n5378, new_n5379, new_n5380, new_n5381, new_n5382, new_n5383,
    new_n5384, new_n5385, new_n5386_1, new_n5387, new_n5388, new_n5389,
    new_n5390, new_n5391, new_n5392, new_n5393, new_n5394, new_n5395,
    new_n5396, new_n5397, new_n5398, new_n5399_1, new_n5400_1, new_n5401,
    new_n5402, new_n5403_1, new_n5404, new_n5405, new_n5406, new_n5407,
    new_n5408, new_n5409, new_n5410, new_n5411, new_n5412, new_n5413,
    new_n5414, new_n5415, new_n5417, new_n5418, new_n5419, new_n5420,
    new_n5421, new_n5422, new_n5423, new_n5424, new_n5425, new_n5426,
    new_n5427, new_n5428, new_n5429, new_n5430_1, new_n5431, new_n5432,
    new_n5433, new_n5434, new_n5435, new_n5436, new_n5437, new_n5438_1,
    new_n5439_1, new_n5440, new_n5441, new_n5442, new_n5443_1, new_n5444,
    new_n5445, new_n5446, new_n5447, new_n5448, new_n5449, new_n5450,
    new_n5451_1, new_n5452, new_n5453, new_n5454, new_n5455, new_n5456,
    new_n5457, new_n5458, new_n5459, new_n5460, new_n5461, new_n5462,
    new_n5463, new_n5464, new_n5465, new_n5466, new_n5467, new_n5468,
    new_n5469, new_n5470, new_n5471, new_n5472_1, new_n5473, new_n5474,
    new_n5475, new_n5476, new_n5477, new_n5478, new_n5479, new_n5480,
    new_n5481, new_n5482, new_n5483, new_n5484, new_n5485_1, new_n5486,
    new_n5487, new_n5488, new_n5489, new_n5490, new_n5491, new_n5492,
    new_n5493, new_n5494, new_n5495, new_n5496, new_n5497, new_n5498,
    new_n5499, new_n5500, new_n5501, new_n5502, new_n5503, new_n5504,
    new_n5505, new_n5506, new_n5507, new_n5508, new_n5509, new_n5510,
    new_n5511, new_n5512, new_n5513, new_n5514, new_n5515, new_n5516,
    new_n5517_1, new_n5518, new_n5519, new_n5520, new_n5521_1, new_n5522,
    new_n5523, new_n5524_1, new_n5525, new_n5526, new_n5527, new_n5528,
    new_n5529, new_n5530, new_n5531, new_n5532_1, new_n5533, new_n5534,
    new_n5535, new_n5536, new_n5537, new_n5538, new_n5539, new_n5540,
    new_n5541, new_n5542, new_n5543, new_n5544, new_n5545, new_n5546,
    new_n5547, new_n5548, new_n5549, new_n5550, new_n5551, new_n5552,
    new_n5553, new_n5554, new_n5555, new_n5556, new_n5557, new_n5558,
    new_n5559, new_n5560, new_n5561, new_n5562, new_n5563, new_n5564_1,
    new_n5565, new_n5566, new_n5567, new_n5568, new_n5569, new_n5570,
    new_n5571, new_n5572, new_n5573, new_n5574, new_n5575, new_n5576,
    new_n5577, new_n5578, new_n5579_1, new_n5580, new_n5581, new_n5582,
    new_n5583, new_n5584, new_n5585, new_n5586, new_n5587, new_n5588,
    new_n5589, new_n5590, new_n5591, new_n5592, new_n5593_1, new_n5594,
    new_n5595, new_n5596, new_n5597, new_n5598, new_n5599, new_n5600,
    new_n5601, new_n5602, new_n5603_1, new_n5604, new_n5605_1, new_n5606,
    new_n5607, new_n5608, new_n5609_1, new_n5610, new_n5611, new_n5612,
    new_n5613, new_n5614, new_n5615, new_n5616, new_n5617, new_n5618,
    new_n5619, new_n5620, new_n5621, new_n5622, new_n5623, new_n5624,
    new_n5625, new_n5626, new_n5627, new_n5628, new_n5629, new_n5630,
    new_n5631, new_n5632, new_n5633, new_n5634_1, new_n5635, new_n5636,
    new_n5637, new_n5638, new_n5639, new_n5640, new_n5641, new_n5642,
    new_n5643_1, new_n5644, new_n5645, new_n5646, new_n5647, new_n5648,
    new_n5649, new_n5650, new_n5651, new_n5652, new_n5653, new_n5654,
    new_n5655, new_n5656, new_n5657, new_n5658, new_n5659, new_n5660,
    new_n5661, new_n5662, new_n5663, new_n5664, new_n5665, new_n5666,
    new_n5667, new_n5668, new_n5669, new_n5670, new_n5671, new_n5672,
    new_n5673, new_n5674, new_n5675, new_n5676, new_n5677, new_n5678,
    new_n5679, new_n5680_1, new_n5681, new_n5682, new_n5683, new_n5684,
    new_n5685, new_n5686, new_n5687_1, new_n5688, new_n5689, new_n5690,
    new_n5691, new_n5692, new_n5693, new_n5694, new_n5695, new_n5696_1,
    new_n5697, new_n5698, new_n5699, new_n5700_1, new_n5701, new_n5702,
    new_n5703, new_n5704_1, new_n5705, new_n5706, new_n5707, new_n5708,
    new_n5709, new_n5710, new_n5711, new_n5712, new_n5713, new_n5714,
    new_n5715, new_n5716, new_n5717, new_n5718, new_n5719, new_n5720,
    new_n5721, new_n5722, new_n5723, new_n5724, new_n5725, new_n5726,
    new_n5727, new_n5728, new_n5729, new_n5730, new_n5731, new_n5732_1,
    new_n5733, new_n5734, new_n5735, new_n5736, new_n5737, new_n5738,
    new_n5739, new_n5740, new_n5741, new_n5742_1, new_n5743, new_n5744,
    new_n5745, new_n5746, new_n5747, new_n5748, new_n5749, new_n5750,
    new_n5751, new_n5752_1, new_n5753, new_n5754, new_n5755, new_n5757,
    new_n5758, new_n5759, new_n5760, new_n5761, new_n5762, new_n5763,
    new_n5764, new_n5765_1, new_n5766, new_n5767, new_n5768, new_n5769,
    new_n5770, new_n5771, new_n5772, new_n5773, new_n5774, new_n5775,
    new_n5776_1, new_n5777, new_n5778, new_n5779, new_n5780, new_n5781,
    new_n5782_1, new_n5783, new_n5784, new_n5785, new_n5786, new_n5787,
    new_n5788, new_n5789, new_n5790, new_n5791, new_n5792, new_n5793,
    new_n5794, new_n5795, new_n5796, new_n5797, new_n5798, new_n5799,
    new_n5800, new_n5801, new_n5802, new_n5803, new_n5804, new_n5805,
    new_n5806, new_n5807, new_n5808, new_n5809, new_n5810, new_n5811,
    new_n5812, new_n5813, new_n5814, new_n5815, new_n5816, new_n5817,
    new_n5818, new_n5819, new_n5820, new_n5821, new_n5822_1, new_n5823,
    new_n5824, new_n5825, new_n5826, new_n5827, new_n5828, new_n5829,
    new_n5830, new_n5831, new_n5832, new_n5833_1, new_n5834_1, new_n5835,
    new_n5836, new_n5837, new_n5838, new_n5839, new_n5840_1, new_n5841_1,
    new_n5842_1, new_n5843, new_n5844, new_n5845, new_n5846, new_n5847,
    new_n5848, new_n5849, new_n5850_1, new_n5851, new_n5852, new_n5853,
    new_n5854, new_n5855, new_n5856, new_n5857, new_n5859, new_n5860,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882_1, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903_1, new_n5904_1, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911_1, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934, new_n5935, new_n5936_1, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5943_1, new_n5944,
    new_n5945, new_n5946, new_n5947, new_n5948, new_n5949, new_n5950,
    new_n5951, new_n5952, new_n5953, new_n5954, new_n5955, new_n5956,
    new_n5957, new_n5958, new_n5959, new_n5960, new_n5961, new_n5962,
    new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968,
    new_n5969, new_n5970, new_n5971, new_n5972, new_n5973, new_n5974,
    new_n5975, new_n5976, new_n5977, new_n5978, new_n5979, new_n5980_1,
    new_n5981, new_n5982, new_n5983, new_n5984, new_n5985, new_n5986,
    new_n5987, new_n5988, new_n5989, new_n5990, new_n5991, new_n5992,
    new_n5993, new_n5994, new_n5995, new_n5996, new_n5997, new_n5998,
    new_n5999, new_n6000, new_n6001, new_n6002, new_n6003, new_n6004,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012_1, new_n6013, new_n6014, new_n6015, new_n6016, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022_1, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031_1, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044_1, new_n6045, new_n6046_1, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084_1, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104_1, new_n6105_1, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160_1, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171_1, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183_1, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189_1, new_n6190, new_n6191,
    new_n6192, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204_1, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218_1, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223_1, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233_1,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245_1,
    new_n6246, new_n6247, new_n6248_1, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254, new_n6255, new_n6256_1, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271_1, new_n6272, new_n6273, new_n6274, new_n6275,
    new_n6276_1, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281,
    new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287,
    new_n6288, new_n6289, new_n6290, new_n6291, new_n6292, new_n6293,
    new_n6294, new_n6295, new_n6296, new_n6297, new_n6298, new_n6299,
    new_n6300, new_n6301, new_n6302, new_n6303, new_n6304, new_n6305,
    new_n6306, new_n6307, new_n6308_1, new_n6309, new_n6310, new_n6311_1,
    new_n6312, new_n6313, new_n6314, new_n6315, new_n6316, new_n6317,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323_1, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330_1,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339_1, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354_1,
    new_n6355, new_n6356_1, new_n6357, new_n6358, new_n6359, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369_1, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375_1, new_n6376, new_n6377, new_n6378,
    new_n6379_1, new_n6380, new_n6381_1, new_n6382, new_n6383_1, new_n6384,
    new_n6385_1, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397_1, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407_1, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427_1, new_n6428, new_n6429, new_n6430, new_n6431_1, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437_1, new_n6438,
    new_n6439, new_n6440, new_n6441, new_n6442, new_n6443, new_n6444,
    new_n6445, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456_1,
    new_n6457_1, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465_1, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470_1, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476_1, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485_1, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502_1, new_n6503, new_n6504,
    new_n6505, new_n6506_1, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513_1, new_n6514_1, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6527, new_n6528,
    new_n6529, new_n6530, new_n6531, new_n6532, new_n6533, new_n6534,
    new_n6535, new_n6536, new_n6537, new_n6538, new_n6539, new_n6540,
    new_n6541, new_n6542_1, new_n6543, new_n6544, new_n6545, new_n6546,
    new_n6547, new_n6548, new_n6549, new_n6550, new_n6551, new_n6552,
    new_n6553, new_n6554, new_n6555, new_n6556_1, new_n6557, new_n6558_1,
    new_n6559, new_n6560_1, new_n6561, new_n6562, new_n6563, new_n6564,
    new_n6565, new_n6566, new_n6567_1, new_n6568, new_n6569, new_n6570,
    new_n6571, new_n6572, new_n6573, new_n6574, new_n6575, new_n6576_1,
    new_n6577, new_n6578, new_n6579, new_n6580, new_n6581, new_n6582,
    new_n6583, new_n6584, new_n6585, new_n6586, new_n6587_1, new_n6588,
    new_n6589, new_n6590_1, new_n6591, new_n6592, new_n6593, new_n6594,
    new_n6595, new_n6596_1, new_n6597, new_n6598, new_n6599, new_n6600,
    new_n6601, new_n6602, new_n6603, new_n6604, new_n6605, new_n6606,
    new_n6607, new_n6608, new_n6609, new_n6610, new_n6611_1, new_n6612_1,
    new_n6613, new_n6614, new_n6615, new_n6616, new_n6617, new_n6618,
    new_n6619, new_n6620, new_n6621, new_n6622, new_n6623, new_n6624,
    new_n6625, new_n6626, new_n6627, new_n6628_1, new_n6629, new_n6630_1,
    new_n6631_1, new_n6632, new_n6633, new_n6634_1, new_n6635, new_n6636,
    new_n6637, new_n6638, new_n6639, new_n6640, new_n6641, new_n6642,
    new_n6643, new_n6644, new_n6645, new_n6646, new_n6647, new_n6648,
    new_n6649, new_n6650, new_n6651, new_n6652_1, new_n6653, new_n6654,
    new_n6655_1, new_n6656, new_n6657, new_n6658, new_n6659_1, new_n6660,
    new_n6661, new_n6662, new_n6663, new_n6664, new_n6665, new_n6666,
    new_n6667, new_n6668, new_n6669_1, new_n6670, new_n6671_1, new_n6672,
    new_n6673_1, new_n6674_1, new_n6675, new_n6676, new_n6677, new_n6678,
    new_n6679, new_n6680, new_n6681, new_n6682, new_n6683, new_n6684_1,
    new_n6685, new_n6686, new_n6687, new_n6688, new_n6689, new_n6690,
    new_n6691_1, new_n6692, new_n6693, new_n6694, new_n6695, new_n6696,
    new_n6697, new_n6698, new_n6699, new_n6700, new_n6701, new_n6702,
    new_n6703, new_n6704, new_n6705, new_n6706_1, new_n6707_1, new_n6708,
    new_n6709, new_n6710, new_n6711, new_n6712, new_n6713, new_n6714,
    new_n6715, new_n6716, new_n6717, new_n6718, new_n6719, new_n6720,
    new_n6722, new_n6723, new_n6724, new_n6725, new_n6726, new_n6727,
    new_n6728, new_n6729_1, new_n6730, new_n6731, new_n6732, new_n6733,
    new_n6734, new_n6735, new_n6736_1, new_n6737, new_n6738, new_n6739,
    new_n6740, new_n6741, new_n6742, new_n6743, new_n6744, new_n6745,
    new_n6746, new_n6747, new_n6748, new_n6749, new_n6750, new_n6751,
    new_n6752, new_n6753, new_n6754, new_n6755, new_n6756, new_n6757,
    new_n6758, new_n6759, new_n6760, new_n6761, new_n6762, new_n6763,
    new_n6764, new_n6766, new_n6767, new_n6768, new_n6769, new_n6770,
    new_n6771, new_n6772, new_n6773_1, new_n6775_1, new_n6777, new_n6778,
    new_n6779, new_n6780, new_n6781, new_n6782, new_n6783, new_n6784,
    new_n6785_1, new_n6786, new_n6787, new_n6788, new_n6789, new_n6790_1,
    new_n6791_1, new_n6792, new_n6793, new_n6794_1, new_n6795, new_n6796,
    new_n6797, new_n6798, new_n6799, new_n6800, new_n6801, new_n6802_1,
    new_n6803, new_n6804, new_n6805, new_n6806, new_n6807, new_n6808,
    new_n6809, new_n6810, new_n6811, new_n6812, new_n6813, new_n6814_1,
    new_n6815, new_n6816, new_n6818, new_n6819, new_n6820, new_n6821,
    new_n6822, new_n6823, new_n6824, new_n6825, new_n6826_1, new_n6827,
    new_n6828, new_n6829, new_n6830, new_n6831, new_n6832, new_n6833,
    new_n6834, new_n6835_1, new_n6836, new_n6837, new_n6838, new_n6839,
    new_n6840, new_n6841, new_n6842, new_n6843, new_n6844, new_n6845,
    new_n6846, new_n6847, new_n6848, new_n6849, new_n6850, new_n6851,
    new_n6852, new_n6853_1, new_n6854, new_n6855, new_n6856, new_n6857,
    new_n6858, new_n6859, new_n6863_1, new_n6864, new_n6865, new_n6866,
    new_n6867_1, new_n6868, new_n6869, new_n6870, new_n6871, new_n6872,
    new_n6873, new_n6874, new_n6875, new_n6876, new_n6877, new_n6878,
    new_n6879, new_n6880, new_n6881, new_n6882, new_n6883, new_n6884,
    new_n6885, new_n6886, new_n6887, new_n6888, new_n6889, new_n6890,
    new_n6891, new_n6892, new_n6893, new_n6894, new_n6895, new_n6896,
    new_n6897, new_n6898, new_n6899, new_n6900, new_n6901, new_n6902,
    new_n6903, new_n6904, new_n6905, new_n6906, new_n6907, new_n6908,
    new_n6909, new_n6910, new_n6911, new_n6912, new_n6913, new_n6914,
    new_n6915, new_n6916, new_n6917, new_n6918, new_n6919, new_n6920,
    new_n6921, new_n6922, new_n6923, new_n6924, new_n6925, new_n6926,
    new_n6927, new_n6928, new_n6929, new_n6930, new_n6931, new_n6932,
    new_n6933, new_n6934, new_n6935, new_n6936, new_n6937, new_n6938,
    new_n6939, new_n6940, new_n6941, new_n6942, new_n6943, new_n6944,
    new_n6945, new_n6946, new_n6947, new_n6948, new_n6949, new_n6950,
    new_n6951, new_n6952, new_n6953, new_n6954, new_n6955, new_n6956,
    new_n6957, new_n6958, new_n6959, new_n6960, new_n6961, new_n6962,
    new_n6963, new_n6964, new_n6965_1, new_n6966, new_n6967_1, new_n6968,
    new_n6969, new_n6970, new_n6971_1, new_n6972, new_n6973, new_n6974,
    new_n6975_1, new_n6976, new_n6977, new_n6978, new_n6979, new_n6980,
    new_n6981, new_n6982, new_n6983_1, new_n6984, new_n6985_1, new_n6986,
    new_n6987, new_n6988, new_n6989, new_n6990, new_n6991, new_n6992,
    new_n6993, new_n6994, new_n6995, new_n6996, new_n6997, new_n6998_1,
    new_n6999, new_n7000, new_n7001, new_n7002, new_n7003, new_n7004,
    new_n7005, new_n7006, new_n7007, new_n7008, new_n7009, new_n7010,
    new_n7011, new_n7012, new_n7013, new_n7014, new_n7015, new_n7016,
    new_n7017, new_n7018, new_n7019, new_n7020, new_n7021, new_n7022,
    new_n7023, new_n7024, new_n7025, new_n7026_1, new_n7027, new_n7028,
    new_n7029, new_n7030, new_n7031, new_n7032_1, new_n7033, new_n7034,
    new_n7035, new_n7036, new_n7037, new_n7038_1, new_n7039, new_n7040,
    new_n7041, new_n7042, new_n7043, new_n7044, new_n7045, new_n7046,
    new_n7047, new_n7048, new_n7049, new_n7050, new_n7051, new_n7052,
    new_n7053, new_n7054, new_n7055, new_n7056, new_n7057_1, new_n7058,
    new_n7059, new_n7060, new_n7061, new_n7062, new_n7063, new_n7064,
    new_n7065, new_n7066, new_n7067, new_n7068, new_n7069, new_n7070,
    new_n7071, new_n7072, new_n7073, new_n7074, new_n7075, new_n7076,
    new_n7077, new_n7078, new_n7079_1, new_n7080, new_n7081, new_n7082,
    new_n7083, new_n7084, new_n7085, new_n7086, new_n7087, new_n7088,
    new_n7089, new_n7090, new_n7091, new_n7092, new_n7093, new_n7094,
    new_n7095, new_n7096, new_n7097, new_n7098, new_n7099_1, new_n7100,
    new_n7101, new_n7102, new_n7103, new_n7104, new_n7105, new_n7106,
    new_n7107, new_n7108, new_n7109, new_n7110, new_n7111, new_n7112,
    new_n7113, new_n7114, new_n7115, new_n7116, new_n7117, new_n7118,
    new_n7119, new_n7120, new_n7121, new_n7122, new_n7123, new_n7124,
    new_n7125, new_n7126, new_n7127, new_n7128, new_n7129, new_n7130,
    new_n7131, new_n7132, new_n7133, new_n7134, new_n7135, new_n7136,
    new_n7137, new_n7138, new_n7139_1, new_n7140, new_n7141, new_n7142,
    new_n7143, new_n7144, new_n7145, new_n7146, new_n7147, new_n7148,
    new_n7149_1, new_n7150, new_n7151, new_n7152, new_n7153, new_n7154,
    new_n7155, new_n7156, new_n7157, new_n7158, new_n7159, new_n7160,
    new_n7161, new_n7162, new_n7163, new_n7164, new_n7165, new_n7166,
    new_n7167, new_n7168, new_n7169, new_n7170, new_n7171, new_n7172,
    new_n7173, new_n7174, new_n7175, new_n7176, new_n7177, new_n7178,
    new_n7179, new_n7180, new_n7181, new_n7182, new_n7183, new_n7184,
    new_n7185, new_n7186, new_n7187, new_n7188, new_n7189, new_n7190_1,
    new_n7191, new_n7192, new_n7193, new_n7194, new_n7195, new_n7196,
    new_n7197, new_n7198, new_n7200, new_n7201, new_n7202, new_n7203,
    new_n7204, new_n7205, new_n7206, new_n7207, new_n7208, new_n7209,
    new_n7210, new_n7211, new_n7212, new_n7213, new_n7214, new_n7215,
    new_n7216, new_n7217, new_n7218, new_n7219, new_n7220, new_n7221,
    new_n7222, new_n7223, new_n7224, new_n7225, new_n7226, new_n7227,
    new_n7228, new_n7229_1, new_n7230_1, new_n7231, new_n7232, new_n7233_1,
    new_n7234, new_n7235, new_n7236_1, new_n7237, new_n7238, new_n7239,
    new_n7240, new_n7241, new_n7242, new_n7243, new_n7244, new_n7245,
    new_n7246, new_n7247, new_n7248, new_n7249, new_n7250, new_n7251,
    new_n7252, new_n7253_1, new_n7254, new_n7255, new_n7256_1, new_n7257,
    new_n7258, new_n7259, new_n7260, new_n7261, new_n7262, new_n7263,
    new_n7264, new_n7265, new_n7266, new_n7267, new_n7268_1, new_n7269,
    new_n7270, new_n7271, new_n7272, new_n7273, new_n7274, new_n7275,
    new_n7276, new_n7277_1, new_n7278, new_n7279, new_n7280_1, new_n7281,
    new_n7282, new_n7283, new_n7284, new_n7285, new_n7286, new_n7287,
    new_n7288, new_n7289, new_n7290, new_n7291, new_n7292, new_n7293,
    new_n7294, new_n7295, new_n7296, new_n7297, new_n7298_1, new_n7299,
    new_n7300, new_n7301, new_n7302, new_n7303, new_n7304, new_n7305_1,
    new_n7306, new_n7307, new_n7308_1, new_n7309, new_n7310, new_n7311,
    new_n7312, new_n7313_1, new_n7314, new_n7315, new_n7316, new_n7317,
    new_n7318, new_n7319, new_n7320, new_n7321, new_n7322, new_n7323,
    new_n7324, new_n7325, new_n7326, new_n7327, new_n7328, new_n7329,
    new_n7330_1, new_n7331, new_n7332, new_n7333, new_n7334, new_n7335_1,
    new_n7336, new_n7337, new_n7338, new_n7339_1, new_n7340, new_n7341,
    new_n7342, new_n7343, new_n7344, new_n7345, new_n7346_1, new_n7347,
    new_n7348, new_n7349_1, new_n7350, new_n7351, new_n7352, new_n7353,
    new_n7354, new_n7355, new_n7356, new_n7357, new_n7358, new_n7359,
    new_n7360, new_n7361, new_n7362, new_n7363_1, new_n7364, new_n7365,
    new_n7366, new_n7367, new_n7368, new_n7369, new_n7370, new_n7371,
    new_n7372, new_n7373, new_n7374, new_n7375, new_n7376, new_n7377_1,
    new_n7378, new_n7379, new_n7380, new_n7381, new_n7382, new_n7383,
    new_n7384, new_n7385, new_n7386, new_n7387, new_n7388, new_n7389,
    new_n7390_1, new_n7391, new_n7392, new_n7393, new_n7394, new_n7395,
    new_n7396, new_n7397, new_n7398, new_n7399, new_n7400, new_n7401,
    new_n7402, new_n7403_1, new_n7404, new_n7405, new_n7406, new_n7407,
    new_n7408_1, new_n7409, new_n7410, new_n7411, new_n7412, new_n7413,
    new_n7414, new_n7415, new_n7416, new_n7417, new_n7418, new_n7419,
    new_n7420, new_n7421_1, new_n7422, new_n7423, new_n7424, new_n7425,
    new_n7426, new_n7427, new_n7428_1, new_n7429, new_n7430, new_n7431,
    new_n7432_1, new_n7433, new_n7434, new_n7435, new_n7436, new_n7437_1,
    new_n7438, new_n7439, new_n7440, new_n7441, new_n7442, new_n7443,
    new_n7444, new_n7445, new_n7446, new_n7447, new_n7448, new_n7449,
    new_n7450, new_n7451, new_n7452, new_n7453, new_n7454, new_n7455,
    new_n7456, new_n7457, new_n7458, new_n7459, new_n7460_1, new_n7461,
    new_n7462, new_n7463, new_n7464, new_n7465, new_n7466, new_n7467,
    new_n7468, new_n7469, new_n7470, new_n7471, new_n7472, new_n7473,
    new_n7474, new_n7475_1, new_n7476, new_n7477_1, new_n7478, new_n7479,
    new_n7480, new_n7481, new_n7482, new_n7483, new_n7484, new_n7485,
    new_n7486, new_n7487, new_n7488, new_n7489, new_n7490, new_n7491,
    new_n7492, new_n7493, new_n7494, new_n7495, new_n7496, new_n7497,
    new_n7498, new_n7499, new_n7500, new_n7501, new_n7502, new_n7503,
    new_n7504, new_n7505, new_n7506, new_n7507_1, new_n7508, new_n7509,
    new_n7510, new_n7511, new_n7512, new_n7513, new_n7514_1, new_n7515,
    new_n7516, new_n7517, new_n7519, new_n7520, new_n7521, new_n7522,
    new_n7523, new_n7524_1, new_n7525, new_n7526, new_n7527, new_n7528,
    new_n7529, new_n7530, new_n7531, new_n7532, new_n7533, new_n7534,
    new_n7535, new_n7536, new_n7537, new_n7538, new_n7539, new_n7540,
    new_n7541, new_n7542, new_n7543, new_n7544, new_n7545, new_n7546,
    new_n7547, new_n7548, new_n7549, new_n7550, new_n7551, new_n7552,
    new_n7553, new_n7554, new_n7555, new_n7556, new_n7557, new_n7558_1,
    new_n7559, new_n7560, new_n7561, new_n7562, new_n7563, new_n7564,
    new_n7565, new_n7566_1, new_n7567, new_n7568, new_n7569_1, new_n7570,
    new_n7571, new_n7572_1, new_n7573, new_n7574, new_n7575_1, new_n7576,
    new_n7577, new_n7578, new_n7579, new_n7580, new_n7581, new_n7582,
    new_n7583, new_n7584, new_n7585_1, new_n7586, new_n7587, new_n7588_1,
    new_n7589, new_n7590, new_n7591, new_n7592, new_n7593_1, new_n7594,
    new_n7595, new_n7596, new_n7597, new_n7598_1, new_n7599, new_n7600,
    new_n7601, new_n7602, new_n7603, new_n7604, new_n7605, new_n7606,
    new_n7607_1, new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612,
    new_n7613, new_n7614, new_n7615, new_n7616_1, new_n7617, new_n7618,
    new_n7619, new_n7620, new_n7621, new_n7622, new_n7623, new_n7624,
    new_n7625, new_n7626, new_n7627, new_n7628, new_n7629, new_n7630_1,
    new_n7631, new_n7632, new_n7633, new_n7634, new_n7635, new_n7636,
    new_n7637, new_n7638, new_n7639, new_n7640, new_n7641, new_n7642,
    new_n7643_1, new_n7644, new_n7645, new_n7646, new_n7647_1, new_n7648,
    new_n7649, new_n7650, new_n7651, new_n7652, new_n7653, new_n7654,
    new_n7655, new_n7656, new_n7657_1, new_n7658, new_n7659, new_n7660,
    new_n7661, new_n7662, new_n7663, new_n7664, new_n7665, new_n7666,
    new_n7667, new_n7668, new_n7669, new_n7670_1, new_n7671, new_n7672,
    new_n7673, new_n7674_1, new_n7675, new_n7676, new_n7677, new_n7678_1,
    new_n7679_1, new_n7680, new_n7681, new_n7682, new_n7683, new_n7684,
    new_n7685, new_n7686_1, new_n7687, new_n7688, new_n7689, new_n7690,
    new_n7691, new_n7692_1, new_n7693_1, new_n7694, new_n7695, new_n7696,
    new_n7697, new_n7698_1, new_n7699, new_n7700, new_n7701, new_n7702,
    new_n7703, new_n7704, new_n7705, new_n7706, new_n7707, new_n7708_1,
    new_n7709, new_n7710, new_n7711, new_n7712, new_n7713, new_n7714,
    new_n7715, new_n7716, new_n7717, new_n7718, new_n7719, new_n7720,
    new_n7721_1, new_n7722, new_n7723, new_n7724, new_n7725, new_n7726,
    new_n7727, new_n7729, new_n7730, new_n7731_1, new_n7733, new_n7734,
    new_n7735, new_n7736, new_n7737, new_n7738, new_n7739, new_n7740,
    new_n7741, new_n7742, new_n7743, new_n7744, new_n7745, new_n7746,
    new_n7747, new_n7748, new_n7749, new_n7750, new_n7751_1, new_n7752,
    new_n7753, new_n7754, new_n7755, new_n7756, new_n7757, new_n7758,
    new_n7759_1, new_n7760, new_n7761, new_n7762, new_n7763, new_n7764,
    new_n7765, new_n7766, new_n7767, new_n7768, new_n7769_1, new_n7770,
    new_n7771, new_n7772, new_n7773_1, new_n7774, new_n7775, new_n7776,
    new_n7777, new_n7778, new_n7779, new_n7780_1, new_n7781, new_n7782,
    new_n7783, new_n7784, new_n7785, new_n7786, new_n7787, new_n7788_1,
    new_n7789, new_n7790, new_n7791, new_n7792, new_n7793, new_n7794_1,
    new_n7795, new_n7796, new_n7797, new_n7798, new_n7799, new_n7800,
    new_n7801, new_n7802, new_n7803, new_n7804, new_n7805, new_n7806,
    new_n7807, new_n7808, new_n7809, new_n7810, new_n7811_1, new_n7812,
    new_n7813, new_n7814, new_n7815, new_n7816, new_n7817, new_n7818,
    new_n7819, new_n7820, new_n7821, new_n7822, new_n7823, new_n7824,
    new_n7825, new_n7826, new_n7827, new_n7828, new_n7829, new_n7830_1,
    new_n7831, new_n7832, new_n7833, new_n7834_1, new_n7835, new_n7836,
    new_n7837, new_n7838, new_n7839, new_n7840, new_n7841_1, new_n7842,
    new_n7843, new_n7844, new_n7845, new_n7846, new_n7847, new_n7848,
    new_n7849, new_n7851, new_n7852, new_n7853, new_n7854, new_n7855,
    new_n7856, new_n7857, new_n7858, new_n7859, new_n7860, new_n7861,
    new_n7862, new_n7863, new_n7864, new_n7865, new_n7866, new_n7867,
    new_n7868, new_n7869, new_n7870, new_n7871, new_n7872, new_n7873,
    new_n7874, new_n7875, new_n7876_1, new_n7877, new_n7878, new_n7879,
    new_n7880, new_n7881, new_n7882, new_n7883, new_n7884_1, new_n7885,
    new_n7886, new_n7887, new_n7888, new_n7889, new_n7890, new_n7891,
    new_n7892, new_n7893, new_n7894, new_n7895, new_n7896, new_n7897,
    new_n7898, new_n7899, new_n7900, new_n7901, new_n7902, new_n7903,
    new_n7904, new_n7905, new_n7906, new_n7907, new_n7908, new_n7909,
    new_n7910, new_n7911, new_n7912, new_n7913, new_n7914, new_n7915,
    new_n7916, new_n7917_1, new_n7918, new_n7919, new_n7920, new_n7921,
    new_n7922, new_n7923, new_n7924, new_n7925, new_n7926, new_n7927,
    new_n7928, new_n7929, new_n7930, new_n7932, new_n7933, new_n7934,
    new_n7935, new_n7936, new_n7937_1, new_n7938, new_n7939, new_n7940,
    new_n7941, new_n7942, new_n7943_1, new_n7944, new_n7945, new_n7946,
    new_n7947, new_n7948, new_n7949_1, new_n7950_1, new_n7951, new_n7952,
    new_n7953, new_n7954, new_n7955, new_n7956, new_n7957, new_n7958,
    new_n7959_1, new_n7960, new_n7961, new_n7962, new_n7963_1, new_n7964,
    new_n7965, new_n7966, new_n7967, new_n7968_1, new_n7969, new_n7970,
    new_n7971, new_n7972, new_n7973, new_n7974, new_n7975, new_n7976,
    new_n7977, new_n7978, new_n7979, new_n7980, new_n7981, new_n7982,
    new_n7983, new_n7984, new_n7985, new_n7986, new_n7987, new_n7988,
    new_n7989, new_n7990, new_n7991, new_n7992_1, new_n7993, new_n7994,
    new_n7995, new_n7996, new_n7997, new_n7998, new_n7999_1, new_n8000,
    new_n8001, new_n8002, new_n8003, new_n8004, new_n8005, new_n8006_1,
    new_n8007, new_n8008, new_n8009, new_n8010, new_n8011, new_n8012,
    new_n8013, new_n8014, new_n8015, new_n8016, new_n8017, new_n8018,
    new_n8019, new_n8020, new_n8021, new_n8022, new_n8023, new_n8024,
    new_n8025, new_n8026, new_n8027_1, new_n8028, new_n8029, new_n8030,
    new_n8031_1, new_n8032, new_n8033, new_n8034, new_n8035, new_n8036,
    new_n8037, new_n8038, new_n8039, new_n8040, new_n8041, new_n8042_1,
    new_n8043, new_n8044, new_n8045, new_n8046, new_n8047, new_n8048,
    new_n8049, new_n8050, new_n8051, new_n8052_1, new_n8053, new_n8054,
    new_n8055, new_n8056, new_n8057, new_n8058, new_n8059, new_n8060,
    new_n8061, new_n8062, new_n8063, new_n8064, new_n8065, new_n8066,
    new_n8067_1, new_n8068, new_n8069, new_n8070, new_n8071, new_n8072,
    new_n8073, new_n8074, new_n8075, new_n8076, new_n8077, new_n8078,
    new_n8079, new_n8080, new_n8081, new_n8082, new_n8083, new_n8084,
    new_n8085, new_n8086, new_n8087, new_n8088, new_n8089, new_n8090,
    new_n8091, new_n8092, new_n8093, new_n8094, new_n8095_1, new_n8096,
    new_n8097, new_n8098, new_n8099, new_n8100, new_n8101, new_n8102,
    new_n8103_1, new_n8104, new_n8105, new_n8106, new_n8107, new_n8108,
    new_n8109_1, new_n8110, new_n8111, new_n8112, new_n8113, new_n8114,
    new_n8115, new_n8116, new_n8117, new_n8118, new_n8119, new_n8120,
    new_n8121, new_n8122, new_n8123, new_n8124, new_n8125, new_n8126,
    new_n8127_1, new_n8128, new_n8129, new_n8130_1, new_n8131, new_n8132,
    new_n8133, new_n8134, new_n8135_1, new_n8136, new_n8137, new_n8138,
    new_n8139_1, new_n8140, new_n8141, new_n8142, new_n8143, new_n8144,
    new_n8145, new_n8146, new_n8147, new_n8148_1, new_n8149_1, new_n8150,
    new_n8151, new_n8152, new_n8153, new_n8154, new_n8155, new_n8156,
    new_n8157, new_n8158, new_n8159_1, new_n8160, new_n8161, new_n8162,
    new_n8163, new_n8164, new_n8165, new_n8166, new_n8167, new_n8168,
    new_n8169, new_n8170, new_n8171, new_n8172, new_n8173, new_n8174,
    new_n8175, new_n8176, new_n8177, new_n8178, new_n8179_1, new_n8180,
    new_n8181, new_n8182, new_n8183, new_n8184, new_n8185, new_n8186,
    new_n8187, new_n8188, new_n8189, new_n8190, new_n8191, new_n8192,
    new_n8193, new_n8194_1, new_n8195, new_n8196, new_n8197, new_n8198,
    new_n8200, new_n8201, new_n8202, new_n8203, new_n8204, new_n8205,
    new_n8206, new_n8207, new_n8208, new_n8209, new_n8210, new_n8211,
    new_n8212, new_n8213, new_n8214, new_n8215_1, new_n8216, new_n8217,
    new_n8218, new_n8219, new_n8220, new_n8221, new_n8222, new_n8223,
    new_n8224, new_n8225, new_n8226, new_n8227, new_n8228, new_n8229,
    new_n8230, new_n8231, new_n8232, new_n8233, new_n8234, new_n8235,
    new_n8236, new_n8237, new_n8238, new_n8239, new_n8240, new_n8241,
    new_n8242, new_n8243, new_n8244_1, new_n8245, new_n8246, new_n8247,
    new_n8248, new_n8249, new_n8250, new_n8251, new_n8252, new_n8253,
    new_n8254, new_n8255_1, new_n8256_1, new_n8257, new_n8258, new_n8259_1,
    new_n8260, new_n8261, new_n8262, new_n8263, new_n8264, new_n8265,
    new_n8266, new_n8267_1, new_n8268, new_n8269, new_n8270, new_n8271,
    new_n8272, new_n8273, new_n8274, new_n8275, new_n8276_1, new_n8277,
    new_n8278, new_n8279, new_n8280, new_n8281, new_n8282, new_n8283,
    new_n8284, new_n8285_1, new_n8286, new_n8287, new_n8288_1, new_n8289,
    new_n8290, new_n8291, new_n8292, new_n8293, new_n8294, new_n8295,
    new_n8296, new_n8297, new_n8298, new_n8299, new_n8300, new_n8301,
    new_n8302, new_n8303, new_n8304, new_n8305_1, new_n8306_1, new_n8307,
    new_n8308, new_n8309_1, new_n8310, new_n8311, new_n8312, new_n8313,
    new_n8314, new_n8315, new_n8316, new_n8317, new_n8318, new_n8319,
    new_n8320_1, new_n8321_1, new_n8322, new_n8323, new_n8324_1, new_n8325,
    new_n8326, new_n8327, new_n8328, new_n8329, new_n8330, new_n8331,
    new_n8332, new_n8333, new_n8334, new_n8335, new_n8336, new_n8337,
    new_n8338, new_n8339_1, new_n8340, new_n8341, new_n8342, new_n8343,
    new_n8344, new_n8345, new_n8346, new_n8347, new_n8348, new_n8349,
    new_n8350, new_n8351, new_n8352, new_n8353, new_n8354, new_n8355,
    new_n8356, new_n8357, new_n8358, new_n8359, new_n8360, new_n8361,
    new_n8362, new_n8363_1, new_n8364, new_n8365, new_n8366, new_n8367,
    new_n8368, new_n8369, new_n8370, new_n8371, new_n8372, new_n8373,
    new_n8374, new_n8375, new_n8376_1, new_n8377, new_n8378, new_n8379,
    new_n8380, new_n8381_1, new_n8382, new_n8383, new_n8384, new_n8385,
    new_n8386, new_n8387, new_n8388, new_n8389, new_n8390, new_n8391,
    new_n8392, new_n8393, new_n8394, new_n8395, new_n8396, new_n8397,
    new_n8398, new_n8399_1, new_n8400, new_n8401, new_n8402, new_n8403,
    new_n8404, new_n8405_1, new_n8406, new_n8407, new_n8408_1, new_n8409,
    new_n8410, new_n8411, new_n8412, new_n8413, new_n8414, new_n8415,
    new_n8416, new_n8417_1, new_n8418, new_n8419, new_n8420, new_n8421,
    new_n8422, new_n8423, new_n8424, new_n8425, new_n8426, new_n8427,
    new_n8428, new_n8429, new_n8430, new_n8431, new_n8432_1, new_n8433,
    new_n8434, new_n8435, new_n8436, new_n8437, new_n8438, new_n8439_1,
    new_n8440, new_n8441, new_n8442, new_n8443, new_n8444, new_n8445,
    new_n8446, new_n8447, new_n8448, new_n8449, new_n8450, new_n8451,
    new_n8452, new_n8453_1, new_n8454, new_n8455, new_n8456, new_n8457,
    new_n8458, new_n8459, new_n8460, new_n8461, new_n8462, new_n8463,
    new_n8464, new_n8465, new_n8466, new_n8467, new_n8468, new_n8469,
    new_n8470, new_n8471, new_n8472, new_n8473, new_n8474, new_n8475,
    new_n8476, new_n8477, new_n8478, new_n8479, new_n8480_1, new_n8481,
    new_n8482, new_n8483, new_n8484, new_n8485, new_n8486, new_n8487,
    new_n8488, new_n8490, new_n8491, new_n8492, new_n8493, new_n8494,
    new_n8495, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505_1, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510_1, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519_1,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526_1, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535_1, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550_1, new_n8551, new_n8552, new_n8553, new_n8554, new_n8555,
    new_n8556, new_n8557, new_n8558, new_n8559, new_n8560, new_n8561,
    new_n8562, new_n8563_1, new_n8564, new_n8565, new_n8566, new_n8567,
    new_n8568, new_n8569, new_n8570, new_n8571, new_n8572, new_n8573,
    new_n8574, new_n8575, new_n8576, new_n8577, new_n8578, new_n8579,
    new_n8580, new_n8581_1, new_n8582, new_n8583, new_n8584, new_n8585,
    new_n8586, new_n8587, new_n8588, new_n8589, new_n8590, new_n8591,
    new_n8592, new_n8593, new_n8594_1, new_n8595, new_n8596, new_n8597,
    new_n8598, new_n8599, new_n8600, new_n8601, new_n8602, new_n8603,
    new_n8604, new_n8605, new_n8606, new_n8607, new_n8608_1, new_n8609,
    new_n8610, new_n8611, new_n8612, new_n8613, new_n8614_1, new_n8615,
    new_n8616, new_n8617, new_n8618, new_n8619, new_n8620_1, new_n8621,
    new_n8622, new_n8623, new_n8624, new_n8625, new_n8626, new_n8627,
    new_n8628, new_n8629, new_n8630, new_n8631, new_n8632, new_n8633,
    new_n8634, new_n8635, new_n8636, new_n8637_1, new_n8638_1, new_n8639,
    new_n8640, new_n8641, new_n8642, new_n8643, new_n8644, new_n8645,
    new_n8646, new_n8647, new_n8648, new_n8649, new_n8650, new_n8651,
    new_n8652, new_n8653, new_n8654, new_n8655, new_n8656_1, new_n8657,
    new_n8658, new_n8659, new_n8660, new_n8661, new_n8662_1, new_n8663,
    new_n8664, new_n8665, new_n8666, new_n8667, new_n8668, new_n8669,
    new_n8670, new_n8671, new_n8672, new_n8673, new_n8674, new_n8675,
    new_n8676, new_n8677, new_n8678_1, new_n8679, new_n8680, new_n8681,
    new_n8682, new_n8683, new_n8684, new_n8685, new_n8686, new_n8687_1,
    new_n8688, new_n8689, new_n8690, new_n8691, new_n8692, new_n8693,
    new_n8694_1, new_n8695, new_n8696, new_n8697, new_n8698, new_n8699,
    new_n8700, new_n8701, new_n8702, new_n8703, new_n8704, new_n8705,
    new_n8706, new_n8707, new_n8708, new_n8709, new_n8710, new_n8711,
    new_n8712, new_n8713, new_n8714, new_n8715, new_n8716_1, new_n8717,
    new_n8718, new_n8719, new_n8720, new_n8721_1, new_n8722, new_n8723,
    new_n8724, new_n8725, new_n8726, new_n8727, new_n8728, new_n8729,
    new_n8730, new_n8731, new_n8732, new_n8733, new_n8734, new_n8735,
    new_n8736, new_n8737, new_n8738, new_n8739, new_n8740, new_n8741,
    new_n8742, new_n8743, new_n8744_1, new_n8745_1, new_n8746, new_n8747,
    new_n8748, new_n8749, new_n8750, new_n8751, new_n8752, new_n8753,
    new_n8754, new_n8755, new_n8756, new_n8757, new_n8758, new_n8759,
    new_n8760, new_n8761, new_n8762, new_n8763, new_n8764, new_n8765,
    new_n8766, new_n8767, new_n8768, new_n8769, new_n8770, new_n8771,
    new_n8772, new_n8773, new_n8774, new_n8775, new_n8776, new_n8777,
    new_n8778, new_n8779, new_n8780, new_n8781, new_n8782_1, new_n8783,
    new_n8784, new_n8785, new_n8786, new_n8787, new_n8789, new_n8790,
    new_n8791, new_n8792, new_n8793, new_n8794, new_n8795, new_n8796,
    new_n8797, new_n8798, new_n8799, new_n8800, new_n8801, new_n8802,
    new_n8803_1, new_n8804, new_n8805, new_n8806_1, new_n8807, new_n8808,
    new_n8809_1, new_n8810, new_n8811, new_n8812, new_n8813, new_n8814,
    new_n8815, new_n8816, new_n8817, new_n8818, new_n8819, new_n8820,
    new_n8821_1, new_n8822, new_n8823, new_n8824_1, new_n8825, new_n8826,
    new_n8827_1, new_n8828, new_n8829, new_n8830, new_n8831, new_n8832,
    new_n8833, new_n8834, new_n8835, new_n8836, new_n8837, new_n8838,
    new_n8839, new_n8840, new_n8841, new_n8842, new_n8843, new_n8844,
    new_n8845, new_n8846, new_n8847, new_n8848, new_n8849_1, new_n8850,
    new_n8851, new_n8852, new_n8853, new_n8854, new_n8855, new_n8856_1,
    new_n8857, new_n8858, new_n8859, new_n8860, new_n8861_1, new_n8862_1,
    new_n8863, new_n8864, new_n8865, new_n8866, new_n8867, new_n8868,
    new_n8869_1, new_n8870, new_n8871, new_n8872, new_n8873, new_n8874,
    new_n8875, new_n8876, new_n8877, new_n8878, new_n8879, new_n8880,
    new_n8881, new_n8882, new_n8883, new_n8884_1, new_n8885, new_n8886,
    new_n8887, new_n8888, new_n8889, new_n8890, new_n8891, new_n8892,
    new_n8893, new_n8894, new_n8895, new_n8896, new_n8897, new_n8898,
    new_n8899, new_n8900, new_n8901, new_n8902, new_n8903, new_n8904,
    new_n8905, new_n8906, new_n8907, new_n8908, new_n8909_1, new_n8910,
    new_n8911_1, new_n8912, new_n8913, new_n8914, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920_1, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943_1, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964_1,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971_1, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982_1,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993_1, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003_1, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012_1,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9030, new_n9031,
    new_n9032_1, new_n9033, new_n9034, new_n9035, new_n9036, new_n9037,
    new_n9038, new_n9039, new_n9040, new_n9041, new_n9042_1, new_n9043,
    new_n9044, new_n9045, new_n9046_1, new_n9047_1, new_n9048, new_n9049,
    new_n9050, new_n9051, new_n9052, new_n9053, new_n9054, new_n9055,
    new_n9056, new_n9057, new_n9058, new_n9059, new_n9060, new_n9061,
    new_n9062, new_n9063, new_n9064, new_n9065, new_n9066, new_n9067,
    new_n9068, new_n9069, new_n9070, new_n9071, new_n9072, new_n9073,
    new_n9074, new_n9075, new_n9076, new_n9077, new_n9078, new_n9079,
    new_n9080, new_n9081, new_n9082, new_n9083, new_n9084, new_n9085,
    new_n9086, new_n9087, new_n9088, new_n9089, new_n9090_1, new_n9091,
    new_n9092, new_n9093, new_n9094, new_n9095, new_n9096, new_n9097,
    new_n9098, new_n9099, new_n9100, new_n9101, new_n9102, new_n9103,
    new_n9104_1, new_n9105, new_n9106, new_n9107, new_n9108, new_n9109,
    new_n9110, new_n9111, new_n9112, new_n9113, new_n9114, new_n9115,
    new_n9116, new_n9117, new_n9118, new_n9119, new_n9120, new_n9121,
    new_n9122, new_n9123, new_n9124, new_n9125, new_n9126, new_n9127,
    new_n9128, new_n9129_1, new_n9130, new_n9131, new_n9132, new_n9133,
    new_n9134, new_n9135, new_n9136, new_n9137, new_n9138, new_n9139,
    new_n9140, new_n9141, new_n9142, new_n9143, new_n9144, new_n9145,
    new_n9146_1, new_n9147, new_n9148, new_n9149, new_n9150, new_n9151,
    new_n9152, new_n9153, new_n9154, new_n9155, new_n9156, new_n9157,
    new_n9158, new_n9159, new_n9160, new_n9161, new_n9162, new_n9163,
    new_n9164_1, new_n9165, new_n9166_1, new_n9167, new_n9168, new_n9169,
    new_n9170, new_n9171, new_n9172_1, new_n9173, new_n9174, new_n9175,
    new_n9176, new_n9177, new_n9178, new_n9179, new_n9180, new_n9181,
    new_n9182_1, new_n9183, new_n9184, new_n9185, new_n9186, new_n9187,
    new_n9188, new_n9189, new_n9190, new_n9191_1, new_n9192, new_n9193,
    new_n9194, new_n9195, new_n9196, new_n9197, new_n9198, new_n9199,
    new_n9200, new_n9201, new_n9202, new_n9203, new_n9204, new_n9205,
    new_n9206, new_n9207, new_n9208, new_n9209, new_n9210, new_n9211,
    new_n9212, new_n9213, new_n9214, new_n9215, new_n9216, new_n9217_1,
    new_n9218, new_n9219, new_n9220_1, new_n9221, new_n9222, new_n9223,
    new_n9224, new_n9225, new_n9226, new_n9227, new_n9228, new_n9229,
    new_n9230, new_n9231, new_n9232, new_n9233, new_n9234, new_n9235,
    new_n9236, new_n9237, new_n9238, new_n9239, new_n9240, new_n9241,
    new_n9242, new_n9243, new_n9244, new_n9245, new_n9246_1, new_n9247,
    new_n9248, new_n9249, new_n9250, new_n9251_1, new_n9252, new_n9253,
    new_n9254, new_n9255, new_n9256, new_n9257, new_n9258, new_n9259_1,
    new_n9260, new_n9261_1, new_n9262, new_n9263, new_n9264, new_n9265,
    new_n9266, new_n9267, new_n9268, new_n9269, new_n9270, new_n9271,
    new_n9272, new_n9273, new_n9274, new_n9275, new_n9276, new_n9277,
    new_n9278, new_n9279, new_n9280, new_n9281, new_n9282, new_n9283,
    new_n9284, new_n9285, new_n9286, new_n9287_1, new_n9288, new_n9289,
    new_n9290, new_n9291, new_n9292, new_n9293, new_n9294, new_n9295,
    new_n9296, new_n9297, new_n9298, new_n9299, new_n9300, new_n9301,
    new_n9302, new_n9303, new_n9304, new_n9305, new_n9306, new_n9307,
    new_n9308_1, new_n9309, new_n9310, new_n9311, new_n9312, new_n9313,
    new_n9314, new_n9315, new_n9316, new_n9317, new_n9318_1, new_n9319,
    new_n9320, new_n9321, new_n9322, new_n9323_1, new_n9324, new_n9325,
    new_n9326, new_n9327, new_n9328, new_n9329, new_n9330, new_n9331,
    new_n9332, new_n9333, new_n9334, new_n9335, new_n9336, new_n9337,
    new_n9338, new_n9339, new_n9340, new_n9341, new_n9342, new_n9343,
    new_n9344_1, new_n9345, new_n9346, new_n9347, new_n9348, new_n9349,
    new_n9350, new_n9351, new_n9352, new_n9353, new_n9354, new_n9355,
    new_n9356, new_n9357, new_n9358, new_n9359, new_n9360, new_n9361,
    new_n9362, new_n9363, new_n9364_1, new_n9365, new_n9366, new_n9367,
    new_n9368, new_n9369, new_n9370, new_n9371_1, new_n9372_1, new_n9373,
    new_n9374, new_n9375, new_n9376, new_n9377, new_n9378, new_n9379,
    new_n9380_1, new_n9381, new_n9382_1, new_n9383, new_n9384, new_n9385,
    new_n9386, new_n9387, new_n9388, new_n9389, new_n9390, new_n9391,
    new_n9392, new_n9393, new_n9394, new_n9396_1, new_n9397, new_n9398,
    new_n9399_1, new_n9400, new_n9401, new_n9402, new_n9403_1, new_n9404,
    new_n9405, new_n9406, new_n9407, new_n9408, new_n9409, new_n9410,
    new_n9411, new_n9412, new_n9413, new_n9414, new_n9415, new_n9416,
    new_n9417, new_n9418, new_n9419_1, new_n9420, new_n9421, new_n9422,
    new_n9423_1, new_n9424, new_n9425, new_n9426, new_n9427, new_n9428,
    new_n9429, new_n9430_1, new_n9431, new_n9432, new_n9433, new_n9434,
    new_n9435_1, new_n9436, new_n9437, new_n9438, new_n9439, new_n9440,
    new_n9441, new_n9442, new_n9443, new_n9444, new_n9445_1, new_n9446,
    new_n9447, new_n9448, new_n9449, new_n9450, new_n9451_1, new_n9452,
    new_n9453, new_n9454, new_n9455, new_n9456, new_n9457, new_n9458_1,
    new_n9459_1, new_n9460_1, new_n9461, new_n9462, new_n9463, new_n9464,
    new_n9465, new_n9466, new_n9467, new_n9468, new_n9469, new_n9470,
    new_n9471, new_n9472, new_n9473, new_n9474, new_n9475, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493_1, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507_1, new_n9508_1, new_n9509, new_n9510, new_n9511, new_n9512_1,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552_1, new_n9553, new_n9554_1,
    new_n9555, new_n9556_1, new_n9557_1, new_n9558_1, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9568, new_n9569, new_n9570, new_n9571, new_n9572,
    new_n9573, new_n9574, new_n9575, new_n9576, new_n9577, new_n9578,
    new_n9579, new_n9580, new_n9581, new_n9582, new_n9583, new_n9584,
    new_n9585, new_n9586, new_n9587, new_n9588, new_n9589, new_n9590,
    new_n9591, new_n9592, new_n9593, new_n9594, new_n9595, new_n9596,
    new_n9597, new_n9598_1, new_n9599, new_n9600, new_n9601, new_n9602,
    new_n9603, new_n9604, new_n9605, new_n9606, new_n9607, new_n9608,
    new_n9609, new_n9610, new_n9611, new_n9612, new_n9613, new_n9614,
    new_n9615, new_n9616_1, new_n9617, new_n9618, new_n9619, new_n9620,
    new_n9621, new_n9622_1, new_n9623, new_n9624, new_n9625, new_n9626_1,
    new_n9627, new_n9628, new_n9629, new_n9630, new_n9631, new_n9632,
    new_n9633_1, new_n9634, new_n9635_1, new_n9636, new_n9637, new_n9638,
    new_n9639, new_n9640, new_n9641, new_n9642, new_n9643, new_n9644,
    new_n9645, new_n9646_1, new_n9647, new_n9648_1, new_n9649, new_n9650,
    new_n9651, new_n9652, new_n9653, new_n9654, new_n9655_1, new_n9656,
    new_n9657, new_n9658, new_n9659, new_n9660, new_n9661, new_n9662,
    new_n9663, new_n9664, new_n9665, new_n9666, new_n9667, new_n9668,
    new_n9669, new_n9670, new_n9671, new_n9672, new_n9673, new_n9674,
    new_n9675, new_n9676, new_n9677, new_n9678, new_n9679, new_n9680,
    new_n9681, new_n9682, new_n9683, new_n9684, new_n9685, new_n9686,
    new_n9687, new_n9688, new_n9689_1, new_n9690, new_n9691, new_n9692,
    new_n9693, new_n9694, new_n9695_1, new_n9696, new_n9697, new_n9698,
    new_n9699_1, new_n9700, new_n9701, new_n9702, new_n9703, new_n9704,
    new_n9705, new_n9706, new_n9707, new_n9708, new_n9709, new_n9710,
    new_n9711, new_n9712, new_n9713, new_n9714, new_n9715, new_n9716,
    new_n9717, new_n9718, new_n9719, new_n9720, new_n9721, new_n9722,
    new_n9723, new_n9724, new_n9725, new_n9726_1, new_n9727, new_n9728,
    new_n9729, new_n9730, new_n9731, new_n9732, new_n9733, new_n9734,
    new_n9735, new_n9736, new_n9737, new_n9738, new_n9739, new_n9740,
    new_n9741, new_n9742, new_n9743, new_n9744, new_n9745, new_n9746,
    new_n9747, new_n9748, new_n9749, new_n9752, new_n9753_1, new_n9754,
    new_n9755, new_n9756, new_n9757, new_n9758, new_n9759, new_n9760,
    new_n9761_1, new_n9762, new_n9763_1, new_n9764, new_n9765, new_n9766,
    new_n9767_1, new_n9768, new_n9769, new_n9770, new_n9771_1, new_n9772,
    new_n9773, new_n9774, new_n9775, new_n9776, new_n9777, new_n9778_1,
    new_n9779, new_n9780, new_n9781, new_n9782, new_n9783_1, new_n9784,
    new_n9785, new_n9786, new_n9787, new_n9788, new_n9789, new_n9790,
    new_n9791, new_n9792, new_n9793, new_n9794, new_n9795, new_n9796,
    new_n9797, new_n9798, new_n9799, new_n9800, new_n9801, new_n9802,
    new_n9803_1, new_n9804, new_n9805, new_n9806, new_n9807, new_n9808,
    new_n9809, new_n9810, new_n9811, new_n9812, new_n9813, new_n9814,
    new_n9815, new_n9816, new_n9817, new_n9818, new_n9819, new_n9820,
    new_n9821, new_n9822, new_n9823, new_n9824, new_n9825, new_n9826,
    new_n9827, new_n9828, new_n9829, new_n9830, new_n9831, new_n9832_1,
    new_n9833_1, new_n9834, new_n9835, new_n9836, new_n9837, new_n9838_1,
    new_n9839, new_n9840, new_n9841, new_n9842, new_n9843, new_n9844,
    new_n9845, new_n9846, new_n9847, new_n9848, new_n9849, new_n9850,
    new_n9851, new_n9852, new_n9853, new_n9854, new_n9855, new_n9856,
    new_n9857, new_n9858, new_n9859, new_n9860, new_n9861, new_n9862,
    new_n9863, new_n9864, new_n9865, new_n9866, new_n9867_1, new_n9868,
    new_n9869, new_n9870, new_n9871, new_n9872_1, new_n9873, new_n9874,
    new_n9875, new_n9876, new_n9877, new_n9878, new_n9879, new_n9880,
    new_n9881, new_n9882, new_n9883, new_n9884, new_n9885, new_n9886,
    new_n9887, new_n9888, new_n9889, new_n9890_1, new_n9891, new_n9892,
    new_n9893, new_n9894, new_n9895, new_n9896, new_n9897, new_n9898,
    new_n9899, new_n9900, new_n9901, new_n9902, new_n9903, new_n9904,
    new_n9905, new_n9906, new_n9907, new_n9908, new_n9909, new_n9910,
    new_n9911, new_n9912, new_n9913, new_n9914, new_n9915, new_n9916,
    new_n9917_1, new_n9918, new_n9919_1, new_n9920, new_n9921, new_n9922,
    new_n9923, new_n9924, new_n9925, new_n9926_1, new_n9927, new_n9928,
    new_n9929, new_n9930, new_n9931, new_n9932, new_n9933, new_n9934_1,
    new_n9935, new_n9936, new_n9937, new_n9938_1, new_n9939, new_n9940,
    new_n9941, new_n9942_1, new_n9943, new_n9944, new_n9945, new_n9946_1,
    new_n9947, new_n9948, new_n9949, new_n9950, new_n9951, new_n9952,
    new_n9953, new_n9954, new_n9955, new_n9956, new_n9957, new_n9958,
    new_n9959, new_n9960, new_n9961, new_n9962, new_n9963, new_n9964,
    new_n9965, new_n9966, new_n9967_1, new_n9968_1, new_n9969, new_n9970,
    new_n9971, new_n9972, new_n9973, new_n9974, new_n9975, new_n9976,
    new_n9977, new_n9978, new_n9979, new_n9980, new_n9981, new_n9982,
    new_n9983, new_n9984, new_n9985, new_n9986, new_n9987, new_n9988,
    new_n9989, new_n9990, new_n9991, new_n9992, new_n9993, new_n9994,
    new_n9995, new_n9996, new_n9997, new_n9998, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009_1, new_n10010_1, new_n10011, new_n10012,
    new_n10013, new_n10014, new_n10015, new_n10016, new_n10017_1,
    new_n10018_1, new_n10019_1, new_n10020, new_n10021_1, new_n10022,
    new_n10023, new_n10024, new_n10025, new_n10026, new_n10027, new_n10028,
    new_n10029, new_n10030, new_n10031, new_n10032, new_n10033, new_n10034,
    new_n10035, new_n10036, new_n10037, new_n10038, new_n10039, new_n10040,
    new_n10041, new_n10042, new_n10043, new_n10044, new_n10045, new_n10046,
    new_n10047, new_n10049, new_n10050, new_n10051, new_n10052,
    new_n10053_1, new_n10054, new_n10055_1, new_n10056, new_n10057_1,
    new_n10058, new_n10059, new_n10060, new_n10061, new_n10062, new_n10063,
    new_n10064, new_n10065, new_n10066, new_n10067, new_n10068, new_n10069,
    new_n10070, new_n10071, new_n10072, new_n10073, new_n10074, new_n10075,
    new_n10076, new_n10077, new_n10078, new_n10079, new_n10080, new_n10081,
    new_n10082, new_n10083, new_n10084, new_n10085, new_n10086, new_n10087,
    new_n10088, new_n10089, new_n10090, new_n10091, new_n10092, new_n10093,
    new_n10094, new_n10095, new_n10096_1, new_n10097, new_n10098,
    new_n10099, new_n10100, new_n10101_1, new_n10102, new_n10103,
    new_n10104, new_n10106, new_n10107, new_n10108, new_n10109, new_n10110,
    new_n10111_1, new_n10112, new_n10113, new_n10114, new_n10115,
    new_n10116, new_n10117_1, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125_1,
    new_n10126, new_n10127, new_n10128, new_n10129, new_n10130, new_n10131,
    new_n10132, new_n10133, new_n10134, new_n10135, new_n10136, new_n10137,
    new_n10138, new_n10139, new_n10140, new_n10141, new_n10142, new_n10143,
    new_n10144, new_n10145, new_n10146, new_n10147, new_n10148, new_n10149,
    new_n10150, new_n10151, new_n10152, new_n10153, new_n10154, new_n10155,
    new_n10156, new_n10157, new_n10158_1, new_n10159, new_n10160,
    new_n10161, new_n10162, new_n10163, new_n10164, new_n10165_1,
    new_n10166, new_n10167, new_n10168, new_n10169, new_n10170, new_n10171,
    new_n10172, new_n10173, new_n10174, new_n10175, new_n10176, new_n10177,
    new_n10178, new_n10179, new_n10180, new_n10181, new_n10182, new_n10183,
    new_n10184, new_n10185, new_n10186, new_n10187, new_n10188, new_n10189,
    new_n10190, new_n10191, new_n10192, new_n10193, new_n10194, new_n10195,
    new_n10196, new_n10197, new_n10198, new_n10199, new_n10200,
    new_n10201_1, new_n10202, new_n10203, new_n10204, new_n10205,
    new_n10206, new_n10207, new_n10208, new_n10209, new_n10210, new_n10211,
    new_n10212, new_n10213, new_n10214, new_n10215, new_n10216, new_n10217,
    new_n10218, new_n10219, new_n10220, new_n10221, new_n10222, new_n10223,
    new_n10224, new_n10226, new_n10227, new_n10228, new_n10229, new_n10230,
    new_n10231, new_n10232, new_n10233, new_n10234, new_n10235,
    new_n10236_1, new_n10237, new_n10238, new_n10239_1, new_n10240,
    new_n10241, new_n10242, new_n10243, new_n10244_1, new_n10245,
    new_n10246, new_n10247, new_n10248, new_n10249, new_n10250_1,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261_1,
    new_n10262_1, new_n10263, new_n10264, new_n10265, new_n10266,
    new_n10267, new_n10268, new_n10269, new_n10270, new_n10271, new_n10272,
    new_n10273, new_n10274, new_n10275_1, new_n10276, new_n10277,
    new_n10278, new_n10279, new_n10280, new_n10281, new_n10282, new_n10283,
    new_n10284, new_n10285, new_n10286, new_n10287_1, new_n10288,
    new_n10289, new_n10290, new_n10291, new_n10292, new_n10293, new_n10294,
    new_n10295_1, new_n10296, new_n10297, new_n10298, new_n10299,
    new_n10300, new_n10301, new_n10302, new_n10303, new_n10304, new_n10305,
    new_n10306, new_n10307, new_n10308, new_n10309, new_n10310, new_n10311,
    new_n10312, new_n10313, new_n10314, new_n10315, new_n10316, new_n10317,
    new_n10318, new_n10319, new_n10320, new_n10321_1, new_n10322,
    new_n10324, new_n10325, new_n10326_1, new_n10327_1, new_n10328,
    new_n10329, new_n10330_1, new_n10331, new_n10332, new_n10333,
    new_n10334, new_n10335, new_n10336, new_n10337, new_n10338, new_n10339,
    new_n10340_1, new_n10341, new_n10342, new_n10343, new_n10344,
    new_n10345_1, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356_1, new_n10357, new_n10358, new_n10359, new_n10360,
    new_n10361, new_n10362, new_n10363, new_n10364, new_n10365, new_n10366,
    new_n10367, new_n10368, new_n10369, new_n10370, new_n10371,
    new_n10372_1, new_n10373, new_n10374, new_n10375, new_n10376,
    new_n10377, new_n10378, new_n10379, new_n10380, new_n10381, new_n10382,
    new_n10383, new_n10384, new_n10385_1, new_n10386, new_n10387_1,
    new_n10388_1, new_n10389, new_n10390_1, new_n10391, new_n10392,
    new_n10393, new_n10394, new_n10395, new_n10396, new_n10397, new_n10398,
    new_n10399, new_n10400, new_n10401, new_n10402, new_n10403,
    new_n10404_1, new_n10405_1, new_n10406, new_n10407, new_n10408,
    new_n10409_1, new_n10410, new_n10411_1, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420_1, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432_1, new_n10433, new_n10434, new_n10435,
    new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476, new_n10477,
    new_n10478, new_n10479, new_n10480, new_n10481, new_n10482, new_n10483,
    new_n10484_1, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489_1, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10504, new_n10505,
    new_n10506, new_n10507, new_n10508, new_n10509, new_n10510, new_n10511,
    new_n10512, new_n10513, new_n10514_1, new_n10515, new_n10516,
    new_n10517, new_n10518, new_n10519, new_n10520, new_n10521, new_n10522,
    new_n10523, new_n10524, new_n10525_1, new_n10526, new_n10527,
    new_n10528, new_n10529, new_n10530, new_n10531, new_n10532, new_n10533,
    new_n10534, new_n10535, new_n10536, new_n10537, new_n10538, new_n10539,
    new_n10540_1, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561_1,
    new_n10562, new_n10563, new_n10564_1, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577_1,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588_1,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593_1,
    new_n10594, new_n10595_1, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611_1, new_n10612, new_n10613, new_n10614_1, new_n10615,
    new_n10616, new_n10617_1, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628_1, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647_1, new_n10648,
    new_n10649, new_n10650_1, new_n10651, new_n10652, new_n10653_1,
    new_n10654, new_n10655, new_n10656, new_n10657, new_n10658, new_n10659,
    new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665,
    new_n10666, new_n10668, new_n10669, new_n10670, new_n10671, new_n10672,
    new_n10673, new_n10674, new_n10676, new_n10677, new_n10678, new_n10679,
    new_n10680, new_n10681, new_n10682, new_n10683, new_n10684, new_n10685,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692_1, new_n10693, new_n10694_1, new_n10695, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701_1,
    new_n10702, new_n10703, new_n10704, new_n10705, new_n10706, new_n10707,
    new_n10708, new_n10709, new_n10710_1, new_n10711, new_n10712_1,
    new_n10713, new_n10714, new_n10715, new_n10716, new_n10717, new_n10718,
    new_n10719, new_n10720, new_n10721, new_n10722, new_n10723, new_n10724,
    new_n10725, new_n10726, new_n10727, new_n10728, new_n10729, new_n10730,
    new_n10731, new_n10732, new_n10733, new_n10734, new_n10735, new_n10736,
    new_n10737, new_n10738, new_n10739_1, new_n10740, new_n10741,
    new_n10742, new_n10743, new_n10744, new_n10745, new_n10746, new_n10747,
    new_n10748, new_n10749, new_n10750, new_n10751, new_n10752, new_n10753,
    new_n10754, new_n10755, new_n10756_1, new_n10757, new_n10758,
    new_n10759, new_n10760, new_n10761, new_n10762, new_n10763_1,
    new_n10764, new_n10765, new_n10766, new_n10767, new_n10768, new_n10769,
    new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775_1, new_n10776, new_n10777, new_n10778, new_n10779,
    new_n10780_1, new_n10781, new_n10782, new_n10783, new_n10784,
    new_n10785, new_n10786, new_n10787, new_n10788, new_n10789, new_n10790,
    new_n10791, new_n10792_1, new_n10793, new_n10794, new_n10795,
    new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807,
    new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817_1, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834_1, new_n10835,
    new_n10836, new_n10837, new_n10838, new_n10839, new_n10840, new_n10841,
    new_n10842, new_n10843, new_n10844, new_n10845, new_n10846, new_n10847,
    new_n10848, new_n10849, new_n10850, new_n10851_1, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10868, new_n10869, new_n10870, new_n10871,
    new_n10872, new_n10873, new_n10874_1, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923,
    new_n10924_1, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943_1, new_n10944, new_n10945,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961_1, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005_1, new_n11006, new_n11007, new_n11008, new_n11009,
    new_n11010, new_n11011_1, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023_1, new_n11024, new_n11025_1,
    new_n11026, new_n11027, new_n11028, new_n11029, new_n11030, new_n11031,
    new_n11032, new_n11033, new_n11034, new_n11035, new_n11036, new_n11037,
    new_n11038, new_n11039, new_n11040, new_n11041, new_n11042, new_n11043,
    new_n11044_1, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056_1, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063_1, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078_1, new_n11079, new_n11082, new_n11084,
    new_n11086, new_n11087, new_n11088, new_n11089, new_n11090, new_n11091,
    new_n11092, new_n11093, new_n11094_1, new_n11095, new_n11096,
    new_n11097, new_n11098, new_n11099, new_n11100, new_n11101_1,
    new_n11102, new_n11103_1, new_n11104, new_n11105, new_n11106,
    new_n11107, new_n11108, new_n11109, new_n11110, new_n11111, new_n11112,
    new_n11113, new_n11114, new_n11115, new_n11116, new_n11117, new_n11118,
    new_n11119, new_n11120_1, new_n11121_1, new_n11122, new_n11123,
    new_n11124, new_n11125, new_n11126, new_n11127_1, new_n11128,
    new_n11129, new_n11130, new_n11131, new_n11132_1, new_n11133,
    new_n11134_1, new_n11135, new_n11136, new_n11137, new_n11138_1,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153, new_n11154, new_n11155, new_n11156,
    new_n11157, new_n11158, new_n11159, new_n11160, new_n11161, new_n11162,
    new_n11163, new_n11164, new_n11165, new_n11166, new_n11167, new_n11168,
    new_n11169, new_n11170, new_n11171, new_n11172, new_n11173, new_n11174,
    new_n11175, new_n11176, new_n11177, new_n11178, new_n11179, new_n11180,
    new_n11181, new_n11182_1, new_n11183, new_n11184_1, new_n11185,
    new_n11186, new_n11187, new_n11188, new_n11189, new_n11190, new_n11191,
    new_n11192_1, new_n11193, new_n11194, new_n11195, new_n11196,
    new_n11197, new_n11198, new_n11199, new_n11200, new_n11201_1,
    new_n11202, new_n11203, new_n11204, new_n11205, new_n11206, new_n11207,
    new_n11208, new_n11209, new_n11210, new_n11211, new_n11212, new_n11213,
    new_n11214, new_n11215, new_n11216, new_n11217, new_n11218, new_n11219,
    new_n11220_1, new_n11221, new_n11222, new_n11223_1, new_n11224,
    new_n11225, new_n11226, new_n11227, new_n11228, new_n11229, new_n11230,
    new_n11231, new_n11232, new_n11233, new_n11234_1, new_n11235,
    new_n11236, new_n11237, new_n11238, new_n11239, new_n11240, new_n11241,
    new_n11242, new_n11243, new_n11244, new_n11245_1, new_n11246,
    new_n11247, new_n11248, new_n11249, new_n11250, new_n11251, new_n11252,
    new_n11253, new_n11254, new_n11255, new_n11256, new_n11257, new_n11258,
    new_n11259, new_n11260, new_n11261_1, new_n11262, new_n11263,
    new_n11264, new_n11265, new_n11266_1, new_n11267, new_n11268,
    new_n11269, new_n11270, new_n11271, new_n11272, new_n11273_1,
    new_n11274, new_n11275_1, new_n11276, new_n11277, new_n11278,
    new_n11279, new_n11280, new_n11281, new_n11282, new_n11283, new_n11284,
    new_n11285, new_n11286, new_n11287, new_n11288, new_n11289,
    new_n11290_1, new_n11291, new_n11292, new_n11293, new_n11295,
    new_n11296, new_n11297, new_n11298, new_n11299, new_n11300, new_n11301,
    new_n11302_1, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313_1, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323,
    new_n11324, new_n11325_1, new_n11326_1, new_n11327, new_n11328,
    new_n11329, new_n11330_1, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345,
    new_n11346, new_n11347_1, new_n11348_1, new_n11349, new_n11350,
    new_n11351, new_n11352_1, new_n11353, new_n11354, new_n11355,
    new_n11356_1, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375_1, new_n11376, new_n11377,
    new_n11378, new_n11379_1, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386_1, new_n11387,
    new_n11388, new_n11389, new_n11390, new_n11391_1, new_n11392,
    new_n11393, new_n11394, new_n11395, new_n11396, new_n11397,
    new_n11398_1, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403_1, new_n11404, new_n11405, new_n11406, new_n11407,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11417, new_n11419_1, new_n11420,
    new_n11421, new_n11422, new_n11423, new_n11424_1, new_n11425,
    new_n11426, new_n11427, new_n11428, new_n11429, new_n11430, new_n11431,
    new_n11432, new_n11433, new_n11434, new_n11435, new_n11436, new_n11437,
    new_n11438, new_n11439_1, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455_1, new_n11456, new_n11457, new_n11458, new_n11459,
    new_n11460, new_n11461, new_n11462_1, new_n11463, new_n11464,
    new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470_1, new_n11471, new_n11472_1, new_n11473_1, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479_1,
    new_n11480, new_n11481_1, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486_1, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496_1, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503_1, new_n11504, new_n11505,
    new_n11506_1, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515_1,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536, new_n11537, new_n11538_1,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548_1, new_n11550,
    new_n11551, new_n11552, new_n11553, new_n11554, new_n11555, new_n11556,
    new_n11557, new_n11558, new_n11559, new_n11560, new_n11561, new_n11562,
    new_n11563, new_n11564_1, new_n11565, new_n11566_1, new_n11567,
    new_n11568, new_n11569, new_n11570, new_n11571, new_n11572, new_n11573,
    new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579_1, new_n11580_1, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11587, new_n11588, new_n11589,
    new_n11590, new_n11591_1, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607_1, new_n11608, new_n11609, new_n11610, new_n11611,
    new_n11612, new_n11613, new_n11614, new_n11615_1, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630_1, new_n11631, new_n11632, new_n11633,
    new_n11634, new_n11635, new_n11636, new_n11637, new_n11638, new_n11639,
    new_n11640, new_n11641, new_n11642, new_n11643, new_n11644, new_n11645,
    new_n11646, new_n11647_1, new_n11648, new_n11649, new_n11650,
    new_n11651, new_n11652, new_n11653, new_n11654, new_n11655, new_n11656,
    new_n11657, new_n11658, new_n11659, new_n11660, new_n11661, new_n11662,
    new_n11663, new_n11664, new_n11665, new_n11666, new_n11667_1,
    new_n11668, new_n11669, new_n11670, new_n11671, new_n11672, new_n11673,
    new_n11674_1, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682_1, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706, new_n11707,
    new_n11708, new_n11709, new_n11710_1, new_n11712_1, new_n11714,
    new_n11715, new_n11716, new_n11717, new_n11719, new_n11720, new_n11721,
    new_n11722, new_n11723, new_n11724_1, new_n11725, new_n11726,
    new_n11727, new_n11728, new_n11729, new_n11730, new_n11731, new_n11732,
    new_n11733, new_n11734, new_n11735, new_n11736_1, new_n11737,
    new_n11738, new_n11739, new_n11740, new_n11741_1, new_n11743,
    new_n11744, new_n11745, new_n11746, new_n11747, new_n11748,
    new_n11749_1, new_n11750, new_n11751, new_n11752, new_n11753,
    new_n11754, new_n11755, new_n11757, new_n11758, new_n11759, new_n11760,
    new_n11761, new_n11762, new_n11763, new_n11764, new_n11765, new_n11766,
    new_n11767, new_n11768, new_n11769, new_n11770_1, new_n11771_1,
    new_n11772, new_n11773, new_n11774, new_n11775_1, new_n11776,
    new_n11777, new_n11778, new_n11779, new_n11780, new_n11781, new_n11782,
    new_n11783, new_n11784, new_n11785, new_n11786, new_n11787, new_n11788,
    new_n11789, new_n11790, new_n11791, new_n11792, new_n11793, new_n11794,
    new_n11795, new_n11796, new_n11797, new_n11798, new_n11799, new_n11800,
    new_n11801, new_n11802, new_n11803, new_n11804, new_n11805, new_n11806,
    new_n11807, new_n11808, new_n11809, new_n11810, new_n11811, new_n11812,
    new_n11813, new_n11814, new_n11815, new_n11816, new_n11817,
    new_n11818_1, new_n11819, new_n11820, new_n11821, new_n11822,
    new_n11823, new_n11824, new_n11825, new_n11826, new_n11827, new_n11828,
    new_n11829, new_n11830, new_n11831, new_n11832, new_n11833, new_n11834,
    new_n11835, new_n11836, new_n11837_1, new_n11838, new_n11839,
    new_n11840, new_n11841_1, new_n11842_1, new_n11843_1, new_n11844,
    new_n11845, new_n11846, new_n11847, new_n11848, new_n11849, new_n11850,
    new_n11851, new_n11852, new_n11853, new_n11854, new_n11855, new_n11856,
    new_n11857, new_n11858, new_n11859, new_n11860, new_n11861, new_n11862,
    new_n11863, new_n11864, new_n11865, new_n11866, new_n11867, new_n11868,
    new_n11869, new_n11870, new_n11871, new_n11872, new_n11873, new_n11874,
    new_n11875, new_n11876, new_n11877, new_n11878, new_n11879, new_n11880,
    new_n11881, new_n11882, new_n11883, new_n11884, new_n11885, new_n11886,
    new_n11887, new_n11888, new_n11889, new_n11890, new_n11891, new_n11892,
    new_n11893, new_n11894, new_n11895, new_n11896, new_n11897,
    new_n11898_1, new_n11899, new_n11900, new_n11901, new_n11902,
    new_n11903, new_n11904, new_n11905_1, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917, new_n11918, new_n11919,
    new_n11920, new_n11921, new_n11922, new_n11923, new_n11924, new_n11925,
    new_n11926_1, new_n11927, new_n11928, new_n11929, new_n11930,
    new_n11931, new_n11932, new_n11933, new_n11934, new_n11935, new_n11936,
    new_n11937, new_n11938, new_n11939, new_n11940, new_n11941, new_n11942,
    new_n11943, new_n11944, new_n11945, new_n11946, new_n11947, new_n11948,
    new_n11949, new_n11950, new_n11951, new_n11952, new_n11953, new_n11954,
    new_n11955, new_n11956, new_n11957, new_n11958, new_n11959, new_n11960,
    new_n11961, new_n11962, new_n11963, new_n11964, new_n11965_1,
    new_n11966, new_n11967, new_n11968, new_n11969, new_n11970, new_n11971,
    new_n11972, new_n11973, new_n11974, new_n11975, new_n11976, new_n11977,
    new_n11978, new_n11979, new_n11980_1, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11998, new_n11999,
    new_n12000_1, new_n12001, new_n12002, new_n12003_1, new_n12004,
    new_n12005, new_n12006, new_n12007, new_n12008, new_n12009, new_n12010,
    new_n12011_1, new_n12012, new_n12013, new_n12014, new_n12015,
    new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021,
    new_n12022, new_n12023, new_n12024, new_n12025, new_n12026, new_n12027,
    new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033,
    new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039,
    new_n12040, new_n12041, new_n12042, new_n12043, new_n12044, new_n12045,
    new_n12046, new_n12047, new_n12048, new_n12049, new_n12050, new_n12051,
    new_n12052, new_n12053, new_n12054, new_n12055, new_n12056, new_n12057,
    new_n12058, new_n12059, new_n12060, new_n12061, new_n12062, new_n12063,
    new_n12064, new_n12065, new_n12066, new_n12067, new_n12068, new_n12069,
    new_n12070, new_n12071, new_n12072_1, new_n12073, new_n12074,
    new_n12075, new_n12076, new_n12077, new_n12078, new_n12079, new_n12080,
    new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086,
    new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092,
    new_n12093, new_n12095, new_n12096, new_n12097, new_n12098, new_n12099,
    new_n12100, new_n12101, new_n12102, new_n12103, new_n12104, new_n12105,
    new_n12106, new_n12107, new_n12108, new_n12109, new_n12110, new_n12111,
    new_n12112, new_n12113_1, new_n12114, new_n12115, new_n12116,
    new_n12117, new_n12118, new_n12119, new_n12120, new_n12121_1,
    new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127,
    new_n12128, new_n12129, new_n12130, new_n12131_1, new_n12132,
    new_n12133, new_n12134, new_n12135, new_n12136, new_n12137, new_n12138,
    new_n12139, new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145, new_n12146_1, new_n12147, new_n12148, new_n12149,
    new_n12150, new_n12151, new_n12152_1, new_n12153_1, new_n12154,
    new_n12155, new_n12156, new_n12157_1, new_n12158_1, new_n12159,
    new_n12160, new_n12161_1, new_n12162, new_n12163, new_n12164,
    new_n12165, new_n12166, new_n12167, new_n12168, new_n12169, new_n12170,
    new_n12171, new_n12172, new_n12173, new_n12174, new_n12175, new_n12176,
    new_n12177, new_n12178, new_n12179_1, new_n12180, new_n12181,
    new_n12182, new_n12183, new_n12184, new_n12185, new_n12186, new_n12187,
    new_n12188, new_n12189, new_n12190, new_n12191, new_n12192_1,
    new_n12193, new_n12194, new_n12195, new_n12196, new_n12197, new_n12198,
    new_n12199, new_n12200, new_n12201, new_n12202, new_n12203, new_n12204,
    new_n12205, new_n12206, new_n12207, new_n12208, new_n12209_1,
    new_n12210, new_n12211, new_n12212, new_n12213, new_n12214, new_n12215,
    new_n12216, new_n12217, new_n12218, new_n12219, new_n12220, new_n12221,
    new_n12222, new_n12223_1, new_n12224, new_n12225_1, new_n12226,
    new_n12227, new_n12228_1, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235_1, new_n12236,
    new_n12237, new_n12238, new_n12239, new_n12240, new_n12241, new_n12242,
    new_n12243, new_n12244, new_n12245, new_n12246, new_n12247, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299, new_n12300, new_n12301,
    new_n12302_1, new_n12303, new_n12304_1, new_n12305, new_n12306,
    new_n12307, new_n12308, new_n12309, new_n12310, new_n12311, new_n12312,
    new_n12313, new_n12314, new_n12316, new_n12317, new_n12318, new_n12319,
    new_n12320, new_n12321, new_n12322, new_n12323, new_n12324_1,
    new_n12325_1, new_n12326, new_n12327, new_n12328, new_n12329_1,
    new_n12330_1, new_n12331, new_n12332, new_n12333, new_n12334,
    new_n12335, new_n12336, new_n12337, new_n12338, new_n12339, new_n12340,
    new_n12341_1, new_n12342, new_n12343, new_n12344, new_n12345,
    new_n12346_1, new_n12347, new_n12348, new_n12349_1, new_n12350,
    new_n12351, new_n12352, new_n12353, new_n12354, new_n12355, new_n12356,
    new_n12357, new_n12358, new_n12359, new_n12360, new_n12361, new_n12362,
    new_n12363, new_n12364_1, new_n12365, new_n12366, new_n12367,
    new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373,
    new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380_1, new_n12381, new_n12382, new_n12383_1, new_n12384_1,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397_1, new_n12398_1, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408_1, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446_1, new_n12447,
    new_n12448, new_n12449_1, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461_1, new_n12462_1, new_n12463,
    new_n12464, new_n12465, new_n12466, new_n12467_1, new_n12468,
    new_n12469_1, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495_1, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507_1,
    new_n12508, new_n12509, new_n12510, new_n12511, new_n12512, new_n12513,
    new_n12514, new_n12515_1, new_n12516_1, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540_1, new_n12541,
    new_n12542, new_n12543, new_n12544, new_n12545_1, new_n12546_1,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552_1, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561,
    new_n12562_1, new_n12563, new_n12564, new_n12565, new_n12566_1,
    new_n12567, new_n12568, new_n12569_1, new_n12570, new_n12571,
    new_n12572, new_n12573, new_n12574, new_n12575, new_n12576, new_n12577,
    new_n12578, new_n12579, new_n12580, new_n12581, new_n12582, new_n12583,
    new_n12584, new_n12585, new_n12586, new_n12587_1, new_n12588,
    new_n12589, new_n12590, new_n12591, new_n12592, new_n12593_1,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607_1, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620_1, new_n12621_1,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626_1,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648, new_n12649, new_n12650_1,
    new_n12651, new_n12652, new_n12653, new_n12654_1, new_n12655,
    new_n12656, new_n12657_1, new_n12658, new_n12659, new_n12660,
    new_n12661, new_n12662, new_n12663, new_n12664, new_n12665_1,
    new_n12666, new_n12667, new_n12668, new_n12669, new_n12670_1,
    new_n12671, new_n12672, new_n12673, new_n12674, new_n12675, new_n12676,
    new_n12677, new_n12678, new_n12679, new_n12680, new_n12681, new_n12682,
    new_n12683, new_n12684, new_n12685, new_n12686, new_n12687, new_n12688,
    new_n12689, new_n12690, new_n12691, new_n12692, new_n12693, new_n12694,
    new_n12695, new_n12696, new_n12697, new_n12698, new_n12699, new_n12700,
    new_n12701, new_n12702_1, new_n12703, new_n12704, new_n12705,
    new_n12706, new_n12707_1, new_n12708, new_n12709, new_n12710,
    new_n12711, new_n12712, new_n12713, new_n12714, new_n12715, new_n12716,
    new_n12717, new_n12718, new_n12719, new_n12720, new_n12721, new_n12722,
    new_n12723, new_n12724, new_n12725_1, new_n12726, new_n12727_1,
    new_n12728, new_n12729, new_n12730, new_n12731, new_n12732, new_n12733,
    new_n12734, new_n12735, new_n12736, new_n12737, new_n12738, new_n12739,
    new_n12740_1, new_n12741, new_n12743, new_n12744, new_n12745,
    new_n12746_1, new_n12747, new_n12748, new_n12749, new_n12750,
    new_n12751, new_n12752, new_n12753, new_n12754, new_n12755,
    new_n12756_1, new_n12757, new_n12758, new_n12759, new_n12760,
    new_n12761, new_n12762, new_n12763, new_n12764, new_n12765, new_n12766,
    new_n12767, new_n12768, new_n12769, new_n12770, new_n12771, new_n12772,
    new_n12773, new_n12774, new_n12775, new_n12776, new_n12777, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783_1,
    new_n12784, new_n12785, new_n12786, new_n12787, new_n12788, new_n12789,
    new_n12790, new_n12791, new_n12792, new_n12793, new_n12794, new_n12795,
    new_n12796, new_n12797, new_n12798, new_n12799, new_n12800,
    new_n12801_1, new_n12802, new_n12803, new_n12804, new_n12805,
    new_n12806, new_n12807, new_n12808, new_n12809, new_n12810,
    new_n12811_1, new_n12812_1, new_n12813, new_n12814, new_n12815,
    new_n12816_1, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821_1, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12837,
    new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843_1, new_n12844, new_n12845, new_n12846, new_n12847,
    new_n12848, new_n12849, new_n12850, new_n12851, new_n12852, new_n12853,
    new_n12854, new_n12855, new_n12856, new_n12857, new_n12858, new_n12859,
    new_n12860, new_n12861_1, new_n12862, new_n12863, new_n12864_1,
    new_n12865_1, new_n12866, new_n12867, new_n12868, new_n12870_1,
    new_n12871_1, new_n12872, new_n12873_1, new_n12874, new_n12875_1,
    new_n12876, new_n12877, new_n12878, new_n12879, new_n12880, new_n12881,
    new_n12882, new_n12883, new_n12884, new_n12885, new_n12886, new_n12887,
    new_n12888, new_n12889, new_n12890, new_n12891, new_n12892_1,
    new_n12893, new_n12894, new_n12895, new_n12896, new_n12897, new_n12898,
    new_n12899, new_n12900_1, new_n12901, new_n12902, new_n12903,
    new_n12904_1, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917_1, new_n12918, new_n12919,
    new_n12920, new_n12921, new_n12922, new_n12923, new_n12924, new_n12925,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941_1, new_n12942_1,
    new_n12943, new_n12944, new_n12945, new_n12946, new_n12947, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956_1, new_n12957, new_n12958, new_n12959,
    new_n12960, new_n12961, new_n12962, new_n12963, new_n12964, new_n12965,
    new_n12966, new_n12967, new_n12968, new_n12969, new_n12970, new_n12971,
    new_n12972, new_n12973, new_n12974, new_n12975, new_n12976, new_n12977,
    new_n12978_1, new_n12979, new_n12980_1, new_n12981, new_n12982,
    new_n12983, new_n12984, new_n12985_1, new_n12986, new_n12987_1,
    new_n12988, new_n12989, new_n12990, new_n12991, new_n12992_1,
    new_n12993, new_n12994, new_n12995, new_n12996, new_n12997, new_n12998,
    new_n12999, new_n13000, new_n13001, new_n13002, new_n13003, new_n13004,
    new_n13005_1, new_n13006, new_n13007, new_n13008, new_n13009,
    new_n13010, new_n13011, new_n13012, new_n13013, new_n13014, new_n13015,
    new_n13016, new_n13017, new_n13018, new_n13019, new_n13020, new_n13021,
    new_n13022, new_n13023, new_n13024, new_n13025, new_n13026_1,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043_1,
    new_n13044_1, new_n13045, new_n13046, new_n13047, new_n13048_1,
    new_n13049, new_n13050, new_n13051, new_n13052, new_n13053,
    new_n13054_1, new_n13055, new_n13056, new_n13057, new_n13058,
    new_n13059, new_n13060, new_n13061, new_n13062, new_n13063, new_n13064,
    new_n13065, new_n13066, new_n13067, new_n13068, new_n13069, new_n13070,
    new_n13071, new_n13073, new_n13074_1, new_n13076, new_n13077,
    new_n13078, new_n13079, new_n13080, new_n13081, new_n13082_1,
    new_n13083, new_n13084, new_n13085, new_n13086, new_n13087, new_n13088,
    new_n13089, new_n13090, new_n13091, new_n13092, new_n13093, new_n13094,
    new_n13095, new_n13096_1, new_n13097, new_n13098, new_n13099,
    new_n13100, new_n13101, new_n13102, new_n13103, new_n13104, new_n13105,
    new_n13106, new_n13107, new_n13108, new_n13109, new_n13110_1,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115,
    new_n13116_1, new_n13117, new_n13118, new_n13119, new_n13120,
    new_n13121, new_n13122_1, new_n13123, new_n13124, new_n13125,
    new_n13126, new_n13127, new_n13128, new_n13129, new_n13130, new_n13131,
    new_n13132, new_n13133, new_n13134, new_n13135, new_n13136,
    new_n13137_1, new_n13138, new_n13139, new_n13140, new_n13141_1,
    new_n13142, new_n13143, new_n13144_1, new_n13145, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168_1, new_n13169,
    new_n13170, new_n13171, new_n13172, new_n13173, new_n13174, new_n13175,
    new_n13176, new_n13177, new_n13178, new_n13179, new_n13180, new_n13181,
    new_n13182, new_n13183, new_n13184, new_n13185, new_n13186, new_n13187,
    new_n13188, new_n13189, new_n13190_1, new_n13191, new_n13192,
    new_n13193, new_n13194, new_n13195, new_n13196, new_n13197,
    new_n13199_1, new_n13200, new_n13201, new_n13202, new_n13203,
    new_n13204_1, new_n13205, new_n13206, new_n13207, new_n13208,
    new_n13209_1, new_n13210, new_n13211, new_n13212, new_n13213,
    new_n13214, new_n13215, new_n13216, new_n13217, new_n13218, new_n13219,
    new_n13220, new_n13221, new_n13222, new_n13223, new_n13224, new_n13225,
    new_n13226, new_n13227, new_n13228, new_n13229, new_n13230, new_n13231,
    new_n13232, new_n13233, new_n13234, new_n13235, new_n13236, new_n13237,
    new_n13238, new_n13239, new_n13240, new_n13241, new_n13242, new_n13243,
    new_n13244, new_n13245, new_n13246, new_n13247, new_n13248, new_n13249,
    new_n13250, new_n13251, new_n13252, new_n13253, new_n13254, new_n13255,
    new_n13256, new_n13257, new_n13258, new_n13259, new_n13260, new_n13261,
    new_n13262, new_n13263_1, new_n13264, new_n13265, new_n13266,
    new_n13267, new_n13268, new_n13269, new_n13270_1, new_n13271,
    new_n13272, new_n13273_1, new_n13274, new_n13275, new_n13276,
    new_n13277, new_n13278, new_n13279, new_n13280, new_n13281, new_n13282,
    new_n13283, new_n13284, new_n13285_1, new_n13286, new_n13287,
    new_n13288, new_n13289, new_n13290, new_n13291, new_n13292, new_n13293,
    new_n13294, new_n13295, new_n13296, new_n13297, new_n13298, new_n13299,
    new_n13300, new_n13301, new_n13302, new_n13303, new_n13304, new_n13305,
    new_n13306, new_n13307, new_n13308, new_n13309, new_n13310, new_n13311,
    new_n13312, new_n13313, new_n13314, new_n13315, new_n13316, new_n13317,
    new_n13318, new_n13319_1, new_n13320, new_n13321, new_n13322,
    new_n13323, new_n13324, new_n13325, new_n13326, new_n13327, new_n13328,
    new_n13329, new_n13330, new_n13331, new_n13332, new_n13333_1,
    new_n13334, new_n13335, new_n13336, new_n13337, new_n13338_1,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13346, new_n13347, new_n13348, new_n13349, new_n13350,
    new_n13351, new_n13352, new_n13353, new_n13354, new_n13355, new_n13356,
    new_n13357, new_n13358, new_n13359, new_n13360, new_n13361, new_n13362,
    new_n13363, new_n13364, new_n13365, new_n13366, new_n13367_1,
    new_n13368, new_n13369, new_n13370, new_n13371, new_n13372, new_n13373,
    new_n13374, new_n13375, new_n13376, new_n13377, new_n13378, new_n13379,
    new_n13380, new_n13381, new_n13382, new_n13383, new_n13384, new_n13385,
    new_n13386, new_n13387, new_n13388, new_n13389, new_n13390, new_n13391,
    new_n13392, new_n13393, new_n13394, new_n13395, new_n13396, new_n13397,
    new_n13398, new_n13399, new_n13400, new_n13401, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407_1, new_n13408,
    new_n13409_1, new_n13410, new_n13411, new_n13412, new_n13413,
    new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419_1, new_n13420, new_n13421, new_n13422, new_n13423,
    new_n13424_1, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453_1, new_n13454, new_n13455, new_n13456_1, new_n13457_1,
    new_n13458, new_n13459, new_n13460_1, new_n13462, new_n13463,
    new_n13464, new_n13465, new_n13466, new_n13467, new_n13468, new_n13469,
    new_n13470, new_n13471, new_n13472, new_n13473, new_n13474, new_n13475,
    new_n13476, new_n13477_1, new_n13478, new_n13479, new_n13480,
    new_n13481, new_n13482, new_n13483, new_n13484_1, new_n13485,
    new_n13486_1, new_n13487_1, new_n13488, new_n13489, new_n13490_1,
    new_n13491, new_n13492, new_n13493, new_n13494_1, new_n13495,
    new_n13496, new_n13497, new_n13498, new_n13499, new_n13500_1,
    new_n13501_1, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506_1, new_n13507, new_n13508, new_n13509, new_n13510,
    new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13533, new_n13534, new_n13535,
    new_n13536, new_n13537, new_n13538, new_n13539, new_n13540, new_n13542,
    new_n13543, new_n13544, new_n13545, new_n13546, new_n13547,
    new_n13548_1, new_n13549_1, new_n13550, new_n13551_1, new_n13552,
    new_n13553, new_n13554, new_n13555, new_n13556, new_n13557, new_n13558,
    new_n13559, new_n13560, new_n13561, new_n13562, new_n13563, new_n13564,
    new_n13565, new_n13566, new_n13567, new_n13568, new_n13569, new_n13570,
    new_n13571, new_n13572, new_n13573, new_n13574, new_n13575, new_n13576,
    new_n13577, new_n13578, new_n13579, new_n13580, new_n13581, new_n13582,
    new_n13583, new_n13584, new_n13585, new_n13586, new_n13587, new_n13588,
    new_n13589, new_n13590, new_n13591, new_n13592, new_n13593, new_n13594,
    new_n13595, new_n13596, new_n13597, new_n13598, new_n13599, new_n13600,
    new_n13601, new_n13602_1, new_n13603, new_n13604, new_n13605,
    new_n13606, new_n13607, new_n13608, new_n13609, new_n13610, new_n13611,
    new_n13612, new_n13613, new_n13614, new_n13615, new_n13616, new_n13617,
    new_n13618, new_n13619, new_n13620, new_n13621, new_n13622, new_n13623,
    new_n13624, new_n13625, new_n13626_1, new_n13627, new_n13628,
    new_n13629, new_n13630, new_n13631, new_n13632, new_n13633, new_n13634,
    new_n13635, new_n13636, new_n13637, new_n13638, new_n13639, new_n13640,
    new_n13641, new_n13642, new_n13643, new_n13644, new_n13645, new_n13646,
    new_n13647, new_n13648, new_n13649, new_n13650, new_n13651, new_n13652,
    new_n13653, new_n13654, new_n13655, new_n13656, new_n13657, new_n13658,
    new_n13659, new_n13660, new_n13661, new_n13662, new_n13663, new_n13664,
    new_n13665, new_n13666, new_n13667, new_n13668_1, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677_1, new_n13678, new_n13679, new_n13680,
    new_n13681, new_n13682, new_n13683_1, new_n13684, new_n13685,
    new_n13686, new_n13687, new_n13688, new_n13689, new_n13690, new_n13691,
    new_n13692, new_n13693, new_n13694, new_n13695, new_n13696, new_n13697,
    new_n13698, new_n13699, new_n13700, new_n13701, new_n13702, new_n13703,
    new_n13704, new_n13705, new_n13706, new_n13707, new_n13708_1,
    new_n13710_1, new_n13713, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719_1, new_n13720, new_n13721, new_n13722_1,
    new_n13723, new_n13724, new_n13725, new_n13726, new_n13727, new_n13728,
    new_n13729, new_n13730, new_n13731, new_n13732, new_n13733, new_n13734,
    new_n13735, new_n13736, new_n13737, new_n13738, new_n13739, new_n13740,
    new_n13741, new_n13742, new_n13743, new_n13744, new_n13745, new_n13746,
    new_n13747, new_n13748, new_n13749, new_n13750, new_n13751, new_n13752,
    new_n13753, new_n13754_1, new_n13755, new_n13756, new_n13757,
    new_n13758, new_n13759, new_n13760, new_n13761, new_n13762, new_n13763,
    new_n13764_1, new_n13765, new_n13766, new_n13767, new_n13768,
    new_n13769, new_n13770, new_n13771, new_n13772, new_n13773, new_n13774,
    new_n13775_1, new_n13776, new_n13777, new_n13778, new_n13779,
    new_n13780, new_n13781_1, new_n13782, new_n13783_1, new_n13784,
    new_n13785, new_n13786, new_n13787, new_n13788, new_n13789, new_n13790,
    new_n13791, new_n13792, new_n13793, new_n13794, new_n13795, new_n13796,
    new_n13797, new_n13798_1, new_n13799, new_n13800, new_n13801,
    new_n13802, new_n13803, new_n13804, new_n13805, new_n13806, new_n13807,
    new_n13808, new_n13809, new_n13810, new_n13811, new_n13812, new_n13813,
    new_n13814, new_n13815, new_n13816, new_n13817, new_n13818, new_n13819,
    new_n13820, new_n13821, new_n13822, new_n13823, new_n13824, new_n13825,
    new_n13826, new_n13827, new_n13828, new_n13829, new_n13830, new_n13831,
    new_n13832, new_n13833, new_n13834, new_n13835_1, new_n13836,
    new_n13837, new_n13838, new_n13839, new_n13840, new_n13841, new_n13842,
    new_n13843, new_n13844, new_n13845, new_n13846, new_n13847, new_n13848,
    new_n13849, new_n13850_1, new_n13851_1, new_n13852, new_n13853,
    new_n13854, new_n13855, new_n13856, new_n13857, new_n13858, new_n13859,
    new_n13860, new_n13861, new_n13862, new_n13863, new_n13864, new_n13865,
    new_n13866, new_n13867, new_n13868, new_n13869, new_n13870, new_n13871,
    new_n13872, new_n13873, new_n13874, new_n13875, new_n13876, new_n13877,
    new_n13878, new_n13879, new_n13880, new_n13881, new_n13882, new_n13883,
    new_n13884, new_n13885, new_n13886, new_n13887, new_n13888, new_n13889,
    new_n13890, new_n13891, new_n13892, new_n13893, new_n13894, new_n13895,
    new_n13897, new_n13898, new_n13899, new_n13900, new_n13901, new_n13902,
    new_n13903, new_n13904, new_n13905, new_n13906, new_n13907, new_n13908,
    new_n13909, new_n13910, new_n13911, new_n13912_1, new_n13913,
    new_n13914_1, new_n13915, new_n13916, new_n13917, new_n13918,
    new_n13919, new_n13920, new_n13921, new_n13922_1, new_n13923_1,
    new_n13924, new_n13925, new_n13926, new_n13927, new_n13928, new_n13929,
    new_n13930, new_n13931, new_n13932, new_n13933, new_n13934, new_n13935,
    new_n13936, new_n13937, new_n13938, new_n13939, new_n13940, new_n13941,
    new_n13942, new_n13943, new_n13944, new_n13945, new_n13946, new_n13947,
    new_n13948, new_n13949, new_n13950, new_n13951_1, new_n13952,
    new_n13953, new_n13954, new_n13955, new_n13956, new_n13957, new_n13958,
    new_n13959, new_n13960, new_n13961, new_n13962, new_n13963, new_n13964,
    new_n13965, new_n13966, new_n13967, new_n13968, new_n13969, new_n13970,
    new_n13971, new_n13972, new_n13973, new_n13974, new_n13975, new_n13976,
    new_n13977, new_n13978, new_n13979, new_n13980, new_n13981, new_n13982,
    new_n13983, new_n13984, new_n13985, new_n13986, new_n13987, new_n13988,
    new_n13989, new_n13990, new_n13991, new_n13992, new_n13993, new_n13994,
    new_n13995, new_n13996, new_n13997, new_n13998, new_n13999, new_n14000,
    new_n14001, new_n14002, new_n14003, new_n14004_1, new_n14005,
    new_n14006, new_n14007, new_n14008, new_n14009, new_n14010, new_n14011,
    new_n14012, new_n14013, new_n14014, new_n14015, new_n14016, new_n14017,
    new_n14018, new_n14019, new_n14020, new_n14021, new_n14022, new_n14023,
    new_n14024, new_n14025, new_n14026, new_n14027, new_n14028, new_n14029,
    new_n14030, new_n14031, new_n14032, new_n14033, new_n14034, new_n14035,
    new_n14036_1, new_n14037, new_n14038, new_n14039, new_n14040,
    new_n14041, new_n14042, new_n14043, new_n14044, new_n14045, new_n14046,
    new_n14047, new_n14048, new_n14049, new_n14050, new_n14051, new_n14052,
    new_n14053, new_n14054, new_n14055, new_n14056, new_n14057, new_n14058,
    new_n14059_1, new_n14060, new_n14061, new_n14062, new_n14063,
    new_n14064, new_n14065, new_n14066, new_n14067, new_n14068, new_n14069,
    new_n14070, new_n14071_1, new_n14072, new_n14073, new_n14074,
    new_n14075, new_n14076, new_n14077, new_n14078, new_n14079, new_n14080,
    new_n14081_1, new_n14082, new_n14083, new_n14084, new_n14085,
    new_n14086, new_n14087, new_n14088, new_n14089, new_n14090_1,
    new_n14091, new_n14092, new_n14093, new_n14094, new_n14095_1,
    new_n14096, new_n14097, new_n14098, new_n14099, new_n14100, new_n14101,
    new_n14102, new_n14103, new_n14104, new_n14105, new_n14106,
    new_n14107_1, new_n14108, new_n14109, new_n14110, new_n14111,
    new_n14112, new_n14113, new_n14114, new_n14115, new_n14116, new_n14117,
    new_n14118, new_n14119, new_n14120, new_n14121_1, new_n14122,
    new_n14123, new_n14124, new_n14125, new_n14126_1, new_n14127,
    new_n14128, new_n14129, new_n14130_1, new_n14131, new_n14132,
    new_n14133, new_n14134, new_n14135, new_n14136_1, new_n14137,
    new_n14138, new_n14139, new_n14140, new_n14141, new_n14142, new_n14143,
    new_n14144, new_n14145, new_n14146, new_n14147_1, new_n14148_1,
    new_n14149, new_n14150, new_n14151, new_n14152, new_n14153, new_n14154,
    new_n14155, new_n14156, new_n14157, new_n14159, new_n14162, new_n14163,
    new_n14164, new_n14165, new_n14166, new_n14167, new_n14168, new_n14169,
    new_n14170, new_n14171, new_n14172, new_n14173, new_n14175, new_n14178,
    new_n14179, new_n14180, new_n14181, new_n14182, new_n14183, new_n14184,
    new_n14185, new_n14186, new_n14187, new_n14188, new_n14189,
    new_n14190_1, new_n14191, new_n14192, new_n14193, new_n14194,
    new_n14195, new_n14196, new_n14197, new_n14198, new_n14199, new_n14200,
    new_n14201, new_n14202, new_n14203, new_n14204, new_n14205, new_n14206,
    new_n14207, new_n14210, new_n14211_1, new_n14212, new_n14213,
    new_n14214, new_n14215, new_n14216, new_n14217, new_n14218, new_n14219,
    new_n14220, new_n14221, new_n14222_1, new_n14223, new_n14224,
    new_n14225, new_n14226, new_n14227, new_n14228, new_n14229,
    new_n14230_1, new_n14231, new_n14232, new_n14233, new_n14234,
    new_n14235, new_n14236, new_n14237, new_n14238, new_n14239, new_n14240,
    new_n14241, new_n14242, new_n14243, new_n14244, new_n14245, new_n14246,
    new_n14247, new_n14248, new_n14249, new_n14250, new_n14251, new_n14252,
    new_n14253, new_n14254, new_n14255, new_n14256, new_n14257, new_n14258,
    new_n14259, new_n14260, new_n14261, new_n14262, new_n14263, new_n14264,
    new_n14265, new_n14266, new_n14267_1, new_n14268, new_n14269,
    new_n14270, new_n14271_1, new_n14272, new_n14273, new_n14274,
    new_n14275_1, new_n14276, new_n14277_1, new_n14278, new_n14279,
    new_n14280, new_n14281, new_n14282, new_n14283, new_n14284, new_n14285,
    new_n14286, new_n14287, new_n14288, new_n14289, new_n14290, new_n14291,
    new_n14292, new_n14293, new_n14294_1, new_n14295, new_n14296,
    new_n14297, new_n14298, new_n14299, new_n14300, new_n14301, new_n14302,
    new_n14303, new_n14304, new_n14305, new_n14306, new_n14307, new_n14308,
    new_n14309, new_n14310_1, new_n14311, new_n14312, new_n14313,
    new_n14314, new_n14315, new_n14316, new_n14317, new_n14318, new_n14319,
    new_n14320, new_n14321, new_n14322, new_n14323_1, new_n14324,
    new_n14325, new_n14326_1, new_n14327, new_n14328, new_n14329,
    new_n14330, new_n14331, new_n14332, new_n14333, new_n14334, new_n14335,
    new_n14336, new_n14337, new_n14338, new_n14339, new_n14340, new_n14341,
    new_n14342_1, new_n14343, new_n14344, new_n14345_1, new_n14346,
    new_n14347, new_n14348, new_n14349, new_n14350, new_n14351, new_n14352,
    new_n14353_1, new_n14354, new_n14355, new_n14356, new_n14357,
    new_n14358, new_n14359, new_n14360, new_n14361, new_n14362, new_n14363,
    new_n14364_1, new_n14365, new_n14366, new_n14367, new_n14368,
    new_n14369, new_n14370, new_n14371, new_n14372, new_n14373, new_n14374,
    new_n14375_1, new_n14376, new_n14377, new_n14378, new_n14379,
    new_n14380, new_n14381, new_n14382, new_n14383, new_n14384, new_n14385,
    new_n14386, new_n14387, new_n14388, new_n14389, new_n14390, new_n14391,
    new_n14392, new_n14393, new_n14394, new_n14395, new_n14396, new_n14397,
    new_n14398, new_n14399, new_n14401, new_n14403, new_n14404, new_n14405,
    new_n14406, new_n14407, new_n14408, new_n14409, new_n14410, new_n14411,
    new_n14412_1, new_n14413, new_n14414_1, new_n14415, new_n14416,
    new_n14417, new_n14418, new_n14419, new_n14420, new_n14421, new_n14422,
    new_n14423, new_n14424, new_n14425, new_n14426, new_n14427, new_n14428,
    new_n14429, new_n14430, new_n14431, new_n14432, new_n14433, new_n14434,
    new_n14435, new_n14436, new_n14437, new_n14438, new_n14439,
    new_n14440_1, new_n14441, new_n14442, new_n14443, new_n14444,
    new_n14445, new_n14446, new_n14447, new_n14448, new_n14449, new_n14450,
    new_n14451, new_n14452, new_n14453, new_n14454, new_n14455, new_n14456,
    new_n14457_1, new_n14458, new_n14459, new_n14460, new_n14461,
    new_n14462, new_n14463, new_n14464_1, new_n14465, new_n14466,
    new_n14467, new_n14468, new_n14469, new_n14470, new_n14471_1,
    new_n14472, new_n14473, new_n14474, new_n14475_1, new_n14476,
    new_n14477, new_n14478, new_n14479, new_n14480, new_n14481, new_n14482,
    new_n14483, new_n14484, new_n14485, new_n14486, new_n14487, new_n14488,
    new_n14489, new_n14490, new_n14491, new_n14492, new_n14493, new_n14494,
    new_n14495, new_n14496, new_n14497, new_n14498, new_n14499, new_n14500,
    new_n14501, new_n14502, new_n14503, new_n14504, new_n14505, new_n14506,
    new_n14507, new_n14508, new_n14509, new_n14510_1, new_n14511,
    new_n14512, new_n14513, new_n14514, new_n14515, new_n14516, new_n14517,
    new_n14518, new_n14519, new_n14520, new_n14521, new_n14522, new_n14523,
    new_n14524, new_n14525, new_n14526, new_n14527, new_n14528, new_n14529,
    new_n14530, new_n14531, new_n14532, new_n14533, new_n14534, new_n14535,
    new_n14536, new_n14537, new_n14538, new_n14539, new_n14540,
    new_n14541_1, new_n14542, new_n14543, new_n14545, new_n14546_1,
    new_n14547_1, new_n14548, new_n14549, new_n14550, new_n14551,
    new_n14552, new_n14553, new_n14554, new_n14555, new_n14556, new_n14557,
    new_n14558, new_n14559, new_n14560, new_n14561, new_n14562, new_n14563,
    new_n14564, new_n14565, new_n14566, new_n14567, new_n14568, new_n14569,
    new_n14570_1, new_n14571, new_n14572, new_n14573, new_n14574,
    new_n14575_1, new_n14576_1, new_n14577, new_n14578, new_n14579,
    new_n14580, new_n14581, new_n14582, new_n14583, new_n14584, new_n14585,
    new_n14586, new_n14587, new_n14588, new_n14589, new_n14590, new_n14591,
    new_n14592, new_n14593_1, new_n14594, new_n14595, new_n14596,
    new_n14597, new_n14598, new_n14599, new_n14600, new_n14601, new_n14602,
    new_n14603_1, new_n14604, new_n14605, new_n14606, new_n14607,
    new_n14608, new_n14609, new_n14610, new_n14611, new_n14612, new_n14613,
    new_n14614, new_n14615, new_n14616, new_n14617, new_n14618, new_n14619,
    new_n14620, new_n14621, new_n14622, new_n14623, new_n14624, new_n14625,
    new_n14626, new_n14627, new_n14628, new_n14629, new_n14630, new_n14631,
    new_n14632, new_n14633_1, new_n14634, new_n14635, new_n14636_1,
    new_n14637, new_n14638, new_n14639, new_n14640, new_n14641, new_n14642,
    new_n14643, new_n14644, new_n14645, new_n14646, new_n14647, new_n14648,
    new_n14649, new_n14650, new_n14651, new_n14652, new_n14653, new_n14654,
    new_n14655, new_n14656, new_n14657, new_n14658, new_n14659, new_n14660,
    new_n14661, new_n14662, new_n14663, new_n14664, new_n14665, new_n14666,
    new_n14667, new_n14668, new_n14669, new_n14670, new_n14671, new_n14672,
    new_n14673, new_n14674, new_n14675, new_n14676, new_n14677, new_n14678,
    new_n14679, new_n14680_1, new_n14681, new_n14682, new_n14683,
    new_n14685, new_n14686, new_n14687, new_n14688, new_n14689, new_n14690,
    new_n14691, new_n14692_1, new_n14693, new_n14694, new_n14695,
    new_n14696, new_n14697, new_n14698, new_n14699, new_n14700,
    new_n14701_1, new_n14702_1, new_n14703, new_n14704_1, new_n14705,
    new_n14706, new_n14707, new_n14708, new_n14709, new_n14710, new_n14711,
    new_n14712, new_n14713, new_n14714, new_n14715, new_n14716, new_n14717,
    new_n14718, new_n14719, new_n14720, new_n14721, new_n14722, new_n14723,
    new_n14724, new_n14725, new_n14727, new_n14730, new_n14731, new_n14732,
    new_n14733, new_n14734_1, new_n14735, new_n14736, new_n14737,
    new_n14738, new_n14739, new_n14740, new_n14741, new_n14742, new_n14743,
    new_n14744, new_n14745, new_n14746_1, new_n14747, new_n14748,
    new_n14749, new_n14750, new_n14751, new_n14752, new_n14753, new_n14754,
    new_n14755, new_n14756, new_n14757, new_n14758, new_n14759, new_n14760,
    new_n14761, new_n14762, new_n14763_1, new_n14764, new_n14765,
    new_n14766, new_n14767, new_n14768, new_n14769, new_n14770, new_n14771,
    new_n14772_1, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14778, new_n14779, new_n14780, new_n14781, new_n14782,
    new_n14783, new_n14784, new_n14785, new_n14786, new_n14787, new_n14788,
    new_n14789, new_n14790_1, new_n14791, new_n14792, new_n14793,
    new_n14794, new_n14795, new_n14796, new_n14797, new_n14798, new_n14799,
    new_n14800, new_n14801_1, new_n14802, new_n14803, new_n14804,
    new_n14805, new_n14806, new_n14807, new_n14808, new_n14809, new_n14810,
    new_n14811, new_n14812, new_n14813, new_n14816, new_n14817, new_n14818,
    new_n14819_1, new_n14820, new_n14821, new_n14822, new_n14823,
    new_n14824, new_n14825, new_n14826_1, new_n14827_1, new_n14828,
    new_n14829, new_n14830, new_n14831, new_n14832, new_n14833, new_n14834,
    new_n14835, new_n14836, new_n14837, new_n14838, new_n14839_1,
    new_n14840, new_n14841, new_n14842, new_n14843, new_n14844, new_n14845,
    new_n14846, new_n14847, new_n14848, new_n14849_1, new_n14850,
    new_n14851, new_n14852, new_n14853, new_n14854, new_n14855, new_n14856,
    new_n14857, new_n14858, new_n14859, new_n14860, new_n14861, new_n14862,
    new_n14863, new_n14864, new_n14865, new_n14866, new_n14867, new_n14868,
    new_n14869, new_n14870, new_n14871, new_n14872, new_n14873, new_n14874,
    new_n14875, new_n14876, new_n14877, new_n14878, new_n14879, new_n14880,
    new_n14881, new_n14882, new_n14883, new_n14884, new_n14885, new_n14886,
    new_n14887, new_n14888, new_n14889, new_n14890, new_n14891_1,
    new_n14892, new_n14893, new_n14894, new_n14895, new_n14896, new_n14897,
    new_n14898, new_n14899_1, new_n14900, new_n14901, new_n14902,
    new_n14903, new_n14904, new_n14905, new_n14906, new_n14907, new_n14908,
    new_n14909, new_n14910, new_n14911, new_n14912, new_n14913, new_n14914,
    new_n14915, new_n14916, new_n14917, new_n14918, new_n14919, new_n14920,
    new_n14921, new_n14922, new_n14923, new_n14924, new_n14925, new_n14926,
    new_n14927, new_n14928, new_n14929, new_n14930, new_n14931_1,
    new_n14932, new_n14933, new_n14934, new_n14935, new_n14936, new_n14937,
    new_n14938, new_n14939, new_n14940, new_n14941, new_n14942, new_n14943,
    new_n14944_1, new_n14945, new_n14946, new_n14947, new_n14948,
    new_n14949, new_n14950, new_n14951, new_n14952, new_n14953,
    new_n14954_1, new_n14955, new_n14956, new_n14957, new_n14958,
    new_n14959, new_n14960, new_n14961, new_n14962, new_n14963, new_n14964,
    new_n14965, new_n14966, new_n14967, new_n14968, new_n14969, new_n14970,
    new_n14971, new_n14972, new_n14973, new_n14974, new_n14975, new_n14976,
    new_n14977_1, new_n14978, new_n14979, new_n14980, new_n14981,
    new_n14982, new_n14983, new_n14984, new_n14985, new_n14986, new_n14987,
    new_n14988, new_n14989_1, new_n14990, new_n14991, new_n14992,
    new_n14993, new_n14994, new_n14995, new_n14996, new_n14997, new_n14998,
    new_n14999, new_n15000, new_n15001, new_n15002_1, new_n15003,
    new_n15004_1, new_n15005, new_n15006, new_n15007, new_n15008,
    new_n15009, new_n15010, new_n15011_1, new_n15012, new_n15013,
    new_n15014, new_n15015, new_n15016, new_n15017, new_n15018,
    new_n15019_1, new_n15020, new_n15021, new_n15022, new_n15023,
    new_n15024, new_n15025, new_n15026, new_n15027, new_n15028, new_n15029,
    new_n15030, new_n15031_1, new_n15032, new_n15033_1, new_n15034,
    new_n15035, new_n15036, new_n15037, new_n15038, new_n15039, new_n15040,
    new_n15041, new_n15042, new_n15043, new_n15044, new_n15045, new_n15046,
    new_n15047, new_n15048, new_n15049, new_n15050, new_n15051,
    new_n15052_1, new_n15053_1, new_n15054, new_n15055, new_n15056,
    new_n15057, new_n15058, new_n15059, new_n15060, new_n15061, new_n15062,
    new_n15063, new_n15064, new_n15065, new_n15066, new_n15067, new_n15068,
    new_n15069, new_n15070, new_n15071, new_n15072, new_n15073, new_n15074,
    new_n15075, new_n15076, new_n15077_1, new_n15078, new_n15079,
    new_n15080, new_n15081, new_n15082_1, new_n15083, new_n15084,
    new_n15085, new_n15086, new_n15087, new_n15088, new_n15089, new_n15090,
    new_n15091, new_n15092, new_n15093, new_n15094_1, new_n15095,
    new_n15097, new_n15099, new_n15100, new_n15101, new_n15102, new_n15103,
    new_n15104, new_n15105, new_n15106, new_n15107, new_n15108, new_n15109,
    new_n15110, new_n15111, new_n15112, new_n15113, new_n15114, new_n15115,
    new_n15116, new_n15117, new_n15118_1, new_n15119, new_n15120,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128_1, new_n15129, new_n15130, new_n15131,
    new_n15133, new_n15134, new_n15135, new_n15136, new_n15137, new_n15138,
    new_n15139_1, new_n15140, new_n15141, new_n15142, new_n15143,
    new_n15144, new_n15145_1, new_n15146_1, new_n15147, new_n15148,
    new_n15149, new_n15150, new_n15151, new_n15152, new_n15153, new_n15154,
    new_n15155, new_n15156, new_n15157, new_n15158, new_n15159, new_n15160,
    new_n15161, new_n15162, new_n15163, new_n15164, new_n15165_1,
    new_n15166, new_n15167_1, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175,
    new_n15176_1, new_n15177, new_n15178, new_n15179, new_n15180_1,
    new_n15181, new_n15182_1, new_n15183, new_n15184, new_n15185,
    new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191,
    new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197,
    new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203,
    new_n15204, new_n15205_1, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230_1, new_n15231,
    new_n15232, new_n15233, new_n15234, new_n15235, new_n15236, new_n15237,
    new_n15238, new_n15239, new_n15240, new_n15241_1, new_n15242,
    new_n15243, new_n15244, new_n15245, new_n15246, new_n15247, new_n15248,
    new_n15249, new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15255_1, new_n15256, new_n15257, new_n15258_1, new_n15259,
    new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265,
    new_n15266, new_n15267, new_n15268, new_n15269, new_n15270,
    new_n15271_1, new_n15272, new_n15273, new_n15274, new_n15275_1,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289_1, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300_1, new_n15301, new_n15302, new_n15303,
    new_n15304, new_n15305, new_n15306, new_n15307_1, new_n15308,
    new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314,
    new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320,
    new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326,
    new_n15327_1, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332_1, new_n15333, new_n15334, new_n15335, new_n15336,
    new_n15337, new_n15338, new_n15339, new_n15340, new_n15341, new_n15342,
    new_n15343, new_n15344, new_n15345_1, new_n15346, new_n15347,
    new_n15348, new_n15349, new_n15350, new_n15351, new_n15352,
    new_n15353_1, new_n15354, new_n15355, new_n15356, new_n15357,
    new_n15358, new_n15359, new_n15360, new_n15361, new_n15362, new_n15363,
    new_n15364, new_n15365, new_n15366_1, new_n15367, new_n15368,
    new_n15369, new_n15370, new_n15371, new_n15372, new_n15373, new_n15374,
    new_n15375, new_n15376, new_n15377, new_n15378_1, new_n15379,
    new_n15380, new_n15381, new_n15382_1, new_n15383, new_n15384,
    new_n15385, new_n15386, new_n15387, new_n15388, new_n15389, new_n15390,
    new_n15391, new_n15392, new_n15393, new_n15394, new_n15395, new_n15396,
    new_n15397, new_n15398, new_n15399, new_n15400, new_n15401, new_n15402,
    new_n15403, new_n15404, new_n15405, new_n15406, new_n15407_1,
    new_n15408, new_n15409, new_n15410, new_n15411, new_n15412, new_n15413,
    new_n15414, new_n15415, new_n15416, new_n15417, new_n15418, new_n15419,
    new_n15420, new_n15421, new_n15422, new_n15423, new_n15424_1,
    new_n15425, new_n15426, new_n15427, new_n15428_1, new_n15429,
    new_n15430, new_n15431, new_n15432, new_n15433, new_n15434,
    new_n15435_1, new_n15436, new_n15437, new_n15438_1, new_n15439,
    new_n15440, new_n15441, new_n15442, new_n15443, new_n15444, new_n15445,
    new_n15446, new_n15447, new_n15448, new_n15449, new_n15450, new_n15451,
    new_n15452, new_n15453, new_n15454, new_n15455, new_n15456, new_n15457,
    new_n15458, new_n15459, new_n15460, new_n15461, new_n15462, new_n15463,
    new_n15464, new_n15465_1, new_n15466, new_n15467_1, new_n15468,
    new_n15469, new_n15470_1, new_n15471, new_n15472, new_n15473,
    new_n15474, new_n15475, new_n15476, new_n15477_1, new_n15478,
    new_n15479, new_n15480, new_n15481_1, new_n15482, new_n15483,
    new_n15484, new_n15485, new_n15486, new_n15487, new_n15488, new_n15489,
    new_n15490_1, new_n15491, new_n15492, new_n15493, new_n15494,
    new_n15495, new_n15496_1, new_n15497, new_n15498, new_n15499,
    new_n15500, new_n15501_1, new_n15502, new_n15503, new_n15504,
    new_n15505, new_n15506_1, new_n15507, new_n15508_1, new_n15509,
    new_n15510, new_n15511, new_n15512, new_n15513, new_n15514, new_n15515,
    new_n15516, new_n15517, new_n15518, new_n15519, new_n15520, new_n15522,
    new_n15524, new_n15525, new_n15526, new_n15527, new_n15528, new_n15529,
    new_n15530, new_n15531, new_n15532, new_n15533, new_n15534, new_n15535,
    new_n15536, new_n15537, new_n15538, new_n15539_1, new_n15540,
    new_n15541, new_n15542, new_n15543, new_n15544, new_n15545,
    new_n15546_1, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555_1,
    new_n15556, new_n15557, new_n15558_1, new_n15559_1, new_n15560,
    new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566,
    new_n15567, new_n15568, new_n15569, new_n15570_1, new_n15571,
    new_n15572, new_n15573_1, new_n15574, new_n15575, new_n15576,
    new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582,
    new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588_1, new_n15589, new_n15590_1, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597,
    new_n15598_1, new_n15599, new_n15600, new_n15601, new_n15602_1,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613,
    new_n15614_1, new_n15616, new_n15619, new_n15621, new_n15622,
    new_n15623, new_n15624, new_n15625, new_n15626, new_n15627, new_n15628,
    new_n15629, new_n15630, new_n15631, new_n15632, new_n15633, new_n15634,
    new_n15635, new_n15636_1, new_n15637, new_n15638, new_n15639,
    new_n15640, new_n15642, new_n15644, new_n15646, new_n15647, new_n15648,
    new_n15649, new_n15650, new_n15651, new_n15652_1, new_n15653,
    new_n15654, new_n15655, new_n15656, new_n15657, new_n15658, new_n15659,
    new_n15660, new_n15661, new_n15662_1, new_n15663, new_n15664,
    new_n15665, new_n15666, new_n15667, new_n15668, new_n15669, new_n15670,
    new_n15671, new_n15672, new_n15673, new_n15674, new_n15675, new_n15676,
    new_n15677, new_n15678, new_n15679, new_n15680, new_n15681, new_n15684,
    new_n15686, new_n15687, new_n15688, new_n15689, new_n15690, new_n15691,
    new_n15692, new_n15693, new_n15694, new_n15695, new_n15696, new_n15697,
    new_n15698, new_n15699, new_n15700, new_n15701, new_n15702, new_n15703,
    new_n15704, new_n15705, new_n15706, new_n15707, new_n15708, new_n15709,
    new_n15710, new_n15711, new_n15712, new_n15713, new_n15714, new_n15715,
    new_n15716_1, new_n15717, new_n15718, new_n15719, new_n15720,
    new_n15721, new_n15722, new_n15724, new_n15725, new_n15726, new_n15727,
    new_n15728, new_n15729, new_n15730, new_n15731, new_n15732, new_n15733,
    new_n15734, new_n15735, new_n15736, new_n15737, new_n15738, new_n15739,
    new_n15740, new_n15741, new_n15742, new_n15743_1, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749_1,
    new_n15750, new_n15751, new_n15752, new_n15753, new_n15754, new_n15755,
    new_n15756, new_n15757, new_n15758, new_n15759, new_n15760,
    new_n15761_1, new_n15762_1, new_n15763, new_n15764, new_n15766_1,
    new_n15768, new_n15770, new_n15771, new_n15772, new_n15773, new_n15774,
    new_n15775, new_n15776, new_n15777, new_n15778, new_n15779,
    new_n15780_1, new_n15781, new_n15782, new_n15783, new_n15784,
    new_n15785, new_n15786, new_n15787, new_n15788, new_n15789, new_n15790,
    new_n15791, new_n15792, new_n15793_1, new_n15794, new_n15795,
    new_n15796, new_n15797, new_n15798, new_n15799, new_n15800, new_n15801,
    new_n15802, new_n15803, new_n15804, new_n15805, new_n15806, new_n15807,
    new_n15808, new_n15809, new_n15810, new_n15811, new_n15812_1,
    new_n15813, new_n15814, new_n15815_1, new_n15816_1, new_n15817,
    new_n15818, new_n15819, new_n15820, new_n15821, new_n15822, new_n15823,
    new_n15824, new_n15825, new_n15826, new_n15827, new_n15828, new_n15829,
    new_n15830, new_n15831_1, new_n15832, new_n15833, new_n15834,
    new_n15835, new_n15836, new_n15837, new_n15838, new_n15839, new_n15840,
    new_n15841, new_n15842, new_n15843, new_n15844, new_n15845,
    new_n15846_1, new_n15847, new_n15850, new_n15851, new_n15852,
    new_n15853, new_n15854, new_n15855, new_n15856, new_n15857, new_n15858,
    new_n15859_1, new_n15860, new_n15861, new_n15862, new_n15863,
    new_n15864, new_n15865, new_n15866, new_n15867, new_n15868,
    new_n15869_1, new_n15870, new_n15871, new_n15872, new_n15873,
    new_n15874, new_n15875, new_n15876, new_n15877, new_n15878, new_n15879,
    new_n15880, new_n15881, new_n15882, new_n15883, new_n15884_1,
    new_n15885_1, new_n15886, new_n15887, new_n15888, new_n15889_1,
    new_n15890, new_n15891, new_n15892, new_n15893, new_n15894, new_n15895,
    new_n15896, new_n15897, new_n15898, new_n15899, new_n15900, new_n15901,
    new_n15902, new_n15903, new_n15904, new_n15905, new_n15906, new_n15907,
    new_n15908, new_n15909, new_n15910, new_n15911, new_n15912, new_n15913,
    new_n15914, new_n15915, new_n15916, new_n15917_1, new_n15918_1,
    new_n15919, new_n15920, new_n15921, new_n15922_1, new_n15923,
    new_n15924, new_n15925, new_n15926, new_n15927, new_n15928, new_n15929,
    new_n15930, new_n15931, new_n15932, new_n15933, new_n15934, new_n15935,
    new_n15936_1, new_n15937, new_n15938, new_n15939, new_n15940,
    new_n15941, new_n15942, new_n15943, new_n15944, new_n15945, new_n15946,
    new_n15947_1, new_n15948, new_n15949, new_n15950, new_n15951,
    new_n15952, new_n15953, new_n15954, new_n15955, new_n15956_1,
    new_n15957, new_n15958_1, new_n15959, new_n15960, new_n15961,
    new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967_1, new_n15968, new_n15969, new_n15970, new_n15971,
    new_n15972, new_n15973, new_n15974, new_n15975, new_n15976, new_n15977,
    new_n15978, new_n15979_1, new_n15980, new_n15981, new_n15982,
    new_n15983, new_n15984, new_n15985, new_n15986_1, new_n15988,
    new_n15989, new_n15990, new_n15991, new_n15992, new_n15993, new_n15994,
    new_n15995, new_n15996, new_n15997, new_n15998, new_n15999, new_n16000,
    new_n16001, new_n16002, new_n16003, new_n16004, new_n16005, new_n16006,
    new_n16007, new_n16008, new_n16009, new_n16010, new_n16011, new_n16012,
    new_n16013_1, new_n16014, new_n16015, new_n16016, new_n16017,
    new_n16018, new_n16019, new_n16020, new_n16021, new_n16022, new_n16023,
    new_n16024, new_n16025, new_n16026, new_n16027, new_n16028,
    new_n16029_1, new_n16030, new_n16031, new_n16032, new_n16033,
    new_n16034, new_n16035, new_n16036, new_n16037, new_n16038, new_n16039,
    new_n16040, new_n16041, new_n16042, new_n16043, new_n16044, new_n16045,
    new_n16046, new_n16047, new_n16048, new_n16049, new_n16050, new_n16051,
    new_n16052, new_n16053, new_n16054, new_n16055, new_n16056, new_n16057,
    new_n16058, new_n16059, new_n16060_1, new_n16061, new_n16062_1,
    new_n16063, new_n16064, new_n16065, new_n16066, new_n16067,
    new_n16068_1, new_n16069, new_n16070, new_n16071, new_n16072,
    new_n16073, new_n16074, new_n16075, new_n16076, new_n16077, new_n16078,
    new_n16079, new_n16080_1, new_n16081, new_n16082, new_n16083,
    new_n16084, new_n16085, new_n16086, new_n16087, new_n16088, new_n16089,
    new_n16090, new_n16091, new_n16092, new_n16093, new_n16094, new_n16095,
    new_n16096, new_n16097, new_n16098_1, new_n16099, new_n16100,
    new_n16101, new_n16102, new_n16103, new_n16104, new_n16105, new_n16106,
    new_n16107, new_n16108, new_n16109, new_n16110_1, new_n16111,
    new_n16112, new_n16113, new_n16114, new_n16115, new_n16116, new_n16117,
    new_n16118, new_n16119, new_n16120, new_n16121, new_n16122, new_n16123,
    new_n16124, new_n16125, new_n16126, new_n16127, new_n16128, new_n16129,
    new_n16130, new_n16131, new_n16132, new_n16133, new_n16134, new_n16135,
    new_n16136, new_n16138, new_n16139, new_n16140, new_n16141,
    new_n16142_1, new_n16143, new_n16144, new_n16145, new_n16146,
    new_n16147, new_n16148, new_n16149, new_n16150, new_n16151, new_n16152,
    new_n16153, new_n16154, new_n16155, new_n16156, new_n16157,
    new_n16158_1, new_n16159, new_n16160, new_n16161, new_n16162,
    new_n16163, new_n16164, new_n16165, new_n16166, new_n16167_1,
    new_n16168, new_n16169, new_n16170, new_n16171, new_n16172, new_n16173,
    new_n16174, new_n16175, new_n16176, new_n16177, new_n16178, new_n16179,
    new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185_1, new_n16186, new_n16187, new_n16188, new_n16189,
    new_n16190, new_n16191, new_n16192, new_n16193, new_n16194, new_n16195,
    new_n16196_1, new_n16197, new_n16198, new_n16199, new_n16200,
    new_n16201, new_n16202, new_n16203, new_n16204, new_n16205,
    new_n16206_1, new_n16207, new_n16208, new_n16210, new_n16212,
    new_n16213, new_n16214, new_n16215_1, new_n16216, new_n16217_1,
    new_n16218_1, new_n16219_1, new_n16220, new_n16221, new_n16222,
    new_n16223_1, new_n16224, new_n16225, new_n16226, new_n16227,
    new_n16228, new_n16230_1, new_n16231, new_n16232, new_n16233,
    new_n16234, new_n16235, new_n16236, new_n16237, new_n16238, new_n16239,
    new_n16240, new_n16241, new_n16242, new_n16243_1, new_n16244,
    new_n16245, new_n16246, new_n16247_1, new_n16248, new_n16249,
    new_n16250, new_n16251, new_n16252, new_n16253, new_n16254, new_n16255,
    new_n16256, new_n16257, new_n16258, new_n16259, new_n16260, new_n16261,
    new_n16262, new_n16263, new_n16264, new_n16265, new_n16266, new_n16267,
    new_n16268, new_n16269, new_n16270, new_n16271, new_n16272, new_n16273,
    new_n16274, new_n16275_1, new_n16276, new_n16277, new_n16278,
    new_n16279_1, new_n16280, new_n16281, new_n16282, new_n16283,
    new_n16284, new_n16285, new_n16286, new_n16287, new_n16288, new_n16289,
    new_n16290, new_n16291, new_n16292, new_n16293, new_n16294, new_n16295,
    new_n16296, new_n16297, new_n16298, new_n16299, new_n16300, new_n16301,
    new_n16302, new_n16303, new_n16304, new_n16305, new_n16306, new_n16307,
    new_n16308, new_n16309, new_n16310, new_n16311, new_n16312, new_n16313,
    new_n16314, new_n16315, new_n16316, new_n16317, new_n16318, new_n16319,
    new_n16320, new_n16321, new_n16322_1, new_n16323, new_n16324,
    new_n16325, new_n16326, new_n16327_1, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350_1, new_n16351, new_n16352,
    new_n16353, new_n16354, new_n16355, new_n16356, new_n16357, new_n16358,
    new_n16359, new_n16360, new_n16361, new_n16362, new_n16363, new_n16364,
    new_n16365, new_n16366, new_n16367_1, new_n16368, new_n16369,
    new_n16370, new_n16371, new_n16372, new_n16373, new_n16374, new_n16375,
    new_n16376_1, new_n16377, new_n16378, new_n16379_1, new_n16380,
    new_n16381, new_n16382, new_n16383, new_n16384, new_n16385, new_n16386,
    new_n16387, new_n16388, new_n16389, new_n16390, new_n16391, new_n16392,
    new_n16393, new_n16394, new_n16395, new_n16396_1, new_n16397,
    new_n16398_1, new_n16399, new_n16400, new_n16401, new_n16402,
    new_n16403, new_n16404, new_n16405, new_n16406_1, new_n16407_1,
    new_n16408, new_n16409, new_n16410, new_n16411, new_n16412, new_n16413,
    new_n16414, new_n16415, new_n16416, new_n16417, new_n16418,
    new_n16419_1, new_n16420, new_n16421, new_n16422, new_n16423,
    new_n16424_1, new_n16425, new_n16426, new_n16429, new_n16430,
    new_n16431, new_n16432, new_n16433_1, new_n16434, new_n16435,
    new_n16436, new_n16437, new_n16438, new_n16439_1, new_n16440_1,
    new_n16441, new_n16442, new_n16443, new_n16444, new_n16445_1,
    new_n16446, new_n16447, new_n16448, new_n16449, new_n16450, new_n16451,
    new_n16452, new_n16453, new_n16454, new_n16455, new_n16456, new_n16457,
    new_n16458, new_n16459, new_n16460_1, new_n16461, new_n16462,
    new_n16463, new_n16464, new_n16465, new_n16466, new_n16467, new_n16468,
    new_n16469, new_n16470, new_n16471, new_n16472, new_n16473, new_n16474,
    new_n16475, new_n16476_1, new_n16477, new_n16478, new_n16479,
    new_n16480, new_n16481_1, new_n16482_1, new_n16483, new_n16484,
    new_n16485, new_n16486, new_n16487, new_n16488, new_n16489, new_n16490,
    new_n16491, new_n16492, new_n16493_1, new_n16494, new_n16495,
    new_n16496, new_n16497, new_n16498, new_n16499, new_n16500, new_n16501,
    new_n16502_1, new_n16503, new_n16504, new_n16505, new_n16506_1,
    new_n16507_1, new_n16508, new_n16509, new_n16510, new_n16511,
    new_n16512, new_n16513, new_n16514, new_n16515, new_n16516_1,
    new_n16517_1, new_n16518, new_n16519, new_n16520, new_n16521_1,
    new_n16522, new_n16523, new_n16524_1, new_n16525, new_n16526,
    new_n16527_1, new_n16528, new_n16529, new_n16530, new_n16531,
    new_n16533, new_n16534, new_n16535, new_n16536, new_n16537, new_n16538,
    new_n16539, new_n16540, new_n16543, new_n16544_1, new_n16545,
    new_n16546, new_n16547, new_n16548, new_n16549, new_n16550, new_n16551,
    new_n16552, new_n16553, new_n16554_1, new_n16555, new_n16556,
    new_n16557, new_n16558, new_n16559, new_n16560, new_n16561, new_n16562,
    new_n16563, new_n16564, new_n16565, new_n16566, new_n16567, new_n16568,
    new_n16569, new_n16570, new_n16571, new_n16572, new_n16573, new_n16574,
    new_n16575, new_n16576, new_n16577, new_n16578, new_n16579, new_n16580,
    new_n16581, new_n16582, new_n16583_1, new_n16584_1, new_n16585,
    new_n16586, new_n16587, new_n16588, new_n16589_1, new_n16590,
    new_n16591, new_n16592, new_n16593, new_n16594, new_n16595,
    new_n16596_1, new_n16597, new_n16598, new_n16599, new_n16600,
    new_n16601, new_n16602, new_n16603, new_n16604, new_n16605, new_n16606,
    new_n16607, new_n16608_1, new_n16609, new_n16610, new_n16611,
    new_n16612, new_n16613, new_n16614, new_n16615, new_n16616,
    new_n16617_1, new_n16618, new_n16619, new_n16620, new_n16621,
    new_n16622, new_n16623, new_n16624, new_n16625, new_n16626, new_n16627,
    new_n16628, new_n16629, new_n16630_1, new_n16631, new_n16632,
    new_n16633, new_n16634, new_n16635, new_n16636, new_n16637, new_n16638,
    new_n16639, new_n16640_1, new_n16641, new_n16642, new_n16643,
    new_n16644, new_n16645, new_n16646, new_n16647, new_n16648, new_n16649,
    new_n16650, new_n16651, new_n16652, new_n16653, new_n16654, new_n16655,
    new_n16657, new_n16658, new_n16659, new_n16660, new_n16661, new_n16662,
    new_n16663, new_n16664, new_n16665, new_n16666, new_n16667, new_n16668,
    new_n16669, new_n16670, new_n16671, new_n16672, new_n16673,
    new_n16674_1, new_n16675, new_n16676, new_n16677, new_n16678,
    new_n16679, new_n16680, new_n16681, new_n16682_1, new_n16683,
    new_n16684_1, new_n16685, new_n16686, new_n16687, new_n16688_1,
    new_n16689, new_n16690, new_n16691, new_n16692, new_n16693, new_n16694,
    new_n16695, new_n16696, new_n16697, new_n16698, new_n16699, new_n16700,
    new_n16701, new_n16702, new_n16703, new_n16704, new_n16705, new_n16706,
    new_n16707, new_n16708, new_n16709, new_n16710, new_n16711, new_n16712,
    new_n16713, new_n16714, new_n16715, new_n16716, new_n16717, new_n16718,
    new_n16719, new_n16720, new_n16721, new_n16722_1, new_n16723,
    new_n16724, new_n16725, new_n16726, new_n16727, new_n16728, new_n16729,
    new_n16730, new_n16731, new_n16732, new_n16733_1, new_n16734,
    new_n16735, new_n16736, new_n16737, new_n16738, new_n16739, new_n16740,
    new_n16741, new_n16742, new_n16743_1, new_n16744, new_n16745,
    new_n16746, new_n16747, new_n16748, new_n16749, new_n16750, new_n16751,
    new_n16752, new_n16753, new_n16754, new_n16755, new_n16756, new_n16757,
    new_n16758, new_n16759, new_n16760, new_n16761, new_n16762, new_n16763,
    new_n16764, new_n16765, new_n16766, new_n16767, new_n16768, new_n16769,
    new_n16770, new_n16771, new_n16772, new_n16773, new_n16774, new_n16775,
    new_n16776, new_n16777, new_n16778, new_n16779, new_n16780, new_n16781,
    new_n16782, new_n16783, new_n16784, new_n16785, new_n16786, new_n16787,
    new_n16788, new_n16789, new_n16790, new_n16791, new_n16792, new_n16793,
    new_n16794, new_n16795, new_n16796, new_n16797, new_n16798_1,
    new_n16799, new_n16800, new_n16801, new_n16802, new_n16803, new_n16804,
    new_n16805, new_n16806, new_n16807, new_n16808, new_n16809, new_n16810,
    new_n16811, new_n16812_1, new_n16813, new_n16814, new_n16815,
    new_n16816, new_n16817, new_n16818_1, new_n16820, new_n16822,
    new_n16823, new_n16824_1, new_n16825, new_n16826, new_n16827,
    new_n16828, new_n16829, new_n16830, new_n16831, new_n16832, new_n16833,
    new_n16834_1, new_n16835, new_n16836, new_n16837_1, new_n16838,
    new_n16839, new_n16840, new_n16841_1, new_n16842, new_n16843,
    new_n16844, new_n16845, new_n16846, new_n16847, new_n16848, new_n16849,
    new_n16850, new_n16851, new_n16852, new_n16853, new_n16854, new_n16855,
    new_n16856, new_n16857, new_n16858, new_n16859, new_n16860, new_n16861,
    new_n16862, new_n16863, new_n16864, new_n16865, new_n16866, new_n16867,
    new_n16868, new_n16869, new_n16870, new_n16871, new_n16872, new_n16873,
    new_n16874, new_n16875, new_n16876, new_n16877, new_n16879, new_n16881,
    new_n16882, new_n16883, new_n16884, new_n16885_1, new_n16886,
    new_n16887, new_n16888, new_n16889, new_n16890, new_n16891, new_n16892,
    new_n16893, new_n16894, new_n16895, new_n16896, new_n16897, new_n16898,
    new_n16899, new_n16900, new_n16901, new_n16902, new_n16903, new_n16904,
    new_n16905_1, new_n16906, new_n16907, new_n16908, new_n16909,
    new_n16910, new_n16911_1, new_n16912, new_n16913, new_n16914,
    new_n16915, new_n16916, new_n16917, new_n16918, new_n16919, new_n16920,
    new_n16921, new_n16922, new_n16923, new_n16924, new_n16925, new_n16926,
    new_n16927, new_n16928, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951_1, new_n16952, new_n16953, new_n16954_1, new_n16955,
    new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961,
    new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967,
    new_n16968_1, new_n16969, new_n16970, new_n16971_1, new_n16972,
    new_n16973, new_n16974, new_n16975, new_n16976, new_n16977, new_n16978,
    new_n16979, new_n16980, new_n16981, new_n16982, new_n16983, new_n16984,
    new_n16985, new_n16986, new_n16987, new_n16988_1, new_n16989_1,
    new_n16990, new_n16991, new_n16992, new_n16993, new_n16994_1,
    new_n16995, new_n16996, new_n16997, new_n16998, new_n16999, new_n17000,
    new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006_1, new_n17007, new_n17008, new_n17009, new_n17010,
    new_n17011, new_n17012, new_n17013, new_n17014, new_n17015, new_n17016,
    new_n17017, new_n17018, new_n17019, new_n17020, new_n17021, new_n17022,
    new_n17023, new_n17024, new_n17025, new_n17026, new_n17027, new_n17028,
    new_n17029, new_n17030, new_n17031, new_n17032, new_n17033, new_n17034,
    new_n17035_1, new_n17036, new_n17037_1, new_n17038, new_n17039,
    new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17046,
    new_n17047, new_n17048, new_n17049, new_n17050, new_n17051, new_n17052,
    new_n17053, new_n17054, new_n17055, new_n17056, new_n17057, new_n17058,
    new_n17059, new_n17060, new_n17061, new_n17062, new_n17063, new_n17064,
    new_n17065, new_n17066, new_n17067, new_n17068_1, new_n17069_1,
    new_n17070_1, new_n17071, new_n17072, new_n17073, new_n17074,
    new_n17075_1, new_n17076, new_n17077_1, new_n17078, new_n17079,
    new_n17080, new_n17081, new_n17082, new_n17083, new_n17084_1,
    new_n17085, new_n17086, new_n17088, new_n17089, new_n17090_1,
    new_n17091, new_n17092, new_n17093, new_n17094, new_n17095_1,
    new_n17096, new_n17097, new_n17098, new_n17099, new_n17100, new_n17101,
    new_n17102, new_n17103, new_n17104_1, new_n17105, new_n17106_1,
    new_n17107, new_n17108, new_n17109, new_n17110, new_n17111, new_n17112,
    new_n17113, new_n17114, new_n17115, new_n17116, new_n17117, new_n17118,
    new_n17119_1, new_n17120, new_n17121, new_n17122, new_n17123,
    new_n17124, new_n17125, new_n17126, new_n17127, new_n17128, new_n17129,
    new_n17130_1, new_n17131, new_n17132, new_n17133, new_n17134,
    new_n17135, new_n17136, new_n17137, new_n17138_1, new_n17139,
    new_n17140, new_n17141, new_n17142, new_n17143, new_n17144, new_n17145,
    new_n17146, new_n17147, new_n17148, new_n17149, new_n17150, new_n17151,
    new_n17152, new_n17153, new_n17154, new_n17155, new_n17156, new_n17157,
    new_n17158, new_n17159, new_n17160, new_n17161, new_n17162,
    new_n17163_1, new_n17164, new_n17165, new_n17166, new_n17167,
    new_n17168_1, new_n17169, new_n17170, new_n17171, new_n17172,
    new_n17173, new_n17174, new_n17175, new_n17176, new_n17177, new_n17178,
    new_n17179, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184,
    new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190,
    new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196,
    new_n17197, new_n17198, new_n17199, new_n17200, new_n17201,
    new_n17202_1, new_n17203, new_n17204, new_n17205, new_n17206,
    new_n17207, new_n17208, new_n17209, new_n17210, new_n17211, new_n17212,
    new_n17213, new_n17214, new_n17215, new_n17216, new_n17217, new_n17218,
    new_n17219_1, new_n17220, new_n17221, new_n17222, new_n17223,
    new_n17224, new_n17225, new_n17226, new_n17227, new_n17228, new_n17229,
    new_n17230, new_n17231, new_n17232_1, new_n17233, new_n17234,
    new_n17235, new_n17236_1, new_n17237, new_n17238, new_n17239,
    new_n17240, new_n17241, new_n17242, new_n17243_1, new_n17244,
    new_n17245, new_n17246, new_n17247, new_n17248, new_n17249,
    new_n17250_1, new_n17251_1, new_n17252, new_n17253, new_n17254,
    new_n17255, new_n17256, new_n17257, new_n17258, new_n17259, new_n17260,
    new_n17261, new_n17262, new_n17263_1, new_n17264, new_n17265,
    new_n17266, new_n17267, new_n17268, new_n17269, new_n17270, new_n17271,
    new_n17272, new_n17273, new_n17274, new_n17275, new_n17276, new_n17277,
    new_n17278, new_n17279, new_n17280, new_n17281, new_n17282, new_n17283,
    new_n17284, new_n17285_1, new_n17286, new_n17287, new_n17288,
    new_n17289, new_n17290, new_n17291, new_n17292, new_n17293, new_n17294,
    new_n17295, new_n17296, new_n17297, new_n17298, new_n17299, new_n17300,
    new_n17301, new_n17302_1, new_n17303, new_n17304, new_n17305,
    new_n17306, new_n17307, new_n17308, new_n17309, new_n17310, new_n17311,
    new_n17312, new_n17313, new_n17314, new_n17315, new_n17316, new_n17317,
    new_n17318, new_n17319, new_n17320_1, new_n17321, new_n17322,
    new_n17323, new_n17324, new_n17325, new_n17326, new_n17327, new_n17328,
    new_n17329, new_n17330, new_n17331, new_n17332, new_n17333, new_n17334,
    new_n17335, new_n17336, new_n17338, new_n17339, new_n17340, new_n17341,
    new_n17342, new_n17343, new_n17344_1, new_n17345, new_n17346,
    new_n17347, new_n17348, new_n17349, new_n17350, new_n17351_1,
    new_n17352, new_n17353, new_n17354, new_n17355, new_n17356, new_n17357,
    new_n17358, new_n17359_1, new_n17360, new_n17361, new_n17362,
    new_n17363, new_n17364, new_n17365, new_n17366, new_n17367, new_n17368,
    new_n17369, new_n17370, new_n17371, new_n17372, new_n17373, new_n17374,
    new_n17375, new_n17376, new_n17377, new_n17378, new_n17379, new_n17380,
    new_n17381, new_n17382, new_n17383, new_n17384, new_n17385, new_n17386,
    new_n17387_1, new_n17388, new_n17389, new_n17390, new_n17391_1,
    new_n17392_1, new_n17393, new_n17394, new_n17395, new_n17396,
    new_n17397, new_n17398, new_n17399, new_n17400, new_n17401, new_n17402,
    new_n17403, new_n17404, new_n17405, new_n17406, new_n17407, new_n17408,
    new_n17409, new_n17410, new_n17411, new_n17412, new_n17413, new_n17414,
    new_n17415, new_n17416, new_n17417, new_n17418, new_n17419, new_n17420,
    new_n17421_1, new_n17422, new_n17423, new_n17424, new_n17425,
    new_n17426, new_n17427, new_n17428, new_n17429, new_n17430, new_n17431,
    new_n17432_1, new_n17433, new_n17434, new_n17435, new_n17436_1,
    new_n17437, new_n17438, new_n17439, new_n17440_1, new_n17441,
    new_n17442, new_n17443, new_n17444, new_n17445, new_n17446, new_n17447,
    new_n17448, new_n17449, new_n17450_1, new_n17451, new_n17452,
    new_n17453, new_n17454, new_n17455, new_n17456, new_n17457,
    new_n17458_1, new_n17459, new_n17460, new_n17461_1, new_n17462,
    new_n17463, new_n17464, new_n17465, new_n17466_1, new_n17467,
    new_n17468, new_n17469, new_n17470, new_n17471, new_n17472, new_n17473,
    new_n17474, new_n17475, new_n17476, new_n17477, new_n17478, new_n17479,
    new_n17480, new_n17481, new_n17482, new_n17483, new_n17484, new_n17485,
    new_n17486, new_n17487, new_n17488, new_n17489, new_n17490, new_n17491,
    new_n17492, new_n17493_1, new_n17494, new_n17495, new_n17496,
    new_n17497, new_n17498, new_n17499, new_n17500_1, new_n17501,
    new_n17502, new_n17503, new_n17504, new_n17505, new_n17506, new_n17507,
    new_n17508, new_n17509, new_n17510, new_n17511, new_n17512, new_n17513,
    new_n17514, new_n17515, new_n17516, new_n17517, new_n17518, new_n17519,
    new_n17520, new_n17521, new_n17522, new_n17523, new_n17524_1,
    new_n17525, new_n17526, new_n17527, new_n17528, new_n17529_1,
    new_n17530, new_n17531, new_n17532, new_n17533, new_n17534, new_n17535,
    new_n17536, new_n17537, new_n17538, new_n17539, new_n17540, new_n17541,
    new_n17542, new_n17543, new_n17544, new_n17545, new_n17546, new_n17547,
    new_n17548, new_n17549, new_n17550, new_n17551, new_n17552, new_n17553,
    new_n17554, new_n17555, new_n17556, new_n17557_1, new_n17558,
    new_n17559, new_n17560, new_n17561, new_n17562, new_n17563, new_n17565,
    new_n17566, new_n17567, new_n17568, new_n17569, new_n17570, new_n17571,
    new_n17572, new_n17573, new_n17574, new_n17575, new_n17576, new_n17577,
    new_n17578, new_n17579, new_n17580, new_n17581, new_n17582,
    new_n17583_1, new_n17584, new_n17585, new_n17586, new_n17587,
    new_n17588, new_n17589, new_n17590, new_n17591, new_n17592_1,
    new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17598,
    new_n17599, new_n17600, new_n17601, new_n17602, new_n17603, new_n17604,
    new_n17605, new_n17606, new_n17607, new_n17608, new_n17609, new_n17610,
    new_n17611, new_n17612, new_n17613, new_n17614, new_n17615, new_n17616,
    new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17622,
    new_n17623, new_n17624, new_n17625, new_n17626, new_n17627, new_n17628,
    new_n17629, new_n17630, new_n17631, new_n17632, new_n17633, new_n17634,
    new_n17635, new_n17636, new_n17637, new_n17638_1, new_n17639,
    new_n17640, new_n17641, new_n17642, new_n17643, new_n17644, new_n17645,
    new_n17646, new_n17647, new_n17648, new_n17649, new_n17650, new_n17651,
    new_n17652, new_n17653, new_n17654, new_n17655, new_n17656, new_n17657,
    new_n17658, new_n17659, new_n17660, new_n17661, new_n17662, new_n17663,
    new_n17664_1, new_n17665, new_n17666, new_n17667, new_n17668,
    new_n17669, new_n17670, new_n17671, new_n17672, new_n17673, new_n17674,
    new_n17675, new_n17676, new_n17677, new_n17678, new_n17679, new_n17680,
    new_n17681, new_n17682, new_n17683, new_n17684, new_n17685, new_n17686,
    new_n17687_1, new_n17688, new_n17689, new_n17690, new_n17691,
    new_n17692, new_n17693, new_n17694, new_n17695, new_n17696, new_n17697,
    new_n17698, new_n17699, new_n17700, new_n17701, new_n17702, new_n17703,
    new_n17704, new_n17705, new_n17706, new_n17707, new_n17708, new_n17709,
    new_n17710, new_n17711, new_n17712, new_n17713, new_n17714, new_n17715,
    new_n17716, new_n17717, new_n17718, new_n17719, new_n17720,
    new_n17721_1, new_n17722, new_n17723, new_n17724, new_n17725,
    new_n17726, new_n17727, new_n17728, new_n17729, new_n17730, new_n17731,
    new_n17732, new_n17733, new_n17734, new_n17735_1, new_n17736,
    new_n17737, new_n17738_1, new_n17739, new_n17740, new_n17741,
    new_n17742, new_n17743, new_n17744, new_n17745, new_n17746_1,
    new_n17747, new_n17748, new_n17749_1, new_n17750, new_n17751,
    new_n17752, new_n17753, new_n17754, new_n17755, new_n17756, new_n17757,
    new_n17759, new_n17760, new_n17761, new_n17762, new_n17763, new_n17764,
    new_n17765, new_n17766, new_n17767, new_n17768, new_n17769, new_n17770,
    new_n17771, new_n17772, new_n17773, new_n17774, new_n17775, new_n17776,
    new_n17777, new_n17778, new_n17779, new_n17780, new_n17781, new_n17782,
    new_n17783, new_n17784_1, new_n17785, new_n17786, new_n17787,
    new_n17788, new_n17789, new_n17790, new_n17791, new_n17792, new_n17793,
    new_n17794, new_n17795, new_n17796, new_n17797, new_n17798, new_n17799,
    new_n17800, new_n17801, new_n17802, new_n17803, new_n17804, new_n17805,
    new_n17806, new_n17807, new_n17808, new_n17809, new_n17810, new_n17811,
    new_n17812, new_n17813, new_n17814, new_n17815, new_n17816, new_n17817,
    new_n17818, new_n17819, new_n17820_1, new_n17821, new_n17822,
    new_n17823, new_n17824, new_n17825, new_n17826, new_n17827, new_n17828,
    new_n17829, new_n17830, new_n17831, new_n17832, new_n17833, new_n17834,
    new_n17835, new_n17836, new_n17837, new_n17838, new_n17839, new_n17840,
    new_n17841, new_n17842, new_n17843, new_n17844, new_n17845, new_n17846,
    new_n17847, new_n17848, new_n17849, new_n17850, new_n17851, new_n17852,
    new_n17853, new_n17854, new_n17855_1, new_n17856, new_n17857,
    new_n17858, new_n17859, new_n17860, new_n17861, new_n17862, new_n17863,
    new_n17864, new_n17865, new_n17866, new_n17867, new_n17868, new_n17869,
    new_n17870, new_n17871, new_n17872, new_n17873, new_n17874, new_n17875,
    new_n17876, new_n17877_1, new_n17878, new_n17879, new_n17880,
    new_n17881, new_n17882, new_n17883, new_n17884, new_n17885, new_n17886,
    new_n17887, new_n17889_1, new_n17890, new_n17891, new_n17892,
    new_n17893, new_n17894, new_n17895, new_n17896, new_n17897, new_n17898,
    new_n17899, new_n17900, new_n17901, new_n17902, new_n17903, new_n17904,
    new_n17905, new_n17906, new_n17907, new_n17908, new_n17909, new_n17910,
    new_n17911_1, new_n17912_1, new_n17913, new_n17914, new_n17915,
    new_n17916, new_n17917, new_n17918, new_n17919, new_n17920, new_n17921,
    new_n17922, new_n17923, new_n17924, new_n17925, new_n17926,
    new_n17927_1, new_n17928, new_n17929, new_n17930, new_n17931_1,
    new_n17932, new_n17933, new_n17934, new_n17935, new_n17936, new_n17937,
    new_n17938, new_n17939, new_n17940, new_n17941, new_n17942, new_n17943,
    new_n17944, new_n17945, new_n17946, new_n17947, new_n17948_1,
    new_n17949, new_n17950, new_n17951, new_n17952, new_n17953,
    new_n17954_1, new_n17955, new_n17956_1, new_n17957, new_n17958,
    new_n17959_1, new_n17960, new_n17961, new_n17963_1, new_n17965,
    new_n17966, new_n17967, new_n17968_1, new_n17969, new_n17970,
    new_n17971, new_n17972, new_n17973, new_n17974, new_n17975,
    new_n17976_1, new_n17977, new_n17978, new_n17979, new_n17980,
    new_n17981, new_n17982, new_n17983, new_n17984, new_n17985, new_n17986,
    new_n17987, new_n17988, new_n17989, new_n17990, new_n17991, new_n17992,
    new_n17993, new_n17994, new_n17995, new_n17996, new_n17997,
    new_n17998_1, new_n17999, new_n18000, new_n18001, new_n18002,
    new_n18003, new_n18004, new_n18005, new_n18006, new_n18007, new_n18008,
    new_n18009, new_n18010, new_n18011, new_n18012, new_n18013, new_n18014,
    new_n18015, new_n18016, new_n18017, new_n18018, new_n18019, new_n18020,
    new_n18021, new_n18022, new_n18023, new_n18024, new_n18025_1,
    new_n18026, new_n18027, new_n18028, new_n18029, new_n18030, new_n18031,
    new_n18032, new_n18033, new_n18034, new_n18035_1, new_n18036,
    new_n18037, new_n18038, new_n18039, new_n18040, new_n18041, new_n18042,
    new_n18043_1, new_n18044, new_n18045_1, new_n18046, new_n18047,
    new_n18048, new_n18049, new_n18050, new_n18051, new_n18052, new_n18053,
    new_n18054, new_n18055, new_n18056, new_n18057, new_n18058,
    new_n18059_1, new_n18060, new_n18061_1, new_n18062, new_n18063,
    new_n18064, new_n18065, new_n18066, new_n18067, new_n18068, new_n18069,
    new_n18070, new_n18071_1, new_n18072, new_n18073, new_n18074,
    new_n18075, new_n18076, new_n18077, new_n18078, new_n18079, new_n18080,
    new_n18081, new_n18082, new_n18083, new_n18084, new_n18085, new_n18086,
    new_n18087, new_n18088, new_n18089, new_n18090, new_n18091, new_n18092,
    new_n18093, new_n18094, new_n18095, new_n18096, new_n18097, new_n18098,
    new_n18099, new_n18100, new_n18101, new_n18102, new_n18103, new_n18104,
    new_n18105_1, new_n18106, new_n18107, new_n18108, new_n18109,
    new_n18110, new_n18111, new_n18112, new_n18113, new_n18114, new_n18115,
    new_n18116, new_n18117, new_n18118, new_n18119, new_n18120, new_n18121,
    new_n18122, new_n18123, new_n18124, new_n18125, new_n18126, new_n18127,
    new_n18128, new_n18129, new_n18130, new_n18131, new_n18132, new_n18133,
    new_n18134, new_n18135, new_n18136, new_n18137, new_n18138, new_n18139,
    new_n18140, new_n18141, new_n18142, new_n18143_1, new_n18144,
    new_n18145_1, new_n18146, new_n18147, new_n18148, new_n18149,
    new_n18150, new_n18151_1, new_n18152_1, new_n18153, new_n18154,
    new_n18155, new_n18156, new_n18157_1, new_n18158, new_n18159,
    new_n18160, new_n18161, new_n18163, new_n18164, new_n18165, new_n18166,
    new_n18167, new_n18168, new_n18169, new_n18170, new_n18171_1,
    new_n18172, new_n18173, new_n18174, new_n18175, new_n18176, new_n18177,
    new_n18178, new_n18179, new_n18180, new_n18181, new_n18182, new_n18183,
    new_n18184, new_n18185, new_n18186, new_n18187, new_n18188, new_n18189,
    new_n18190, new_n18191, new_n18192, new_n18193_1, new_n18194,
    new_n18195, new_n18196, new_n18197, new_n18198, new_n18199, new_n18200,
    new_n18201, new_n18202, new_n18203, new_n18204, new_n18205, new_n18206,
    new_n18207, new_n18208, new_n18209, new_n18210, new_n18211, new_n18212,
    new_n18213, new_n18214, new_n18215, new_n18216, new_n18217, new_n18218,
    new_n18219, new_n18220, new_n18221, new_n18222, new_n18223, new_n18224,
    new_n18225, new_n18226, new_n18227_1, new_n18228, new_n18229,
    new_n18230, new_n18231, new_n18232_1, new_n18233, new_n18234,
    new_n18235, new_n18236, new_n18237, new_n18238_1, new_n18239,
    new_n18240, new_n18241_1, new_n18242, new_n18243, new_n18244,
    new_n18245, new_n18246, new_n18247, new_n18248, new_n18249, new_n18250,
    new_n18251, new_n18252, new_n18253, new_n18254_1, new_n18255,
    new_n18256, new_n18257, new_n18258, new_n18259, new_n18260, new_n18261,
    new_n18262, new_n18263, new_n18264, new_n18265, new_n18266, new_n18267,
    new_n18268, new_n18269, new_n18270, new_n18271, new_n18272, new_n18273,
    new_n18274_1, new_n18275, new_n18276, new_n18277, new_n18278,
    new_n18279, new_n18280, new_n18281, new_n18282, new_n18283, new_n18284,
    new_n18285, new_n18286, new_n18287, new_n18288_1, new_n18289,
    new_n18290_1, new_n18291, new_n18292, new_n18298, new_n18300,
    new_n18302, new_n18303, new_n18304_1, new_n18306, new_n18307,
    new_n18308, new_n18309, new_n18310_1, new_n18311_1, new_n18312,
    new_n18313, new_n18314, new_n18315, new_n18316, new_n18317, new_n18318,
    new_n18319, new_n18320, new_n18321, new_n18322, new_n18323_1,
    new_n18324, new_n18325, new_n18326, new_n18327, new_n18328, new_n18329,
    new_n18330, new_n18331, new_n18332_1, new_n18333, new_n18334,
    new_n18335, new_n18336, new_n18337, new_n18338, new_n18339, new_n18340,
    new_n18341, new_n18342, new_n18343_1, new_n18346, new_n18347,
    new_n18348, new_n18349, new_n18350_1, new_n18351, new_n18352,
    new_n18353, new_n18354, new_n18355, new_n18356, new_n18357, new_n18358,
    new_n18359, new_n18360, new_n18361, new_n18362_1, new_n18363,
    new_n18364, new_n18365, new_n18366, new_n18367, new_n18368, new_n18369,
    new_n18370, new_n18371, new_n18372, new_n18373, new_n18374, new_n18375,
    new_n18376, new_n18377_1, new_n18378, new_n18379, new_n18380,
    new_n18381, new_n18382, new_n18383, new_n18384, new_n18385, new_n18386,
    new_n18387, new_n18388, new_n18389, new_n18390, new_n18391, new_n18392,
    new_n18393, new_n18394, new_n18395, new_n18396, new_n18397, new_n18398,
    new_n18399, new_n18400, new_n18401, new_n18402, new_n18403, new_n18404,
    new_n18405_1, new_n18406, new_n18407, new_n18408, new_n18409_1,
    new_n18410, new_n18411, new_n18412, new_n18413, new_n18414_1,
    new_n18415, new_n18416, new_n18417, new_n18418_1, new_n18419,
    new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425,
    new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431,
    new_n18434, new_n18436, new_n18439_1, new_n18440, new_n18441,
    new_n18442, new_n18443, new_n18444_1, new_n18445_1, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451,
    new_n18452_1, new_n18453, new_n18454, new_n18455, new_n18456,
    new_n18457, new_n18458, new_n18459, new_n18460, new_n18461, new_n18462,
    new_n18463, new_n18464, new_n18465, new_n18466, new_n18467_1,
    new_n18468, new_n18469, new_n18470, new_n18471, new_n18472, new_n18473,
    new_n18474, new_n18475, new_n18476, new_n18477, new_n18478, new_n18479,
    new_n18480, new_n18481, new_n18482_1, new_n18483_1, new_n18484,
    new_n18485, new_n18486, new_n18487, new_n18488, new_n18489, new_n18490,
    new_n18491, new_n18492, new_n18493, new_n18494, new_n18495,
    new_n18496_1, new_n18497, new_n18498, new_n18499, new_n18500,
    new_n18501, new_n18502, new_n18503, new_n18504, new_n18505, new_n18506,
    new_n18507, new_n18508, new_n18509_1, new_n18510, new_n18511,
    new_n18512, new_n18513_1, new_n18514, new_n18515_1, new_n18516,
    new_n18517, new_n18518, new_n18519, new_n18520, new_n18521, new_n18522,
    new_n18523, new_n18524, new_n18525, new_n18526, new_n18527, new_n18528,
    new_n18529, new_n18530, new_n18531, new_n18532, new_n18533, new_n18534,
    new_n18535, new_n18536, new_n18537_1, new_n18538, new_n18539,
    new_n18540, new_n18541, new_n18542, new_n18543, new_n18544, new_n18545,
    new_n18546, new_n18547, new_n18548, new_n18549, new_n18550, new_n18551,
    new_n18552, new_n18553, new_n18554, new_n18555, new_n18556, new_n18557,
    new_n18558_1, new_n18559, new_n18560, new_n18561, new_n18562,
    new_n18563, new_n18564, new_n18565, new_n18566, new_n18567, new_n18568,
    new_n18569, new_n18570, new_n18571, new_n18572_1, new_n18573,
    new_n18574_1, new_n18575, new_n18576_1, new_n18577, new_n18578_1,
    new_n18579, new_n18580, new_n18581, new_n18582_1, new_n18583_1,
    new_n18584_1, new_n18585, new_n18586, new_n18587, new_n18588,
    new_n18589, new_n18590, new_n18591, new_n18592, new_n18593, new_n18594,
    new_n18595, new_n18596, new_n18597, new_n18598, new_n18599, new_n18600,
    new_n18601, new_n18602, new_n18603, new_n18604, new_n18605, new_n18606,
    new_n18607, new_n18609, new_n18611, new_n18612, new_n18613, new_n18614,
    new_n18615, new_n18616, new_n18617, new_n18618, new_n18619, new_n18620,
    new_n18621, new_n18622, new_n18623, new_n18624, new_n18625, new_n18626,
    new_n18627, new_n18628, new_n18629, new_n18630, new_n18631, new_n18632,
    new_n18633, new_n18634, new_n18635_1, new_n18636, new_n18637,
    new_n18638, new_n18639, new_n18640, new_n18641, new_n18642, new_n18643,
    new_n18644, new_n18645, new_n18646, new_n18647, new_n18648,
    new_n18649_1, new_n18650, new_n18651, new_n18652, new_n18653_1,
    new_n18654, new_n18655, new_n18656, new_n18657, new_n18658, new_n18659,
    new_n18660, new_n18661, new_n18662, new_n18663, new_n18664, new_n18665,
    new_n18666, new_n18667, new_n18668, new_n18669, new_n18670, new_n18671,
    new_n18672, new_n18673, new_n18674, new_n18675, new_n18676, new_n18677,
    new_n18678, new_n18679_1, new_n18680, new_n18681, new_n18682,
    new_n18683, new_n18684, new_n18685, new_n18686, new_n18687, new_n18688,
    new_n18689, new_n18690_1, new_n18691, new_n18692, new_n18694,
    new_n18695, new_n18696, new_n18697, new_n18698, new_n18699, new_n18700,
    new_n18701, new_n18702, new_n18703, new_n18704, new_n18705, new_n18706,
    new_n18707, new_n18708_1, new_n18709, new_n18710, new_n18711,
    new_n18712, new_n18713, new_n18714, new_n18715, new_n18716, new_n18717,
    new_n18718, new_n18719, new_n18720, new_n18721_1, new_n18722,
    new_n18723, new_n18724, new_n18725_1, new_n18726, new_n18727,
    new_n18728, new_n18729, new_n18730, new_n18731, new_n18732, new_n18733,
    new_n18735, new_n18737_1, new_n18738, new_n18739, new_n18740,
    new_n18741, new_n18742, new_n18743, new_n18744, new_n18745_1,
    new_n18746, new_n18747, new_n18748, new_n18749, new_n18750,
    new_n18751_1, new_n18752, new_n18753, new_n18754, new_n18755,
    new_n18756, new_n18757, new_n18758, new_n18759, new_n18760, new_n18761,
    new_n18762, new_n18763, new_n18764, new_n18765, new_n18766, new_n18767,
    new_n18768, new_n18769, new_n18770, new_n18771, new_n18772, new_n18773,
    new_n18774, new_n18775, new_n18776, new_n18777, new_n18778, new_n18779,
    new_n18780_1, new_n18781, new_n18782_1, new_n18783, new_n18784,
    new_n18786, new_n18787, new_n18788, new_n18789, new_n18790, new_n18791,
    new_n18792, new_n18793, new_n18794, new_n18795, new_n18796, new_n18797,
    new_n18798, new_n18799, new_n18800, new_n18801, new_n18802_1,
    new_n18803, new_n18804, new_n18805, new_n18806, new_n18807, new_n18808,
    new_n18809, new_n18810, new_n18811, new_n18812, new_n18813, new_n18814,
    new_n18815, new_n18816, new_n18817, new_n18818, new_n18819, new_n18820,
    new_n18821, new_n18822, new_n18823, new_n18824, new_n18825, new_n18826,
    new_n18827, new_n18828, new_n18829, new_n18830_1, new_n18831_1,
    new_n18832, new_n18833, new_n18835, new_n18836, new_n18837, new_n18838,
    new_n18839, new_n18840, new_n18841, new_n18842, new_n18843_1,
    new_n18844, new_n18845, new_n18846, new_n18847, new_n18848, new_n18849,
    new_n18850, new_n18851, new_n18852, new_n18853, new_n18854, new_n18855,
    new_n18856, new_n18857, new_n18858_1, new_n18859_1, new_n18860,
    new_n18861, new_n18862, new_n18863, new_n18864_1, new_n18865_1,
    new_n18866, new_n18867, new_n18868, new_n18869, new_n18870, new_n18871,
    new_n18872, new_n18873, new_n18874, new_n18875, new_n18876, new_n18877,
    new_n18878, new_n18879, new_n18880_1, new_n18881, new_n18882,
    new_n18883, new_n18884, new_n18885, new_n18886_1, new_n18887_1,
    new_n18888, new_n18889, new_n18890, new_n18891, new_n18892, new_n18893,
    new_n18894, new_n18895, new_n18896, new_n18897, new_n18898, new_n18899,
    new_n18900, new_n18901_1, new_n18902, new_n18903, new_n18904,
    new_n18905, new_n18906, new_n18907_1, new_n18908, new_n18909,
    new_n18910, new_n18911, new_n18912, new_n18913, new_n18914, new_n18915,
    new_n18916, new_n18917, new_n18918, new_n18919_1, new_n18920,
    new_n18921, new_n18922, new_n18923, new_n18924, new_n18925,
    new_n18926_1, new_n18927, new_n18928, new_n18929, new_n18930,
    new_n18931, new_n18932, new_n18933, new_n18934, new_n18935, new_n18936,
    new_n18937, new_n18938, new_n18939, new_n18940_1, new_n18941,
    new_n18942, new_n18943, new_n18944, new_n18945_1, new_n18946,
    new_n18947, new_n18948, new_n18949, new_n18950, new_n18951, new_n18952,
    new_n18953, new_n18954, new_n18955, new_n18956, new_n18957, new_n18958,
    new_n18959, new_n18960, new_n18961, new_n18962_1, new_n18963,
    new_n18964, new_n18965, new_n18966, new_n18967, new_n18968, new_n18969,
    new_n18970_1, new_n18971, new_n18972, new_n18973, new_n18974,
    new_n18975, new_n18976, new_n18977_1, new_n18978, new_n18979,
    new_n18980, new_n18981, new_n18982_1, new_n18983, new_n18984,
    new_n18985, new_n18986, new_n18987, new_n18988, new_n18989, new_n18990,
    new_n18991, new_n18992, new_n18993, new_n18994, new_n18995, new_n18996,
    new_n18997, new_n18998, new_n18999_1, new_n19000, new_n19001,
    new_n19002, new_n19003, new_n19004, new_n19005_1, new_n19006,
    new_n19007, new_n19008, new_n19009, new_n19010, new_n19011, new_n19012,
    new_n19013, new_n19014, new_n19015, new_n19016, new_n19017, new_n19018,
    new_n19019, new_n19020, new_n19021, new_n19022, new_n19023, new_n19024,
    new_n19025, new_n19026, new_n19027, new_n19028, new_n19029, new_n19030,
    new_n19031, new_n19032, new_n19033_1, new_n19034, new_n19035,
    new_n19036, new_n19037, new_n19038, new_n19039, new_n19040, new_n19041,
    new_n19042_1, new_n19043, new_n19044_1, new_n19045, new_n19046,
    new_n19047, new_n19048, new_n19049, new_n19050, new_n19051, new_n19052,
    new_n19054, new_n19057, new_n19059, new_n19060, new_n19061, new_n19062,
    new_n19063, new_n19064, new_n19065, new_n19066, new_n19067, new_n19068,
    new_n19069, new_n19070, new_n19071, new_n19072, new_n19073, new_n19074,
    new_n19075, new_n19076, new_n19077, new_n19078, new_n19079, new_n19082,
    new_n19083, new_n19084, new_n19085, new_n19086, new_n19087, new_n19088,
    new_n19089, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19106,
    new_n19107_1, new_n19108, new_n19109, new_n19110, new_n19111,
    new_n19112, new_n19113, new_n19114, new_n19115, new_n19116_1,
    new_n19117, new_n19118, new_n19119, new_n19120, new_n19121, new_n19122,
    new_n19123, new_n19124, new_n19125_1, new_n19126, new_n19127,
    new_n19128, new_n19129, new_n19130, new_n19131, new_n19132, new_n19133,
    new_n19134, new_n19135, new_n19136, new_n19137, new_n19138, new_n19139,
    new_n19140, new_n19141_1, new_n19142, new_n19143, new_n19144_1,
    new_n19145, new_n19146, new_n19147, new_n19148, new_n19149, new_n19150,
    new_n19151, new_n19152, new_n19153, new_n19154, new_n19155, new_n19156,
    new_n19157, new_n19158, new_n19159, new_n19160, new_n19161, new_n19162,
    new_n19163_1, new_n19164_1, new_n19165, new_n19166, new_n19167,
    new_n19168, new_n19169, new_n19170, new_n19171, new_n19172, new_n19173,
    new_n19174_1, new_n19175, new_n19176_1, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19187, new_n19188, new_n19189, new_n19190,
    new_n19191, new_n19192, new_n19193, new_n19194, new_n19195,
    new_n19196_1, new_n19197, new_n19198, new_n19199, new_n19200,
    new_n19201, new_n19202_1, new_n19203, new_n19204, new_n19205,
    new_n19206, new_n19207, new_n19208, new_n19209, new_n19210, new_n19211,
    new_n19212, new_n19213, new_n19214, new_n19215, new_n19216, new_n19217,
    new_n19218, new_n19219, new_n19220_1, new_n19221_1, new_n19222,
    new_n19223_1, new_n19224_1, new_n19225, new_n19226, new_n19227,
    new_n19228_1, new_n19229, new_n19230, new_n19231, new_n19234_1,
    new_n19235, new_n19236, new_n19237, new_n19238, new_n19239, new_n19240,
    new_n19241, new_n19242, new_n19243, new_n19244_1, new_n19245,
    new_n19246, new_n19247, new_n19248, new_n19249, new_n19250, new_n19251,
    new_n19252, new_n19253, new_n19254, new_n19255, new_n19256, new_n19257,
    new_n19258, new_n19259, new_n19260, new_n19262, new_n19263, new_n19264,
    new_n19265, new_n19266, new_n19267, new_n19268, new_n19269,
    new_n19270_1, new_n19271, new_n19272, new_n19273, new_n19274,
    new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280,
    new_n19281, new_n19282_1, new_n19283, new_n19284, new_n19285,
    new_n19286, new_n19287, new_n19288, new_n19289, new_n19290, new_n19291,
    new_n19292, new_n19293, new_n19296, new_n19297, new_n19298, new_n19299,
    new_n19300, new_n19301, new_n19302, new_n19303, new_n19304, new_n19305,
    new_n19306, new_n19307, new_n19308, new_n19309, new_n19310, new_n19311,
    new_n19312, new_n19313, new_n19314_1, new_n19315_1, new_n19316,
    new_n19317, new_n19318, new_n19319, new_n19320, new_n19321, new_n19322,
    new_n19323_1, new_n19324, new_n19325, new_n19326, new_n19327_1,
    new_n19328, new_n19329, new_n19330, new_n19331, new_n19332,
    new_n19333_1, new_n19334, new_n19335, new_n19336, new_n19337,
    new_n19338, new_n19339, new_n19340, new_n19341, new_n19342, new_n19343,
    new_n19344, new_n19345, new_n19346, new_n19347, new_n19348_1,
    new_n19349, new_n19350, new_n19351, new_n19353, new_n19354_1,
    new_n19355, new_n19356, new_n19357_1, new_n19358, new_n19359,
    new_n19360, new_n19361_1, new_n19362, new_n19363, new_n19364,
    new_n19365, new_n19366, new_n19367_1, new_n19368, new_n19369,
    new_n19370, new_n19371, new_n19372, new_n19373, new_n19374, new_n19375,
    new_n19376, new_n19377, new_n19378, new_n19379, new_n19380, new_n19381,
    new_n19382, new_n19383, new_n19384, new_n19385_1, new_n19386,
    new_n19387, new_n19388, new_n19389_1, new_n19390, new_n19391,
    new_n19392, new_n19393, new_n19394, new_n19395, new_n19396, new_n19397,
    new_n19398, new_n19399, new_n19400, new_n19401_1, new_n19402,
    new_n19403, new_n19404, new_n19405, new_n19406, new_n19407, new_n19408,
    new_n19409, new_n19410, new_n19411, new_n19412, new_n19413,
    new_n19414_1, new_n19415, new_n19416, new_n19417, new_n19418,
    new_n19419, new_n19420, new_n19421, new_n19422, new_n19423,
    new_n19424_1, new_n19425, new_n19426, new_n19427, new_n19428,
    new_n19429, new_n19430, new_n19431, new_n19432, new_n19433, new_n19434,
    new_n19435, new_n19436, new_n19437, new_n19438, new_n19439, new_n19440,
    new_n19441, new_n19442, new_n19443, new_n19444, new_n19445, new_n19446,
    new_n19447, new_n19448, new_n19449, new_n19450_1, new_n19451,
    new_n19452, new_n19453, new_n19454_1, new_n19455, new_n19456,
    new_n19457, new_n19458_1, new_n19459, new_n19460, new_n19461,
    new_n19462, new_n19463, new_n19464, new_n19465, new_n19466,
    new_n19467_1, new_n19468, new_n19469, new_n19470, new_n19471,
    new_n19472_1, new_n19473, new_n19474, new_n19475, new_n19476,
    new_n19477_1, new_n19478, new_n19479, new_n19480, new_n19481,
    new_n19482, new_n19483, new_n19484, new_n19485, new_n19486, new_n19487,
    new_n19488, new_n19489, new_n19490, new_n19491, new_n19492, new_n19493,
    new_n19494_1, new_n19495, new_n19496_1, new_n19497, new_n19498,
    new_n19499, new_n19500, new_n19501, new_n19502, new_n19503, new_n19504,
    new_n19505, new_n19506, new_n19507, new_n19508, new_n19509, new_n19510,
    new_n19511, new_n19512, new_n19513, new_n19514_1, new_n19515_1,
    new_n19516, new_n19517, new_n19518, new_n19519, new_n19520, new_n19521,
    new_n19522, new_n19523_1, new_n19524, new_n19525, new_n19526,
    new_n19527, new_n19528, new_n19529, new_n19530, new_n19531_1,
    new_n19532, new_n19533, new_n19534, new_n19535, new_n19536, new_n19537,
    new_n19538, new_n19539_1, new_n19540, new_n19541, new_n19542,
    new_n19543, new_n19544, new_n19545, new_n19546, new_n19547, new_n19548,
    new_n19549, new_n19550, new_n19551, new_n19552, new_n19553, new_n19554,
    new_n19555, new_n19556, new_n19557, new_n19558, new_n19559, new_n19560,
    new_n19561, new_n19562, new_n19563, new_n19564, new_n19565, new_n19566,
    new_n19567, new_n19568, new_n19569, new_n19570_1, new_n19571,
    new_n19572, new_n19573, new_n19574, new_n19575_1, new_n19576,
    new_n19577, new_n19578, new_n19579, new_n19581, new_n19582, new_n19583,
    new_n19584_1, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602_1, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608_1, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617_1, new_n19618_1, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623_1, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641_1, new_n19642, new_n19643,
    new_n19644, new_n19645, new_n19646, new_n19647, new_n19648_1,
    new_n19649, new_n19650, new_n19651, new_n19652_1, new_n19653,
    new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659,
    new_n19660, new_n19661, new_n19662, new_n19663, new_n19664_1,
    new_n19665, new_n19666, new_n19667, new_n19668, new_n19669, new_n19670,
    new_n19671, new_n19672, new_n19673, new_n19674, new_n19675, new_n19676,
    new_n19677, new_n19678, new_n19679, new_n19680_1, new_n19681,
    new_n19682, new_n19683, new_n19684, new_n19685, new_n19686, new_n19687,
    new_n19688, new_n19689, new_n19690, new_n19691, new_n19692, new_n19693,
    new_n19694, new_n19695, new_n19696, new_n19697, new_n19698, new_n19699,
    new_n19700, new_n19701_1, new_n19702, new_n19703, new_n19704,
    new_n19705, new_n19706, new_n19707, new_n19708, new_n19709, new_n19710,
    new_n19711, new_n19712, new_n19713, new_n19714, new_n19715, new_n19716,
    new_n19717, new_n19718, new_n19719, new_n19722, new_n19723, new_n19724,
    new_n19725, new_n19726, new_n19727, new_n19728, new_n19729, new_n19730,
    new_n19731, new_n19732, new_n19733, new_n19734, new_n19735,
    new_n19736_1, new_n19737, new_n19738, new_n19739, new_n19740,
    new_n19741, new_n19742, new_n19743, new_n19744, new_n19745, new_n19746,
    new_n19747, new_n19748, new_n19749_1, new_n19750, new_n19751,
    new_n19752, new_n19753, new_n19754, new_n19755, new_n19756_1,
    new_n19757, new_n19758, new_n19759, new_n19760, new_n19761, new_n19762,
    new_n19763, new_n19764, new_n19765, new_n19766, new_n19767_1,
    new_n19768, new_n19769, new_n19770_1, new_n19771, new_n19772,
    new_n19773, new_n19774, new_n19775, new_n19776, new_n19777, new_n19778,
    new_n19779, new_n19780_1, new_n19781, new_n19782, new_n19783,
    new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789_1, new_n19790, new_n19791, new_n19792_1, new_n19793,
    new_n19794, new_n19795, new_n19796, new_n19797, new_n19798_1,
    new_n19799, new_n19800, new_n19801, new_n19802, new_n19803_1,
    new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809,
    new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815,
    new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821,
    new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827,
    new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833,
    new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839,
    new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845,
    new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851,
    new_n19852, new_n19854, new_n19855, new_n19856, new_n19857, new_n19858,
    new_n19859, new_n19860, new_n19861, new_n19862, new_n19863, new_n19864,
    new_n19865, new_n19866, new_n19867, new_n19868, new_n19869, new_n19870,
    new_n19871, new_n19872, new_n19873_1, new_n19874, new_n19875,
    new_n19876, new_n19877, new_n19878, new_n19879, new_n19880, new_n19881,
    new_n19882, new_n19883, new_n19884, new_n19885, new_n19886, new_n19887,
    new_n19888, new_n19889, new_n19890, new_n19891, new_n19892, new_n19893,
    new_n19894, new_n19895, new_n19896, new_n19897, new_n19898, new_n19899,
    new_n19900, new_n19901, new_n19902, new_n19903, new_n19904,
    new_n19905_1, new_n19906, new_n19907, new_n19908, new_n19909_1,
    new_n19910, new_n19911_1, new_n19912, new_n19913, new_n19914,
    new_n19915, new_n19916_1, new_n19917, new_n19918, new_n19919,
    new_n19920, new_n19921, new_n19923_1, new_n19924, new_n19925,
    new_n19926, new_n19927, new_n19928, new_n19929, new_n19930_1,
    new_n19931, new_n19932, new_n19933, new_n19934, new_n19935, new_n19936,
    new_n19937, new_n19938, new_n19939, new_n19940, new_n19941_1,
    new_n19942, new_n19943, new_n19944, new_n19945, new_n19946, new_n19947,
    new_n19948, new_n19949, new_n19950, new_n19951, new_n19952, new_n19953,
    new_n19954, new_n19955, new_n19956, new_n19957, new_n19958, new_n19959,
    new_n19961, new_n19963, new_n19964, new_n19965, new_n19966, new_n19967,
    new_n19968_1, new_n19969, new_n19970, new_n19971, new_n19972,
    new_n19973, new_n19974, new_n19975, new_n19976, new_n19977, new_n19978,
    new_n19979, new_n19980, new_n19981, new_n19982, new_n19983, new_n19984,
    new_n19985, new_n19986, new_n19987, new_n19988_1, new_n19989,
    new_n19990, new_n19991, new_n19992, new_n19993, new_n19994, new_n19995,
    new_n19996, new_n19997, new_n19998, new_n19999, new_n20000, new_n20001,
    new_n20002, new_n20003, new_n20004_1, new_n20005, new_n20006,
    new_n20007, new_n20008, new_n20009, new_n20010, new_n20011, new_n20012,
    new_n20013_1, new_n20014, new_n20015, new_n20016, new_n20017_1,
    new_n20018, new_n20019, new_n20020, new_n20021, new_n20022, new_n20023,
    new_n20024, new_n20025, new_n20026, new_n20027, new_n20028, new_n20029,
    new_n20030, new_n20031, new_n20032, new_n20033_1, new_n20034,
    new_n20035, new_n20036_1, new_n20037, new_n20038, new_n20039,
    new_n20040_1, new_n20041, new_n20042, new_n20043, new_n20044,
    new_n20045, new_n20046, new_n20047, new_n20048, new_n20049, new_n20050,
    new_n20051, new_n20052, new_n20053, new_n20054, new_n20055, new_n20057,
    new_n20060, new_n20061_1, new_n20062, new_n20063, new_n20064,
    new_n20065, new_n20066, new_n20067, new_n20068, new_n20069_1,
    new_n20070, new_n20071, new_n20072, new_n20073, new_n20074, new_n20075,
    new_n20076, new_n20077_1, new_n20079, new_n20082, new_n20083,
    new_n20084, new_n20085, new_n20086_1, new_n20087, new_n20088,
    new_n20089, new_n20090, new_n20091, new_n20092, new_n20093, new_n20094,
    new_n20095, new_n20096_1, new_n20097, new_n20098, new_n20099,
    new_n20100, new_n20101, new_n20102, new_n20103_1, new_n20104,
    new_n20105, new_n20106, new_n20107, new_n20108, new_n20109, new_n20110,
    new_n20111, new_n20112, new_n20113, new_n20114, new_n20115, new_n20116,
    new_n20119, new_n20120, new_n20121, new_n20122, new_n20123, new_n20124,
    new_n20125, new_n20126_1, new_n20127, new_n20128, new_n20129,
    new_n20130, new_n20131, new_n20132, new_n20133, new_n20134, new_n20135,
    new_n20136, new_n20137, new_n20138_1, new_n20139, new_n20140,
    new_n20141, new_n20142, new_n20143, new_n20144, new_n20145, new_n20146,
    new_n20147, new_n20148, new_n20149_1, new_n20150, new_n20151_1,
    new_n20152, new_n20153, new_n20154, new_n20155, new_n20156, new_n20157,
    new_n20158, new_n20159, new_n20160, new_n20161, new_n20162, new_n20163,
    new_n20164, new_n20165, new_n20166, new_n20167, new_n20168,
    new_n20169_1, new_n20170, new_n20171, new_n20172, new_n20173,
    new_n20174, new_n20175, new_n20176, new_n20177, new_n20178,
    new_n20179_1, new_n20180, new_n20181, new_n20182, new_n20183,
    new_n20184, new_n20185, new_n20186, new_n20187_1, new_n20188,
    new_n20189, new_n20190, new_n20191, new_n20192, new_n20193, new_n20194,
    new_n20195, new_n20196, new_n20197, new_n20198, new_n20199, new_n20200,
    new_n20201, new_n20202, new_n20203, new_n20204, new_n20205, new_n20206,
    new_n20207, new_n20208, new_n20209, new_n20210, new_n20211, new_n20212,
    new_n20213_1, new_n20214, new_n20215, new_n20216, new_n20217,
    new_n20218, new_n20219, new_n20220, new_n20221, new_n20222, new_n20223,
    new_n20224, new_n20225, new_n20226, new_n20227, new_n20228, new_n20229,
    new_n20230, new_n20231, new_n20232, new_n20233, new_n20234,
    new_n20235_1, new_n20236, new_n20237, new_n20238, new_n20239,
    new_n20240, new_n20241, new_n20242, new_n20243, new_n20244, new_n20245,
    new_n20247, new_n20250_1, new_n20251, new_n20252, new_n20253,
    new_n20254, new_n20255, new_n20256, new_n20257, new_n20258,
    new_n20259_1, new_n20260, new_n20261, new_n20262, new_n20263,
    new_n20264, new_n20265, new_n20266, new_n20267, new_n20268, new_n20269,
    new_n20270, new_n20271, new_n20272, new_n20273, new_n20274, new_n20275,
    new_n20276, new_n20277, new_n20278, new_n20279_1, new_n20280,
    new_n20281, new_n20282, new_n20283, new_n20284, new_n20285, new_n20286,
    new_n20287_1, new_n20288, new_n20289, new_n20290, new_n20291,
    new_n20292, new_n20293, new_n20294, new_n20295, new_n20296, new_n20297,
    new_n20298, new_n20299, new_n20300, new_n20301_1, new_n20302,
    new_n20303, new_n20304, new_n20305, new_n20306, new_n20307, new_n20308,
    new_n20309, new_n20310, new_n20311, new_n20312, new_n20313, new_n20314,
    new_n20315, new_n20316, new_n20317, new_n20318, new_n20319, new_n20320,
    new_n20321, new_n20322, new_n20323, new_n20324, new_n20325, new_n20326,
    new_n20327, new_n20328, new_n20329, new_n20330_1, new_n20331,
    new_n20332, new_n20333_1, new_n20334, new_n20335, new_n20336,
    new_n20337, new_n20338, new_n20339, new_n20340, new_n20341, new_n20342,
    new_n20343, new_n20344, new_n20345, new_n20346, new_n20347, new_n20348,
    new_n20349_1, new_n20350, new_n20351, new_n20352, new_n20353,
    new_n20354, new_n20355_1, new_n20356, new_n20357, new_n20358,
    new_n20359_1, new_n20360, new_n20361, new_n20362, new_n20363,
    new_n20364, new_n20365, new_n20366_1, new_n20367, new_n20368,
    new_n20369, new_n20370, new_n20371, new_n20372, new_n20373, new_n20374,
    new_n20375, new_n20376, new_n20377, new_n20378, new_n20379, new_n20380,
    new_n20381, new_n20382, new_n20383, new_n20384, new_n20385_1,
    new_n20386, new_n20387, new_n20388_1, new_n20389, new_n20390,
    new_n20391, new_n20392, new_n20393, new_n20394, new_n20395, new_n20396,
    new_n20397, new_n20398, new_n20399, new_n20400, new_n20401,
    new_n20402_1, new_n20403_1, new_n20404, new_n20405, new_n20406,
    new_n20407, new_n20408, new_n20409_1, new_n20410, new_n20411_1,
    new_n20412, new_n20413, new_n20414, new_n20415, new_n20416, new_n20417,
    new_n20418, new_n20420, new_n20421, new_n20422, new_n20423,
    new_n20424_1, new_n20425, new_n20426, new_n20427, new_n20428,
    new_n20429_1, new_n20430, new_n20431, new_n20432, new_n20433,
    new_n20434, new_n20435, new_n20436_1, new_n20437, new_n20438,
    new_n20440, new_n20441_1, new_n20442, new_n20443, new_n20444,
    new_n20445_1, new_n20446, new_n20447, new_n20448, new_n20449,
    new_n20450_1, new_n20451, new_n20452, new_n20453, new_n20454,
    new_n20455_1, new_n20456, new_n20457, new_n20458, new_n20459,
    new_n20460, new_n20461, new_n20462, new_n20463, new_n20464, new_n20465,
    new_n20466, new_n20467, new_n20468, new_n20469, new_n20470_1,
    new_n20471, new_n20472, new_n20473, new_n20474, new_n20475, new_n20476,
    new_n20477, new_n20478_1, new_n20479, new_n20480, new_n20481,
    new_n20482, new_n20483, new_n20485, new_n20486, new_n20487, new_n20488,
    new_n20489_1, new_n20490_1, new_n20491, new_n20492, new_n20493,
    new_n20494, new_n20495_1, new_n20496, new_n20497, new_n20498,
    new_n20499, new_n20500, new_n20501, new_n20502, new_n20503, new_n20504,
    new_n20505, new_n20506, new_n20507, new_n20508, new_n20509, new_n20510,
    new_n20511, new_n20512, new_n20513, new_n20514, new_n20515_1,
    new_n20516, new_n20517, new_n20518, new_n20519, new_n20520, new_n20521,
    new_n20522, new_n20523, new_n20524, new_n20525, new_n20526, new_n20527,
    new_n20528, new_n20529, new_n20530, new_n20532, new_n20533_1,
    new_n20534, new_n20535, new_n20536, new_n20537, new_n20538, new_n20539,
    new_n20540, new_n20541, new_n20542, new_n20543, new_n20544, new_n20545,
    new_n20546, new_n20547, new_n20548, new_n20549, new_n20550, new_n20551,
    new_n20552, new_n20553, new_n20554, new_n20555, new_n20556, new_n20557,
    new_n20558, new_n20559, new_n20560, new_n20561, new_n20562, new_n20563,
    new_n20564, new_n20565, new_n20566, new_n20567, new_n20568, new_n20569,
    new_n20570, new_n20571, new_n20572, new_n20573, new_n20574, new_n20576,
    new_n20578, new_n20579, new_n20580, new_n20581, new_n20582_1,
    new_n20583, new_n20584, new_n20585, new_n20586, new_n20587, new_n20588,
    new_n20589, new_n20590_1, new_n20591, new_n20592, new_n20593,
    new_n20594, new_n20595, new_n20596, new_n20597, new_n20598, new_n20599,
    new_n20600, new_n20601, new_n20602_1, new_n20604_1, new_n20605,
    new_n20606, new_n20607, new_n20608, new_n20609_1, new_n20610,
    new_n20611, new_n20612, new_n20613, new_n20614, new_n20615, new_n20616,
    new_n20617, new_n20618, new_n20619, new_n20620, new_n20621, new_n20622,
    new_n20623_1, new_n20624, new_n20625, new_n20626, new_n20627,
    new_n20628, new_n20629_1, new_n20630, new_n20631, new_n20632,
    new_n20633, new_n20634, new_n20635, new_n20636, new_n20637, new_n20638,
    new_n20639, new_n20640, new_n20641, new_n20642, new_n20643, new_n20644,
    new_n20645, new_n20646, new_n20647, new_n20648, new_n20649, new_n20650,
    new_n20651, new_n20652, new_n20653, new_n20654, new_n20655, new_n20656,
    new_n20657, new_n20658_1, new_n20659, new_n20660, new_n20661_1,
    new_n20662, new_n20663, new_n20664, new_n20665, new_n20666, new_n20667,
    new_n20668, new_n20669, new_n20670, new_n20671, new_n20672,
    new_n20673_1, new_n20674, new_n20675, new_n20676, new_n20677,
    new_n20678_1, new_n20679, new_n20680_1, new_n20681, new_n20682,
    new_n20683, new_n20684, new_n20685_1, new_n20686, new_n20687,
    new_n20688, new_n20689, new_n20690, new_n20691_1, new_n20692,
    new_n20693, new_n20694, new_n20695, new_n20696_1, new_n20697,
    new_n20698, new_n20699, new_n20701, new_n20702, new_n20703,
    new_n20704_1, new_n20705_1, new_n20706, new_n20707, new_n20708,
    new_n20709_1, new_n20710, new_n20711, new_n20712, new_n20713_1,
    new_n20714, new_n20715, new_n20716, new_n20717, new_n20718, new_n20719,
    new_n20720, new_n20721, new_n20722_1, new_n20723_1, new_n20724,
    new_n20725, new_n20726, new_n20727, new_n20728, new_n20729, new_n20730,
    new_n20731, new_n20732, new_n20733, new_n20734, new_n20735, new_n20736,
    new_n20737, new_n20738, new_n20739, new_n20740, new_n20741, new_n20742,
    new_n20743, new_n20744, new_n20745, new_n20746, new_n20747,
    new_n20748_1, new_n20749, new_n20750, new_n20751, new_n20752,
    new_n20753, new_n20754, new_n20755, new_n20756, new_n20757, new_n20758,
    new_n20759, new_n20760, new_n20761_1, new_n20762, new_n20763,
    new_n20764, new_n20765, new_n20766, new_n20767, new_n20768, new_n20769,
    new_n20770, new_n20771, new_n20772, new_n20773, new_n20774_1,
    new_n20775, new_n20776, new_n20777, new_n20778, new_n20779, new_n20780,
    new_n20781, new_n20782, new_n20783, new_n20784, new_n20785, new_n20786,
    new_n20787, new_n20788_1, new_n20789, new_n20790, new_n20791,
    new_n20792, new_n20793, new_n20794_1, new_n20795_1, new_n20796,
    new_n20797, new_n20798, new_n20799, new_n20800, new_n20801, new_n20802,
    new_n20803_1, new_n20804, new_n20805, new_n20806, new_n20807,
    new_n20808, new_n20809, new_n20810, new_n20811, new_n20812, new_n20813,
    new_n20814, new_n20815, new_n20816, new_n20817, new_n20818, new_n20819,
    new_n20820, new_n20821, new_n20822, new_n20823, new_n20824, new_n20825,
    new_n20826_1, new_n20827, new_n20828, new_n20829, new_n20830,
    new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20836,
    new_n20837, new_n20838, new_n20839, new_n20840, new_n20841, new_n20842,
    new_n20843, new_n20844, new_n20845, new_n20846, new_n20847, new_n20848,
    new_n20849, new_n20850, new_n20851, new_n20852, new_n20853, new_n20854,
    new_n20855, new_n20856, new_n20857, new_n20858, new_n20859, new_n20860,
    new_n20861, new_n20862, new_n20863, new_n20864, new_n20865, new_n20866,
    new_n20867, new_n20868, new_n20869_1, new_n20870, new_n20871,
    new_n20872, new_n20873, new_n20874, new_n20875, new_n20876, new_n20877,
    new_n20878, new_n20879_1, new_n20880, new_n20881, new_n20882,
    new_n20883, new_n20884, new_n20885, new_n20886, new_n20887, new_n20888,
    new_n20889, new_n20890, new_n20891, new_n20892, new_n20893, new_n20894,
    new_n20895, new_n20896, new_n20897, new_n20899, new_n20900, new_n20901,
    new_n20902, new_n20903, new_n20904, new_n20905, new_n20906, new_n20907,
    new_n20908, new_n20909, new_n20910, new_n20911, new_n20912, new_n20913,
    new_n20914, new_n20915_1, new_n20916, new_n20917, new_n20918,
    new_n20919, new_n20920, new_n20921, new_n20922, new_n20925, new_n20926,
    new_n20927, new_n20928, new_n20929_1, new_n20930, new_n20931,
    new_n20932, new_n20933, new_n20934, new_n20935_1, new_n20936_1,
    new_n20937, new_n20938, new_n20940, new_n20942, new_n20945,
    new_n20946_1, new_n20947, new_n20948, new_n20949, new_n20950,
    new_n20951, new_n20952, new_n20953, new_n20954, new_n20955, new_n20956,
    new_n20957, new_n20958, new_n20962, new_n20964, new_n20966, new_n20968,
    new_n20969, new_n20970, new_n20971, new_n20972, new_n20973, new_n20974,
    new_n20975, new_n20976, new_n20977, new_n20978, new_n20979, new_n20980,
    new_n20981, new_n20982, new_n20983, new_n20984, new_n20985,
    new_n20986_1, new_n20987, new_n20988, new_n20989, new_n20990,
    new_n20991, new_n20992, new_n20993, new_n20994, new_n20995, new_n20996,
    new_n20997, new_n20998, new_n20999, new_n21000, new_n21001, new_n21002,
    new_n21003, new_n21004, new_n21005, new_n21006, new_n21007,
    new_n21008_1, new_n21009, new_n21010, new_n21011, new_n21012,
    new_n21013, new_n21014, new_n21015, new_n21016, new_n21017_1,
    new_n21018, new_n21019, new_n21020, new_n21021, new_n21022, new_n21023,
    new_n21024, new_n21025, new_n21026, new_n21027, new_n21028, new_n21029,
    new_n21030, new_n21031, new_n21032, new_n21033, new_n21034_1,
    new_n21035, new_n21036, new_n21037, new_n21038, new_n21039, new_n21040,
    new_n21041, new_n21042, new_n21043, new_n21044, new_n21045,
    new_n21046_1, new_n21047, new_n21048, new_n21049, new_n21050,
    new_n21051, new_n21052, new_n21053, new_n21054, new_n21055, new_n21056,
    new_n21057, new_n21058, new_n21059, new_n21060, new_n21061,
    new_n21062_1, new_n21063, new_n21064, new_n21065, new_n21066,
    new_n21067, new_n21068, new_n21069, new_n21070, new_n21071, new_n21072,
    new_n21073, new_n21074, new_n21075, new_n21076, new_n21077,
    new_n21078_1, new_n21079, new_n21080, new_n21081, new_n21082,
    new_n21083, new_n21084, new_n21085, new_n21086, new_n21087, new_n21088,
    new_n21089, new_n21090, new_n21091, new_n21092, new_n21093_1,
    new_n21095_1, new_n21096, new_n21097, new_n21098, new_n21099,
    new_n21100, new_n21101, new_n21102, new_n21103, new_n21104, new_n21105,
    new_n21106, new_n21107, new_n21108, new_n21109, new_n21110, new_n21111,
    new_n21112, new_n21113, new_n21114, new_n21115, new_n21116, new_n21117,
    new_n21118, new_n21119, new_n21120, new_n21121, new_n21122,
    new_n21123_1, new_n21124, new_n21125, new_n21126, new_n21127,
    new_n21128, new_n21129, new_n21130, new_n21131, new_n21132, new_n21133,
    new_n21134_1, new_n21135, new_n21136, new_n21137, new_n21138_1,
    new_n21139, new_n21140, new_n21141, new_n21142, new_n21143, new_n21144,
    new_n21145, new_n21146, new_n21148, new_n21149, new_n21150, new_n21151,
    new_n21152, new_n21153, new_n21154_1, new_n21155, new_n21156,
    new_n21157_1, new_n21158, new_n21159, new_n21160, new_n21161,
    new_n21162, new_n21163, new_n21164, new_n21165, new_n21166, new_n21167,
    new_n21168_1, new_n21169, new_n21170, new_n21171, new_n21172,
    new_n21173_1, new_n21174, new_n21175, new_n21176_1, new_n21177,
    new_n21178, new_n21179, new_n21180, new_n21181, new_n21182_1,
    new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193_1,
    new_n21194, new_n21195, new_n21196, new_n21197, new_n21198, new_n21199,
    new_n21200, new_n21201, new_n21202, new_n21203_1, new_n21204,
    new_n21205, new_n21206, new_n21207, new_n21208, new_n21209, new_n21210,
    new_n21211, new_n21212, new_n21213, new_n21214, new_n21215, new_n21216,
    new_n21217, new_n21218, new_n21219, new_n21220, new_n21221,
    new_n21222_1, new_n21223, new_n21224, new_n21225_1, new_n21226_1,
    new_n21227, new_n21228, new_n21229, new_n21230, new_n21231, new_n21232,
    new_n21233, new_n21234, new_n21235, new_n21236, new_n21237,
    new_n21238_1, new_n21239, new_n21240, new_n21241, new_n21242,
    new_n21243, new_n21244, new_n21245, new_n21246, new_n21247, new_n21248,
    new_n21249, new_n21250, new_n21251, new_n21252, new_n21253,
    new_n21254_1, new_n21255, new_n21256, new_n21257, new_n21258,
    new_n21259, new_n21260, new_n21261, new_n21262, new_n21263, new_n21264,
    new_n21265, new_n21266, new_n21267, new_n21268, new_n21269, new_n21270,
    new_n21271, new_n21272, new_n21273, new_n21274, new_n21275,
    new_n21276_1, new_n21277, new_n21278, new_n21279, new_n21280,
    new_n21281, new_n21282, new_n21283, new_n21284, new_n21285, new_n21286,
    new_n21287_1, new_n21288, new_n21289, new_n21290, new_n21291,
    new_n21292, new_n21293, new_n21294, new_n21295, new_n21296, new_n21297,
    new_n21298_1, new_n21299, new_n21300, new_n21301, new_n21302_1,
    new_n21303, new_n21304, new_n21305, new_n21306, new_n21307, new_n21308,
    new_n21309, new_n21310, new_n21311, new_n21312, new_n21313, new_n21314,
    new_n21315, new_n21316, new_n21317_1, new_n21318, new_n21319,
    new_n21320, new_n21321, new_n21322, new_n21323, new_n21324, new_n21325,
    new_n21326, new_n21327, new_n21328, new_n21329, new_n21331, new_n21332,
    new_n21333, new_n21334, new_n21335, new_n21336, new_n21337, new_n21338,
    new_n21339, new_n21340, new_n21341, new_n21342, new_n21343, new_n21344,
    new_n21345, new_n21346, new_n21347, new_n21348, new_n21349_1,
    new_n21350, new_n21351, new_n21352, new_n21353, new_n21354, new_n21355,
    new_n21356, new_n21357, new_n21358, new_n21359, new_n21360, new_n21361,
    new_n21362, new_n21363, new_n21364, new_n21365_1, new_n21366,
    new_n21367_1, new_n21368, new_n21369, new_n21370, new_n21371,
    new_n21372, new_n21373, new_n21374, new_n21375, new_n21376, new_n21377,
    new_n21378, new_n21379, new_n21380, new_n21381, new_n21382, new_n21383,
    new_n21384, new_n21385, new_n21388, new_n21389, new_n21390, new_n21391,
    new_n21392, new_n21393, new_n21394, new_n21395, new_n21396_1,
    new_n21397, new_n21398_1, new_n21399_1, new_n21400, new_n21401,
    new_n21402, new_n21403, new_n21404_1, new_n21405, new_n21406,
    new_n21407, new_n21408, new_n21409, new_n21411, new_n21413, new_n21414,
    new_n21415, new_n21416, new_n21417, new_n21418, new_n21419, new_n21420,
    new_n21423, new_n21425, new_n21426, new_n21427, new_n21428, new_n21429,
    new_n21430, new_n21431, new_n21432, new_n21433, new_n21434, new_n21435,
    new_n21436, new_n21437, new_n21438, new_n21439, new_n21440, new_n21441,
    new_n21442, new_n21443, new_n21444, new_n21445, new_n21446_1,
    new_n21447, new_n21448, new_n21449, new_n21450, new_n21451, new_n21452,
    new_n21453, new_n21454, new_n21455, new_n21456, new_n21457, new_n21458,
    new_n21459, new_n21460, new_n21461, new_n21462, new_n21463, new_n21464,
    new_n21465, new_n21466, new_n21467, new_n21468, new_n21469, new_n21470,
    new_n21471_1, new_n21472_1, new_n21473, new_n21474, new_n21475,
    new_n21476, new_n21477, new_n21478, new_n21479, new_n21480, new_n21481,
    new_n21482, new_n21483, new_n21484, new_n21485, new_n21486, new_n21487,
    new_n21488, new_n21489_1, new_n21491, new_n21493, new_n21494,
    new_n21495, new_n21496, new_n21497, new_n21498, new_n21499, new_n21500,
    new_n21501, new_n21502, new_n21503, new_n21504, new_n21505, new_n21506,
    new_n21507, new_n21508, new_n21509, new_n21510, new_n21511, new_n21512,
    new_n21513, new_n21514, new_n21515, new_n21516, new_n21517, new_n21518,
    new_n21519, new_n21520, new_n21521, new_n21522, new_n21523, new_n21524,
    new_n21525_1, new_n21526, new_n21527, new_n21528, new_n21529,
    new_n21530, new_n21531, new_n21532, new_n21533, new_n21534, new_n21535,
    new_n21536, new_n21537, new_n21538_1, new_n21539, new_n21540,
    new_n21541, new_n21542, new_n21543, new_n21544, new_n21545, new_n21546,
    new_n21547, new_n21548, new_n21549_1, new_n21550, new_n21551,
    new_n21552, new_n21553, new_n21554, new_n21555, new_n21556, new_n21557,
    new_n21558, new_n21559, new_n21560, new_n21561, new_n21562, new_n21563,
    new_n21564, new_n21565, new_n21566, new_n21567, new_n21568, new_n21569,
    new_n21570, new_n21571, new_n21572, new_n21573, new_n21574, new_n21575,
    new_n21576, new_n21577, new_n21578, new_n21579, new_n21580, new_n21581,
    new_n21582, new_n21583, new_n21584, new_n21585, new_n21586, new_n21587,
    new_n21588, new_n21589, new_n21590, new_n21591, new_n21592, new_n21593,
    new_n21594, new_n21595, new_n21596, new_n21597, new_n21598,
    new_n21599_1, new_n21600, new_n21601, new_n21602, new_n21603,
    new_n21604, new_n21605, new_n21606, new_n21607, new_n21608, new_n21610,
    new_n21611, new_n21612, new_n21613, new_n21614, new_n21615_1,
    new_n21616, new_n21617, new_n21618, new_n21619, new_n21620, new_n21621,
    new_n21622, new_n21623, new_n21624, new_n21625, new_n21626, new_n21627,
    new_n21628_1, new_n21629, new_n21630, new_n21631, new_n21632,
    new_n21633, new_n21634, new_n21635, new_n21636, new_n21637_1,
    new_n21638, new_n21639, new_n21640, new_n21641, new_n21642, new_n21643,
    new_n21644, new_n21645_1, new_n21646, new_n21647, new_n21648,
    new_n21649_1, new_n21650, new_n21651, new_n21652, new_n21653,
    new_n21654_1, new_n21655, new_n21656, new_n21657, new_n21658,
    new_n21659, new_n21660, new_n21661, new_n21662, new_n21663, new_n21664,
    new_n21665_1, new_n21667, new_n21668, new_n21669, new_n21670,
    new_n21671, new_n21672, new_n21673, new_n21674_1, new_n21675,
    new_n21676, new_n21677, new_n21678, new_n21679, new_n21680_1,
    new_n21681, new_n21682, new_n21683, new_n21684, new_n21685_1,
    new_n21686, new_n21687_1, new_n21688, new_n21689, new_n21690,
    new_n21691, new_n21692, new_n21693, new_n21694, new_n21695, new_n21696,
    new_n21697, new_n21698, new_n21699, new_n21700, new_n21701, new_n21702,
    new_n21703, new_n21704, new_n21705, new_n21706, new_n21707, new_n21708,
    new_n21709, new_n21710, new_n21711, new_n21712, new_n21713, new_n21714,
    new_n21715, new_n21716, new_n21717_1, new_n21718, new_n21719_1,
    new_n21720, new_n21721, new_n21722, new_n21723, new_n21724, new_n21725,
    new_n21726, new_n21727, new_n21728, new_n21729, new_n21730, new_n21731,
    new_n21732, new_n21733, new_n21734, new_n21735_1, new_n21736,
    new_n21737, new_n21738, new_n21739, new_n21740, new_n21741, new_n21742,
    new_n21743, new_n21744, new_n21745, new_n21746, new_n21747, new_n21748,
    new_n21749_1, new_n21750_1, new_n21751, new_n21752, new_n21753_1,
    new_n21754, new_n21755, new_n21759, new_n21762, new_n21763, new_n21764,
    new_n21765_1, new_n21766, new_n21767, new_n21768, new_n21769,
    new_n21770, new_n21771, new_n21772, new_n21773, new_n21774, new_n21775,
    new_n21776, new_n21777, new_n21778, new_n21779_1, new_n21780,
    new_n21781, new_n21782, new_n21783, new_n21784_1, new_n21785,
    new_n21786, new_n21787, new_n21788, new_n21789, new_n21790, new_n21791,
    new_n21792, new_n21793, new_n21794, new_n21795, new_n21796, new_n21797,
    new_n21798, new_n21799, new_n21800_1, new_n21801, new_n21802,
    new_n21803, new_n21804, new_n21805, new_n21806, new_n21807, new_n21808,
    new_n21809, new_n21810, new_n21811, new_n21812, new_n21813, new_n21814,
    new_n21815, new_n21816, new_n21817, new_n21818, new_n21819,
    new_n21820_1, new_n21821, new_n21822, new_n21823, new_n21824,
    new_n21825, new_n21826, new_n21827, new_n21828, new_n21829, new_n21830,
    new_n21831, new_n21832_1, new_n21833, new_n21834, new_n21835,
    new_n21836, new_n21837, new_n21838, new_n21839_1, new_n21840,
    new_n21841, new_n21842, new_n21843, new_n21844, new_n21845, new_n21846,
    new_n21847, new_n21848, new_n21849, new_n21850, new_n21851, new_n21854,
    new_n21855, new_n21856, new_n21857, new_n21858, new_n21859, new_n21860,
    new_n21861, new_n21862, new_n21863, new_n21864, new_n21865, new_n21866,
    new_n21867, new_n21868, new_n21869, new_n21870, new_n21871, new_n21872,
    new_n21873, new_n21874_1, new_n21875, new_n21876, new_n21877,
    new_n21878, new_n21879, new_n21880, new_n21881, new_n21882, new_n21883,
    new_n21884, new_n21885, new_n21888, new_n21889, new_n21890, new_n21891,
    new_n21892, new_n21893, new_n21894, new_n21895, new_n21896, new_n21897,
    new_n21898_1, new_n21899, new_n21900, new_n21901, new_n21902,
    new_n21903, new_n21904, new_n21905_1, new_n21906, new_n21907,
    new_n21908, new_n21909, new_n21910, new_n21911, new_n21913,
    new_n21915_1, new_n21917, new_n21920, new_n21921, new_n21922,
    new_n21923, new_n21924, new_n21925, new_n21926, new_n21927, new_n21928,
    new_n21929, new_n21930, new_n21931, new_n21932, new_n21933,
    new_n21934_1, new_n21935, new_n21936, new_n21937, new_n21938,
    new_n21939, new_n21940, new_n21941, new_n21942, new_n21943_1,
    new_n21944, new_n21945, new_n21946, new_n21947, new_n21948, new_n21949,
    new_n21950, new_n21951, new_n21952, new_n21953, new_n21954, new_n21955,
    new_n21956, new_n21957_1, new_n21958, new_n21959, new_n21960_1,
    new_n21961, new_n21962, new_n21963, new_n21964, new_n21965, new_n21966,
    new_n21967, new_n21968, new_n21969, new_n21970, new_n21971, new_n21972,
    new_n21973, new_n21974, new_n21975, new_n21976_1, new_n21977,
    new_n21978, new_n21979, new_n21980, new_n21981_1, new_n21982,
    new_n21983, new_n21984, new_n21985, new_n21986_1, new_n21987,
    new_n21988, new_n21989, new_n21990, new_n21991, new_n21992,
    new_n21993_1, new_n21994, new_n21995, new_n21996, new_n21997_1,
    new_n21998, new_n21999, new_n22000, new_n22001, new_n22002, new_n22003,
    new_n22004, new_n22005, new_n22006, new_n22007, new_n22008, new_n22009,
    new_n22010, new_n22011, new_n22012, new_n22013, new_n22014, new_n22015,
    new_n22016_1, new_n22017, new_n22018, new_n22019, new_n22020,
    new_n22021, new_n22022, new_n22023, new_n22024, new_n22025, new_n22026,
    new_n22027_1, new_n22028, new_n22029, new_n22030, new_n22031,
    new_n22032, new_n22033, new_n22034, new_n22035, new_n22036, new_n22037,
    new_n22038, new_n22039, new_n22040, new_n22041, new_n22042,
    new_n22043_1, new_n22044, new_n22045, new_n22046, new_n22047,
    new_n22048, new_n22049, new_n22050_1, new_n22051, new_n22052,
    new_n22053, new_n22054, new_n22055, new_n22056, new_n22059, new_n22061,
    new_n22062, new_n22063_1, new_n22064, new_n22065, new_n22066,
    new_n22067, new_n22068_1, new_n22069, new_n22070, new_n22071,
    new_n22072_1, new_n22073, new_n22074, new_n22075, new_n22076_1,
    new_n22077, new_n22078, new_n22079, new_n22080, new_n22081, new_n22082,
    new_n22083, new_n22084, new_n22085, new_n22086, new_n22087, new_n22088,
    new_n22089, new_n22090_1, new_n22091, new_n22092, new_n22094,
    new_n22098, new_n22101, new_n22102, new_n22103, new_n22104, new_n22105,
    new_n22106, new_n22107_1, new_n22108, new_n22109, new_n22110,
    new_n22111, new_n22112, new_n22113_1, new_n22114, new_n22115,
    new_n22116, new_n22117, new_n22118, new_n22119, new_n22120, new_n22121,
    new_n22122, new_n22123, new_n22124_1, new_n22125, new_n22126_1,
    new_n22127, new_n22128, new_n22129, new_n22130_1, new_n22131,
    new_n22132, new_n22133, new_n22134, new_n22135, new_n22136, new_n22137,
    new_n22138, new_n22139, new_n22140, new_n22141, new_n22142, new_n22143,
    new_n22144_1, new_n22145, new_n22146, new_n22147, new_n22148,
    new_n22149, new_n22150_1, new_n22151, new_n22152, new_n22153,
    new_n22154, new_n22155, new_n22156, new_n22157_1, new_n22158,
    new_n22159, new_n22160, new_n22161, new_n22162, new_n22163, new_n22164,
    new_n22165, new_n22166, new_n22167, new_n22168, new_n22169, new_n22170,
    new_n22171, new_n22172, new_n22173_1, new_n22174, new_n22175,
    new_n22176, new_n22177, new_n22178, new_n22179, new_n22180, new_n22181,
    new_n22182, new_n22183, new_n22184, new_n22185, new_n22186, new_n22187,
    new_n22188, new_n22189, new_n22190, new_n22191, new_n22192, new_n22193,
    new_n22194, new_n22195, new_n22196, new_n22197, new_n22198_1,
    new_n22199, new_n22200, new_n22201_1, new_n22204, new_n22205,
    new_n22206, new_n22207, new_n22208, new_n22209, new_n22210, new_n22211,
    new_n22212, new_n22213_1, new_n22214, new_n22215, new_n22216,
    new_n22217, new_n22218, new_n22219, new_n22220, new_n22221, new_n22222,
    new_n22223, new_n22224, new_n22225, new_n22226, new_n22227, new_n22228,
    new_n22229, new_n22230, new_n22231, new_n22232, new_n22233, new_n22234,
    new_n22235, new_n22236, new_n22237, new_n22238, new_n22239, new_n22240,
    new_n22241, new_n22242, new_n22243, new_n22244, new_n22245, new_n22246,
    new_n22247, new_n22248, new_n22249, new_n22250, new_n22251, new_n22252,
    new_n22253_1, new_n22254, new_n22255, new_n22256, new_n22257,
    new_n22258, new_n22259, new_n22260, new_n22261, new_n22262, new_n22263,
    new_n22264, new_n22265, new_n22266, new_n22267, new_n22268, new_n22269,
    new_n22270_1, new_n22271, new_n22272, new_n22273, new_n22274_1,
    new_n22275, new_n22276, new_n22277, new_n22278, new_n22279, new_n22280,
    new_n22281, new_n22282, new_n22283_1, new_n22284, new_n22285,
    new_n22286, new_n22287, new_n22288, new_n22289, new_n22290_1,
    new_n22291, new_n22292, new_n22293, new_n22294, new_n22295, new_n22296,
    new_n22297, new_n22298, new_n22299, new_n22300, new_n22301, new_n22302,
    new_n22303, new_n22304, new_n22305, new_n22306, new_n22307,
    new_n22309_1, new_n22310, new_n22311_1, new_n22312, new_n22313,
    new_n22314, new_n22315, new_n22316, new_n22317_1, new_n22318,
    new_n22319, new_n22320, new_n22321, new_n22322, new_n22323, new_n22324,
    new_n22325, new_n22326, new_n22327, new_n22328, new_n22329, new_n22330,
    new_n22331, new_n22332_1, new_n22333, new_n22334, new_n22335_1,
    new_n22336, new_n22337, new_n22338, new_n22339, new_n22340,
    new_n22341_1, new_n22342, new_n22343, new_n22344, new_n22345,
    new_n22346, new_n22347, new_n22348, new_n22349, new_n22350, new_n22351,
    new_n22352, new_n22353_1, new_n22354, new_n22355, new_n22356,
    new_n22357, new_n22358_1, new_n22359_1, new_n22360, new_n22361,
    new_n22362, new_n22363, new_n22364, new_n22365, new_n22366, new_n22367,
    new_n22368, new_n22370, new_n22371, new_n22372, new_n22373, new_n22374,
    new_n22375, new_n22376, new_n22377, new_n22378, new_n22379_1,
    new_n22380, new_n22381, new_n22382, new_n22383, new_n22384, new_n22385,
    new_n22386, new_n22387, new_n22388, new_n22389, new_n22390, new_n22391,
    new_n22392, new_n22393, new_n22394, new_n22395, new_n22396, new_n22397,
    new_n22398, new_n22399, new_n22400, new_n22401, new_n22402, new_n22403,
    new_n22404, new_n22405, new_n22406, new_n22407, new_n22408, new_n22409,
    new_n22410, new_n22411, new_n22412, new_n22413, new_n22414, new_n22415,
    new_n22416, new_n22417, new_n22418, new_n22420, new_n22424, new_n22425,
    new_n22426, new_n22427, new_n22428, new_n22429, new_n22430, new_n22431,
    new_n22432, new_n22433_1, new_n22434, new_n22435, new_n22436,
    new_n22437, new_n22438, new_n22439, new_n22440, new_n22441,
    new_n22442_1, new_n22445, new_n22447, new_n22449, new_n22450,
    new_n22451, new_n22452, new_n22453, new_n22454, new_n22455, new_n22456,
    new_n22457, new_n22458, new_n22459, new_n22460, new_n22461, new_n22462,
    new_n22463, new_n22464, new_n22465, new_n22466, new_n22467_1,
    new_n22468, new_n22469, new_n22470_1, new_n22471, new_n22472,
    new_n22473, new_n22474, new_n22475, new_n22476, new_n22477, new_n22478,
    new_n22479, new_n22480, new_n22481, new_n22482, new_n22483,
    new_n22484_1, new_n22485, new_n22486, new_n22487, new_n22488,
    new_n22489_1, new_n22490, new_n22491, new_n22492_1, new_n22493,
    new_n22494_1, new_n22495, new_n22496, new_n22497, new_n22498,
    new_n22499, new_n22500, new_n22501, new_n22502, new_n22503, new_n22504,
    new_n22505, new_n22506, new_n22507, new_n22508, new_n22509, new_n22510,
    new_n22511, new_n22512, new_n22513, new_n22515, new_n22516, new_n22517,
    new_n22518, new_n22519, new_n22520, new_n22521, new_n22522, new_n22523,
    new_n22524, new_n22525, new_n22526, new_n22527, new_n22528, new_n22529,
    new_n22530, new_n22532, new_n22533_1, new_n22534, new_n22535,
    new_n22536, new_n22537, new_n22538, new_n22539, new_n22540, new_n22541,
    new_n22542, new_n22543, new_n22544, new_n22545, new_n22546, new_n22547,
    new_n22548, new_n22549, new_n22550, new_n22554_1, new_n22555,
    new_n22556, new_n22557, new_n22558, new_n22559, new_n22560, new_n22561,
    new_n22562, new_n22563, new_n22564, new_n22565, new_n22566, new_n22567,
    new_n22568, new_n22569, new_n22570, new_n22571, new_n22572, new_n22573,
    new_n22575, new_n22576, new_n22577, new_n22578, new_n22579, new_n22580,
    new_n22581, new_n22582, new_n22583, new_n22584_1, new_n22585,
    new_n22586, new_n22587, new_n22588_1, new_n22589_1, new_n22590,
    new_n22591_1, new_n22592, new_n22593, new_n22594, new_n22595,
    new_n22596, new_n22597_1, new_n22598, new_n22599, new_n22600,
    new_n22601, new_n22602, new_n22603, new_n22604, new_n22605, new_n22606,
    new_n22607, new_n22608, new_n22609, new_n22610, new_n22611, new_n22612,
    new_n22613, new_n22614, new_n22615, new_n22616, new_n22617, new_n22618,
    new_n22619_1, new_n22620_1, new_n22621, new_n22622, new_n22623_1,
    new_n22624, new_n22625, new_n22626_1, new_n22627, new_n22628,
    new_n22629, new_n22630, new_n22631_1, new_n22632, new_n22633,
    new_n22634, new_n22635, new_n22636, new_n22637, new_n22638, new_n22639,
    new_n22640, new_n22641, new_n22642, new_n22643, new_n22644, new_n22645,
    new_n22646, new_n22647, new_n22648, new_n22649, new_n22650, new_n22652,
    new_n22653, new_n22654, new_n22655, new_n22656, new_n22657, new_n22658,
    new_n22659, new_n22660_1, new_n22661, new_n22662, new_n22663,
    new_n22664, new_n22666, new_n22667, new_n22668, new_n22669, new_n22670,
    new_n22671, new_n22672, new_n22673, new_n22674, new_n22675, new_n22676,
    new_n22677, new_n22678, new_n22679, new_n22680, new_n22681, new_n22682,
    new_n22683, new_n22684, new_n22685, new_n22686, new_n22687, new_n22688,
    new_n22689, new_n22690, new_n22691, new_n22692, new_n22693, new_n22694,
    new_n22695, new_n22696, new_n22697_1, new_n22698, new_n22699,
    new_n22700, new_n22701, new_n22702, new_n22703, new_n22704, new_n22705,
    new_n22706, new_n22707, new_n22708, new_n22709, new_n22710, new_n22711,
    new_n22712, new_n22713, new_n22714_1, new_n22715, new_n22716,
    new_n22717, new_n22718, new_n22719, new_n22720, new_n22721, new_n22722,
    new_n22723, new_n22724, new_n22725, new_n22726, new_n22727, new_n22728,
    new_n22729, new_n22730, new_n22731, new_n22732, new_n22733, new_n22734,
    new_n22735, new_n22736, new_n22737, new_n22738, new_n22739, new_n22740,
    new_n22741, new_n22742, new_n22743, new_n22744, new_n22745, new_n22746,
    new_n22747, new_n22748, new_n22749, new_n22750, new_n22751, new_n22752,
    new_n22753, new_n22754, new_n22755, new_n22756, new_n22757, new_n22758,
    new_n22759, new_n22760, new_n22761_1, new_n22762, new_n22763,
    new_n22764_1, new_n22765, new_n22766, new_n22767, new_n22768,
    new_n22769, new_n22770, new_n22771, new_n22772, new_n22773, new_n22774,
    new_n22775, new_n22776, new_n22777, new_n22778, new_n22779_1,
    new_n22780, new_n22781, new_n22782, new_n22783, new_n22784, new_n22785,
    new_n22786, new_n22787_1, new_n22788, new_n22789, new_n22790,
    new_n22791, new_n22792, new_n22793_1, new_n22794, new_n22795,
    new_n22796, new_n22797, new_n22798, new_n22799, new_n22800, new_n22801,
    new_n22802, new_n22803, new_n22804, new_n22805, new_n22806, new_n22807,
    new_n22808, new_n22809, new_n22810, new_n22811, new_n22812, new_n22813,
    new_n22814, new_n22815, new_n22816, new_n22817, new_n22818,
    new_n22819_1, new_n22820, new_n22821, new_n22822, new_n22823,
    new_n22824, new_n22825, new_n22826, new_n22827, new_n22828, new_n22829,
    new_n22830, new_n22831, new_n22832, new_n22833, new_n22834, new_n22835,
    new_n22836, new_n22837, new_n22838, new_n22839, new_n22840, new_n22841,
    new_n22842, new_n22843_1, new_n22844, new_n22845, new_n22846,
    new_n22847, new_n22848, new_n22849, new_n22850, new_n22851, new_n22852,
    new_n22853, new_n22854, new_n22855, new_n22856, new_n22857,
    new_n22858_1, new_n22859, new_n22860, new_n22861, new_n22862,
    new_n22863, new_n22864, new_n22865, new_n22866, new_n22867, new_n22868,
    new_n22869, new_n22870_1, new_n22871_1, new_n22872, new_n22873,
    new_n22874, new_n22875, new_n22876, new_n22877, new_n22878,
    new_n22879_1, new_n22880, new_n22881, new_n22882, new_n22883,
    new_n22884, new_n22885, new_n22886, new_n22887, new_n22888, new_n22889,
    new_n22890, new_n22891_1, new_n22892, new_n22893, new_n22894,
    new_n22895, new_n22896, new_n22897_1, new_n22898, new_n22899,
    new_n22900, new_n22901, new_n22902, new_n22903_1, new_n22904,
    new_n22905, new_n22906, new_n22907_1, new_n22908, new_n22909,
    new_n22910_1, new_n22911, new_n22912, new_n22913, new_n22914_1,
    new_n22915, new_n22916, new_n22917, new_n22918_1, new_n22921,
    new_n22922, new_n22923, new_n22924, new_n22925, new_n22926, new_n22927,
    new_n22928, new_n22929, new_n22930, new_n22931, new_n22932, new_n22933,
    new_n22934, new_n22935, new_n22936, new_n22937, new_n22938,
    new_n22939_1, new_n22940, new_n22941, new_n22942, new_n22943,
    new_n22944, new_n22945, new_n22946, new_n22947, new_n22948, new_n22949,
    new_n22950, new_n22951, new_n22952, new_n22953, new_n22954, new_n22955,
    new_n22956, new_n22957, new_n22958, new_n22959, new_n22961, new_n22962,
    new_n22963, new_n22964, new_n22965, new_n22966, new_n22967, new_n22968,
    new_n22969, new_n22970, new_n22971, new_n22972, new_n22973, new_n22974,
    new_n22975, new_n22976, new_n22977, new_n22979, new_n22981, new_n22982,
    new_n22983, new_n22984, new_n22985, new_n22986, new_n22988, new_n22992,
    new_n22993, new_n22994, new_n22995, new_n22996, new_n22997,
    new_n22998_1, new_n22999, new_n23000, new_n23001, new_n23002,
    new_n23003, new_n23004, new_n23005, new_n23006_1, new_n23007_1,
    new_n23008, new_n23009_1, new_n23010, new_n23011, new_n23012,
    new_n23013, new_n23014_1, new_n23015, new_n23016, new_n23017,
    new_n23018, new_n23019, new_n23020, new_n23021, new_n23022, new_n23023,
    new_n23024, new_n23025, new_n23026, new_n23027, new_n23028, new_n23029,
    new_n23030, new_n23031, new_n23032, new_n23033, new_n23034,
    new_n23035_1, new_n23036, new_n23037, new_n23038, new_n23039_1,
    new_n23040, new_n23041, new_n23042, new_n23043, new_n23044, new_n23045,
    new_n23046, new_n23047_1, new_n23048, new_n23049, new_n23050,
    new_n23051, new_n23052, new_n23053, new_n23054, new_n23055, new_n23056,
    new_n23057, new_n23058_1, new_n23059, new_n23060, new_n23061,
    new_n23062, new_n23063, new_n23064, new_n23065_1, new_n23066_1,
    new_n23067_1, new_n23068_1, new_n23069, new_n23070, new_n23071,
    new_n23072, new_n23073, new_n23074, new_n23075, new_n23076, new_n23077,
    new_n23078, new_n23079, new_n23080, new_n23081, new_n23082, new_n23083,
    new_n23084, new_n23085, new_n23086, new_n23087, new_n23088, new_n23089,
    new_n23090, new_n23091, new_n23092, new_n23093, new_n23094, new_n23095,
    new_n23096, new_n23097, new_n23098, new_n23099, new_n23100, new_n23101,
    new_n23102, new_n23103, new_n23104, new_n23105, new_n23106, new_n23107,
    new_n23108, new_n23109, new_n23110, new_n23111, new_n23113, new_n23115,
    new_n23116, new_n23117, new_n23118, new_n23119, new_n23120_1,
    new_n23121, new_n23122, new_n23123, new_n23124, new_n23125, new_n23126,
    new_n23127, new_n23128, new_n23129, new_n23130, new_n23131, new_n23132,
    new_n23133, new_n23135, new_n23136, new_n23137, new_n23138, new_n23139,
    new_n23140, new_n23141, new_n23142, new_n23143, new_n23144, new_n23145,
    new_n23146_1, new_n23147, new_n23148, new_n23149, new_n23150,
    new_n23151, new_n23152, new_n23153, new_n23154, new_n23155, new_n23156,
    new_n23157, new_n23158, new_n23159, new_n23160_1, new_n23161,
    new_n23162, new_n23163, new_n23164, new_n23165, new_n23166_1,
    new_n23167, new_n23168, new_n23169, new_n23170, new_n23171, new_n23172,
    new_n23173, new_n23174, new_n23175, new_n23176, new_n23177, new_n23178,
    new_n23179, new_n23180, new_n23181, new_n23182, new_n23183, new_n23184,
    new_n23185, new_n23186, new_n23187, new_n23188, new_n23189, new_n23190,
    new_n23191, new_n23192, new_n23193, new_n23195, new_n23197, new_n23198,
    new_n23199, new_n23200_1, new_n23201, new_n23202, new_n23203,
    new_n23204, new_n23205, new_n23206, new_n23207, new_n23208, new_n23209,
    new_n23210, new_n23211, new_n23212, new_n23213, new_n23214, new_n23215,
    new_n23216, new_n23217, new_n23218, new_n23219, new_n23220, new_n23221,
    new_n23222, new_n23223, new_n23224, new_n23225, new_n23226, new_n23227,
    new_n23228, new_n23229, new_n23230, new_n23231, new_n23232, new_n23233,
    new_n23234, new_n23235, new_n23236, new_n23238_1, new_n23239,
    new_n23240, new_n23241, new_n23242, new_n23243, new_n23244, new_n23245,
    new_n23246, new_n23247_1, new_n23248_1, new_n23249, new_n23250_1,
    new_n23251, new_n23252, new_n23253, new_n23254, new_n23255, new_n23256,
    new_n23257, new_n23258, new_n23259, new_n23260, new_n23261, new_n23262,
    new_n23263, new_n23264, new_n23265, new_n23266, new_n23267, new_n23268,
    new_n23269, new_n23270_1, new_n23271, new_n23272_1, new_n23273,
    new_n23274, new_n23275, new_n23276, new_n23277, new_n23278, new_n23279,
    new_n23281, new_n23283, new_n23285, new_n23286, new_n23287,
    new_n23289_1, new_n23290, new_n23291, new_n23292, new_n23293,
    new_n23294, new_n23295, new_n23296, new_n23297, new_n23298, new_n23299,
    new_n23300, new_n23301, new_n23302, new_n23303, new_n23304_1,
    new_n23305_1, new_n23306, new_n23307, new_n23308, new_n23309,
    new_n23310, new_n23312, new_n23315, new_n23317, new_n23318, new_n23319,
    new_n23320, new_n23321, new_n23322, new_n23323, new_n23324, new_n23325,
    new_n23326, new_n23327, new_n23328, new_n23329, new_n23330, new_n23331,
    new_n23332, new_n23333_1, new_n23334, new_n23335, new_n23336,
    new_n23337, new_n23338, new_n23339, new_n23340, new_n23341_1,
    new_n23342_1, new_n23343, new_n23344, new_n23345, new_n23346,
    new_n23347, new_n23348, new_n23349, new_n23350, new_n23351, new_n23352,
    new_n23353, new_n23354, new_n23355_1, new_n23356, new_n23357,
    new_n23358, new_n23359, new_n23360, new_n23361, new_n23362, new_n23363,
    new_n23364, new_n23365, new_n23366, new_n23367, new_n23368,
    new_n23369_1, new_n23370, new_n23371_1, new_n23372, new_n23373,
    new_n23374, new_n23375, new_n23376, new_n23377, new_n23378, new_n23379,
    new_n23380, new_n23381, new_n23382, new_n23383, new_n23384, new_n23385,
    new_n23386, new_n23387, new_n23388, new_n23389, new_n23390, new_n23391,
    new_n23392, new_n23393, new_n23394, new_n23395, new_n23396, new_n23397,
    new_n23398, new_n23399, new_n23400, new_n23401_1, new_n23402,
    new_n23403, new_n23404, new_n23405, new_n23406, new_n23407, new_n23408,
    new_n23409, new_n23410, new_n23411, new_n23412, new_n23413,
    new_n23414_1, new_n23415, new_n23416, new_n23417, new_n23418,
    new_n23419, new_n23420, new_n23421, new_n23423, new_n23426, new_n23428,
    new_n23430_1, new_n23431, new_n23432, new_n23433_1, new_n23434_1,
    new_n23435, new_n23436, new_n23437, new_n23438, new_n23439, new_n23440,
    new_n23441, new_n23442, new_n23443, new_n23444, new_n23445, new_n23446,
    new_n23447, new_n23448, new_n23449, new_n23450_1, new_n23451,
    new_n23452, new_n23453, new_n23454, new_n23455, new_n23457, new_n23458,
    new_n23459, new_n23460, new_n23461, new_n23462, new_n23463_1,
    new_n23464, new_n23465, new_n23466, new_n23467, new_n23468, new_n23469,
    new_n23470, new_n23471_1, new_n23472, new_n23473, new_n23474,
    new_n23475, new_n23476, new_n23477, new_n23478, new_n23479,
    new_n23480_1, new_n23481, new_n23482, new_n23483, new_n23484,
    new_n23485, new_n23486, new_n23487, new_n23488, new_n23489, new_n23490,
    new_n23491, new_n23492, new_n23493_1, new_n23494, new_n23495,
    new_n23496, new_n23497, new_n23498, new_n23499, new_n23500, new_n23501,
    new_n23502, new_n23503, new_n23504, new_n23505, new_n23506, new_n23507,
    new_n23508, new_n23509, new_n23510, new_n23511, new_n23512,
    new_n23513_1, new_n23514, new_n23515, new_n23516, new_n23517,
    new_n23518, new_n23519, new_n23520, new_n23521, new_n23522, new_n23523,
    new_n23524, new_n23525, new_n23526, new_n23527, new_n23528,
    new_n23529_1, new_n23530, new_n23531, new_n23532, new_n23533,
    new_n23534, new_n23535, new_n23536, new_n23537, new_n23538, new_n23539,
    new_n23540, new_n23541_1, new_n23542, new_n23543, new_n23544,
    new_n23545, new_n23546_1, new_n23547, new_n23552, new_n23553,
    new_n23554, new_n23555, new_n23556, new_n23557, new_n23558, new_n23559,
    new_n23560, new_n23561, new_n23562, new_n23563, new_n23564, new_n23565,
    new_n23566, new_n23567, new_n23568, new_n23569, new_n23570, new_n23571,
    new_n23572, new_n23573, new_n23574, new_n23575, new_n23576, new_n23577,
    new_n23578, new_n23579, new_n23580, new_n23581, new_n23582, new_n23583,
    new_n23584, new_n23585_1, new_n23586_1, new_n23587, new_n23588_1,
    new_n23589, new_n23590, new_n23591, new_n23592, new_n23593, new_n23594,
    new_n23595, new_n23596, new_n23597, new_n23598, new_n23599, new_n23600,
    new_n23601, new_n23602, new_n23603, new_n23604, new_n23605, new_n23606,
    new_n23607, new_n23608, new_n23609, new_n23610, new_n23611, new_n23612,
    new_n23613, new_n23614, new_n23615, new_n23616, new_n23617, new_n23618,
    new_n23619_1, new_n23620, new_n23621, new_n23622, new_n23623,
    new_n23624_1, new_n23625, new_n23626, new_n23627, new_n23628_1,
    new_n23629, new_n23630, new_n23631, new_n23632, new_n23633, new_n23634,
    new_n23635, new_n23636, new_n23637_1, new_n23638, new_n23639,
    new_n23640, new_n23641, new_n23642, new_n23643, new_n23644, new_n23645,
    new_n23646, new_n23647, new_n23648, new_n23649, new_n23650, new_n23651,
    new_n23652, new_n23653, new_n23654, new_n23655, new_n23658, new_n23659,
    new_n23660, new_n23661, new_n23662, new_n23663_1, new_n23664,
    new_n23665, new_n23666, new_n23667, new_n23668, new_n23669_1,
    new_n23670, new_n23671, new_n23672, new_n23673, new_n23674, new_n23675,
    new_n23676, new_n23677, new_n23678, new_n23679, new_n23680, new_n23681,
    new_n23682, new_n23683, new_n23684_1, new_n23685, new_n23686,
    new_n23687, new_n23688, new_n23689, new_n23690_1, new_n23691,
    new_n23692, new_n23693, new_n23694, new_n23695, new_n23696,
    new_n23697_1, new_n23698, new_n23699, new_n23700, new_n23701,
    new_n23702, new_n23703, new_n23704, new_n23705, new_n23706, new_n23707,
    new_n23708, new_n23709, new_n23710, new_n23711, new_n23712, new_n23713,
    new_n23714_1, new_n23715, new_n23716, new_n23717_1, new_n23718,
    new_n23719_1, new_n23720, new_n23721, new_n23722, new_n23723,
    new_n23724, new_n23725, new_n23726, new_n23727, new_n23728, new_n23729,
    new_n23730, new_n23731, new_n23733, new_n23735, new_n23736, new_n23737,
    new_n23738, new_n23739, new_n23740, new_n23741, new_n23742, new_n23743,
    new_n23744, new_n23745, new_n23746, new_n23747, new_n23748_1,
    new_n23749, new_n23750, new_n23751, new_n23752, new_n23753, new_n23754,
    new_n23755_1, new_n23756, new_n23757, new_n23758, new_n23760,
    new_n23761, new_n23762, new_n23763, new_n23764, new_n23765, new_n23766,
    new_n23767, new_n23768, new_n23769, new_n23770, new_n23771, new_n23772,
    new_n23773, new_n23774, new_n23775_1, new_n23776, new_n23777,
    new_n23778, new_n23779, new_n23780, new_n23782, new_n23783, new_n23784,
    new_n23785, new_n23786, new_n23787, new_n23788, new_n23789, new_n23790,
    new_n23791, new_n23792, new_n23793, new_n23794, new_n23795, new_n23796,
    new_n23797, new_n23798, new_n23799, new_n23800, new_n23801, new_n23802,
    new_n23803, new_n23804, new_n23805, new_n23806, new_n23807, new_n23808,
    new_n23809, new_n23810, new_n23811, new_n23812, new_n23813, new_n23814,
    new_n23815, new_n23816, new_n23817, new_n23818, new_n23819, new_n23820,
    new_n23821, new_n23822, new_n23823, new_n23824, new_n23825, new_n23826,
    new_n23827, new_n23828, new_n23829, new_n23830, new_n23831_1,
    new_n23832, new_n23833, new_n23834, new_n23835, new_n23836, new_n23839,
    new_n23841, new_n23842_1, new_n23843, new_n23844, new_n23845,
    new_n23846, new_n23847, new_n23848, new_n23849_1, new_n23850,
    new_n23851, new_n23852, new_n23853, new_n23854, new_n23855,
    new_n23856_1, new_n23857, new_n23858, new_n23859, new_n23860,
    new_n23861, new_n23862, new_n23863, new_n23864, new_n23865, new_n23866,
    new_n23867, new_n23868, new_n23869, new_n23870, new_n23871, new_n23872,
    new_n23873, new_n23874, new_n23875, new_n23876, new_n23877, new_n23878,
    new_n23879, new_n23880, new_n23881, new_n23882, new_n23883_1,
    new_n23884, new_n23885, new_n23886, new_n23887, new_n23888_1,
    new_n23889, new_n23890, new_n23891, new_n23892, new_n23893, new_n23894,
    new_n23895_1, new_n23896, new_n23897, new_n23898, new_n23899_1,
    new_n23900, new_n23901, new_n23903_1, new_n23904, new_n23905,
    new_n23906, new_n23907, new_n23908, new_n23909, new_n23910, new_n23911,
    new_n23912_1, new_n23913_1, new_n23914, new_n23915, new_n23916,
    new_n23917, new_n23918, new_n23919, new_n23920, new_n23921, new_n23922,
    new_n23923_1, new_n23924_1, new_n23925, new_n23926, new_n23927,
    new_n23928, new_n23929, new_n23930, new_n23931, new_n23932, new_n23933,
    new_n23934, new_n23935_1, new_n23937, new_n23938, new_n23939,
    new_n23940, new_n23941, new_n23942_1, new_n23943, new_n23944,
    new_n23945, new_n23946, new_n23947, new_n23948, new_n23949, new_n23950,
    new_n23951, new_n23952, new_n23953, new_n23954_1, new_n23955,
    new_n23956, new_n23958_1, new_n23961, new_n23963, new_n23964,
    new_n23965, new_n23966, new_n23967, new_n23968, new_n23969, new_n23970,
    new_n23971, new_n23972, new_n23973, new_n23974_1, new_n23977,
    new_n23978, new_n23979, new_n23980, new_n23981, new_n23982, new_n23983,
    new_n23984, new_n23985, new_n23986_1, new_n23987, new_n23988,
    new_n23989, new_n23990, new_n23991, new_n23992, new_n23993, new_n23994,
    new_n23995, new_n23996, new_n23997, new_n23998, new_n23999, new_n24000,
    new_n24001, new_n24002_1, new_n24003, new_n24004_1, new_n24005,
    new_n24006, new_n24007, new_n24008, new_n24009, new_n24010, new_n24011,
    new_n24012, new_n24013, new_n24014, new_n24015, new_n24016, new_n24017,
    new_n24018, new_n24019, new_n24020, new_n24021, new_n24022, new_n24023,
    new_n24024, new_n24025, new_n24026, new_n24027, new_n24028, new_n24029,
    new_n24030, new_n24031, new_n24032_1, new_n24033, new_n24034,
    new_n24035, new_n24036, new_n24037, new_n24038, new_n24039_1,
    new_n24040, new_n24041, new_n24042, new_n24043, new_n24044, new_n24045,
    new_n24046, new_n24047, new_n24048_1, new_n24049, new_n24050,
    new_n24051, new_n24052_1, new_n24053, new_n24054, new_n24055,
    new_n24056, new_n24057, new_n24058, new_n24059, new_n24060, new_n24061,
    new_n24062, new_n24064, new_n24068, new_n24069, new_n24070, new_n24071,
    new_n24072, new_n24073, new_n24074, new_n24075, new_n24076, new_n24077,
    new_n24078, new_n24079, new_n24080, new_n24081, new_n24082, new_n24083,
    new_n24084, new_n24085_1, new_n24086, new_n24087, new_n24088,
    new_n24089, new_n24090, new_n24091, new_n24092_1, new_n24093_1,
    new_n24096_1, new_n24098, new_n24099, new_n24100, new_n24101,
    new_n24102, new_n24103, new_n24104, new_n24105_1, new_n24106,
    new_n24107, new_n24108, new_n24109, new_n24110, new_n24111, new_n24112,
    new_n24113, new_n24114, new_n24115, new_n24116, new_n24117, new_n24118,
    new_n24119_1, new_n24120, new_n24121, new_n24122, new_n24123,
    new_n24124, new_n24125, new_n24126, new_n24127, new_n24128,
    new_n24129_1, new_n24130, new_n24131, new_n24132, new_n24133_1,
    new_n24134, new_n24135, new_n24136, new_n24137, new_n24138, new_n24139,
    new_n24140, new_n24141_1, new_n24142, new_n24143, new_n24144,
    new_n24145_1, new_n24146_1, new_n24147, new_n24148, new_n24149,
    new_n24150_1, new_n24151, new_n24152, new_n24153, new_n24154,
    new_n24155_1, new_n24156, new_n24157, new_n24158, new_n24159,
    new_n24160_1, new_n24161, new_n24162, new_n24163, new_n24164,
    new_n24165, new_n24166, new_n24167_1, new_n24168, new_n24169,
    new_n24170_1, new_n24171, new_n24172_1, new_n24173, new_n24174,
    new_n24175, new_n24176, new_n24177_1, new_n24178, new_n24179,
    new_n24180, new_n24181, new_n24182, new_n24183, new_n24184, new_n24185,
    new_n24186, new_n24187, new_n24188, new_n24189, new_n24190, new_n24191,
    new_n24192, new_n24193, new_n24194, new_n24195, new_n24196_1,
    new_n24197, new_n24198, new_n24199, new_n24200, new_n24201, new_n24202,
    new_n24203, new_n24204, new_n24205, new_n24206, new_n24207, new_n24208,
    new_n24209, new_n24210, new_n24211, new_n24212, new_n24213, new_n24214,
    new_n24215, new_n24216, new_n24217, new_n24218, new_n24219, new_n24220,
    new_n24221, new_n24222, new_n24224, new_n24226, new_n24228_1,
    new_n24231, new_n24234, new_n24235, new_n24236, new_n24237, new_n24238,
    new_n24239, new_n24240, new_n24241, new_n24242, new_n24243, new_n24244,
    new_n24245, new_n24246, new_n24247, new_n24248, new_n24249, new_n24250,
    new_n24251, new_n24252, new_n24253, new_n24254, new_n24255, new_n24256,
    new_n24257, new_n24258_1, new_n24259, new_n24260_1, new_n24261,
    new_n24262, new_n24263, new_n24264, new_n24265, new_n24266, new_n24267,
    new_n24268, new_n24269, new_n24270, new_n24271, new_n24272, new_n24273,
    new_n24274, new_n24275, new_n24276, new_n24277, new_n24278_1,
    new_n24279, new_n24280, new_n24281, new_n24282, new_n24283, new_n24286,
    new_n24288, new_n24289_1, new_n24290, new_n24291, new_n24292,
    new_n24293, new_n24294, new_n24295, new_n24296, new_n24297_1,
    new_n24298, new_n24299, new_n24300, new_n24301, new_n24302, new_n24303,
    new_n24304, new_n24305, new_n24306, new_n24307_1, new_n24308,
    new_n24309, new_n24310, new_n24311, new_n24312, new_n24313, new_n24314,
    new_n24315, new_n24316, new_n24317, new_n24318, new_n24319_1,
    new_n24320, new_n24321, new_n24322, new_n24323_1, new_n24324,
    new_n24325, new_n24326, new_n24327_1, new_n24328, new_n24329,
    new_n24330, new_n24331, new_n24332, new_n24333, new_n24334, new_n24335,
    new_n24336, new_n24337, new_n24338, new_n24339, new_n24340, new_n24341,
    new_n24342_1, new_n24343, new_n24344, new_n24345_1, new_n24346,
    new_n24347_1, new_n24348, new_n24349, new_n24350, new_n24351,
    new_n24352, new_n24353, new_n24354, new_n24355, new_n24356, new_n24357,
    new_n24358, new_n24359, new_n24360, new_n24361, new_n24362, new_n24363,
    new_n24364, new_n24365, new_n24366, new_n24367, new_n24368, new_n24369,
    new_n24370, new_n24371, new_n24372, new_n24373_1, new_n24374_1,
    new_n24375, new_n24376, new_n24377, new_n24378, new_n24379, new_n24380,
    new_n24381, new_n24382, new_n24383, new_n24384, new_n24385, new_n24386,
    new_n24387, new_n24388, new_n24389, new_n24390, new_n24391, new_n24392,
    new_n24393, new_n24394, new_n24395, new_n24396, new_n24397, new_n24398,
    new_n24400, new_n24401, new_n24402, new_n24403, new_n24404, new_n24405,
    new_n24406_1, new_n24407, new_n24408, new_n24409, new_n24411,
    new_n24413, new_n24415_1, new_n24416, new_n24417, new_n24418,
    new_n24419, new_n24420, new_n24421_1, new_n24422, new_n24423,
    new_n24424, new_n24425, new_n24426, new_n24427, new_n24428, new_n24429,
    new_n24430, new_n24431_1, new_n24432, new_n24433, new_n24434,
    new_n24435, new_n24436, new_n24437, new_n24438, new_n24439, new_n24440,
    new_n24441, new_n24442, new_n24443, new_n24444, new_n24445, new_n24446,
    new_n24447, new_n24448, new_n24449, new_n24451, new_n24452, new_n24453,
    new_n24454, new_n24455, new_n24456, new_n24457, new_n24458, new_n24459,
    new_n24460, new_n24461, new_n24462, new_n24463, new_n24464, new_n24465,
    new_n24466, new_n24467, new_n24468, new_n24469, new_n24470, new_n24471,
    new_n24472_1, new_n24473, new_n24474, new_n24475, new_n24476_1,
    new_n24477, new_n24478, new_n24479, new_n24480, new_n24481, new_n24482,
    new_n24483_1, new_n24484, new_n24485_1, new_n24486, new_n24487,
    new_n24488, new_n24489, new_n24490, new_n24491, new_n24492, new_n24493,
    new_n24494, new_n24495, new_n24496, new_n24497, new_n24498, new_n24499,
    new_n24500, new_n24501_1, new_n24502, new_n24503, new_n24504,
    new_n24505, new_n24506, new_n24507, new_n24508, new_n24509, new_n24510,
    new_n24511, new_n24512_1, new_n24513, new_n24514, new_n24515,
    new_n24516, new_n24517, new_n24518, new_n24519, new_n24520, new_n24521,
    new_n24522, new_n24523, new_n24524, new_n24525, new_n24526, new_n24527,
    new_n24528, new_n24529, new_n24530, new_n24531, new_n24532, new_n24533,
    new_n24534, new_n24535, new_n24536, new_n24538, new_n24539, new_n24542,
    new_n24543, new_n24544, new_n24545, new_n24546, new_n24547, new_n24548,
    new_n24549, new_n24550, new_n24551, new_n24552, new_n24553, new_n24554,
    new_n24555, new_n24556, new_n24557, new_n24558_1, new_n24559,
    new_n24560, new_n24561, new_n24562, new_n24563, new_n24564, new_n24565,
    new_n24566, new_n24567, new_n24568, new_n24569, new_n24570, new_n24571,
    new_n24572, new_n24573, new_n24574, new_n24575, new_n24576_1,
    new_n24577, new_n24578, new_n24579_1, new_n24580, new_n24581,
    new_n24582, new_n24583, new_n24584, new_n24585, new_n24586, new_n24587,
    new_n24588, new_n24589, new_n24590, new_n24591, new_n24592, new_n24593,
    new_n24594, new_n24595, new_n24596, new_n24597, new_n24598, new_n24599,
    new_n24600, new_n24601, new_n24602_1, new_n24603, new_n24604_1,
    new_n24605, new_n24606, new_n24607, new_n24608, new_n24609, new_n24610,
    new_n24611, new_n24612, new_n24613, new_n24614, new_n24615, new_n24616,
    new_n24617, new_n24618_1, new_n24619, new_n24620_1, new_n24621,
    new_n24622, new_n24623, new_n24624, new_n24625, new_n24626_1,
    new_n24627, new_n24628, new_n24629_1, new_n24630, new_n24631,
    new_n24632, new_n24633, new_n24634, new_n24635, new_n24636_1,
    new_n24637, new_n24638_1, new_n24639, new_n24640, new_n24641,
    new_n24642, new_n24643, new_n24644, new_n24645, new_n24646, new_n24647,
    new_n24648, new_n24649, new_n24650, new_n24651, new_n24652, new_n24653,
    new_n24654, new_n24655, new_n24656, new_n24657, new_n24658, new_n24659,
    new_n24660, new_n24661, new_n24662, new_n24663, new_n24664, new_n24665,
    new_n24666, new_n24667, new_n24668, new_n24669, new_n24670, new_n24671,
    new_n24672, new_n24673, new_n24674, new_n24675, new_n24676, new_n24677,
    new_n24678, new_n24679, new_n24680, new_n24681, new_n24682, new_n24683,
    new_n24684, new_n24685, new_n24686, new_n24687, new_n24689, new_n24691,
    new_n24692, new_n24693, new_n24694, new_n24695, new_n24696, new_n24697,
    new_n24698, new_n24699, new_n24700, new_n24701, new_n24702, new_n24703,
    new_n24704, new_n24705, new_n24706, new_n24707, new_n24708, new_n24709,
    new_n24710, new_n24711, new_n24712, new_n24713, new_n24714,
    new_n24715_1, new_n24716, new_n24717, new_n24718, new_n24719,
    new_n24720, new_n24721, new_n24722, new_n24723_1, new_n24724,
    new_n24725, new_n24726, new_n24727, new_n24728, new_n24729, new_n24730,
    new_n24731, new_n24732_1, new_n24733, new_n24734, new_n24735,
    new_n24736, new_n24737, new_n24738, new_n24739, new_n24740, new_n24741,
    new_n24742, new_n24743, new_n24744, new_n24745, new_n24746, new_n24747,
    new_n24748, new_n24749_1, new_n24750, new_n24751, new_n24752,
    new_n24753, new_n24754, new_n24755, new_n24756, new_n24757,
    new_n24758_1, new_n24759, new_n24760, new_n24761, new_n24762,
    new_n24763, new_n24764, new_n24765, new_n24766, new_n24767,
    new_n24768_1, new_n24769, new_n24770, new_n24771, new_n24772,
    new_n24774, new_n24776, new_n24778, new_n24780, new_n24782,
    new_n24784_1, new_n24785, new_n24786_1, new_n24788, new_n24791,
    new_n24792, new_n24793, new_n24794, new_n24795, new_n24796, new_n24797,
    new_n24798, new_n24799, new_n24800, new_n24801, new_n24802, new_n24803,
    new_n24804, new_n24805, new_n24806, new_n24807_1, new_n24808,
    new_n24809, new_n24810, new_n24811, new_n24812, new_n24813, new_n24814,
    new_n24815, new_n24816, new_n24817, new_n24818, new_n24819, new_n24820,
    new_n24821, new_n24822, new_n24823, new_n24824, new_n24825,
    new_n24826_1, new_n24827, new_n24828, new_n24829, new_n24830,
    new_n24831, new_n24832, new_n24833, new_n24834, new_n24835, new_n24836,
    new_n24837, new_n24838, new_n24839, new_n24840_1, new_n24841_1,
    new_n24842, new_n24843, new_n24844, new_n24845, new_n24846, new_n24847,
    new_n24848, new_n24849, new_n24850, new_n24851, new_n24852,
    new_n24853_1, new_n24854, new_n24855, new_n24856, new_n24857_1,
    new_n24858, new_n24859, new_n24860, new_n24861, new_n24862, new_n24863,
    new_n24864, new_n24865, new_n24866, new_n24867, new_n24868, new_n24869,
    new_n24870, new_n24871, new_n24872, new_n24873, new_n24874, new_n24875,
    new_n24876, new_n24877, new_n24878, new_n24879_1, new_n24880,
    new_n24881, new_n24882, new_n24883, new_n24884, new_n24885, new_n24886,
    new_n24887_1, new_n24888, new_n24889, new_n24890, new_n24891,
    new_n24892, new_n24893, new_n24894, new_n24895, new_n24896, new_n24897,
    new_n24898, new_n24899, new_n24900, new_n24901, new_n24902, new_n24903,
    new_n24904, new_n24905, new_n24906, new_n24907, new_n24908, new_n24909,
    new_n24910, new_n24911, new_n24912, new_n24913, new_n24914, new_n24915,
    new_n24916, new_n24917, new_n24918, new_n24919, new_n24920, new_n24921,
    new_n24922, new_n24923, new_n24924, new_n24925, new_n24926, new_n24927,
    new_n24928, new_n24929, new_n24930, new_n24931, new_n24932, new_n24933,
    new_n24934_1, new_n24935, new_n24936, new_n24937_1, new_n24938,
    new_n24939, new_n24940, new_n24941, new_n24942, new_n24943, new_n24944,
    new_n24945, new_n24946, new_n24947, new_n24948, new_n24949, new_n24950,
    new_n24953, new_n24954, new_n24955, new_n24956, new_n24957, new_n24958,
    new_n24959, new_n24960, new_n24961, new_n24962, new_n24963, new_n24964,
    new_n24965, new_n24966, new_n24967, new_n24968, new_n24969, new_n24970,
    new_n24971, new_n24972, new_n24973, new_n24974, new_n24975, new_n24976,
    new_n24977, new_n24978, new_n24979, new_n24980, new_n24981, new_n24982,
    new_n24983, new_n24984, new_n24985, new_n24986, new_n24987, new_n24988,
    new_n24989, new_n24990, new_n24991, new_n24992, new_n24993, new_n24994,
    new_n24995, new_n24996, new_n24997, new_n24998_1, new_n24999,
    new_n25000, new_n25001, new_n25002, new_n25003, new_n25004, new_n25005,
    new_n25006_1, new_n25007, new_n25008, new_n25009, new_n25010,
    new_n25011, new_n25012, new_n25013, new_n25014, new_n25015, new_n25016,
    new_n25017, new_n25018, new_n25019, new_n25020, new_n25021, new_n25022,
    new_n25023_1, new_n25024, new_n25025, new_n25026, new_n25027,
    new_n25028, new_n25029, new_n25030, new_n25031, new_n25032_1,
    new_n25033, new_n25034, new_n25035, new_n25036, new_n25037, new_n25038,
    new_n25039, new_n25040, new_n25041, new_n25042, new_n25043, new_n25044,
    new_n25045, new_n25046, new_n25047, new_n25048, new_n25049, new_n25050,
    new_n25051, new_n25052, new_n25053, new_n25054, new_n25055, new_n25056,
    new_n25057, new_n25058, new_n25059, new_n25060, new_n25061,
    new_n25062_1, new_n25063, new_n25064, new_n25065, new_n25066,
    new_n25067, new_n25068_1, new_n25069, new_n25070, new_n25071,
    new_n25072, new_n25073_1, new_n25075, new_n25077, new_n25079,
    new_n25081, new_n25082, new_n25083_1, new_n25084, new_n25085,
    new_n25086, new_n25087, new_n25088, new_n25089, new_n25090, new_n25091,
    new_n25092, new_n25093, new_n25094_1, new_n25095, new_n25096,
    new_n25097_1, new_n25098, new_n25099, new_n25100, new_n25101,
    new_n25102, new_n25103, new_n25104, new_n25105, new_n25106, new_n25107,
    new_n25108, new_n25109, new_n25110, new_n25111, new_n25112, new_n25113,
    new_n25114, new_n25115, new_n25116, new_n25117, new_n25118,
    new_n25119_1, new_n25120_1, new_n25121, new_n25122, new_n25123,
    new_n25124, new_n25125, new_n25126_1, new_n25127, new_n25128,
    new_n25129, new_n25130, new_n25131, new_n25132, new_n25133_1,
    new_n25134, new_n25135, new_n25136, new_n25137, new_n25138, new_n25139,
    new_n25140, new_n25141, new_n25142, new_n25143, new_n25144, new_n25145,
    new_n25146, new_n25147, new_n25148, new_n25149, new_n25150, new_n25151,
    new_n25152, new_n25153, new_n25154, new_n25155_1, new_n25156,
    new_n25157, new_n25158, new_n25159, new_n25160, new_n25161, new_n25162,
    new_n25163, new_n25164, new_n25165, new_n25166, new_n25167,
    new_n25168_1, new_n25169, new_n25170, new_n25171, new_n25172,
    new_n25173, new_n25174, new_n25175, new_n25176, new_n25177, new_n25178,
    new_n25179, new_n25180, new_n25181_1, new_n25182, new_n25183,
    new_n25184, new_n25185, new_n25186, new_n25187, new_n25188, new_n25189,
    new_n25190, new_n25191, new_n25192, new_n25193, new_n25194, new_n25195,
    new_n25196, new_n25197, new_n25198, new_n25200_1, new_n25201,
    new_n25202, new_n25203, new_n25204, new_n25205, new_n25206, new_n25207,
    new_n25208, new_n25209_1, new_n25210, new_n25212, new_n25213,
    new_n25214, new_n25215_1, new_n25216, new_n25217, new_n25218,
    new_n25219, new_n25220, new_n25221, new_n25222, new_n25223, new_n25224,
    new_n25225, new_n25226, new_n25227, new_n25228, new_n25229, new_n25230,
    new_n25231, new_n25232, new_n25233, new_n25234, new_n25235, new_n25236,
    new_n25237, new_n25238, new_n25241, new_n25246, new_n25247, new_n25248,
    new_n25249, new_n25250, new_n25251, new_n25252, new_n25253,
    new_n25254_1, new_n25255, new_n25256_1, new_n25257, new_n25258,
    new_n25259, new_n25260, new_n25261, new_n25262, new_n25263, new_n25264,
    new_n25265, new_n25270, new_n25272, new_n25275, new_n25277, new_n25279,
    new_n25282, new_n25283, new_n25284, new_n25285, new_n25286, new_n25287,
    new_n25288, new_n25289, new_n25290, new_n25291, new_n25292,
    new_n25293_1, new_n25294, new_n25295, new_n25296_1, new_n25297,
    new_n25298, new_n25299, new_n25300, new_n25301, new_n25302, new_n25303,
    new_n25304, new_n25305, new_n25306, new_n25307, new_n25308, new_n25309,
    new_n25310, new_n25311, new_n25312, new_n25313, new_n25314, new_n25315,
    new_n25316_1, new_n25317, new_n25318, new_n25319, new_n25320,
    new_n25321, new_n25322, new_n25323, new_n25324, new_n25325, new_n25326,
    new_n25327, new_n25329, new_n25330, new_n25331_1, new_n25332_1,
    new_n25333, new_n25334, new_n25335, new_n25336_1, new_n25337_1,
    new_n25338, new_n25339, new_n25340, new_n25341, new_n25342, new_n25343,
    new_n25344, new_n25345_1, new_n25346, new_n25347, new_n25348,
    new_n25349, new_n25350, new_n25351, new_n25352, new_n25353, new_n25354,
    new_n25355, new_n25356_1, new_n25357, new_n25358, new_n25359,
    new_n25360, new_n25361, new_n25362_1, new_n25363, new_n25364,
    new_n25365_1, new_n25366, new_n25367, new_n25368, new_n25369,
    new_n25370_1, new_n25372, new_n25373, new_n25374, new_n25375,
    new_n25376, new_n25377, new_n25378, new_n25379, new_n25380,
    new_n25381_1, new_n25382, new_n25383, new_n25384, new_n25385,
    new_n25386, new_n25387, new_n25388, new_n25389, new_n25390, new_n25391,
    new_n25392, new_n25393, new_n25394, new_n25395, new_n25396, new_n25397,
    new_n25398, new_n25399, new_n25400, new_n25401, new_n25402, new_n25403,
    new_n25404, new_n25405, new_n25406, new_n25407, new_n25408, new_n25409,
    new_n25410, new_n25411, new_n25412_1, new_n25413, new_n25414,
    new_n25415, new_n25416, new_n25417, new_n25418, new_n25419, new_n25420,
    new_n25421, new_n25422, new_n25423, new_n25424, new_n25425, new_n25426,
    new_n25427, new_n25428, new_n25429, new_n25430, new_n25431, new_n25432,
    new_n25433, new_n25434, new_n25435_1, new_n25436, new_n25437,
    new_n25438, new_n25439, new_n25440, new_n25441, new_n25442, new_n25443,
    new_n25444, new_n25445, new_n25446, new_n25447, new_n25448, new_n25449,
    new_n25450, new_n25451, new_n25452, new_n25453, new_n25454, new_n25455,
    new_n25456, new_n25457, new_n25458, new_n25459, new_n25460_1,
    new_n25461, new_n25462, new_n25463, new_n25464_1, new_n25465,
    new_n25466, new_n25467, new_n25468_1, new_n25469, new_n25470,
    new_n25471_1, new_n25472, new_n25473, new_n25474, new_n25475_1,
    new_n25476, new_n25477, new_n25478, new_n25479, new_n25480, new_n25481,
    new_n25482, new_n25483, new_n25484, new_n25485, new_n25486, new_n25487,
    new_n25488, new_n25489, new_n25490, new_n25491, new_n25492, new_n25493,
    new_n25494_1, new_n25495, new_n25496, new_n25497, new_n25498,
    new_n25499_1, new_n25500, new_n25501, new_n25502, new_n25503,
    new_n25504, new_n25505, new_n25506, new_n25507, new_n25508, new_n25509,
    new_n25510, new_n25511, new_n25512, new_n25513_1, new_n25514,
    new_n25515, new_n25516, new_n25517, new_n25518_1, new_n25519,
    new_n25520, new_n25521, new_n25522, new_n25523_1, new_n25524,
    new_n25525, new_n25526, new_n25527, new_n25528, new_n25529, new_n25530,
    new_n25531, new_n25532_1, new_n25533, new_n25534, new_n25535,
    new_n25536, new_n25537, new_n25538, new_n25539_1, new_n25540,
    new_n25541, new_n25542, new_n25543, new_n25544, new_n25545, new_n25546,
    new_n25547, new_n25548, new_n25549, new_n25550_1, new_n25551,
    new_n25552, new_n25553, new_n25554, new_n25555, new_n25556, new_n25557,
    new_n25558, new_n25559, new_n25560, new_n25561, new_n25562, new_n25563,
    new_n25564, new_n25565_1, new_n25566, new_n25567, new_n25568,
    new_n25569, new_n25570, new_n25571, new_n25572, new_n25573, new_n25574,
    new_n25575, new_n25576, new_n25577, new_n25578, new_n25579, new_n25580,
    new_n25581, new_n25582, new_n25583, new_n25584, new_n25585,
    new_n25586_1, new_n25587, new_n25588, new_n25589, new_n25590,
    new_n25593, new_n25595, new_n25597, new_n25598, new_n25599, new_n25600,
    new_n25601, new_n25602, new_n25603, new_n25604, new_n25605, new_n25606,
    new_n25607, new_n25608, new_n25609, new_n25610, new_n25611_1,
    new_n25612, new_n25613, new_n25614_1, new_n25615, new_n25616,
    new_n25617, new_n25618, new_n25619_1, new_n25620, new_n25621,
    new_n25622, new_n25623, new_n25624, new_n25625, new_n25626, new_n25627,
    new_n25628, new_n25629_1, new_n25630, new_n25632, new_n25634,
    new_n25635, new_n25636, new_n25637, new_n25638, new_n25639, new_n25640,
    new_n25641, new_n25642, new_n25643_1, new_n25644, new_n25645,
    new_n25646, new_n25647, new_n25648, new_n25649, new_n25650, new_n25651,
    new_n25652, new_n25653, new_n25654, new_n25655, new_n25656, new_n25657,
    new_n25658, new_n25659, new_n25662, new_n25663, new_n25664,
    new_n25665_1, new_n25666, new_n25667, new_n25668, new_n25670,
    new_n25673, new_n25675, new_n25676, new_n25679, new_n25681, new_n25682,
    new_n25683, new_n25684, new_n25685, new_n25686, new_n25687, new_n25688,
    new_n25689, new_n25690, new_n25691, new_n25692, new_n25693,
    new_n25694_1, new_n25695, new_n25696, new_n25697, new_n25698,
    new_n25699, new_n25700, new_n25701, new_n25704, new_n25706_1,
    new_n25707, new_n25708, new_n25709, new_n25710, new_n25711, new_n25712,
    new_n25713, new_n25714, new_n25715, new_n25716, new_n25717, new_n25718,
    new_n25719_1, new_n25720, new_n25721, new_n25722, new_n25723,
    new_n25725, new_n25726, new_n25727, new_n25728, new_n25729, new_n25730,
    new_n25731, new_n25732, new_n25733, new_n25734, new_n25735, new_n25736,
    new_n25737, new_n25738_1, new_n25739, new_n25740, new_n25741,
    new_n25742, new_n25743, new_n25744, new_n25745, new_n25746, new_n25747,
    new_n25748, new_n25750, new_n25751_1, new_n25752, new_n25753,
    new_n25754, new_n25755, new_n25756_1, new_n25757, new_n25758_1,
    new_n25759, new_n25760, new_n25761, new_n25762, new_n25763, new_n25764,
    new_n25765, new_n25766, new_n25767, new_n25768, new_n25769, new_n25770,
    new_n25771, new_n25772, new_n25773_1, new_n25774, new_n25775,
    new_n25776, new_n25777, new_n25778, new_n25779, new_n25780, new_n25781,
    new_n25782, new_n25783, new_n25784_1, new_n25785, new_n25786,
    new_n25787, new_n25788, new_n25789, new_n25790, new_n25791,
    new_n25792_1, new_n25793, new_n25794, new_n25795, new_n25796,
    new_n25797_1, new_n25798, new_n25799, new_n25800, new_n25802,
    new_n25803, new_n25804, new_n25805, new_n25806, new_n25807, new_n25808,
    new_n25809, new_n25810, new_n25811, new_n25812, new_n25813, new_n25814,
    new_n25815, new_n25816_1, new_n25817, new_n25818, new_n25819,
    new_n25820, new_n25821, new_n25822, new_n25823, new_n25824, new_n25825,
    new_n25826_1, new_n25827, new_n25828, new_n25829, new_n25830,
    new_n25831, new_n25832, new_n25833, new_n25834, new_n25835, new_n25836,
    new_n25837, new_n25838, new_n25839_1, new_n25840_1, new_n25841,
    new_n25842, new_n25843, new_n25844, new_n25845, new_n25846, new_n25847,
    new_n25848, new_n25849, new_n25850, new_n25851, new_n25852, new_n25853,
    new_n25854, new_n25855, new_n25856, new_n25857, new_n25858, new_n25859,
    new_n25860, new_n25861, new_n25862, new_n25863, new_n25864, new_n25865,
    new_n25866, new_n25867, new_n25868, new_n25869, new_n25870, new_n25871,
    new_n25872_1, new_n25873_1, new_n25874, new_n25875, new_n25876,
    new_n25877_1, new_n25878, new_n25879, new_n25880, new_n25881,
    new_n25882, new_n25883, new_n25884, new_n25885, new_n25886, new_n25887,
    new_n25888, new_n25889, new_n25890, new_n25891, new_n25892, new_n25893,
    new_n25894, new_n25895, new_n25896, new_n25897, new_n25898, new_n25899,
    new_n25900, new_n25901, new_n25902, new_n25903, new_n25904, new_n25905,
    new_n25906, new_n25907, new_n25908, new_n25911, new_n25913, new_n25915,
    new_n25916, new_n25917, new_n25918, new_n25919, new_n25920, new_n25921,
    new_n25922, new_n25923_1, new_n25924, new_n25925, new_n25926_1,
    new_n25927, new_n25928, new_n25929, new_n25930, new_n25931, new_n25932,
    new_n25933, new_n25934_1, new_n25935, new_n25936, new_n25937,
    new_n25938_1, new_n25939, new_n25940, new_n25941, new_n25942,
    new_n25943, new_n25944, new_n25945, new_n25946, new_n25947, new_n25948,
    new_n25949, new_n25950, new_n25951, new_n25952, new_n25953, new_n25954,
    new_n25955, new_n25956, new_n25957, new_n25958, new_n25959, new_n25960,
    new_n25961, new_n25962, new_n25963, new_n25964, new_n25965, new_n25966,
    new_n25967, new_n25968, new_n25969, new_n25970, new_n25971,
    new_n25972_1, new_n25973, new_n25974_1, new_n25975, new_n25976,
    new_n25977, new_n25978, new_n25979, new_n25980, new_n25981, new_n25982,
    new_n25983, new_n25984, new_n25985_1, new_n25986, new_n25987,
    new_n25988, new_n25989, new_n25990, new_n25991, new_n25992, new_n25993,
    new_n25994_1, new_n25995, new_n25996, new_n25997, new_n25998,
    new_n25999, new_n26000, new_n26001, new_n26002, new_n26003, new_n26004,
    new_n26005, new_n26006, new_n26007, new_n26008, new_n26009, new_n26010,
    new_n26011, new_n26012, new_n26013, new_n26014, new_n26015, new_n26016,
    new_n26017, new_n26018, new_n26019, new_n26020, new_n26021, new_n26022,
    new_n26023, new_n26024, new_n26025, new_n26026, new_n26027, new_n26028,
    new_n26029, new_n26030, new_n26031, new_n26032, new_n26033, new_n26034,
    new_n26035, new_n26036_1, new_n26037, new_n26038, new_n26039,
    new_n26040, new_n26041, new_n26042, new_n26043, new_n26044, new_n26045,
    new_n26046, new_n26047, new_n26048, new_n26049, new_n26050, new_n26051,
    new_n26052, new_n26053_1, new_n26054_1, new_n26056, new_n26057,
    new_n26059, new_n26062, new_n26064, new_n26067, new_n26068, new_n26069,
    new_n26070, new_n26071, new_n26072, new_n26073, new_n26074, new_n26075,
    new_n26076, new_n26077, new_n26078, new_n26079, new_n26080, new_n26081,
    new_n26082, new_n26083, new_n26084_1, new_n26085, new_n26086,
    new_n26087, new_n26088, new_n26089, new_n26090, new_n26091, new_n26092,
    new_n26093, new_n26094, new_n26095, new_n26096_1, new_n26097,
    new_n26098, new_n26099, new_n26100, new_n26101, new_n26102, new_n26103,
    new_n26104, new_n26105, new_n26106, new_n26107_1, new_n26108,
    new_n26109, new_n26111_1, new_n26112, new_n26113_1, new_n26114,
    new_n26115, new_n26116, new_n26117, new_n26118, new_n26119, new_n26120,
    new_n26121, new_n26122, new_n26123, new_n26124, new_n26125, new_n26126,
    new_n26127, new_n26128, new_n26129, new_n26130, new_n26131, new_n26132,
    new_n26133, new_n26134, new_n26135, new_n26136, new_n26137, new_n26138,
    new_n26139, new_n26140, new_n26141, new_n26142, new_n26143, new_n26144,
    new_n26145, new_n26146, new_n26148, new_n26151, new_n26153, new_n26158,
    new_n26159_1, new_n26160, new_n26161, new_n26162, new_n26163,
    new_n26164, new_n26165, new_n26166, new_n26167_1, new_n26168,
    new_n26169, new_n26170, new_n26171, new_n26172, new_n26173, new_n26174,
    new_n26175, new_n26176, new_n26177, new_n26178, new_n26179_1,
    new_n26180_1, new_n26181, new_n26182, new_n26183, new_n26185,
    new_n26188, new_n26189, new_n26190, new_n26191_1, new_n26192,
    new_n26193, new_n26194, new_n26195, new_n26196, new_n26197, new_n26198,
    new_n26199, new_n26200, new_n26201, new_n26202, new_n26203, new_n26204,
    new_n26205, new_n26206, new_n26207, new_n26208, new_n26209, new_n26210,
    new_n26211, new_n26212, new_n26213, new_n26214, new_n26215, new_n26216,
    new_n26217, new_n26218, new_n26219, new_n26220_1, new_n26221,
    new_n26222, new_n26223, new_n26224_1, new_n26226, new_n26228,
    new_n26229_1, new_n26230, new_n26231, new_n26232, new_n26233,
    new_n26234, new_n26235, new_n26236, new_n26237_1, new_n26238,
    new_n26239, new_n26240, new_n26241, new_n26242, new_n26243, new_n26244,
    new_n26245, new_n26246, new_n26247, new_n26248, new_n26249,
    new_n26250_1, new_n26251, new_n26252, new_n26253, new_n26254,
    new_n26255, new_n26256, new_n26257, new_n26258, new_n26259, new_n26260,
    new_n26261, new_n26262, new_n26263, new_n26264_1, new_n26265,
    new_n26266, new_n26267, new_n26268, new_n26269, new_n26270, new_n26271,
    new_n26272, new_n26273, new_n26274_1, new_n26275, new_n26276,
    new_n26277, new_n26278, new_n26279, new_n26280, new_n26281, new_n26282,
    new_n26283, new_n26284, new_n26285, new_n26286, new_n26287_1,
    new_n26288, new_n26289, new_n26290, new_n26291, new_n26292, new_n26293,
    new_n26294, new_n26295, new_n26296, new_n26297, new_n26298, new_n26299,
    new_n26301, new_n26302, new_n26303, new_n26304, new_n26305, new_n26306,
    new_n26307, new_n26308, new_n26309, new_n26310, new_n26311, new_n26312,
    new_n26313, new_n26314, new_n26315, new_n26316, new_n26317_1,
    new_n26318_1, new_n26319, new_n26320, new_n26321, new_n26322,
    new_n26323, new_n26324, new_n26325, new_n26326, new_n26327, new_n26328,
    new_n26329, new_n26330, new_n26331, new_n26332, new_n26334, new_n26335,
    new_n26337, new_n26338, new_n26339, new_n26340, new_n26341, new_n26342,
    new_n26343, new_n26344, new_n26345, new_n26346, new_n26347, new_n26348,
    new_n26349, new_n26350, new_n26351, new_n26352, new_n26353_1,
    new_n26354, new_n26355, new_n26356, new_n26357, new_n26358, new_n26359,
    new_n26360, new_n26361, new_n26362, new_n26363, new_n26364, new_n26365,
    new_n26366, new_n26367, new_n26368, new_n26369, new_n26370, new_n26371,
    new_n26372, new_n26373, new_n26374, new_n26375_1, new_n26376,
    new_n26377, new_n26378, new_n26379, new_n26380, new_n26383, new_n26384,
    new_n26386, new_n26388, new_n26389, new_n26390, new_n26391, new_n26392,
    new_n26393, new_n26394, new_n26395, new_n26396_1, new_n26397,
    new_n26398, new_n26399, new_n26400, new_n26401, new_n26402, new_n26403,
    new_n26404, new_n26405, new_n26406, new_n26407, new_n26408_1,
    new_n26409, new_n26410, new_n26411, new_n26412, new_n26413, new_n26414,
    new_n26415, new_n26416, new_n26417, new_n26418, new_n26419, new_n26420,
    new_n26421, new_n26422, new_n26423, new_n26424, new_n26425, new_n26426,
    new_n26427, new_n26428, new_n26429_1, new_n26430, new_n26431_1,
    new_n26432, new_n26433, new_n26434, new_n26435, new_n26436,
    new_n26439_1, new_n26440, new_n26441, new_n26442, new_n26443_1,
    new_n26444, new_n26445, new_n26446, new_n26447, new_n26448, new_n26449,
    new_n26450, new_n26451, new_n26452_1, new_n26453, new_n26454,
    new_n26455, new_n26456, new_n26457, new_n26458, new_n26459, new_n26460,
    new_n26463, new_n26466, new_n26468, new_n26470, new_n26472, new_n26473,
    new_n26474, new_n26475, new_n26476, new_n26477, new_n26478, new_n26479,
    new_n26480, new_n26481, new_n26482, new_n26483_1, new_n26484,
    new_n26485, new_n26486, new_n26487, new_n26488, new_n26489, new_n26490,
    new_n26491, new_n26492_1, new_n26493, new_n26494, new_n26495,
    new_n26496, new_n26497, new_n26498, new_n26499, new_n26500, new_n26501,
    new_n26502, new_n26503, new_n26504, new_n26505, new_n26506, new_n26507,
    new_n26508, new_n26509, new_n26510_1, new_n26511, new_n26512_1,
    new_n26513, new_n26514, new_n26515_1, new_n26516, new_n26517,
    new_n26518, new_n26519, new_n26520, new_n26521, new_n26522, new_n26523,
    new_n26524, new_n26525, new_n26526, new_n26527, new_n26528, new_n26529,
    new_n26530, new_n26531, new_n26532, new_n26533, new_n26534, new_n26535,
    new_n26536, new_n26540, new_n26546, new_n26548, new_n26549, new_n26550,
    new_n26551, new_n26552, new_n26553_1, new_n26554, new_n26555,
    new_n26556, new_n26557, new_n26558, new_n26559, new_n26560, new_n26567,
    new_n26570, new_n26573, new_n26578, new_n26580, new_n26582, new_n26583,
    new_n26584, new_n26585, new_n26586, new_n26587, new_n26588, new_n26589,
    new_n26590_1, new_n26591, new_n26592, new_n26593, new_n26594,
    new_n26595, new_n26596, new_n26597, new_n26598_1, new_n26599,
    new_n26600, new_n26601, new_n26602, new_n26603, new_n26604,
    new_n26605_1, new_n26606, new_n26607, new_n26608, new_n26609,
    new_n26610, new_n26611, new_n26613, new_n26614, new_n26615, new_n26616,
    new_n26617, new_n26618, new_n26619, new_n26620, new_n26621, new_n26622,
    new_n26623, new_n26624, new_n26625_1, new_n26626, new_n26627,
    new_n26628, new_n26629, new_n26630, new_n26631, new_n26632, new_n26633,
    new_n26634, new_n26635, new_n26636, new_n26637, new_n26638, new_n26639,
    new_n26640, new_n26641, new_n26642, new_n26644, new_n26645, new_n26646,
    new_n26647, new_n26648, new_n26649, new_n26650, new_n26651, new_n26652,
    new_n26653, new_n26654, new_n26655, new_n26656_1, new_n26657,
    new_n26658, new_n26659, new_n26660_1, new_n26662, new_n26666,
    new_n26667, new_n26668, new_n26669, new_n26670, new_n26671, new_n26672,
    new_n26673, new_n26674_1, new_n26675_1, new_n26676, new_n26677,
    new_n26678, new_n26679, new_n26680, new_n26681_1, new_n26682,
    new_n26683, new_n26684, new_n26685, new_n26686, new_n26687, new_n26688,
    new_n26689, new_n26690, new_n26691, new_n26692, new_n26693, new_n26694,
    new_n26695, new_n26696_1, new_n26697, new_n26701, new_n26705,
    new_n26708, new_n26709, new_n26710, new_n26711, new_n26712, new_n26713,
    new_n26714, new_n26715, new_n26717, new_n26721, new_n26723, new_n26724,
    new_n26725_1, new_n26726, new_n26727_1, new_n26728, new_n26729_1,
    new_n26730, new_n26731, new_n26732, new_n26733, new_n26734, new_n26735,
    new_n26740, new_n26745_1, new_n26747, new_n26748_1, new_n26749,
    new_n26750, new_n26751, new_n26752_1, new_n26753, new_n26754,
    new_n26755, new_n26756, new_n26757, new_n26758, new_n26759, new_n26760,
    new_n26761, new_n26762, new_n26763, new_n26764, new_n26765, new_n26766,
    new_n26767, new_n26768, new_n26769, new_n26770, new_n26771,
    new_n26775_1, new_n26777, new_n26778, new_n26779, new_n26780_1,
    new_n26781, new_n26782, new_n26783, new_n26786, new_n26787, new_n26788,
    new_n26789, new_n26790, new_n26791, new_n26792, new_n26794_1,
    new_n26796, new_n26798, new_n26800, new_n26801_1, new_n26802,
    new_n26803, new_n26804, new_n26805, new_n26806, new_n26807,
    new_n26808_1, new_n26809, new_n26810, new_n26811, new_n26812,
    new_n26813, new_n26814, new_n26815_1, new_n26816, new_n26817,
    new_n26818, new_n26819, new_n26820, new_n26821, new_n26822,
    new_n26823_1, new_n26824, new_n26825, new_n26826, new_n26827,
    new_n26828, new_n26829, new_n26830, new_n26831, new_n26832, new_n26833,
    new_n26834, new_n26835, new_n26836, new_n26837, new_n26838, new_n26839,
    new_n26840, new_n26841, new_n26842, new_n26843, new_n26844, new_n26845,
    new_n26846, new_n26847_1, new_n26848, new_n26849, new_n26850,
    new_n26851, new_n26852, new_n26853, new_n26854, new_n26855, new_n26856,
    new_n26857, new_n26858, new_n26861, new_n26862, new_n26863, new_n26864,
    new_n26865, new_n26866, new_n26867, new_n26868, new_n26869, new_n26870,
    new_n26872, new_n26873, new_n26874, new_n26875, new_n26876, new_n26877,
    new_n26878, new_n26879, new_n26880, new_n26881, new_n26882_1,
    new_n26883, new_n26884, new_n26885, new_n26886, new_n26887, new_n26888,
    new_n26889, new_n26890, new_n26891, new_n26892, new_n26893, new_n26894,
    new_n26895, new_n26896, new_n26897, new_n26898, new_n26901, new_n26906,
    new_n26908, new_n26910, new_n26912, new_n26913_1, new_n26914,
    new_n26915, new_n26916, new_n26917, new_n26918, new_n26919, new_n26920,
    new_n26921_1, new_n26922, new_n26923_1, new_n26924, new_n26925,
    new_n26926, new_n26927, new_n26928, new_n26929_1, new_n26930_1,
    new_n26931, new_n26932, new_n26933, new_n26934, new_n26935, new_n26936,
    new_n26937, new_n26938, new_n26939, new_n26940, new_n26941, new_n26942,
    new_n26943_1, new_n26944, new_n26945, new_n26946, new_n26947,
    new_n26948, new_n26949, new_n26953, new_n26956, new_n26957, new_n26958,
    new_n26959, new_n26960, new_n26961, new_n26964, new_n26970_1,
    new_n26972, new_n26974, new_n26975, new_n26976, new_n26977, new_n26978,
    new_n26979_1, new_n26980, new_n26981, new_n26982, new_n26983,
    new_n26984, new_n26985, new_n26986_1, new_n26987, new_n26988,
    new_n26989, new_n26990, new_n26991, new_n26992, new_n26993, new_n26994,
    new_n26995, new_n26996, new_n26997, new_n26998, new_n26999, new_n27000,
    new_n27001, new_n27002, new_n27003, new_n27004_1, new_n27005,
    new_n27006, new_n27007, new_n27008, new_n27009, new_n27010,
    new_n27011_1, new_n27012, new_n27013, new_n27014, new_n27015,
    new_n27016, new_n27017, new_n27018, new_n27019_1, new_n27020,
    new_n27021, new_n27022, new_n27023, new_n27024, new_n27025, new_n27026,
    new_n27027, new_n27028, new_n27029, new_n27030, new_n27031_1,
    new_n27032, new_n27033, new_n27034, new_n27035, new_n27036,
    new_n27037_1, new_n27038, new_n27039, new_n27040, new_n27041,
    new_n27042, new_n27043, new_n27044, new_n27045, new_n27046, new_n27047,
    new_n27048, new_n27049, new_n27050, new_n27051_1, new_n27052,
    new_n27053, new_n27054, new_n27055, new_n27056, new_n27057, new_n27058,
    new_n27059, new_n27061, new_n27062, new_n27063, new_n27064, new_n27065,
    new_n27066, new_n27067, new_n27068, new_n27069, new_n27070, new_n27071,
    new_n27072_1, new_n27073, new_n27074, new_n27075, new_n27076,
    new_n27077, new_n27078, new_n27079_1, new_n27080, new_n27081,
    new_n27082, new_n27083, new_n27084, new_n27085, new_n27086, new_n27087,
    new_n27088, new_n27089_1, new_n27090, new_n27091, new_n27092,
    new_n27093, new_n27094, new_n27095, new_n27096_1, new_n27097,
    new_n27098, new_n27099, new_n27100, new_n27101, new_n27102, new_n27103,
    new_n27104_1, new_n27105, new_n27106, new_n27107, new_n27108,
    new_n27109, new_n27110_1, new_n27111, new_n27112_1, new_n27113,
    new_n27114, new_n27115, new_n27116, new_n27117, new_n27118, new_n27119,
    new_n27120_1, new_n27121, new_n27122, new_n27123, new_n27124,
    new_n27125, new_n27126, new_n27127, new_n27128, new_n27129,
    new_n27130_1, new_n27131, new_n27132, new_n27133, new_n27134_1,
    new_n27135, new_n27136, new_n27137, new_n27138, new_n27139, new_n27140,
    new_n27141, new_n27142, new_n27143, new_n27144, new_n27147, new_n27148,
    new_n27149, new_n27150, new_n27151, new_n27152, new_n27153, new_n27154,
    new_n27155, new_n27156, new_n27157, new_n27158_1, new_n27159,
    new_n27160, new_n27161, new_n27162, new_n27163_1, new_n27165,
    new_n27166, new_n27169, new_n27172, new_n27173, new_n27174, new_n27175,
    new_n27176, new_n27177, new_n27178, new_n27179, new_n27180, new_n27181,
    new_n27182, new_n27183, new_n27184, new_n27185, new_n27186, new_n27187,
    new_n27188_1, new_n27189, new_n27190, new_n27191, new_n27192,
    new_n27193, new_n27194_1, new_n27195, new_n27196, new_n27197,
    new_n27198, new_n27199, new_n27200, new_n27201, new_n27202, new_n27203,
    new_n27204, new_n27205, new_n27206, new_n27207, new_n27208, new_n27209,
    new_n27210, new_n27211, new_n27212, new_n27213, new_n27214, new_n27215,
    new_n27216, new_n27217, new_n27218, new_n27219, new_n27220, new_n27221,
    new_n27222, new_n27223, new_n27224, new_n27225, new_n27226, new_n27227,
    new_n27228, new_n27229, new_n27230, new_n27231, new_n27232, new_n27233,
    new_n27234, new_n27235, new_n27236, new_n27237, new_n27238, new_n27239,
    new_n27240, new_n27241, new_n27242, new_n27243, new_n27244, new_n27245,
    new_n27246, new_n27247, new_n27248, new_n27249, new_n27250, new_n27251,
    new_n27252, new_n27253, new_n27254, new_n27255, new_n27256, new_n27257,
    new_n27258, new_n27259, new_n27260, new_n27261, new_n27262, new_n27263,
    new_n27264, new_n27265, new_n27266, new_n27268, new_n27269, new_n27270,
    new_n27271, new_n27272, new_n27273, new_n27274, new_n27275, new_n27276,
    new_n27277, new_n27278, new_n27279, new_n27282, new_n27283, new_n27284,
    new_n27285, new_n27286, new_n27287, new_n27288, new_n27292, new_n27295,
    new_n27296, new_n27297, new_n27298, new_n27299, new_n27300, new_n27301,
    new_n27302, new_n27303, new_n27304, new_n27305, new_n27306, new_n27307,
    new_n27308, new_n27309, new_n27310, new_n27311, new_n27312, new_n27313,
    new_n27314, new_n27315, new_n27316, new_n27317, new_n27318, new_n27319,
    new_n27320, new_n27321, new_n27322, new_n27323, new_n27324, new_n27325,
    new_n27326, new_n27327, new_n27328, new_n27329, new_n27330, new_n27331,
    new_n27332, new_n27333, new_n27334, new_n27335, new_n27336, new_n27337,
    new_n27338, new_n27339, new_n27340, new_n27341, new_n27342, new_n27343,
    new_n27344, new_n27345, new_n27346, new_n27347, new_n27348, new_n27349,
    new_n27350, new_n27351, new_n27352, new_n27353, new_n27354, new_n27355,
    new_n27356, new_n27357, new_n27358, new_n27359, new_n27360, new_n27361,
    new_n27362, new_n27363, new_n27364, new_n27365, new_n27366, new_n27367,
    new_n27368, new_n27369, new_n27370, new_n27371, new_n27372, new_n27373,
    new_n27376, new_n27379, new_n27383, new_n27384, new_n27385, new_n27386,
    new_n27387, new_n27388, new_n27390, new_n27392, new_n27395, new_n27396,
    new_n27397, new_n27400, new_n27402, new_n27403, new_n27404, new_n27405,
    new_n27406, new_n27407, new_n27408, new_n27409, new_n27410, new_n27411,
    new_n27412, new_n27413, new_n27414, new_n27415, new_n27416, new_n27417,
    new_n27418, new_n27419, new_n27420, new_n27421, new_n27422, new_n27423,
    new_n27424, new_n27425, new_n27426, new_n27427, new_n27428, new_n27429,
    new_n27430, new_n27431, new_n27432, new_n27433, new_n27434, new_n27435,
    new_n27436, new_n27437, new_n27438, new_n27439, new_n27440, new_n27441,
    new_n27442, new_n27443, new_n27444, new_n27445, new_n27446, new_n27447,
    new_n27448, new_n27449, new_n27450, new_n27451, new_n27452, new_n27453,
    new_n27454, new_n27455, new_n27456, new_n27459, new_n27460, new_n27461,
    new_n27463, new_n27467, new_n27471, new_n27472, new_n27473, new_n27474,
    new_n27475, new_n27476, new_n27477, new_n27478, new_n27479, new_n27480,
    new_n27481, new_n27482, new_n27483, new_n27484, new_n27485, new_n27486,
    new_n27488, new_n27491, new_n27492, new_n27494, new_n27497, new_n27499,
    new_n27503, new_n27504, new_n27505, new_n27506, new_n27507, new_n27508,
    new_n27509, new_n27510, new_n27511, new_n27512, new_n27513, new_n27514,
    new_n27515, new_n27516, new_n27517, new_n27518, new_n27519, new_n27520,
    new_n27521, new_n27522, new_n27524, new_n27525, new_n27526, new_n27527,
    new_n27528, new_n27529, new_n27530, new_n27531, new_n27532, new_n27533,
    new_n27534, new_n27535, new_n27536, new_n27537, new_n27538, new_n27539,
    new_n27540, new_n27541, new_n27542, new_n27543, new_n27544, new_n27545,
    new_n27546, new_n27551, new_n27553, new_n27554, new_n27555, new_n27556,
    new_n27557, new_n27558, new_n27559, new_n27560, new_n27561, new_n27562,
    new_n27563, new_n27564, new_n27565, new_n27566, new_n27567, new_n27568,
    new_n27569, new_n27570, new_n27571, new_n27572, new_n27573, new_n27574,
    new_n27575, new_n27576, new_n27577, new_n27578, new_n27579, new_n27580,
    new_n27581, new_n27582, new_n27583, new_n27584, new_n27585, new_n27586,
    new_n27587, new_n27588, new_n27589, new_n27590, new_n27591, new_n27592,
    new_n27593, new_n27594, new_n27595, new_n27597, new_n27599, new_n27600,
    new_n27601, new_n27602, new_n27603, new_n27604, new_n27605, new_n27606,
    new_n27607, new_n27608, new_n27609, new_n27610, new_n27611, new_n27612,
    new_n27613, new_n27614, new_n27615, new_n27616, new_n27617, new_n27618,
    new_n27619, new_n27620, new_n27621, new_n27622, new_n27623, new_n27624,
    new_n27625, new_n27626, new_n27627, new_n27628, new_n27629, new_n27630,
    new_n27631, new_n27633, new_n27634, new_n27635, new_n27636, new_n27637,
    new_n27638, new_n27639, new_n27640, new_n27641, new_n27642, new_n27643,
    new_n27644, new_n27646, new_n27647, new_n27648, new_n27649, new_n27650,
    new_n27651, new_n27652, new_n27653, new_n27654, new_n27655, new_n27656,
    new_n27657, new_n27658, new_n27659, new_n27660, new_n27663, new_n27665,
    new_n27666, new_n27667, new_n27670, new_n27673, new_n27674, new_n27675,
    new_n27676, new_n27677, new_n27678, new_n27679, new_n27680, new_n27681,
    new_n27682, new_n27683, new_n27684, new_n27685, new_n27686, new_n27687,
    new_n27688, new_n27689, new_n27690, new_n27691, new_n27692, new_n27693,
    new_n27694, new_n27695, new_n27696, new_n27697, new_n27698, new_n27699,
    new_n27700, new_n27701, new_n27702, new_n27703, new_n27704, new_n27705,
    new_n27706, new_n27707, new_n27708, new_n27709, new_n27710, new_n27711,
    new_n27712, new_n27713, new_n27714, new_n27715, new_n27716, new_n27717,
    new_n27718, new_n27719, new_n27720, new_n27721, new_n27722, new_n27723,
    new_n27724, new_n27725, new_n27726, new_n27727, new_n27728, new_n27730,
    new_n27731, new_n27732, new_n27733, new_n27734, new_n27735, new_n27736,
    new_n27737, new_n27738, new_n27739, new_n27740, new_n27741, new_n27742,
    new_n27743, new_n27744, new_n27745, new_n27746, new_n27747, new_n27748,
    new_n27749, new_n27750, new_n27751, new_n27752, new_n27753, new_n27754,
    new_n27755, new_n27756, new_n27757, new_n27758, new_n27759, new_n27760,
    new_n27761, new_n27762, new_n27763, new_n27764, new_n27765, new_n27766,
    new_n27767, new_n27768, new_n27769, new_n27770, new_n27771, new_n27772,
    new_n27773, new_n27774, new_n27775, new_n27776, new_n27777, new_n27778,
    new_n27779, new_n27780, new_n27781, new_n27782, new_n27783, new_n27784,
    new_n27785, new_n27786, new_n27787, new_n27788, new_n27789, new_n27790,
    new_n27791, new_n27792, new_n27793, new_n27794, new_n27795, new_n27796,
    new_n27798, new_n27800, new_n27802, new_n27804, new_n27806, new_n27808,
    new_n27811, new_n27817, new_n27818, new_n27819, new_n27820, new_n27821,
    new_n27822, new_n27824, new_n27827, new_n27829, new_n27831, new_n27832,
    new_n27834, new_n27836, new_n27839, new_n27842, new_n27843, new_n27844,
    new_n27845, new_n27846, new_n27847, new_n27848, new_n27849, new_n27850,
    new_n27851, new_n27852, new_n27853, new_n27854, new_n27855, new_n27856,
    new_n27857, new_n27858, new_n27859, new_n27860, new_n27861, new_n27862,
    new_n27863, new_n27864, new_n27865, new_n27866, new_n27867, new_n27868,
    new_n27869, new_n27870, new_n27871, new_n27872, new_n27873, new_n27874,
    new_n27875, new_n27876, new_n27877, new_n27878, new_n27879, new_n27880,
    new_n27881, new_n27882, new_n27883, new_n27886, new_n27887, new_n27888,
    new_n27889, new_n27890, new_n27891, new_n27892, new_n27893, new_n27894,
    new_n27895, new_n27896, new_n27897, new_n27898, new_n27899, new_n27900,
    new_n27901, new_n27903, new_n27907, new_n27909, new_n27911, new_n27912,
    new_n27913, new_n27914, new_n27915, new_n27916, new_n27917, new_n27918,
    new_n27919, new_n27920, new_n27921, new_n27922, new_n27923, new_n27924,
    new_n27925, new_n27926, new_n27927, new_n27928, new_n27929, new_n27930,
    new_n27931, new_n27932, new_n27933, new_n27934, new_n27935, new_n27936,
    new_n27937, new_n27938, new_n27939, new_n27940, new_n27941, new_n27942,
    new_n27943, new_n27944, new_n27945, new_n27946, new_n27947, new_n27948,
    new_n27949, new_n27950, new_n27951, new_n27952, new_n27953, new_n27954,
    new_n27955, new_n27956, new_n27957, new_n27958, new_n27959, new_n27960,
    new_n27961, new_n27962, new_n27963, new_n27964, new_n27965, new_n27966,
    new_n27967, new_n27968, new_n27969, new_n27970, new_n27971, new_n27972,
    new_n27973, new_n27974, new_n27975, new_n27976, new_n27977, new_n27978,
    new_n27979, new_n27980, new_n27981, new_n27982, new_n27983, new_n27984,
    new_n27985, new_n27986, new_n27987, new_n27988, new_n27989, new_n27990,
    new_n27991, new_n27992, new_n27993, new_n27994, new_n27995, new_n27996,
    new_n27997, new_n27998, new_n27999, new_n28000, new_n28001, new_n28002,
    new_n28003, new_n28004, new_n28005, new_n28006, new_n28007, new_n28008,
    new_n28009, new_n28010, new_n28011, new_n28012, new_n28013, new_n28014,
    new_n28015, new_n28016, new_n28017, new_n28018, new_n28019, new_n28020,
    new_n28021, new_n28022, new_n28023, new_n28024, new_n28025, new_n28026,
    new_n28027, new_n28028, new_n28029, new_n28030, new_n28031, new_n28032,
    new_n28033, new_n28034, new_n28035, new_n28036, new_n28037, new_n28038,
    new_n28039, new_n28040, new_n28041, new_n28042, new_n28043, new_n28044,
    new_n28045, new_n28046, new_n28047, new_n28048, new_n28049, new_n28050,
    new_n28051, new_n28052, new_n28053, new_n28054, new_n28055, new_n28056,
    new_n28057, new_n28058, new_n28059, new_n28060, new_n28061, new_n28062,
    new_n28063, new_n28064, new_n28065, new_n28066, new_n28072, new_n28073,
    new_n28074, new_n28075, new_n28076, new_n28077, new_n28078, new_n28079,
    new_n28080, new_n28081, new_n28082, new_n28083, new_n28084, new_n28085,
    new_n28086, new_n28087, new_n28088, new_n28089, new_n28090, new_n28091,
    new_n28092, new_n28093, new_n28094, new_n28098, new_n28100, new_n28101,
    new_n28102, new_n28103, new_n28104, new_n28105, new_n28106, new_n28107,
    new_n28108, new_n28109, new_n28110, new_n28111, new_n28112, new_n28113,
    new_n28114, new_n28115, new_n28116, new_n28117, new_n28118, new_n28119,
    new_n28120, new_n28121, new_n28122, new_n28123, new_n28124, new_n28125,
    new_n28127, new_n28128, new_n28129, new_n28130, new_n28131, new_n28132,
    new_n28136, new_n28137, new_n28138, new_n28139, new_n28141, new_n28145,
    new_n28148, new_n28149, new_n28152, new_n28154, new_n28155, new_n28156,
    new_n28157, new_n28158, new_n28159, new_n28160, new_n28161, new_n28162,
    new_n28163, new_n28164, new_n28165, new_n28166, new_n28167, new_n28168,
    new_n28169, new_n28170, new_n28171, new_n28172, new_n28173, new_n28174,
    new_n28175, new_n28176, new_n28177, new_n28178, new_n28179, new_n28180,
    new_n28181, new_n28182, new_n28183, new_n28184, new_n28185, new_n28187,
    new_n28189, new_n28191, new_n28193, new_n28196, new_n28198, new_n28202,
    new_n28207, new_n28210, new_n28213, new_n28215, new_n28217, new_n28218,
    new_n28219, new_n28220, new_n28221, new_n28222, new_n28223, new_n28224,
    new_n28225, new_n28226, new_n28227, new_n28228, new_n28229, new_n28230,
    new_n28231, new_n28232, new_n28233, new_n28234, new_n28235, new_n28236,
    new_n28237, new_n28238, new_n28239, new_n28240, new_n28241, new_n28242,
    new_n28243, new_n28244, new_n28245, new_n28246, new_n28247, new_n28248,
    new_n28249, new_n28250, new_n28251, new_n28252, new_n28253, new_n28254,
    new_n28255, new_n28256, new_n28257, new_n28258, new_n28262, new_n28263,
    new_n28266, new_n28268, new_n28270, new_n28271, new_n28272, new_n28273,
    new_n28274, new_n28275, new_n28276, new_n28277, new_n28278, new_n28279,
    new_n28280, new_n28281, new_n28282, new_n28283, new_n28284, new_n28285,
    new_n28286, new_n28287, new_n28291, new_n28292, new_n28293, new_n28296,
    new_n28297, new_n28298, new_n28299, new_n28300, new_n28301, new_n28302,
    new_n28304, new_n28306, new_n28307, new_n28308, new_n28309, new_n28310,
    new_n28311, new_n28312, new_n28313, new_n28314, new_n28315, new_n28316,
    new_n28317, new_n28318, new_n28319, new_n28320, new_n28321, new_n28322,
    new_n28323, new_n28324, new_n28325, new_n28326, new_n28327, new_n28329,
    new_n28331, new_n28332, new_n28333, new_n28334, new_n28335, new_n28336,
    new_n28337, new_n28338, new_n28339, new_n28340, new_n28341, new_n28342,
    new_n28343, new_n28344, new_n28345, new_n28346, new_n28347, new_n28348,
    new_n28349, new_n28350, new_n28351, new_n28352, new_n28353, new_n28354,
    new_n28355, new_n28356, new_n28357, new_n28358, new_n28359, new_n28360,
    new_n28361, new_n28362, new_n28363, new_n28364, new_n28365, new_n28366,
    new_n28367, new_n28368, new_n28369, new_n28370, new_n28371, new_n28372,
    new_n28373, new_n28374, new_n28375, new_n28376, new_n28377, new_n28378,
    new_n28380, new_n28382, new_n28384, new_n28386, new_n28391, new_n28393,
    new_n28396, new_n28399, new_n28407, new_n28408, new_n28412, new_n28413,
    new_n28414, new_n28415, new_n28416, new_n28417, new_n28418, new_n28419,
    new_n28420, new_n28421, new_n28422, new_n28423, new_n28424, new_n28425,
    new_n28426, new_n28427, new_n28430, new_n28431, new_n28432, new_n28433,
    new_n28434, new_n28435, new_n28436, new_n28437, new_n28438, new_n28439,
    new_n28440, new_n28441, new_n28442, new_n28443, new_n28444, new_n28445,
    new_n28446, new_n28447, new_n28448, new_n28449, new_n28450, new_n28451,
    new_n28454, new_n28456, new_n28457, new_n28458, new_n28459, new_n28460,
    new_n28461, new_n28462, new_n28463, new_n28466, new_n28468, new_n28473,
    new_n28474, new_n28475, new_n28476, new_n28477, new_n28478, new_n28479,
    new_n28480, new_n28481, new_n28482, new_n28483, new_n28485, new_n28486,
    new_n28487, new_n28488, new_n28489, new_n28490, new_n28491, new_n28492,
    new_n28493, new_n28494, new_n28495, new_n28496, new_n28497, new_n28498,
    new_n28499, new_n28500, new_n28501, new_n28502, new_n28503, new_n28504,
    new_n28505, new_n28506, new_n28512, new_n28516, new_n28520, new_n28522,
    new_n28524, new_n28526, new_n28528, new_n28531, new_n28534, new_n28536,
    new_n28538, new_n28539, new_n28541, new_n28542, new_n28543, new_n28544,
    new_n28545, new_n28546, new_n28547, new_n28548, new_n28549, new_n28550,
    new_n28551, new_n28552, new_n28553, new_n28554, new_n28555, new_n28556,
    new_n28557, new_n28558, new_n28559, new_n28560, new_n28561, new_n28562,
    new_n28563, new_n28564, new_n28565, new_n28566, new_n28568, new_n28572,
    new_n28573, new_n28574, new_n28575, new_n28576, new_n28578, new_n28581,
    new_n28583, new_n28586, new_n28588, new_n28590, new_n28593, new_n28595,
    new_n28598, new_n28600, new_n28602, new_n28606, new_n28611, new_n28614,
    new_n28618, new_n28619, new_n28620, new_n28621, new_n28622, new_n28623,
    new_n28627, new_n28629, new_n28632, new_n28634, new_n28636, new_n28639,
    new_n28642, new_n28644, new_n28645, new_n28646, new_n28647, new_n28648,
    new_n28649, new_n28650, new_n28654, new_n28655, new_n28656, new_n28657,
    new_n28658, new_n28659, new_n28660, new_n28661, new_n28662, new_n28663,
    new_n28664, new_n28665, new_n28666, new_n28670, new_n28672, new_n28673,
    new_n28674, new_n28675, new_n28676, new_n28677, new_n28678, new_n28679,
    new_n28680, new_n28682, new_n28684, new_n28685, new_n28688, new_n28690,
    new_n28692, new_n28694, new_n28698, new_n28704, new_n28706, new_n28707,
    new_n28708, new_n28709, new_n28710, new_n28713, new_n28714, new_n28715,
    new_n28716, new_n28717, new_n28718, new_n28719, new_n28720, new_n28721,
    new_n28722, new_n28723, new_n28724, new_n28725, new_n28726, new_n28727,
    new_n28728, new_n28729, new_n28732, new_n28733, new_n28734, new_n28736,
    new_n28740, new_n28741, new_n28742, new_n28743, new_n28744, new_n28745,
    new_n28746, new_n28748, new_n28749, new_n28754, new_n28756, new_n28757,
    new_n28761, new_n28769, new_n28771, new_n28773, new_n28774, new_n28775,
    new_n28776, new_n28777, new_n28778, new_n28779, new_n28780, new_n28781,
    new_n28784, new_n28786, new_n28788, new_n28791, new_n28793, new_n28795,
    new_n28796, new_n28797, new_n28798, new_n28799, new_n28800, new_n28801,
    new_n28802, new_n28803, new_n28804, new_n28806, new_n28807, new_n28813,
    new_n28815, new_n28817, new_n28821, new_n28822, new_n28824, new_n28825,
    new_n28826, new_n28827, new_n28828, new_n28829, new_n28830, new_n28831,
    new_n28832, new_n28833, new_n28834, new_n28835, new_n28836, new_n28837,
    new_n28840, new_n28846, new_n28849, new_n28852, new_n28854, new_n28856,
    new_n28858, new_n28860, new_n28862, new_n28864, new_n28865, new_n28866,
    new_n28867, new_n28868, new_n28869, new_n28870, new_n28871, new_n28872,
    new_n28873, new_n28874, new_n28875, new_n28878, new_n28879, new_n28880,
    new_n28881, new_n28882, new_n28883, new_n28884, new_n28885, new_n28886,
    new_n28887, new_n28888, new_n28889, new_n28894, new_n28895, new_n28896,
    new_n28897, new_n28898, new_n28899, new_n28900, new_n28902, new_n28904,
    new_n28905, new_n28906, new_n28907, new_n28908, new_n28909, new_n28912,
    new_n28913, new_n28914, new_n28915, new_n28916, new_n28917, new_n28918,
    new_n28920, new_n28921, new_n28922, new_n28923, new_n28924, new_n28925,
    new_n28926, new_n28927, new_n28928, new_n28929, new_n28930, new_n28931,
    new_n28932, new_n28933, new_n28934, new_n28935, new_n28936, new_n28937,
    new_n28938, new_n28939, new_n28940, new_n28941, new_n28942, new_n28943,
    new_n28944, new_n28945, new_n28946, new_n28947, new_n28948, new_n28952,
    new_n28953, new_n28954, new_n28955, new_n28956, new_n28957, new_n28958,
    new_n28959, new_n28961, new_n28963, new_n28965, new_n28970, new_n28973,
    new_n28976, new_n28979, new_n28980, new_n28986, new_n28988, new_n28993,
    new_n29000, new_n29001, new_n29002, new_n29003, new_n29004, new_n29005,
    new_n29006, new_n29007, new_n29009, new_n29011, new_n29014, new_n29018,
    new_n29020, new_n29022, new_n29026, new_n29032, new_n29034, new_n29040,
    new_n29043, new_n29045, new_n29049, new_n29053, new_n29060, new_n29063,
    new_n29069, new_n29071, new_n29072, new_n29076, new_n29081, new_n29087,
    new_n29089, new_n29090, new_n29091, new_n29092, new_n29093, new_n29094,
    new_n29095, new_n29096, new_n29097, new_n29099, new_n29101, new_n29106,
    new_n29108, new_n29110, new_n29112, new_n29117, new_n29118, new_n29119,
    new_n29120, new_n29121, new_n29122, new_n29123, new_n29124, new_n29125,
    new_n29126, new_n29127, new_n29130, new_n29133, new_n29135, new_n29136,
    new_n29137, new_n29138, new_n29139, new_n29140, new_n29141, new_n29142,
    new_n29145, new_n29146, new_n29149, new_n29151, new_n29154, new_n29155,
    new_n29156, new_n29157, new_n29158, new_n29159, new_n29160, new_n29161,
    new_n29163, new_n29164, new_n29165, new_n29166, new_n29167, new_n29168,
    new_n29169, new_n29170, new_n29171, new_n29172, new_n29173, new_n29174,
    new_n29175, new_n29176, new_n29177, new_n29183, new_n29189, new_n29191,
    new_n29193, new_n29195, new_n29197, new_n29201, new_n29204, new_n29207,
    new_n29208, new_n29209, new_n29210, new_n29213, new_n29215, new_n29218,
    new_n29220, new_n29222, new_n29226, new_n29232, new_n29234, new_n29236,
    new_n29237, new_n29241, new_n29243, new_n29245, new_n29246, new_n29247,
    new_n29249, new_n29253, new_n29260, new_n29261, new_n29262, new_n29266,
    new_n29268, new_n29270, new_n29275, new_n29278, new_n29280, new_n29281,
    new_n29282, new_n29285, new_n29292, new_n29293, new_n29294, new_n29295,
    new_n29296, new_n29297, new_n29298, new_n29299, new_n29300, new_n29301,
    new_n29302, new_n29303, new_n29304, new_n29305, new_n29306, new_n29308,
    new_n29311, new_n29313, new_n29316, new_n29322, new_n29325, new_n29327,
    new_n29328, new_n29329, new_n29330, new_n29331, new_n29332, new_n29333,
    new_n29334, new_n29339, new_n29342, new_n29343, new_n29347, new_n29348,
    new_n29349, new_n29350, new_n29351, new_n29352, new_n29353, new_n29354,
    new_n29355, new_n29356, new_n29357, new_n29358, new_n29359, new_n29361,
    new_n29363, new_n29365, new_n29366, new_n29367, new_n29370, new_n29372,
    new_n29375, new_n29378, new_n29381, new_n29382, new_n29383, new_n29384,
    new_n29385, new_n29388, new_n29390, new_n29393, new_n29396, new_n29397,
    new_n29398, new_n29399, new_n29400, new_n29401, new_n29402, new_n29405,
    new_n29409, new_n29411, new_n29412, new_n29413, new_n29414, new_n29415,
    new_n29416, new_n29417, new_n29418, new_n29420, new_n29425, new_n29426,
    new_n29429, new_n29435, new_n29436, new_n29437, new_n29438, new_n29439,
    new_n29440, new_n29441, new_n29444, new_n29445, new_n29448, new_n29449,
    new_n29450, new_n29451, new_n29452, new_n29453, new_n29454, new_n29458,
    new_n29460, new_n29463, new_n29470, new_n29471, new_n29472, new_n29473,
    new_n29475, new_n29477, new_n29479, new_n29481, new_n29483, new_n29485,
    new_n29488, new_n29490, new_n29493, new_n29494, new_n29495, new_n29498,
    new_n29500, new_n29502, new_n29505, new_n29508, new_n29509, new_n29511,
    new_n29512, new_n29513, new_n29514, new_n29515, new_n29516, new_n29517,
    new_n29519, new_n29524, new_n29525, new_n29526, new_n29528, new_n29529,
    new_n29531, new_n29532, new_n29533, new_n29537, new_n29538, new_n29539,
    new_n29540, new_n29541, new_n29542, new_n29543, new_n29544, new_n29545,
    new_n29546, new_n29547, new_n29548, new_n29549, new_n29550, new_n29551,
    new_n29552, new_n29553, new_n29554, new_n29555, new_n29556, new_n29557,
    new_n29558, new_n29559, new_n29560, new_n29561, new_n29562, new_n29563,
    new_n29565, new_n29567, new_n29569, new_n29571, new_n29572, new_n29573,
    new_n29576, new_n29578, new_n29579, new_n29580, new_n29581, new_n29582,
    new_n29583, new_n29591, new_n29593, new_n29595, new_n29596, new_n29597,
    new_n29598, new_n29599, new_n29600, new_n29602, new_n29609, new_n29615,
    new_n29617, new_n29621, new_n29624, new_n29625, new_n29626, new_n29627,
    new_n29629, new_n29630, new_n29631, new_n29632, new_n29633, new_n29634,
    new_n29635, new_n29637, new_n29643, new_n29645, new_n29649, new_n29651,
    new_n29653, new_n29659, new_n29664, new_n29665, new_n29669, new_n29670,
    new_n29672, new_n29673, new_n29675, new_n29679, new_n29681, new_n29687,
    new_n29688, new_n29689, new_n29690, new_n29691, new_n29692, new_n29693,
    new_n29694, new_n29695, new_n29696, new_n29697, new_n29698, new_n29706,
    new_n29708, new_n29713, new_n29716, new_n29721, new_n29727, new_n29731,
    new_n29732, new_n29735, new_n29742, new_n29743, new_n29748, new_n29752,
    new_n29755, new_n29756, new_n29757, new_n29758, new_n29759, new_n29760,
    new_n29765, new_n29767, new_n29768, new_n29769, new_n29770, new_n29772,
    new_n29774, new_n29775, new_n29777, new_n29781, new_n29783, new_n29787,
    new_n29789, new_n29793, new_n29796, new_n29798, new_n29800, new_n29804,
    new_n29806, new_n29808, new_n29812, new_n29814, new_n29817, new_n29821,
    new_n29824, new_n29826, new_n29830, new_n29836, new_n29840, new_n29842,
    new_n29846, new_n29847, new_n29848, new_n29849, new_n29852, new_n29855,
    new_n29858, new_n29862, new_n29864, new_n29866, new_n29869, new_n29870,
    new_n29877, new_n29880, new_n29883, new_n29885, new_n29889, new_n29893,
    new_n29897, new_n29900, new_n29902, new_n29906, new_n29910, new_n29915,
    new_n29918, new_n29919, new_n29921, new_n29924, new_n29927, new_n29928,
    new_n29929, new_n29930, new_n29931, new_n29932, new_n29933, new_n29934,
    new_n29938, new_n29939, new_n29941, new_n29942, new_n29944, new_n29946,
    new_n29949, new_n29952, new_n29957, new_n29959, new_n29961, new_n29964,
    new_n29965, new_n29966, new_n29967, new_n29969, new_n29971, new_n29974,
    new_n29975, new_n29976, new_n29977, new_n29978, new_n29979, new_n29983,
    new_n29989, new_n29991, new_n29992, new_n29993, new_n29998, new_n29999,
    new_n30002, new_n30004, new_n30007, new_n30009, new_n30013, new_n30015,
    new_n30017, new_n30020, new_n30022, new_n30023, new_n30025, new_n30027,
    new_n30028, new_n30031, new_n30034, new_n30036, new_n30039, new_n30042,
    new_n30044, new_n30045, new_n30046, new_n30047, new_n30048, new_n30049,
    new_n30050, new_n30051, new_n30053, new_n30055, new_n30057, new_n30059,
    new_n30060, new_n30061, new_n30062, new_n30067, new_n30069, new_n30070,
    new_n30072, new_n30073, new_n30074, new_n30075, new_n30076, new_n30077,
    new_n30078, new_n30079, new_n30080, new_n30082, new_n30085, new_n30087,
    new_n30092, new_n30097, new_n30106, new_n30108, new_n30109, new_n30115,
    new_n30119, new_n30120, new_n30122;
not_3  g00000(new_n2349, n9942);
xor_3  g00001(new_n2350, n10739, new_n2349);
not_3  g00002(new_n2351, new_n2350);
not_3  g00003(new_n2352, n25643);
nand_4 g00004(new_n2353, new_n2352, n21753);
not_3  g00005(new_n2354, n21753);
xor_3  g00006(new_n2355_1, n25643, new_n2354);
not_3  g00007(new_n2356, n21832);
nor_4  g00008(new_n2357, new_n2356, n9557);
not_3  g00009(new_n2358, new_n2357);
not_3  g00010(new_n2359, n9557);
xor_3  g00011(new_n2360, n21832, new_n2359);
not_3  g00012(new_n2361_1, n26913);
nor_4  g00013(new_n2362, new_n2361_1, n3136);
not_3  g00014(new_n2363_1, new_n2362);
not_3  g00015(new_n2364, n3136);
xor_3  g00016(new_n2365, n26913, new_n2364);
not_3  g00017(new_n2366, n6385);
nor_4  g00018(new_n2367, n16223, new_n2366);
not_3  g00019(new_n2368, n16223);
nor_4  g00020(new_n2369, new_n2368, n6385);
not_3  g00021(new_n2370, n20138);
nor_4  g00022(new_n2371, new_n2370, n19494);
not_3  g00023(new_n2372, n19494);
nor_4  g00024(new_n2373, n20138, new_n2372);
not_3  g00025(new_n2374_1, n9251);
nor_4  g00026(new_n2375, new_n2374_1, n2387);
not_3  g00027(new_n2376, new_n2375);
nor_4  g00028(new_n2377, new_n2376, new_n2373);
nor_4  g00029(new_n2378, new_n2377, new_n2371);
nor_4  g00030(new_n2379, new_n2378, new_n2369);
nor_4  g00031(new_n2380, new_n2379, new_n2367);
nand_4 g00032(new_n2381, new_n2380, new_n2365);
nand_4 g00033(new_n2382, new_n2381, new_n2363_1);
nand_4 g00034(new_n2383, new_n2382, new_n2360);
nand_4 g00035(new_n2384, new_n2383, new_n2358);
nand_4 g00036(new_n2385, new_n2384, new_n2355_1);
nand_4 g00037(new_n2386, new_n2385, new_n2353);
xor_3  g00038(new_n2387_1, new_n2386, new_n2351);
nand_4 g00039(new_n2388_1, n13781, n5704);
not_3  g00040(new_n2389, n5704);
not_3  g00041(new_n2390, n13781);
nand_4 g00042(new_n2391, new_n2390, new_n2389);
nand_4 g00043(new_n2392, new_n2391, new_n2388_1);
not_3  g00044(new_n2393, new_n2392);
not_3  g00045(new_n2394, new_n2388_1);
xnor_3 g00046(new_n2395, n18409, n11486);
xnor_3 g00047(new_n2396, new_n2395, new_n2394);
nor_4  g00048(new_n2397, new_n2396, new_n2393);
not_3  g00049(new_n2398, new_n2397);
nor_4  g00050(new_n2399, n16722, n13708);
nand_4 g00051(new_n2400, n16722, n13708);
not_3  g00052(new_n2401, new_n2400);
nor_4  g00053(new_n2402, new_n2401, new_n2399);
not_3  g00054(new_n2403, new_n2402);
nor_4  g00055(new_n2404, n18409, n11486);
not_3  g00056(new_n2405, new_n2404);
not_3  g00057(new_n2406, new_n2395);
nand_4 g00058(new_n2407, new_n2406, new_n2388_1);
nand_4 g00059(new_n2408, new_n2407, new_n2405);
xnor_3 g00060(new_n2409_1, new_n2408, new_n2403);
not_3  g00061(new_n2410, new_n2409_1);
nor_4  g00062(new_n2411, new_n2410, new_n2398);
not_3  g00063(new_n2412, new_n2411);
xor_3  g00064(new_n2413, n19911, n3480);
not_3  g00065(new_n2414, new_n2399);
nand_4 g00066(new_n2415, new_n2408, new_n2402);
nand_4 g00067(new_n2416_1, new_n2415, new_n2414);
xnor_3 g00068(new_n2417, new_n2416_1, new_n2413);
nor_4  g00069(new_n2418, new_n2417, new_n2412);
xor_3  g00070(new_n2419, n3018, n2731);
nor_4  g00071(new_n2420_1, n19911, n3480);
not_3  g00072(new_n2421_1, new_n2420_1);
nand_4 g00073(new_n2422, new_n2416_1, new_n2413);
nand_4 g00074(new_n2423, new_n2422, new_n2421_1);
nor_4  g00075(new_n2424, new_n2423, new_n2419);
not_3  g00076(new_n2425, new_n2419);
not_3  g00077(new_n2426, n3480);
xor_3  g00078(new_n2427, n19911, new_n2426);
not_3  g00079(new_n2428, new_n2416_1);
nor_4  g00080(new_n2429, new_n2428, new_n2427);
nor_4  g00081(new_n2430, new_n2429, new_n2420_1);
nor_4  g00082(new_n2431, new_n2430, new_n2425);
nor_4  g00083(new_n2432, new_n2431, new_n2424);
nand_4 g00084(new_n2433, new_n2432, new_n2418);
xor_3  g00085(new_n2434, n26660, n18907);
nor_4  g00086(new_n2435, n3018, n2731);
not_3  g00087(new_n2436, new_n2435);
nand_4 g00088(new_n2437, new_n2423, new_n2419);
nand_4 g00089(new_n2438, new_n2437, new_n2436);
xnor_3 g00090(new_n2439, new_n2438, new_n2434);
nor_4  g00091(new_n2440_1, new_n2439, new_n2433);
xor_3  g00092(new_n2441, n22332, n13783);
not_3  g00093(new_n2442, new_n2441);
not_3  g00094(new_n2443, n18907);
not_3  g00095(new_n2444_1, n26660);
nand_4 g00096(new_n2445, new_n2444_1, new_n2443);
nand_4 g00097(new_n2446, new_n2438, new_n2434);
nand_4 g00098(new_n2447, new_n2446, new_n2445);
xnor_3 g00099(new_n2448, new_n2447, new_n2442);
xnor_3 g00100(new_n2449, new_n2448, new_n2440_1);
xor_3  g00101(new_n2450, n13490, n7751);
nor_4  g00102(new_n2451, n26823, n22660);
not_3  g00103(new_n2452, new_n2451);
xor_3  g00104(new_n2453, n26823, n22660);
nor_4  g00105(new_n2454, n4812, n1777);
not_3  g00106(new_n2455, new_n2454);
nand_4 g00107(new_n2456, n4812, n1777);
not_3  g00108(new_n2457, new_n2456);
nor_4  g00109(new_n2458, new_n2457, new_n2454);
nor_4  g00110(new_n2459, n24278, n8745);
not_3  g00111(new_n2460, new_n2459);
nand_4 g00112(new_n2461, n24278, n8745);
not_3  g00113(new_n2462, new_n2461);
nor_4  g00114(new_n2463, new_n2462, new_n2459);
nor_4  g00115(new_n2464, n24618, n15636);
not_3  g00116(new_n2465, new_n2464);
nand_4 g00117(new_n2466, n24618, n15636);
not_3  g00118(new_n2467, new_n2466);
nor_4  g00119(new_n2468, new_n2467, new_n2464);
nand_4 g00120(new_n2469, n20077, n3952);
not_3  g00121(new_n2470, new_n2469);
nor_4  g00122(new_n2471, n20077, n3952);
nand_4 g00123(new_n2472, n12315, n6794);
nor_4  g00124(new_n2473, new_n2472, new_n2471);
nor_4  g00125(new_n2474, new_n2473, new_n2470);
nand_4 g00126(new_n2475, new_n2474, new_n2468);
nand_4 g00127(new_n2476, new_n2475, new_n2465);
nand_4 g00128(new_n2477, new_n2476, new_n2463);
nand_4 g00129(new_n2478, new_n2477, new_n2460);
nand_4 g00130(new_n2479_1, new_n2478, new_n2458);
nand_4 g00131(new_n2480, new_n2479_1, new_n2455);
nand_4 g00132(new_n2481, new_n2480, new_n2453);
nand_4 g00133(new_n2482, new_n2481, new_n2452);
xnor_3 g00134(new_n2483, new_n2482, new_n2450);
xnor_3 g00135(new_n2484, new_n2483, new_n2449);
not_3  g00136(new_n2485, new_n2484);
xnor_3 g00137(new_n2486, new_n2439, new_n2433);
not_3  g00138(new_n2487, new_n2453);
not_3  g00139(new_n2488, new_n2458);
not_3  g00140(new_n2489, new_n2478);
nor_4  g00141(new_n2490, new_n2489, new_n2488);
nor_4  g00142(new_n2491, new_n2490, new_n2454);
nor_4  g00143(new_n2492, new_n2491, new_n2487);
nor_4  g00144(new_n2493, new_n2480, new_n2453);
nor_4  g00145(new_n2494, new_n2493, new_n2492);
nand_4 g00146(new_n2495, new_n2494, new_n2486);
xnor_3 g00147(new_n2496, new_n2432, new_n2418);
xnor_3 g00148(new_n2497, new_n2478, new_n2488);
nand_4 g00149(new_n2498, new_n2497, new_n2496);
not_3  g00150(new_n2499, new_n2497);
xnor_3 g00151(new_n2500, new_n2499, new_n2496);
xnor_3 g00152(new_n2501, new_n2417, new_n2412);
xnor_3 g00153(new_n2502, new_n2476, new_n2463);
not_3  g00154(new_n2503, new_n2502);
nand_4 g00155(new_n2504, new_n2503, new_n2501);
xnor_3 g00156(new_n2505, new_n2409_1, new_n2397);
not_3  g00157(new_n2506, new_n2505);
xnor_3 g00158(new_n2507, new_n2474, new_n2468);
nor_4  g00159(new_n2508, new_n2507, new_n2506);
not_3  g00160(new_n2509, new_n2508);
not_3  g00161(new_n2510, new_n2507);
xnor_3 g00162(new_n2511, new_n2510, new_n2505);
xnor_3 g00163(new_n2512, n12315, n6794);
nor_4  g00164(new_n2513_1, new_n2512, new_n2392);
xnor_3 g00165(new_n2514, n20077, n3952);
xnor_3 g00166(new_n2515_1, new_n2514, new_n2472);
not_3  g00167(new_n2516, new_n2515_1);
nor_4  g00168(new_n2517, new_n2516, new_n2513_1);
not_3  g00169(new_n2518, new_n2391);
nor_4  g00170(new_n2519, new_n2407, new_n2518);
nor_4  g00171(new_n2520, new_n2519, new_n2397);
not_3  g00172(new_n2521, new_n2513_1);
nor_4  g00173(new_n2522, new_n2514, new_n2521);
nor_4  g00174(new_n2523, new_n2522, new_n2517);
not_3  g00175(new_n2524, new_n2523);
nor_4  g00176(new_n2525, new_n2524, new_n2520);
nor_4  g00177(new_n2526, new_n2525, new_n2517);
nor_4  g00178(new_n2527, new_n2526, new_n2511);
not_3  g00179(new_n2528, new_n2527);
nand_4 g00180(new_n2529, new_n2528, new_n2509);
xnor_3 g00181(new_n2530, new_n2502, new_n2501);
nand_4 g00182(new_n2531, new_n2530, new_n2529);
nand_4 g00183(new_n2532, new_n2531, new_n2504);
nand_4 g00184(new_n2533_1, new_n2532, new_n2500);
nand_4 g00185(new_n2534, new_n2533_1, new_n2498);
xnor_3 g00186(new_n2535_1, new_n2494, new_n2486);
not_3  g00187(new_n2536, new_n2535_1);
nand_4 g00188(new_n2537_1, new_n2536, new_n2534);
nand_4 g00189(new_n2538, new_n2537_1, new_n2495);
xnor_3 g00190(new_n2539, new_n2538, new_n2485);
xnor_3 g00191(new_n2540, new_n2539, new_n2387_1);
xor_3  g00192(new_n2541, new_n2384, new_n2355_1);
xnor_3 g00193(new_n2542, new_n2536, new_n2534);
nor_4  g00194(new_n2543, new_n2542, new_n2541);
not_3  g00195(new_n2544, new_n2543);
xnor_3 g00196(new_n2545, new_n2535_1, new_n2534);
xnor_3 g00197(new_n2546, new_n2545, new_n2541);
xor_3  g00198(new_n2547_1, new_n2382, new_n2360);
xnor_3 g00199(new_n2548, new_n2532, new_n2500);
nor_4  g00200(new_n2549, new_n2548, new_n2547_1);
not_3  g00201(new_n2550, new_n2549);
xnor_3 g00202(new_n2551, new_n2497, new_n2496);
xnor_3 g00203(new_n2552, new_n2532, new_n2551);
xnor_3 g00204(new_n2553_1, new_n2552, new_n2547_1);
xor_3  g00205(new_n2554, n26913, n3136);
xor_3  g00206(new_n2555_1, new_n2380, new_n2554);
not_3  g00207(new_n2556, new_n2555_1);
xnor_3 g00208(new_n2557, new_n2530, new_n2529);
nor_4  g00209(new_n2558, new_n2557, new_n2556);
not_3  g00210(new_n2559, new_n2558);
not_3  g00211(new_n2560_1, new_n2557);
xnor_3 g00212(new_n2561_1, new_n2560_1, new_n2555_1);
not_3  g00213(new_n2562, new_n2561_1);
xnor_3 g00214(new_n2563, new_n2526, new_n2511);
nor_4  g00215(new_n2564, new_n2369, new_n2367);
not_3  g00216(new_n2565, new_n2564);
xor_3  g00217(new_n2566, new_n2565, new_n2378);
not_3  g00218(new_n2567, new_n2566);
nor_4  g00219(new_n2568, new_n2567, new_n2563);
not_3  g00220(new_n2569, new_n2563);
xnor_3 g00221(new_n2570_1, new_n2566, new_n2569);
not_3  g00222(new_n2571, n2387);
xor_3  g00223(new_n2572, n9251, new_n2571);
not_3  g00224(new_n2573_1, new_n2512);
xor_3  g00225(new_n2574, new_n2573_1, new_n2392);
nor_4  g00226(new_n2575, new_n2574, new_n2572);
nor_4  g00227(new_n2576, new_n2373, new_n2371);
xor_3  g00228(new_n2577, new_n2576, new_n2376);
nor_4  g00229(new_n2578_1, new_n2577, new_n2575);
xor_3  g00230(new_n2579, new_n2523, new_n2520);
xnor_3 g00231(new_n2580, new_n2577, new_n2575);
nor_4  g00232(new_n2581, new_n2580, new_n2579);
nor_4  g00233(new_n2582_1, new_n2581, new_n2578_1);
nor_4  g00234(new_n2583, new_n2582_1, new_n2570_1);
nor_4  g00235(new_n2584, new_n2583, new_n2568);
not_3  g00236(new_n2585, new_n2584);
nand_4 g00237(new_n2586, new_n2585, new_n2562);
nand_4 g00238(new_n2587, new_n2586, new_n2559);
nand_4 g00239(new_n2588, new_n2587, new_n2553_1);
nand_4 g00240(new_n2589, new_n2588, new_n2550);
nand_4 g00241(new_n2590, new_n2589, new_n2546);
nand_4 g00242(new_n2591, new_n2590, new_n2544);
xor_3  g00243(n7, new_n2591, new_n2540);
xnor_3 g00244(new_n2593, n3618, n1681);
xor_3  g00245(new_n2594, new_n2593, n4588);
not_3  g00246(new_n2595, new_n2594);
not_3  g00247(new_n2596, n22201);
xor_3  g00248(new_n2597, n22843, n583);
not_3  g00249(new_n2598, new_n2597);
xor_3  g00250(new_n2599, new_n2598, new_n2596);
xor_3  g00251(n50, new_n2599, new_n2595);
not_3  g00252(new_n2601, n21687);
xor_3  g00253(new_n2602_1, n19922, n6773);
not_3  g00254(new_n2603, new_n2602_1);
xor_3  g00255(new_n2604, new_n2603, new_n2601);
xor_3  g00256(new_n2605, n21398, n14090);
nand_4 g00257(new_n2606, new_n2605, n25926);
not_3  g00258(new_n2607, new_n2606);
nor_4  g00259(new_n2608, new_n2605, n25926);
nor_4  g00260(new_n2609, new_n2608, new_n2607);
xor_3  g00261(n55, new_n2609, new_n2604);
not_3  g00262(new_n2611, n25365);
xor_3  g00263(new_n2612, n20040, n9396);
nor_4  g00264(new_n2613, n19531, n1999);
xor_3  g00265(new_n2614, n19531, n1999);
not_3  g00266(new_n2615, new_n2614);
nor_4  g00267(new_n2616, n25168, n18345);
xor_3  g00268(new_n2617, n25168, n18345);
not_3  g00269(new_n2618, new_n2617);
not_3  g00270(new_n2619_1, n9318);
not_3  g00271(new_n2620, n13190);
nand_4 g00272(new_n2621, new_n2620, new_n2619_1);
xor_3  g00273(new_n2622, n13190, n9318);
nor_4  g00274(new_n2623, n19477, n3460);
not_3  g00275(new_n2624, new_n2623);
xor_3  g00276(new_n2625, n19477, n3460);
nor_4  g00277(new_n2626, n11223, n5226);
not_3  g00278(new_n2627, new_n2626);
xor_3  g00279(new_n2628, n11223, n5226);
nor_4  g00280(new_n2629, n17664, n5115);
not_3  g00281(new_n2630, new_n2629);
nand_4 g00282(new_n2631, n17664, n5115);
not_3  g00283(new_n2632, new_n2631);
nor_4  g00284(new_n2633, new_n2632, new_n2629);
nor_4  g00285(new_n2634, n26572, n23369);
not_3  g00286(new_n2635, new_n2634);
nand_4 g00287(new_n2636, n26572, n23369);
not_3  g00288(new_n2637, new_n2636);
nor_4  g00289(new_n2638, new_n2637, new_n2634);
nor_4  g00290(new_n2639, n11667, n1136);
not_3  g00291(new_n2640, new_n2639);
nand_4 g00292(new_n2641, n21398, n19234);
nand_4 g00293(new_n2642, n11667, n1136);
not_3  g00294(new_n2643, new_n2642);
nor_4  g00295(new_n2644, new_n2643, new_n2639);
nand_4 g00296(new_n2645, new_n2644, new_n2641);
nand_4 g00297(new_n2646_1, new_n2645, new_n2640);
nand_4 g00298(new_n2647, new_n2646_1, new_n2638);
nand_4 g00299(new_n2648, new_n2647, new_n2635);
nand_4 g00300(new_n2649, new_n2648, new_n2633);
nand_4 g00301(new_n2650, new_n2649, new_n2630);
nand_4 g00302(new_n2651, new_n2650, new_n2628);
nand_4 g00303(new_n2652, new_n2651, new_n2627);
nand_4 g00304(new_n2653, new_n2652, new_n2625);
nand_4 g00305(new_n2654, new_n2653, new_n2624);
nand_4 g00306(new_n2655, new_n2654, new_n2622);
nand_4 g00307(new_n2656, new_n2655, new_n2621);
not_3  g00308(new_n2657, new_n2656);
nor_4  g00309(new_n2658, new_n2657, new_n2618);
nor_4  g00310(new_n2659_1, new_n2658, new_n2616);
nor_4  g00311(new_n2660, new_n2659_1, new_n2615);
nor_4  g00312(new_n2661_1, new_n2660, new_n2613);
not_3  g00313(new_n2662, new_n2661_1);
nor_4  g00314(new_n2663, new_n2662, new_n2612);
not_3  g00315(new_n2664, new_n2612);
nor_4  g00316(new_n2665, new_n2661_1, new_n2664);
nor_4  g00317(new_n2666, new_n2665, new_n2663);
xnor_3 g00318(new_n2667, new_n2666, new_n2611);
not_3  g00319(new_n2668, new_n2667);
not_3  g00320(new_n2669, n14704);
not_3  g00321(new_n2670, new_n2659_1);
nor_4  g00322(new_n2671, new_n2670, new_n2614);
nor_4  g00323(new_n2672, new_n2671, new_n2660);
nor_4  g00324(new_n2673, new_n2672, new_n2669);
not_3  g00325(new_n2674, new_n2673);
not_3  g00326(new_n2675, new_n2672);
nor_4  g00327(new_n2676, new_n2675, n14704);
nor_4  g00328(new_n2677, new_n2676, new_n2673);
not_3  g00329(new_n2678, n19270);
nor_4  g00330(new_n2679, new_n2656, new_n2617);
nor_4  g00331(new_n2680_1, new_n2679, new_n2658);
nor_4  g00332(new_n2681, new_n2680_1, new_n2678);
not_3  g00333(new_n2682, new_n2681);
xnor_3 g00334(new_n2683, new_n2680_1, new_n2678);
not_3  g00335(new_n2684, new_n2683);
not_3  g00336(new_n2685, n8687);
not_3  g00337(new_n2686, new_n2622);
xnor_3 g00338(new_n2687, new_n2654, new_n2686);
nor_4  g00339(new_n2688, new_n2687, new_n2685);
not_3  g00340(new_n2689, new_n2688);
not_3  g00341(new_n2690, new_n2625);
xnor_3 g00342(new_n2691, new_n2652, new_n2690);
not_3  g00343(new_n2692, new_n2691);
nor_4  g00344(new_n2693_1, new_n2692, n24768);
not_3  g00345(new_n2694, n24768);
nor_4  g00346(new_n2695, new_n2691, new_n2694);
nor_4  g00347(new_n2696, new_n2695, new_n2693_1);
not_3  g00348(new_n2697, new_n2696);
xnor_3 g00349(new_n2698, new_n2650, new_n2628);
nor_4  g00350(new_n2699, new_n2698, n26483);
xnor_3 g00351(new_n2700, new_n2698, n26483);
not_3  g00352(new_n2701, n15979);
not_3  g00353(new_n2702, new_n2633);
xnor_3 g00354(new_n2703_1, new_n2648, new_n2702);
nor_4  g00355(new_n2704, new_n2703_1, new_n2701);
not_3  g00356(new_n2705, new_n2704);
xnor_3 g00357(new_n2706_1, new_n2648, new_n2633);
nor_4  g00358(new_n2707, new_n2706_1, n15979);
nor_4  g00359(new_n2708, new_n2707, new_n2704);
not_3  g00360(new_n2709, n8638);
not_3  g00361(new_n2710, new_n2638);
xnor_3 g00362(new_n2711_1, new_n2646_1, new_n2710);
nor_4  g00363(new_n2712, new_n2711_1, new_n2709);
not_3  g00364(new_n2713, new_n2712);
not_3  g00365(new_n2714, new_n2641);
nand_4 g00366(new_n2715, new_n2642, new_n2640);
xnor_3 g00367(new_n2716, new_n2715, new_n2714);
nor_4  g00368(new_n2717, new_n2716, n16247);
not_3  g00369(new_n2718, new_n2717);
not_3  g00370(new_n2719, n23541);
xnor_3 g00371(new_n2720, n21398, n19234);
nor_4  g00372(new_n2721, new_n2720, new_n2719);
not_3  g00373(new_n2722, new_n2721);
not_3  g00374(new_n2723, n16247);
nor_4  g00375(new_n2724, new_n2715, new_n2714);
nor_4  g00376(new_n2725, new_n2644, new_n2641);
nor_4  g00377(new_n2726, new_n2725, new_n2724);
nor_4  g00378(new_n2727, new_n2726, new_n2723);
nor_4  g00379(new_n2728, new_n2727, new_n2717);
nand_4 g00380(new_n2729, new_n2728, new_n2722);
nand_4 g00381(new_n2730, new_n2729, new_n2718);
xnor_3 g00382(new_n2731_1, new_n2646_1, new_n2638);
nor_4  g00383(new_n2732, new_n2731_1, n8638);
nor_4  g00384(new_n2733, new_n2732, new_n2712);
not_3  g00385(new_n2734, new_n2733);
nor_4  g00386(new_n2735, new_n2734, new_n2730);
not_3  g00387(new_n2736, new_n2735);
nand_4 g00388(new_n2737, new_n2736, new_n2713);
nand_4 g00389(new_n2738, new_n2737, new_n2708);
nand_4 g00390(new_n2739, new_n2738, new_n2705);
nor_4  g00391(new_n2740, new_n2739, new_n2700);
nor_4  g00392(new_n2741, new_n2740, new_n2699);
nor_4  g00393(new_n2742, new_n2741, new_n2697);
nor_4  g00394(new_n2743_1, new_n2742, new_n2693_1);
not_3  g00395(new_n2744, new_n2687);
nor_4  g00396(new_n2745, new_n2744, n8687);
nor_4  g00397(new_n2746, new_n2745, new_n2688);
nand_4 g00398(new_n2747, new_n2746, new_n2743_1);
nand_4 g00399(new_n2748, new_n2747, new_n2689);
nand_4 g00400(new_n2749, new_n2748, new_n2684);
nand_4 g00401(new_n2750, new_n2749, new_n2682);
nand_4 g00402(new_n2751, new_n2750, new_n2677);
nand_4 g00403(new_n2752, new_n2751, new_n2674);
nand_4 g00404(new_n2753, new_n2752, new_n2668);
not_3  g00405(new_n2754, new_n2753);
nor_4  g00406(new_n2755, new_n2752, new_n2668);
nor_4  g00407(new_n2756, new_n2755, new_n2754);
not_3  g00408(new_n2757, n13951);
not_3  g00409(new_n2758, n8439);
not_3  g00410(new_n2759, n5579);
not_3  g00411(new_n2760, n16971);
nor_4  g00412(new_n2761_1, n18151, n11503);
nand_4 g00413(new_n2762, new_n2761_1, new_n2760);
nor_4  g00414(new_n2763, new_n2762, n10411);
not_3  g00415(new_n2764, new_n2763);
nor_4  g00416(new_n2765, new_n2764, n23430);
nand_4 g00417(new_n2766, new_n2765, new_n2759);
nor_4  g00418(new_n2767, new_n2766, n25523);
nand_4 g00419(new_n2768, new_n2767, new_n2758);
nor_4  g00420(new_n2769, new_n2768, n22793);
xor_3  g00421(new_n2770, new_n2769, new_n2757);
not_3  g00422(new_n2771, new_n2770);
xor_3  g00423(new_n2772, n22270, n2944);
not_3  g00424(new_n2773, new_n2772);
nor_4  g00425(new_n2774_1, n8806, n767);
xor_3  g00426(new_n2775, n8806, n767);
not_3  g00427(new_n2776, new_n2775);
nor_4  g00428(new_n2777, n7330, n2479);
xor_3  g00429(new_n2778, n7330, n2479);
not_3  g00430(new_n2779_1, new_n2778);
not_3  g00431(new_n2780, n9372);
not_3  g00432(new_n2781, n22492);
nand_4 g00433(new_n2782, new_n2781, new_n2780);
xor_3  g00434(new_n2783_1, n22492, n9372);
nor_4  g00435(new_n2784, n12821, n6596);
not_3  g00436(new_n2785, new_n2784);
xor_3  g00437(new_n2786, n12821, n6596);
nor_4  g00438(new_n2787, n15289, n3468);
not_3  g00439(new_n2788, new_n2787);
xor_3  g00440(new_n2789, n15289, n3468);
nor_4  g00441(new_n2790, n18558, n6556);
not_3  g00442(new_n2791, new_n2790);
xor_3  g00443(new_n2792, n18558, n6556);
nor_4  g00444(new_n2793, n22871, n7149);
not_3  g00445(new_n2794, new_n2793);
xor_3  g00446(new_n2795, n22871, n7149);
nor_4  g00447(new_n2796, n14275, n14148);
not_3  g00448(new_n2797, new_n2796);
nand_4 g00449(new_n2798, n25023, n1152);
nand_4 g00450(new_n2799, n14275, n14148);
not_3  g00451(new_n2800, new_n2799);
nor_4  g00452(new_n2801, new_n2800, new_n2796);
nand_4 g00453(new_n2802, new_n2801, new_n2798);
nand_4 g00454(new_n2803, new_n2802, new_n2797);
nand_4 g00455(new_n2804, new_n2803, new_n2795);
nand_4 g00456(new_n2805, new_n2804, new_n2794);
nand_4 g00457(new_n2806, new_n2805, new_n2792);
nand_4 g00458(new_n2807, new_n2806, new_n2791);
nand_4 g00459(new_n2808, new_n2807, new_n2789);
nand_4 g00460(new_n2809_1, new_n2808, new_n2788);
nand_4 g00461(new_n2810, new_n2809_1, new_n2786);
nand_4 g00462(new_n2811, new_n2810, new_n2785);
nand_4 g00463(new_n2812, new_n2811, new_n2783_1);
nand_4 g00464(new_n2813, new_n2812, new_n2782);
not_3  g00465(new_n2814, new_n2813);
nor_4  g00466(new_n2815, new_n2814, new_n2779_1);
nor_4  g00467(new_n2816_1, new_n2815, new_n2777);
nor_4  g00468(new_n2817, new_n2816_1, new_n2776);
nor_4  g00469(new_n2818, new_n2817, new_n2774_1);
xnor_3 g00470(new_n2819, new_n2818, new_n2773);
nor_4  g00471(new_n2820, new_n2819, new_n2771);
xnor_3 g00472(new_n2821, new_n2818, new_n2772);
nor_4  g00473(new_n2822, new_n2821, new_n2770);
nor_4  g00474(new_n2823, new_n2822, new_n2820);
not_3  g00475(new_n2824, new_n2823);
xor_3  g00476(new_n2825, new_n2768, n22793);
xnor_3 g00477(new_n2826_1, new_n2816_1, new_n2775);
nand_4 g00478(new_n2827, new_n2826_1, new_n2825);
not_3  g00479(new_n2828, new_n2827);
xnor_3 g00480(new_n2829, new_n2826_1, new_n2825);
xor_3  g00481(new_n2830, new_n2767, new_n2758);
xnor_3 g00482(new_n2831, new_n2813, new_n2778);
not_3  g00483(new_n2832, new_n2831);
nor_4  g00484(new_n2833, new_n2832, new_n2830);
not_3  g00485(new_n2834, new_n2833);
xnor_3 g00486(new_n2835, new_n2831, new_n2830);
xor_3  g00487(new_n2836, new_n2766, n25523);
not_3  g00488(new_n2837, new_n2783_1);
xnor_3 g00489(new_n2838, new_n2811, new_n2837);
nor_4  g00490(new_n2839, new_n2838, new_n2836);
not_3  g00491(new_n2840, new_n2839);
not_3  g00492(new_n2841, new_n2836);
xnor_3 g00493(new_n2842, new_n2811, new_n2783_1);
nor_4  g00494(new_n2843, new_n2842, new_n2841);
nor_4  g00495(new_n2844, new_n2843, new_n2839);
xor_3  g00496(new_n2845, new_n2765, new_n2759);
not_3  g00497(new_n2846, new_n2786);
xnor_3 g00498(new_n2847, new_n2809_1, new_n2846);
nor_4  g00499(new_n2848, new_n2847, new_n2845);
not_3  g00500(new_n2849, new_n2848);
not_3  g00501(new_n2850, new_n2845);
xnor_3 g00502(new_n2851, new_n2809_1, new_n2786);
nor_4  g00503(new_n2852, new_n2851, new_n2850);
nor_4  g00504(new_n2853_1, new_n2852, new_n2848);
not_3  g00505(new_n2854, n23430);
xor_3  g00506(new_n2855, new_n2763, new_n2854);
not_3  g00507(new_n2856, new_n2789);
xnor_3 g00508(new_n2857, new_n2807, new_n2856);
nor_4  g00509(new_n2858_1, new_n2857, new_n2855);
not_3  g00510(new_n2859, new_n2858_1);
not_3  g00511(new_n2860_1, n10411);
xor_3  g00512(new_n2861, new_n2762, new_n2860_1);
xnor_3 g00513(new_n2862, new_n2805, new_n2792);
nand_4 g00514(new_n2863, new_n2862, new_n2861);
not_3  g00515(new_n2864, new_n2863);
nor_4  g00516(new_n2865, new_n2862, new_n2861);
nor_4  g00517(new_n2866, new_n2865, new_n2864);
xor_3  g00518(new_n2867, new_n2761_1, new_n2760);
not_3  g00519(new_n2868, new_n2803);
xnor_3 g00520(new_n2869, new_n2868, new_n2795);
nor_4  g00521(new_n2870, new_n2869, new_n2867);
not_3  g00522(new_n2871, new_n2870);
not_3  g00523(new_n2872, new_n2867);
xnor_3 g00524(new_n2873, new_n2803, new_n2795);
nor_4  g00525(new_n2874, new_n2873, new_n2872);
nor_4  g00526(new_n2875, new_n2874, new_n2870);
xor_3  g00527(new_n2876, n18151, n11503);
not_3  g00528(new_n2877, new_n2802);
nor_4  g00529(new_n2878, new_n2801, new_n2798);
nor_4  g00530(new_n2879, new_n2878, new_n2877);
nor_4  g00531(new_n2880, new_n2879, new_n2876);
not_3  g00532(new_n2881, new_n2880);
not_3  g00533(new_n2882, n18151);
xor_3  g00534(new_n2883, n25023, n1152);
nand_4 g00535(new_n2884, new_n2883, new_n2882);
not_3  g00536(new_n2885, new_n2884);
not_3  g00537(new_n2886_1, new_n2879);
xnor_3 g00538(new_n2887_1, new_n2886_1, new_n2876);
nand_4 g00539(new_n2888, new_n2887_1, new_n2885);
nand_4 g00540(new_n2889, new_n2888, new_n2881);
nand_4 g00541(new_n2890, new_n2889, new_n2875);
nand_4 g00542(new_n2891, new_n2890, new_n2871);
nand_4 g00543(new_n2892, new_n2891, new_n2866);
nand_4 g00544(new_n2893, new_n2892, new_n2863);
not_3  g00545(new_n2894, new_n2855);
xnor_3 g00546(new_n2895, new_n2807, new_n2789);
nor_4  g00547(new_n2896, new_n2895, new_n2894);
nor_4  g00548(new_n2897, new_n2896, new_n2858_1);
nand_4 g00549(new_n2898, new_n2897, new_n2893);
nand_4 g00550(new_n2899, new_n2898, new_n2859);
nand_4 g00551(new_n2900, new_n2899, new_n2853_1);
nand_4 g00552(new_n2901, new_n2900, new_n2849);
nand_4 g00553(new_n2902, new_n2901, new_n2844);
nand_4 g00554(new_n2903, new_n2902, new_n2840);
nand_4 g00555(new_n2904, new_n2903, new_n2835);
nand_4 g00556(new_n2905, new_n2904, new_n2834);
nor_4  g00557(new_n2906, new_n2905, new_n2829);
nor_4  g00558(new_n2907, new_n2906, new_n2828);
xnor_3 g00559(new_n2908, new_n2907, new_n2824);
xnor_3 g00560(new_n2909, new_n2908, new_n2756);
not_3  g00561(new_n2910, new_n2751);
nor_4  g00562(new_n2911, new_n2750, new_n2677);
nor_4  g00563(new_n2912, new_n2911, new_n2910);
not_3  g00564(new_n2913, new_n2912);
xnor_3 g00565(new_n2914, new_n2905, new_n2829);
nor_4  g00566(new_n2915, new_n2914, new_n2913);
xnor_3 g00567(new_n2916, new_n2914, new_n2913);
xnor_3 g00568(new_n2917, new_n2748, new_n2684);
not_3  g00569(new_n2918, new_n2904);
nor_4  g00570(new_n2919, new_n2903, new_n2835);
nor_4  g00571(new_n2920, new_n2919, new_n2918);
nand_4 g00572(new_n2921, new_n2920, new_n2917);
not_3  g00573(new_n2922, new_n2917);
xnor_3 g00574(new_n2923, new_n2920, new_n2922);
xnor_3 g00575(new_n2924, new_n2746, new_n2743_1);
not_3  g00576(new_n2925, new_n2924);
xnor_3 g00577(new_n2926, new_n2901, new_n2844);
nor_4  g00578(new_n2927, new_n2926, new_n2925);
not_3  g00579(new_n2928, new_n2927);
xnor_3 g00580(new_n2929_1, new_n2926, new_n2924);
xnor_3 g00581(new_n2930, new_n2741, new_n2697);
not_3  g00582(new_n2931, new_n2930);
xnor_3 g00583(new_n2932, new_n2899, new_n2853_1);
not_3  g00584(new_n2933, new_n2932);
nor_4  g00585(new_n2934, new_n2933, new_n2931);
xnor_3 g00586(new_n2935, new_n2932, new_n2930);
xnor_3 g00587(new_n2936, new_n2739, new_n2700);
not_3  g00588(new_n2937, new_n2936);
xnor_3 g00589(new_n2938, new_n2857, new_n2855);
xnor_3 g00590(new_n2939, new_n2938, new_n2893);
nand_4 g00591(new_n2940, new_n2939, new_n2937);
xnor_3 g00592(new_n2941, new_n2939, new_n2936);
xnor_3 g00593(new_n2942, new_n2891, new_n2866);
not_3  g00594(new_n2943, new_n2942);
xnor_3 g00595(new_n2944_1, new_n2737, new_n2708);
nand_4 g00596(new_n2945, new_n2944_1, new_n2943);
xnor_3 g00597(new_n2946, new_n2944_1, new_n2942);
xnor_3 g00598(new_n2947, new_n2889, new_n2875);
not_3  g00599(new_n2948_1, new_n2947);
not_3  g00600(new_n2949, new_n2730);
nor_4  g00601(new_n2950, new_n2733, new_n2949);
nor_4  g00602(new_n2951, new_n2950, new_n2735);
not_3  g00603(new_n2952, new_n2951);
nor_4  g00604(new_n2953, new_n2952, new_n2948_1);
xnor_3 g00605(new_n2954, new_n2951, new_n2947);
xnor_3 g00606(new_n2955, new_n2879, new_n2876);
nor_4  g00607(new_n2956, new_n2955, new_n2884);
nor_4  g00608(new_n2957, new_n2887_1, new_n2885);
nor_4  g00609(new_n2958, new_n2957, new_n2956);
xnor_3 g00610(new_n2959, new_n2728, new_n2722);
not_3  g00611(new_n2960, new_n2959);
nand_4 g00612(new_n2961_1, new_n2960, new_n2958);
xor_3  g00613(new_n2962, new_n2720, new_n2719);
xnor_3 g00614(new_n2963, new_n2883, new_n2882);
nand_4 g00615(new_n2964, new_n2963, new_n2962);
xnor_3 g00616(new_n2965, new_n2959, new_n2958);
nand_4 g00617(new_n2966, new_n2965, new_n2964);
nand_4 g00618(new_n2967, new_n2966, new_n2961_1);
nor_4  g00619(new_n2968, new_n2967, new_n2954);
nor_4  g00620(new_n2969, new_n2968, new_n2953);
nand_4 g00621(new_n2970, new_n2969, new_n2946);
nand_4 g00622(new_n2971_1, new_n2970, new_n2945);
nand_4 g00623(new_n2972, new_n2971_1, new_n2941);
nand_4 g00624(new_n2973, new_n2972, new_n2940);
nor_4  g00625(new_n2974, new_n2973, new_n2935);
nor_4  g00626(new_n2975, new_n2974, new_n2934);
nand_4 g00627(new_n2976, new_n2975, new_n2929_1);
nand_4 g00628(new_n2977, new_n2976, new_n2928);
nand_4 g00629(new_n2978_1, new_n2977, new_n2923);
nand_4 g00630(new_n2979_1, new_n2978_1, new_n2921);
nor_4  g00631(new_n2980, new_n2979_1, new_n2916);
nor_4  g00632(new_n2981, new_n2980, new_n2915);
xnor_3 g00633(n108, new_n2981, new_n2909);
not_3  g00634(new_n2983, n767);
xor_3  g00635(new_n2984, n22379, new_n2983);
not_3  g00636(new_n2985_1, n7330);
nand_4 g00637(new_n2986, new_n2985_1, n1662);
not_3  g00638(new_n2987, n1662);
xor_3  g00639(new_n2988, n7330, new_n2987);
not_3  g00640(new_n2989, n12875);
nor_4  g00641(new_n2990, n22492, new_n2989);
not_3  g00642(new_n2991, new_n2990);
xor_3  g00643(new_n2992, n22492, new_n2989);
not_3  g00644(new_n2993, n2035);
nor_4  g00645(new_n2994, n12821, new_n2993);
not_3  g00646(new_n2995, new_n2994);
xor_3  g00647(new_n2996, n12821, new_n2993);
not_3  g00648(new_n2997, n5213);
nor_4  g00649(new_n2998, new_n2997, n3468);
not_3  g00650(new_n2999_1, new_n2998);
not_3  g00651(new_n3000, n3468);
xor_3  g00652(new_n3001, n5213, new_n3000);
not_3  g00653(new_n3002, n4665);
nor_4  g00654(new_n3003, n18558, new_n3002);
xor_3  g00655(new_n3004, n18558, n4665);
not_3  g00656(new_n3005, n7149);
nor_4  g00657(new_n3006, n19005, new_n3005);
not_3  g00658(new_n3007, n19005);
nor_4  g00659(new_n3008, new_n3007, n7149);
not_3  g00660(new_n3009, n14148);
nor_4  g00661(new_n3010_1, new_n3009, n4326);
not_3  g00662(new_n3011, n4326);
nor_4  g00663(new_n3012, n14148, new_n3011);
not_3  g00664(new_n3013, n1152);
nor_4  g00665(new_n3014, n5438, new_n3013);
not_3  g00666(new_n3015, new_n3014);
nor_4  g00667(new_n3016, new_n3015, new_n3012);
nor_4  g00668(new_n3017_1, new_n3016, new_n3010_1);
nor_4  g00669(new_n3018_1, new_n3017_1, new_n3008);
nor_4  g00670(new_n3019, new_n3018_1, new_n3006);
not_3  g00671(new_n3020_1, new_n3019);
nor_4  g00672(new_n3021, new_n3020_1, new_n3004);
nor_4  g00673(new_n3022, new_n3021, new_n3003);
not_3  g00674(new_n3023, new_n3022);
nand_4 g00675(new_n3024, new_n3023, new_n3001);
nand_4 g00676(new_n3025, new_n3024, new_n2999_1);
nand_4 g00677(new_n3026, new_n3025, new_n2996);
nand_4 g00678(new_n3027, new_n3026, new_n2995);
nand_4 g00679(new_n3028, new_n3027, new_n2992);
nand_4 g00680(new_n3029, new_n3028, new_n2991);
nand_4 g00681(new_n3030_1, new_n3029, new_n2988);
nand_4 g00682(new_n3031, new_n3030_1, new_n2986);
xor_3  g00683(new_n3032, new_n3031, new_n2984);
xor_3  g00684(new_n3033, n10763, n6814);
nor_4  g00685(new_n3034, n19701, n7437);
xor_3  g00686(new_n3035, n19701, n7437);
not_3  g00687(new_n3036, new_n3035);
not_3  g00688(new_n3037, n20700);
not_3  g00689(new_n3038, n23529);
nand_4 g00690(new_n3039, new_n3038, new_n3037);
xor_3  g00691(new_n3040, n23529, n20700);
nor_4  g00692(new_n3041, n24620, n7099);
not_3  g00693(new_n3042, new_n3041);
xor_3  g00694(new_n3043, n24620, n7099);
nor_4  g00695(new_n3044, n12811, n5211);
not_3  g00696(new_n3045, new_n3044);
xor_3  g00697(new_n3046, n12811, n5211);
nor_4  g00698(new_n3047, n12956, n1118);
not_3  g00699(new_n3048, new_n3047);
xor_3  g00700(new_n3049, n12956, n1118);
nor_4  g00701(new_n3050, n25974, n18295);
not_3  g00702(new_n3051, new_n3050);
xor_3  g00703(new_n3052, n25974, n18295);
nor_4  g00704(new_n3053, n6502, n1630);
not_3  g00705(new_n3054, new_n3053);
nand_4 g00706(new_n3055, n15780, n1451);
nand_4 g00707(new_n3056, n6502, n1630);
not_3  g00708(new_n3057, new_n3056);
nor_4  g00709(new_n3058, new_n3057, new_n3053);
nand_4 g00710(new_n3059, new_n3058, new_n3055);
nand_4 g00711(new_n3060, new_n3059, new_n3054);
nand_4 g00712(new_n3061, new_n3060, new_n3052);
nand_4 g00713(new_n3062, new_n3061, new_n3051);
nand_4 g00714(new_n3063, new_n3062, new_n3049);
nand_4 g00715(new_n3064, new_n3063, new_n3048);
nand_4 g00716(new_n3065, new_n3064, new_n3046);
nand_4 g00717(new_n3066, new_n3065, new_n3045);
nand_4 g00718(new_n3067_1, new_n3066, new_n3043);
nand_4 g00719(new_n3068, new_n3067_1, new_n3042);
nand_4 g00720(new_n3069, new_n3068, new_n3040);
nand_4 g00721(new_n3070, new_n3069, new_n3039);
not_3  g00722(new_n3071, new_n3070);
nor_4  g00723(new_n3072, new_n3071, new_n3036);
nor_4  g00724(new_n3073, new_n3072, new_n3034);
xnor_3 g00725(new_n3074, new_n3073, new_n3033);
xor_3  g00726(new_n3075, n27089, n12657);
not_3  g00727(new_n3076_1, new_n3075);
nor_4  g00728(new_n3077, n17077, n11841);
xor_3  g00729(new_n3078, n17077, n11841);
not_3  g00730(new_n3079, new_n3078);
not_3  g00731(new_n3080, n10710);
not_3  g00732(new_n3081, n26510);
nand_4 g00733(new_n3082, new_n3081, new_n3080);
xor_3  g00734(new_n3083, n26510, n10710);
nor_4  g00735(new_n3084, n23068, n20929);
not_3  g00736(new_n3085, new_n3084);
xor_3  g00737(new_n3086, n23068, n20929);
nor_4  g00738(new_n3087, n19514, n8006);
not_3  g00739(new_n3088, new_n3087);
xor_3  g00740(new_n3089_1, n19514, n8006);
nor_4  g00741(new_n3090, n25074, n10053);
not_3  g00742(new_n3091, new_n3090);
xor_3  g00743(new_n3092, n25074, n10053);
nor_4  g00744(new_n3093, n16396, n8399);
not_3  g00745(new_n3094, new_n3093);
nand_4 g00746(new_n3095, n16396, n8399);
not_3  g00747(new_n3096, new_n3095);
nor_4  g00748(new_n3097, new_n3096, new_n3093);
nor_4  g00749(new_n3098, n9507, n9399);
not_3  g00750(new_n3099, new_n3098);
nand_4 g00751(new_n3100, n26979, n2088);
nand_4 g00752(new_n3101, n9507, n9399);
not_3  g00753(new_n3102, new_n3101);
nor_4  g00754(new_n3103, new_n3102, new_n3098);
nand_4 g00755(new_n3104, new_n3103, new_n3100);
nand_4 g00756(new_n3105, new_n3104, new_n3099);
nand_4 g00757(new_n3106, new_n3105, new_n3097);
nand_4 g00758(new_n3107, new_n3106, new_n3094);
nand_4 g00759(new_n3108, new_n3107, new_n3092);
nand_4 g00760(new_n3109, new_n3108, new_n3091);
nand_4 g00761(new_n3110, new_n3109, new_n3089_1);
nand_4 g00762(new_n3111, new_n3110, new_n3088);
nand_4 g00763(new_n3112, new_n3111, new_n3086);
nand_4 g00764(new_n3113, new_n3112, new_n3085);
nand_4 g00765(new_n3114, new_n3113, new_n3083);
nand_4 g00766(new_n3115, new_n3114, new_n3082);
not_3  g00767(new_n3116, new_n3115);
nor_4  g00768(new_n3117, new_n3116, new_n3079);
nor_4  g00769(new_n3118, new_n3117, new_n3077);
xnor_3 g00770(new_n3119, new_n3118, new_n3076_1);
xnor_3 g00771(new_n3120, new_n3119, new_n3074);
xnor_3 g00772(new_n3121, new_n3070, new_n3035);
not_3  g00773(new_n3122, new_n3121);
xnor_3 g00774(new_n3123, new_n3115, new_n3078);
nor_4  g00775(new_n3124, new_n3123, new_n3122);
xnor_3 g00776(new_n3125_1, new_n3115, new_n3079);
xnor_3 g00777(new_n3126_1, new_n3125_1, new_n3121);
xnor_3 g00778(new_n3127, new_n3068, new_n3040);
not_3  g00779(new_n3128, new_n3127);
xnor_3 g00780(new_n3129, new_n3113, new_n3083);
nand_4 g00781(new_n3130, new_n3129, new_n3128);
xnor_3 g00782(new_n3131, new_n3129, new_n3127);
xnor_3 g00783(new_n3132, new_n3066, new_n3043);
not_3  g00784(new_n3133, new_n3132);
xnor_3 g00785(new_n3134, new_n3111, new_n3086);
nand_4 g00786(new_n3135, new_n3134, new_n3133);
xnor_3 g00787(new_n3136_1, new_n3134, new_n3132);
xnor_3 g00788(new_n3137, new_n3064, new_n3046);
not_3  g00789(new_n3138, new_n3137);
xnor_3 g00790(new_n3139, new_n3109, new_n3089_1);
nand_4 g00791(new_n3140, new_n3139, new_n3138);
xnor_3 g00792(new_n3141, new_n3139, new_n3137);
not_3  g00793(new_n3142, new_n3049);
xnor_3 g00794(new_n3143, new_n3062, new_n3142);
not_3  g00795(new_n3144, new_n3107);
xnor_3 g00796(new_n3145, new_n3144, new_n3092);
not_3  g00797(new_n3146, new_n3145);
nand_4 g00798(new_n3147, new_n3146, new_n3143);
not_3  g00799(new_n3148, new_n3147);
nor_4  g00800(new_n3149, new_n3146, new_n3143);
nor_4  g00801(new_n3150, new_n3149, new_n3148);
not_3  g00802(new_n3151, new_n3060);
xnor_3 g00803(new_n3152, new_n3151, new_n3052);
not_3  g00804(new_n3153, new_n3106);
nor_4  g00805(new_n3154, new_n3105, new_n3097);
nor_4  g00806(new_n3155, new_n3154, new_n3153);
not_3  g00807(new_n3156, new_n3155);
nor_4  g00808(new_n3157, new_n3156, new_n3152);
xnor_3 g00809(new_n3158, new_n3156, new_n3152);
xnor_3 g00810(new_n3159, new_n3058, new_n3055);
not_3  g00811(new_n3160, new_n3104);
nor_4  g00812(new_n3161_1, new_n3103, new_n3100);
nor_4  g00813(new_n3162, new_n3161_1, new_n3160);
nor_4  g00814(new_n3163, new_n3162, new_n3159);
not_3  g00815(new_n3164_1, new_n3163);
xor_3  g00816(new_n3165, n15780, n1451);
xor_3  g00817(new_n3166, n26979, n2088);
not_3  g00818(new_n3167, new_n3166);
nor_4  g00819(new_n3168, new_n3167, new_n3165);
not_3  g00820(new_n3169, new_n3159);
not_3  g00821(new_n3170, new_n3162);
nor_4  g00822(new_n3171, new_n3170, new_n3169);
nor_4  g00823(new_n3172, new_n3171, new_n3163);
nand_4 g00824(new_n3173, new_n3172, new_n3168);
nand_4 g00825(new_n3174, new_n3173, new_n3164_1);
nor_4  g00826(new_n3175, new_n3174, new_n3158);
nor_4  g00827(new_n3176, new_n3175, new_n3157);
nand_4 g00828(new_n3177, new_n3176, new_n3150);
nand_4 g00829(new_n3178, new_n3177, new_n3147);
nand_4 g00830(new_n3179, new_n3178, new_n3141);
nand_4 g00831(new_n3180, new_n3179, new_n3140);
nand_4 g00832(new_n3181, new_n3180, new_n3136_1);
nand_4 g00833(new_n3182, new_n3181, new_n3135);
nand_4 g00834(new_n3183, new_n3182, new_n3131);
nand_4 g00835(new_n3184, new_n3183, new_n3130);
nor_4  g00836(new_n3185, new_n3184, new_n3126_1);
nor_4  g00837(new_n3186, new_n3185, new_n3124);
xnor_3 g00838(new_n3187, new_n3186, new_n3120);
xnor_3 g00839(new_n3188, new_n3187, new_n3032);
xnor_3 g00840(new_n3189, new_n3029, new_n2988);
nand_4 g00841(new_n3190, new_n3184, new_n3126_1);
not_3  g00842(new_n3191, new_n3190);
nor_4  g00843(new_n3192, new_n3191, new_n3185);
not_3  g00844(new_n3193, new_n3192);
nand_4 g00845(new_n3194, new_n3193, new_n3189);
xnor_3 g00846(new_n3195, new_n3192, new_n3189);
not_3  g00847(new_n3196, new_n2992);
xor_3  g00848(new_n3197, new_n3027, new_n3196);
not_3  g00849(new_n3198, new_n3183);
nor_4  g00850(new_n3199, new_n3182, new_n3131);
nor_4  g00851(new_n3200, new_n3199, new_n3198);
nand_4 g00852(new_n3201, new_n3200, new_n3197);
not_3  g00853(new_n3202, new_n3200);
xnor_3 g00854(new_n3203, new_n3202, new_n3197);
not_3  g00855(new_n3204, new_n2996);
xor_3  g00856(new_n3205, new_n3025, new_n3204);
xnor_3 g00857(new_n3206, new_n3180, new_n3136_1);
not_3  g00858(new_n3207, new_n3206);
nand_4 g00859(new_n3208_1, new_n3207, new_n3205);
xnor_3 g00860(new_n3209, new_n3206, new_n3205);
xor_3  g00861(new_n3210, new_n3022, new_n3001);
xnor_3 g00862(new_n3211, new_n3178, new_n3141);
not_3  g00863(new_n3212, new_n3211);
nand_4 g00864(new_n3213, new_n3212, new_n3210);
xnor_3 g00865(new_n3214, new_n3211, new_n3210);
not_3  g00866(new_n3215, new_n3176);
xnor_3 g00867(new_n3216, new_n3215, new_n3150);
xor_3  g00868(new_n3217, new_n3020_1, new_n3004);
not_3  g00869(new_n3218, new_n3217);
nand_4 g00870(new_n3219_1, new_n3218, new_n3216);
not_3  g00871(new_n3220, new_n3219_1);
nor_4  g00872(new_n3221, new_n3218, new_n3216);
nor_4  g00873(new_n3222, new_n3221, new_n3220);
not_3  g00874(new_n3223, new_n3158);
xnor_3 g00875(new_n3224, new_n3174, new_n3223);
not_3  g00876(new_n3225, new_n3017_1);
nor_4  g00877(new_n3226, new_n3008, new_n3006);
xor_3  g00878(new_n3227, new_n3226, new_n3225);
not_3  g00879(new_n3228_1, new_n3227);
nor_4  g00880(new_n3229, new_n3228_1, new_n3224);
not_3  g00881(new_n3230, new_n3229);
not_3  g00882(new_n3231, new_n3224);
nor_4  g00883(new_n3232, new_n3227, new_n3231);
nor_4  g00884(new_n3233, new_n3232, new_n3229);
xor_3  g00885(new_n3234, n5438, new_n3013);
not_3  g00886(new_n3235_1, new_n3165);
nor_4  g00887(new_n3236, new_n3166, new_n3235_1);
nor_4  g00888(new_n3237, new_n3236, new_n3168);
nor_4  g00889(new_n3238, new_n3237, new_n3234);
nor_4  g00890(new_n3239, new_n3012, new_n3010_1);
xor_3  g00891(new_n3240, new_n3239, new_n3014);
not_3  g00892(new_n3241, new_n3240);
nor_4  g00893(new_n3242, new_n3241, new_n3238);
not_3  g00894(new_n3243, new_n3242);
xnor_3 g00895(new_n3244_1, new_n3172, new_n3168);
not_3  g00896(new_n3245, new_n3244_1);
not_3  g00897(new_n3246, new_n3238);
nor_4  g00898(new_n3247, new_n3240, new_n3246);
nor_4  g00899(new_n3248, new_n3247, new_n3242);
nand_4 g00900(new_n3249, new_n3248, new_n3245);
nand_4 g00901(new_n3250, new_n3249, new_n3243);
nand_4 g00902(new_n3251, new_n3250, new_n3233);
nand_4 g00903(new_n3252, new_n3251, new_n3230);
nand_4 g00904(new_n3253_1, new_n3252, new_n3222);
nand_4 g00905(new_n3254, new_n3253_1, new_n3219_1);
nand_4 g00906(new_n3255, new_n3254, new_n3214);
nand_4 g00907(new_n3256, new_n3255, new_n3213);
nand_4 g00908(new_n3257, new_n3256, new_n3209);
nand_4 g00909(new_n3258, new_n3257, new_n3208_1);
nand_4 g00910(new_n3259, new_n3258, new_n3203);
nand_4 g00911(new_n3260_1, new_n3259, new_n3201);
nand_4 g00912(new_n3261, new_n3260_1, new_n3195);
nand_4 g00913(new_n3262, new_n3261, new_n3194);
not_3  g00914(new_n3263_1, new_n3262);
xor_3  g00915(n142, new_n3263_1, new_n3188);
nor_4  g00916(new_n3265, n7593, n5101);
xor_3  g00917(new_n3266, n7593, n5101);
not_3  g00918(new_n3267, new_n3266);
nor_4  g00919(new_n3268, n16507, n337);
xor_3  g00920(new_n3269, n16507, n337);
not_3  g00921(new_n3270, new_n3269);
nor_4  g00922(new_n3271, n22470, n3228);
xor_3  g00923(new_n3272, n22470, n3228);
not_3  g00924(new_n3273, new_n3272);
not_3  g00925(new_n3274, n5302);
not_3  g00926(new_n3275, n19116);
nand_4 g00927(new_n3276, new_n3275, new_n3274);
xor_3  g00928(new_n3277, n19116, n5302);
nor_4  g00929(new_n3278, n25738, n6861);
not_3  g00930(new_n3279_1, new_n3278);
xor_3  g00931(new_n3280, n25738, n6861);
nor_4  g00932(new_n3281, n21471, n19357);
not_3  g00933(new_n3282, new_n3281);
xor_3  g00934(new_n3283, n21471, n19357);
nor_4  g00935(new_n3284, n18737, n2328);
not_3  g00936(new_n3285, new_n3284);
xor_3  g00937(new_n3286, n18737, n2328);
nor_4  g00938(new_n3287, n15053, n14603);
not_3  g00939(new_n3288, new_n3287);
xor_3  g00940(new_n3289_1, n15053, n14603);
not_3  g00941(new_n3290, n20794);
not_3  g00942(new_n3291, n25471);
nand_4 g00943(new_n3292, new_n3291, new_n3290);
nand_4 g00944(new_n3293, n23333, n16502);
xor_3  g00945(new_n3294, n25471, n20794);
nand_4 g00946(new_n3295, new_n3294, new_n3293);
nand_4 g00947(new_n3296, new_n3295, new_n3292);
nand_4 g00948(new_n3297, new_n3296, new_n3289_1);
nand_4 g00949(new_n3298, new_n3297, new_n3288);
nand_4 g00950(new_n3299, new_n3298, new_n3286);
nand_4 g00951(new_n3300, new_n3299, new_n3285);
nand_4 g00952(new_n3301_1, new_n3300, new_n3283);
nand_4 g00953(new_n3302, new_n3301_1, new_n3282);
nand_4 g00954(new_n3303, new_n3302, new_n3280);
nand_4 g00955(new_n3304, new_n3303, new_n3279_1);
nand_4 g00956(new_n3305, new_n3304, new_n3277);
nand_4 g00957(new_n3306_1, new_n3305, new_n3276);
not_3  g00958(new_n3307, new_n3306_1);
nor_4  g00959(new_n3308, new_n3307, new_n3273);
nor_4  g00960(new_n3309, new_n3308, new_n3271);
nor_4  g00961(new_n3310, new_n3309, new_n3270);
nor_4  g00962(new_n3311, new_n3310, new_n3268);
nor_4  g00963(new_n3312, new_n3311, new_n3267);
nor_4  g00964(new_n3313, new_n3312, new_n3265);
not_3  g00965(new_n3314, n24618);
nor_4  g00966(new_n3315, n12315, n3952);
nand_4 g00967(new_n3316_1, new_n3315, new_n3314);
nor_4  g00968(new_n3317, new_n3316_1, n24278);
not_3  g00969(new_n3318, new_n3317);
nor_4  g00970(new_n3319, new_n3318, n4812);
not_3  g00971(new_n3320_1, new_n3319);
nor_4  g00972(new_n3321, new_n3320_1, n26823);
not_3  g00973(new_n3322, new_n3321);
nor_4  g00974(new_n3323, new_n3322, n7751);
not_3  g00975(new_n3324_1, new_n3323);
nor_4  g00976(new_n3325, new_n3324_1, n20946);
not_3  g00977(new_n3326, new_n3325);
nor_4  g00978(new_n3327, new_n3326, n9967);
not_3  g00979(new_n3328, new_n3327);
nor_4  g00980(new_n3329, new_n3328, n3425);
not_3  g00981(new_n3330, n3425);
xor_3  g00982(new_n3331, new_n3327, new_n3330);
xor_3  g00983(new_n3332_1, n7335, n4319);
nor_4  g00984(new_n3333, n23463, n5696);
xor_3  g00985(new_n3334, n23463, n5696);
not_3  g00986(new_n3335, n13074);
not_3  g00987(new_n3336, n13367);
nand_4 g00988(new_n3337, new_n3336, new_n3335);
xor_3  g00989(new_n3338, n13367, n13074);
nor_4  g00990(new_n3339, n10739, n932);
not_3  g00991(new_n3340_1, new_n3339);
xor_3  g00992(new_n3341, n10739, n932);
nor_4  g00993(new_n3342, n21753, n6691);
not_3  g00994(new_n3343_1, new_n3342);
xor_3  g00995(new_n3344, n21753, n6691);
nor_4  g00996(new_n3345, n21832, n3260);
not_3  g00997(new_n3346, new_n3345);
nand_4 g00998(new_n3347, n21832, n3260);
not_3  g00999(new_n3348, new_n3347);
nor_4  g01000(new_n3349_1, new_n3348, new_n3345);
nor_4  g01001(new_n3350, n26913, n20489);
not_3  g01002(new_n3351, new_n3350);
nand_4 g01003(new_n3352, n26913, n20489);
not_3  g01004(new_n3353, new_n3352);
nor_4  g01005(new_n3354, new_n3353, new_n3350);
nor_4  g01006(new_n3355, n16223, n2355);
not_3  g01007(new_n3356, new_n3355);
nand_4 g01008(new_n3357, n16223, n2355);
not_3  g01009(new_n3358, new_n3357);
nor_4  g01010(new_n3359, new_n3358, new_n3355);
nand_4 g01011(new_n3360, n19494, n11121);
not_3  g01012(new_n3361, new_n3360);
nor_4  g01013(new_n3362, n19494, n11121);
nand_4 g01014(new_n3363, n16217, n2387);
nor_4  g01015(new_n3364, new_n3363, new_n3362);
nor_4  g01016(new_n3365, new_n3364, new_n3361);
nand_4 g01017(new_n3366_1, new_n3365, new_n3359);
nand_4 g01018(new_n3367, new_n3366_1, new_n3356);
nand_4 g01019(new_n3368, new_n3367, new_n3354);
nand_4 g01020(new_n3369, new_n3368, new_n3351);
nand_4 g01021(new_n3370, new_n3369, new_n3349_1);
nand_4 g01022(new_n3371, new_n3370, new_n3346);
nand_4 g01023(new_n3372, new_n3371, new_n3344);
nand_4 g01024(new_n3373, new_n3372, new_n3343_1);
nand_4 g01025(new_n3374, new_n3373, new_n3341);
nand_4 g01026(new_n3375, new_n3374, new_n3340_1);
nand_4 g01027(new_n3376, new_n3375, new_n3338);
nand_4 g01028(new_n3377, new_n3376, new_n3337);
nand_4 g01029(new_n3378, new_n3377, new_n3334);
not_3  g01030(new_n3379, new_n3378);
nor_4  g01031(new_n3380, new_n3379, new_n3333);
xnor_3 g01032(new_n3381, new_n3380, new_n3332_1);
xnor_3 g01033(new_n3382, new_n3381, n5025);
xnor_3 g01034(new_n3383, new_n3377, new_n3334);
not_3  g01035(new_n3384, new_n3383);
nor_4  g01036(new_n3385, new_n3384, n6485);
not_3  g01037(new_n3386, new_n3385);
not_3  g01038(new_n3387, n6485);
nor_4  g01039(new_n3388, new_n3383, new_n3387);
nor_4  g01040(new_n3389, new_n3388, new_n3385);
xnor_3 g01041(new_n3390_1, new_n3375, new_n3338);
not_3  g01042(new_n3391, new_n3390_1);
nor_4  g01043(new_n3392, new_n3391, n26036);
not_3  g01044(new_n3393, new_n3392);
not_3  g01045(new_n3394, n26036);
nor_4  g01046(new_n3395, new_n3390_1, new_n3394);
nor_4  g01047(new_n3396, new_n3395, new_n3392);
xnor_3 g01048(new_n3397, new_n3373, new_n3341);
not_3  g01049(new_n3398, new_n3397);
nor_4  g01050(new_n3399, new_n3398, n19770);
not_3  g01051(new_n3400, new_n3399);
not_3  g01052(new_n3401, n19770);
nor_4  g01053(new_n3402, new_n3397, new_n3401);
nor_4  g01054(new_n3403, new_n3402, new_n3399);
not_3  g01055(new_n3404, new_n3372);
nor_4  g01056(new_n3405, new_n3371, new_n3344);
nor_4  g01057(new_n3406, new_n3405, new_n3404);
nor_4  g01058(new_n3407, new_n3406, n8782);
not_3  g01059(new_n3408, new_n3407);
not_3  g01060(new_n3409, n8782);
xnor_3 g01061(new_n3410, new_n3371, new_n3344);
nor_4  g01062(new_n3411, new_n3410, new_n3409);
nor_4  g01063(new_n3412, new_n3411, new_n3407);
xnor_3 g01064(new_n3413, new_n3369, new_n3349_1);
not_3  g01065(new_n3414, new_n3413);
nor_4  g01066(new_n3415, new_n3414, n8678);
not_3  g01067(new_n3416, new_n3415);
not_3  g01068(new_n3417, n8678);
nor_4  g01069(new_n3418, new_n3413, new_n3417);
nor_4  g01070(new_n3419, new_n3418, new_n3415);
xnor_3 g01071(new_n3420, new_n3367, new_n3354);
not_3  g01072(new_n3421, new_n3420);
nor_4  g01073(new_n3422, new_n3421, n1432);
not_3  g01074(new_n3423, new_n3422);
not_3  g01075(new_n3424, n1432);
nor_4  g01076(new_n3425_1, new_n3420, new_n3424);
nor_4  g01077(new_n3426_1, new_n3425_1, new_n3422);
xnor_3 g01078(new_n3427, new_n3365, new_n3359);
not_3  g01079(new_n3428, new_n3427);
nor_4  g01080(new_n3429, new_n3428, n21599);
not_3  g01081(new_n3430, new_n3429);
not_3  g01082(new_n3431, n21599);
nor_4  g01083(new_n3432, new_n3427, new_n3431);
nor_4  g01084(new_n3433, new_n3432, new_n3429);
not_3  g01085(new_n3434, n25336);
xnor_3 g01086(new_n3435, n16217, n2387);
nor_4  g01087(new_n3436, new_n3435, n11424);
nand_4 g01088(new_n3437, new_n3436, new_n3434);
not_3  g01089(new_n3438, new_n3437);
nor_4  g01090(new_n3439, new_n3436, new_n3434);
nor_4  g01091(new_n3440, new_n3439, new_n3438);
xnor_3 g01092(new_n3441, n19494, n11121);
xnor_3 g01093(new_n3442, new_n3441, new_n3363);
not_3  g01094(new_n3443, new_n3442);
nand_4 g01095(new_n3444, new_n3443, new_n3440);
nand_4 g01096(new_n3445, new_n3444, new_n3437);
nand_4 g01097(new_n3446, new_n3445, new_n3433);
nand_4 g01098(new_n3447, new_n3446, new_n3430);
nand_4 g01099(new_n3448, new_n3447, new_n3426_1);
nand_4 g01100(new_n3449, new_n3448, new_n3423);
nand_4 g01101(new_n3450, new_n3449, new_n3419);
nand_4 g01102(new_n3451_1, new_n3450, new_n3416);
nand_4 g01103(new_n3452, new_n3451_1, new_n3412);
nand_4 g01104(new_n3453, new_n3452, new_n3408);
nand_4 g01105(new_n3454, new_n3453, new_n3403);
nand_4 g01106(new_n3455, new_n3454, new_n3400);
nand_4 g01107(new_n3456, new_n3455, new_n3396);
nand_4 g01108(new_n3457, new_n3456, new_n3393);
nand_4 g01109(new_n3458, new_n3457, new_n3389);
nand_4 g01110(new_n3459_1, new_n3458, new_n3386);
xnor_3 g01111(new_n3460_1, new_n3459_1, new_n3382);
not_3  g01112(new_n3461, new_n3460_1);
nand_4 g01113(new_n3462, new_n3461, new_n3331);
xnor_3 g01114(new_n3463, new_n3460_1, new_n3331);
not_3  g01115(new_n3464, n9967);
xor_3  g01116(new_n3465, new_n3325, new_n3464);
xnor_3 g01117(new_n3466, new_n3457, new_n3389);
nand_4 g01118(new_n3467, new_n3466, new_n3465);
not_3  g01119(new_n3468_1, new_n3465);
xnor_3 g01120(new_n3469, new_n3466, new_n3468_1);
xor_3  g01121(new_n3470, new_n3324_1, n20946);
xnor_3 g01122(new_n3471, new_n3455, new_n3396);
nand_4 g01123(new_n3472, new_n3471, new_n3470);
not_3  g01124(new_n3473, new_n3470);
xnor_3 g01125(new_n3474, new_n3471, new_n3473);
not_3  g01126(new_n3475, n7751);
xor_3  g01127(new_n3476, new_n3321, new_n3475);
xnor_3 g01128(new_n3477, new_n3397, new_n3401);
xnor_3 g01129(new_n3478, new_n3453, new_n3477);
not_3  g01130(new_n3479, new_n3478);
nand_4 g01131(new_n3480_1, new_n3479, new_n3476);
xnor_3 g01132(new_n3481, new_n3478, new_n3476);
not_3  g01133(new_n3482, n26823);
xor_3  g01134(new_n3483, new_n3320_1, new_n3482);
not_3  g01135(new_n3484, new_n3483);
xnor_3 g01136(new_n3485, new_n3451_1, new_n3412);
nand_4 g01137(new_n3486, new_n3485, new_n3484);
xnor_3 g01138(new_n3487, new_n3485, new_n3483);
xor_3  g01139(new_n3488, new_n3317, n4812);
not_3  g01140(new_n3489, new_n3488);
xnor_3 g01141(new_n3490, new_n3449, new_n3419);
nand_4 g01142(new_n3491, new_n3490, new_n3489);
xnor_3 g01143(new_n3492, new_n3490, new_n3488);
xor_3  g01144(new_n3493, new_n3316_1, n24278);
xnor_3 g01145(new_n3494, new_n3447, new_n3426_1);
nand_4 g01146(new_n3495, new_n3494, new_n3493);
not_3  g01147(new_n3496, new_n3493);
xnor_3 g01148(new_n3497, new_n3494, new_n3496);
xor_3  g01149(new_n3498, new_n3315, new_n3314);
xnor_3 g01150(new_n3499, new_n3436, new_n3434);
nor_4  g01151(new_n3500, new_n3442, new_n3499);
nor_4  g01152(new_n3501, new_n3500, new_n3438);
xnor_3 g01153(new_n3502_1, new_n3501, new_n3433);
not_3  g01154(new_n3503, new_n3502_1);
nand_4 g01155(new_n3504, new_n3503, new_n3498);
xnor_3 g01156(new_n3505, new_n3502_1, new_n3498);
not_3  g01157(new_n3506_1, n12315);
not_3  g01158(new_n3507, n11424);
not_3  g01159(new_n3508, new_n3435);
nor_4  g01160(new_n3509, new_n3508, new_n3507);
nor_4  g01161(new_n3510, new_n3509, new_n3436);
nor_4  g01162(new_n3511, new_n3510, new_n3506_1);
not_3  g01163(new_n3512, new_n3511);
nor_4  g01164(new_n3513, new_n3512, n3952);
not_3  g01165(new_n3514, new_n3513);
xnor_3 g01166(new_n3515, new_n3442, new_n3499);
nand_4 g01167(new_n3516_1, n12315, n3952);
not_3  g01168(new_n3517, new_n3516_1);
nor_4  g01169(new_n3518, new_n3517, new_n3315);
nor_4  g01170(new_n3519, new_n3518, new_n3511);
nor_4  g01171(new_n3520, new_n3519, new_n3513);
nand_4 g01172(new_n3521, new_n3520, new_n3515);
nand_4 g01173(new_n3522, new_n3521, new_n3514);
nand_4 g01174(new_n3523, new_n3522, new_n3505);
nand_4 g01175(new_n3524, new_n3523, new_n3504);
nand_4 g01176(new_n3525, new_n3524, new_n3497);
nand_4 g01177(new_n3526, new_n3525, new_n3495);
nand_4 g01178(new_n3527, new_n3526, new_n3492);
nand_4 g01179(new_n3528_1, new_n3527, new_n3491);
nand_4 g01180(new_n3529, new_n3528_1, new_n3487);
nand_4 g01181(new_n3530, new_n3529, new_n3486);
nand_4 g01182(new_n3531, new_n3530, new_n3481);
nand_4 g01183(new_n3532, new_n3531, new_n3480_1);
nand_4 g01184(new_n3533, new_n3532, new_n3474);
nand_4 g01185(new_n3534, new_n3533, new_n3472);
nand_4 g01186(new_n3535, new_n3534, new_n3469);
nand_4 g01187(new_n3536, new_n3535, new_n3467);
nand_4 g01188(new_n3537, new_n3536, new_n3463);
nand_4 g01189(new_n3538, new_n3537, new_n3462);
nor_4  g01190(new_n3539, new_n3381, n5025);
not_3  g01191(new_n3540, new_n3459_1);
nor_4  g01192(new_n3541_1, new_n3540, new_n3382);
nor_4  g01193(new_n3542, new_n3541_1, new_n3539);
nor_4  g01194(new_n3543, n7335, n4319);
not_3  g01195(new_n3544, new_n3332_1);
nor_4  g01196(new_n3545, new_n3380, new_n3544);
nor_4  g01197(new_n3546, new_n3545, new_n3543);
not_3  g01198(new_n3547, new_n3546);
xnor_3 g01199(new_n3548, new_n3547, new_n3542);
not_3  g01200(new_n3549, new_n3548);
nor_4  g01201(new_n3550, new_n3549, new_n3538);
not_3  g01202(new_n3551, new_n3538);
nor_4  g01203(new_n3552, new_n3548, new_n3551);
nor_4  g01204(new_n3553, new_n3552, new_n3550);
xnor_3 g01205(new_n3554, new_n3553, new_n3329);
nand_4 g01206(new_n3555_1, new_n3554, new_n3313);
not_3  g01207(new_n3556, new_n3537);
nor_4  g01208(new_n3557, new_n3536, new_n3463);
nor_4  g01209(new_n3558, new_n3557, new_n3556);
xor_3  g01210(new_n3559, new_n3311, new_n3266);
nor_4  g01211(new_n3560, new_n3559, new_n3558);
xnor_3 g01212(new_n3561_1, new_n3559, new_n3558);
not_3  g01213(new_n3562, new_n3535);
nor_4  g01214(new_n3563_1, new_n3534, new_n3469);
nor_4  g01215(new_n3564, new_n3563_1, new_n3562);
xor_3  g01216(new_n3565, new_n3309, new_n3269);
nor_4  g01217(new_n3566, new_n3565, new_n3564);
xnor_3 g01218(new_n3567, new_n3565, new_n3564);
not_3  g01219(new_n3568, new_n3533);
nor_4  g01220(new_n3569, new_n3532, new_n3474);
nor_4  g01221(new_n3570_1, new_n3569, new_n3568);
xor_3  g01222(new_n3571, new_n3307, new_n3272);
nor_4  g01223(new_n3572, new_n3571, new_n3570_1);
xnor_3 g01224(new_n3573, new_n3571, new_n3570_1);
xnor_3 g01225(new_n3574, new_n3530, new_n3481);
not_3  g01226(new_n3575, new_n3304);
xor_3  g01227(new_n3576, new_n3575, new_n3277);
not_3  g01228(new_n3577, new_n3576);
nand_4 g01229(new_n3578, new_n3577, new_n3574);
not_3  g01230(new_n3579, new_n3578);
nor_4  g01231(new_n3580, new_n3577, new_n3574);
nor_4  g01232(new_n3581, new_n3580, new_n3579);
xnor_3 g01233(new_n3582_1, new_n3528_1, new_n3487);
not_3  g01234(new_n3583, new_n3302);
xor_3  g01235(new_n3584, new_n3583, new_n3280);
not_3  g01236(new_n3585, new_n3584);
nand_4 g01237(new_n3586, new_n3585, new_n3582_1);
xnor_3 g01238(new_n3587, new_n3584, new_n3582_1);
xnor_3 g01239(new_n3588, new_n3526, new_n3492);
not_3  g01240(new_n3589, new_n3300);
xor_3  g01241(new_n3590, new_n3589, new_n3283);
not_3  g01242(new_n3591, new_n3590);
nand_4 g01243(new_n3592, new_n3591, new_n3588);
xnor_3 g01244(new_n3593, new_n3590, new_n3588);
not_3  g01245(new_n3594, new_n3524);
xnor_3 g01246(new_n3595, new_n3594, new_n3497);
not_3  g01247(new_n3596, new_n3286);
not_3  g01248(new_n3597, new_n3298);
xor_3  g01249(new_n3598, new_n3597, new_n3596);
not_3  g01250(new_n3599, new_n3598);
nor_4  g01251(new_n3600, new_n3599, new_n3595);
not_3  g01252(new_n3601, new_n3600);
not_3  g01253(new_n3602, new_n3595);
nor_4  g01254(new_n3603, new_n3598, new_n3602);
nor_4  g01255(new_n3604, new_n3603, new_n3600);
xnor_3 g01256(new_n3605, new_n3522, new_n3505);
xnor_3 g01257(new_n3606, new_n3296, new_n3289_1);
not_3  g01258(new_n3607, new_n3606);
nand_4 g01259(new_n3608, new_n3607, new_n3605);
not_3  g01260(new_n3609, new_n3608);
nor_4  g01261(new_n3610, new_n3607, new_n3605);
nor_4  g01262(new_n3611, new_n3610, new_n3609);
xor_3  g01263(new_n3612, n23333, n16502);
not_3  g01264(new_n3613, new_n3612);
xor_3  g01265(new_n3614, new_n3510, n12315);
nor_4  g01266(new_n3615, new_n3614, new_n3613);
not_3  g01267(new_n3616, new_n3294);
xor_3  g01268(new_n3617_1, new_n3616, new_n3293);
nor_4  g01269(new_n3618_1, new_n3617_1, new_n3615);
not_3  g01270(new_n3619, new_n3618_1);
xnor_3 g01271(new_n3620, new_n3520, new_n3515);
xor_3  g01272(new_n3621, new_n3510, new_n3506_1);
nand_4 g01273(new_n3622, new_n3621, new_n3612);
nor_4  g01274(new_n3623, new_n3622, new_n3616);
nor_4  g01275(new_n3624, new_n3623, new_n3618_1);
nand_4 g01276(new_n3625, new_n3624, new_n3620);
nand_4 g01277(new_n3626, new_n3625, new_n3619);
nand_4 g01278(new_n3627, new_n3626, new_n3611);
nand_4 g01279(new_n3628, new_n3627, new_n3608);
nand_4 g01280(new_n3629, new_n3628, new_n3604);
nand_4 g01281(new_n3630, new_n3629, new_n3601);
nand_4 g01282(new_n3631, new_n3630, new_n3593);
nand_4 g01283(new_n3632, new_n3631, new_n3592);
nand_4 g01284(new_n3633, new_n3632, new_n3587);
nand_4 g01285(new_n3634, new_n3633, new_n3586);
nand_4 g01286(new_n3635, new_n3634, new_n3581);
not_3  g01287(new_n3636, new_n3635);
nor_4  g01288(new_n3637, new_n3636, new_n3579);
nor_4  g01289(new_n3638, new_n3637, new_n3573);
nor_4  g01290(new_n3639, new_n3638, new_n3572);
nor_4  g01291(new_n3640, new_n3639, new_n3567);
nor_4  g01292(new_n3641, new_n3640, new_n3566);
nor_4  g01293(new_n3642_1, new_n3641, new_n3561_1);
nor_4  g01294(new_n3643, new_n3642_1, new_n3560);
not_3  g01295(new_n3644, new_n3313);
xnor_3 g01296(new_n3645, new_n3554, new_n3644);
nand_4 g01297(new_n3646, new_n3645, new_n3643);
nand_4 g01298(new_n3647, new_n3646, new_n3555_1);
not_3  g01299(new_n3648, new_n3550);
not_3  g01300(new_n3649_1, new_n3329);
nand_4 g01301(new_n3650, new_n3547, new_n3542);
xor_3  g01302(new_n3651, new_n3650, new_n3649_1);
nor_4  g01303(new_n3652, new_n3651, new_n3648);
xor_3  g01304(new_n3653, new_n3650, new_n3329);
nor_4  g01305(new_n3654, new_n3653, new_n3551);
nor_4  g01306(new_n3655, new_n3654, new_n3652);
nand_4 g01307(new_n3656, new_n3655, new_n3647);
nor_4  g01308(new_n3657, new_n3650, new_n3329);
and_4  g01309(new_n3658, new_n3657, new_n3551);
xnor_3 g01310(n175, new_n3658, new_n3656);
not_3  g01311(new_n3660, n26180);
not_3  g01312(new_n3661, n25494);
not_3  g01313(new_n3662, n8856);
nor_4  g01314(new_n3663, n20138, n9251);
nand_4 g01315(new_n3664, new_n3663, new_n2366);
nor_4  g01316(new_n3665_1, new_n3664, n3136);
nand_4 g01317(new_n3666, new_n3665_1, new_n2359);
nor_4  g01318(new_n3667, new_n3666, n25643);
nand_4 g01319(new_n3668, new_n3667, new_n2349);
nor_4  g01320(new_n3669, new_n3668, n16482);
not_3  g01321(new_n3670, new_n3669);
nor_4  g01322(new_n3671, new_n3670, n14130);
xor_3  g01323(new_n3672, new_n3671, new_n3662);
not_3  g01324(new_n3673, new_n3672);
nor_4  g01325(new_n3674, new_n3673, new_n3661);
nor_4  g01326(new_n3675, new_n3672, n25494);
nor_4  g01327(new_n3676, new_n3675, new_n3674);
xor_3  g01328(new_n3677, new_n3670, n14130);
nor_4  g01329(new_n3678, new_n3677, n10117);
not_3  g01330(new_n3679_1, new_n3677);
xor_3  g01331(new_n3680, new_n3679_1, n10117);
xor_3  g01332(new_n3681, new_n3668, n16482);
nor_4  g01333(new_n3682, new_n3681, n13460);
not_3  g01334(new_n3683, new_n3681);
xor_3  g01335(new_n3684, new_n3683, n13460);
xor_3  g01336(new_n3685, new_n3667, new_n2349);
nor_4  g01337(new_n3686, new_n3685, n6104);
not_3  g01338(new_n3687, new_n3685);
xor_3  g01339(new_n3688, new_n3687, n6104);
nand_4 g01340(new_n3689, new_n3666, n25643);
not_3  g01341(new_n3690, new_n3689);
nor_4  g01342(new_n3691, new_n3690, new_n3667);
nor_4  g01343(new_n3692, new_n3691, n4119);
not_3  g01344(new_n3693, n4119);
not_3  g01345(new_n3694, new_n3691);
nor_4  g01346(new_n3695, new_n3694, new_n3693);
nor_4  g01347(new_n3696, new_n3695, new_n3692);
not_3  g01348(new_n3697, new_n3696);
xnor_3 g01349(new_n3698, new_n3665_1, n9557);
nor_4  g01350(new_n3699, new_n3698, n14510);
not_3  g01351(new_n3700, n14510);
not_3  g01352(new_n3701, new_n3698);
nor_4  g01353(new_n3702, new_n3701, new_n3700);
nor_4  g01354(new_n3703, new_n3702, new_n3699);
nand_4 g01355(new_n3704, new_n3664, n3136);
not_3  g01356(new_n3705, new_n3704);
nor_4  g01357(new_n3706, new_n3705, new_n3665_1);
nor_4  g01358(new_n3707, new_n3706, n13263);
not_3  g01359(new_n3708, new_n3707);
xnor_3 g01360(new_n3709, new_n3663, n6385);
nor_4  g01361(new_n3710_1, new_n3709, n20455);
not_3  g01362(new_n3711, new_n3710_1);
not_3  g01363(new_n3712, n20455);
not_3  g01364(new_n3713, new_n3709);
nor_4  g01365(new_n3714, new_n3713, new_n3712);
nor_4  g01366(new_n3715, new_n3714, new_n3710_1);
not_3  g01367(new_n3716, n1639);
xnor_3 g01368(new_n3717, n20138, n9251);
nand_4 g01369(new_n3718, new_n3717, new_n3716);
nand_4 g01370(new_n3719, n16968, n9251);
xnor_3 g01371(new_n3720, new_n3717, n1639);
nand_4 g01372(new_n3721, new_n3720, new_n3719);
nand_4 g01373(new_n3722, new_n3721, new_n3718);
nand_4 g01374(new_n3723, new_n3722, new_n3715);
nand_4 g01375(new_n3724, new_n3723, new_n3711);
not_3  g01376(new_n3725_1, n13263);
not_3  g01377(new_n3726, new_n3706);
nor_4  g01378(new_n3727, new_n3726, new_n3725_1);
nor_4  g01379(new_n3728, new_n3727, new_n3707);
nand_4 g01380(new_n3729, new_n3728, new_n3724);
nand_4 g01381(new_n3730, new_n3729, new_n3708);
nand_4 g01382(new_n3731, new_n3730, new_n3703);
not_3  g01383(new_n3732, new_n3731);
nor_4  g01384(new_n3733_1, new_n3732, new_n3699);
nor_4  g01385(new_n3734, new_n3733_1, new_n3697);
nor_4  g01386(new_n3735, new_n3734, new_n3692);
nor_4  g01387(new_n3736, new_n3735, new_n3688);
nor_4  g01388(new_n3737, new_n3736, new_n3686);
nor_4  g01389(new_n3738, new_n3737, new_n3684);
nor_4  g01390(new_n3739, new_n3738, new_n3682);
nor_4  g01391(new_n3740_1, new_n3739, new_n3680);
nor_4  g01392(new_n3741, new_n3740_1, new_n3678);
xnor_3 g01393(new_n3742, new_n3741, new_n3676);
nor_4  g01394(new_n3743, new_n3742, new_n3660);
not_3  g01395(new_n3744, new_n3742);
nor_4  g01396(new_n3745, new_n3744, n26180);
nor_4  g01397(new_n3746, new_n3745, new_n3743);
xnor_3 g01398(new_n3747, new_n3739, new_n3680);
nor_4  g01399(new_n3748, new_n3747, n24004);
not_3  g01400(new_n3749, n24004);
not_3  g01401(new_n3750, new_n3747);
nor_4  g01402(new_n3751, new_n3750, new_n3749);
nor_4  g01403(new_n3752, new_n3751, new_n3748);
not_3  g01404(new_n3753, new_n3752);
not_3  g01405(new_n3754, n12871);
not_3  g01406(new_n3755_1, new_n3737);
xnor_3 g01407(new_n3756, new_n3755_1, new_n3684);
nand_4 g01408(new_n3757, new_n3756, new_n3754);
xnor_3 g01409(new_n3758_1, new_n3756, n12871);
not_3  g01410(new_n3759, new_n3735);
xnor_3 g01411(new_n3760_1, new_n3759, new_n3688);
not_3  g01412(new_n3761, new_n3760_1);
nor_4  g01413(new_n3762, new_n3761, n23304);
not_3  g01414(new_n3763, new_n3762);
not_3  g01415(new_n3764, n23304);
nor_4  g01416(new_n3765, new_n3760_1, new_n3764);
nor_4  g01417(new_n3766, new_n3765, new_n3762);
not_3  g01418(new_n3767, n19361);
not_3  g01419(new_n3768, new_n3733_1);
nor_4  g01420(new_n3769, new_n3768, new_n3696);
nor_4  g01421(new_n3770, new_n3769, new_n3734);
nand_4 g01422(new_n3771, new_n3770, new_n3767);
not_3  g01423(new_n3772, new_n3770);
nor_4  g01424(new_n3773, new_n3772, n19361);
nor_4  g01425(new_n3774, new_n3770, new_n3767);
nor_4  g01426(new_n3775, new_n3774, new_n3773);
xnor_3 g01427(new_n3776, new_n3730, new_n3703);
nor_4  g01428(new_n3777, new_n3776, n1437);
not_3  g01429(new_n3778, new_n3777);
not_3  g01430(new_n3779, n1437);
not_3  g01431(new_n3780, new_n3776);
nor_4  g01432(new_n3781_1, new_n3780, new_n3779);
nor_4  g01433(new_n3782, new_n3781_1, new_n3777);
xnor_3 g01434(new_n3783, new_n3728, new_n3724);
nor_4  g01435(new_n3784, new_n3783, n4722);
not_3  g01436(new_n3785_1, new_n3784);
not_3  g01437(new_n3786, n4722);
not_3  g01438(new_n3787, new_n3783);
nor_4  g01439(new_n3788, new_n3787, new_n3786);
nor_4  g01440(new_n3789, new_n3788, new_n3784);
not_3  g01441(new_n3790, n14633);
xnor_3 g01442(new_n3791, new_n3722, new_n3715);
not_3  g01443(new_n3792, new_n3791);
nor_4  g01444(new_n3793, new_n3792, new_n3790);
nor_4  g01445(new_n3794_1, new_n3791, n14633);
nor_4  g01446(new_n3795_1, new_n3794_1, new_n3793);
not_3  g01447(new_n3796, new_n3795_1);
not_3  g01448(new_n3797, n8721);
xnor_3 g01449(new_n3798, new_n3720, new_n3719);
not_3  g01450(new_n3799, new_n3798);
nor_4  g01451(new_n3800, new_n3799, new_n3797);
xor_3  g01452(new_n3801, n16968, n9251);
nand_4 g01453(new_n3802, new_n3801, n18578);
nor_4  g01454(new_n3803, new_n3798, n8721);
nor_4  g01455(new_n3804, new_n3803, new_n3800);
not_3  g01456(new_n3805, new_n3804);
nor_4  g01457(new_n3806, new_n3805, new_n3802);
nor_4  g01458(new_n3807, new_n3806, new_n3800);
nor_4  g01459(new_n3808, new_n3807, new_n3796);
nor_4  g01460(new_n3809, new_n3808, new_n3793);
nand_4 g01461(new_n3810, new_n3809, new_n3789);
nand_4 g01462(new_n3811, new_n3810, new_n3785_1);
nand_4 g01463(new_n3812, new_n3811, new_n3782);
nand_4 g01464(new_n3813, new_n3812, new_n3778);
nand_4 g01465(new_n3814, new_n3813, new_n3775);
nand_4 g01466(new_n3815, new_n3814, new_n3771);
nand_4 g01467(new_n3816, new_n3815, new_n3766);
nand_4 g01468(new_n3817, new_n3816, new_n3763);
nand_4 g01469(new_n3818, new_n3817, new_n3758_1);
nand_4 g01470(new_n3819, new_n3818, new_n3757);
not_3  g01471(new_n3820, new_n3819);
nor_4  g01472(new_n3821, new_n3820, new_n3753);
nor_4  g01473(new_n3822, new_n3821, new_n3748);
xnor_3 g01474(new_n3823, new_n3822, new_n3746);
not_3  g01475(new_n3824, new_n3823);
not_3  g01476(new_n3825, n2743);
xor_3  g01477(new_n3826, n3506, new_n3825);
not_3  g01478(new_n3827, new_n3826);
not_3  g01479(new_n3828_1, n7026);
nor_4  g01480(new_n3829, n14899, new_n3828_1);
xor_3  g01481(new_n3830, n14899, new_n3828_1);
not_3  g01482(new_n3831, n13719);
or_4   g01483(new_n3832, n18444, new_n3831);
xor_3  g01484(new_n3833, n18444, new_n3831);
not_3  g01485(new_n3834, n24638);
nand_4 g01486(new_n3835, new_n3834, n442);
not_3  g01487(new_n3836, n442);
xor_3  g01488(new_n3837, n24638, new_n3836);
not_3  g01489(new_n3838, n21674);
nand_4 g01490(new_n3839, new_n3838, n9172);
not_3  g01491(new_n3840, n9172);
xor_3  g01492(new_n3841, n21674, new_n3840);
not_3  g01493(new_n3842_1, n4913);
nor_4  g01494(new_n3843, n17251, new_n3842_1);
not_3  g01495(new_n3844, new_n3843);
xor_3  g01496(new_n3845, n17251, new_n3842_1);
not_3  g01497(new_n3846, n604);
nor_4  g01498(new_n3847, n14790, new_n3846);
not_3  g01499(new_n3848, new_n3847);
xor_3  g01500(new_n3849, n14790, new_n3846);
not_3  g01501(new_n3850_1, n10096);
nor_4  g01502(new_n3851, n16824, new_n3850_1);
not_3  g01503(new_n3852, n16824);
nor_4  g01504(new_n3853, new_n3852, n10096);
not_3  g01505(new_n3854, n16994);
nor_4  g01506(new_n3855, new_n3854, n16521);
not_3  g01507(new_n3856, n16521);
nor_4  g01508(new_n3857, n16994, new_n3856);
not_3  g01509(new_n3858, n7139);
nand_4 g01510(new_n3859, n9246, new_n3858);
nor_4  g01511(new_n3860, new_n3859, new_n3857);
nor_4  g01512(new_n3861, new_n3860, new_n3855);
nor_4  g01513(new_n3862, new_n3861, new_n3853);
nor_4  g01514(new_n3863, new_n3862, new_n3851);
nand_4 g01515(new_n3864, new_n3863, new_n3849);
nand_4 g01516(new_n3865, new_n3864, new_n3848);
nand_4 g01517(new_n3866, new_n3865, new_n3845);
nand_4 g01518(new_n3867, new_n3866, new_n3844);
nand_4 g01519(new_n3868, new_n3867, new_n3841);
nand_4 g01520(new_n3869_1, new_n3868, new_n3839);
nand_4 g01521(new_n3870, new_n3869_1, new_n3837);
nand_4 g01522(new_n3871_1, new_n3870, new_n3835);
nand_4 g01523(new_n3872, new_n3871_1, new_n3833);
nand_4 g01524(new_n3873, new_n3872, new_n3832);
nand_4 g01525(new_n3874, new_n3873, new_n3830);
not_3  g01526(new_n3875, new_n3874);
nor_4  g01527(new_n3876, new_n3875, new_n3829);
xor_3  g01528(new_n3877, new_n3876, new_n3827);
nor_4  g01529(new_n3878, n25565, n21993);
not_3  g01530(new_n3879, new_n3878);
nor_4  g01531(new_n3880, new_n3879, n11273);
not_3  g01532(new_n3881, new_n3880);
nor_4  g01533(new_n3882, new_n3881, n22290);
not_3  g01534(new_n3883, new_n3882);
nor_4  g01535(new_n3884, new_n3883, n9598);
not_3  g01536(new_n3885, new_n3884);
nor_4  g01537(new_n3886, new_n3885, n7670);
not_3  g01538(new_n3887, new_n3886);
nor_4  g01539(new_n3888, new_n3887, n13912);
not_3  g01540(new_n3889, new_n3888);
nor_4  g01541(new_n3890, new_n3889, n20213);
not_3  g01542(new_n3891_1, new_n3890);
nor_4  g01543(new_n3892, new_n3891_1, n21489);
not_3  g01544(new_n3893, new_n3892);
xor_3  g01545(new_n3894, new_n3893, n9259);
xnor_3 g01546(new_n3895, new_n3894, new_n3877);
xnor_3 g01547(new_n3896, new_n3873, new_n3830);
not_3  g01548(new_n3897, n21489);
xor_3  g01549(new_n3898, new_n3890, new_n3897);
not_3  g01550(new_n3899, new_n3898);
nor_4  g01551(new_n3900, new_n3899, new_n3896);
not_3  g01552(new_n3901, new_n3896);
xor_3  g01553(new_n3902, new_n3899, new_n3901);
not_3  g01554(new_n3903, new_n3833);
xnor_3 g01555(new_n3904, new_n3871_1, new_n3903);
xor_3  g01556(new_n3905, new_n3889, n20213);
nor_4  g01557(new_n3906, new_n3905, new_n3904);
not_3  g01558(new_n3907, new_n3906);
not_3  g01559(new_n3908, new_n3904);
not_3  g01560(new_n3909_1, new_n3905);
xor_3  g01561(new_n3910, new_n3909_1, new_n3908);
not_3  g01562(new_n3911, new_n3837);
xnor_3 g01563(new_n3912, new_n3869_1, new_n3911);
not_3  g01564(new_n3913, n13912);
xor_3  g01565(new_n3914, new_n3886, new_n3913);
nor_4  g01566(new_n3915, new_n3914, new_n3912);
not_3  g01567(new_n3916, new_n3915);
not_3  g01568(new_n3917, new_n3912);
not_3  g01569(new_n3918_1, new_n3914);
xor_3  g01570(new_n3919, new_n3918_1, new_n3917);
xnor_3 g01571(new_n3920, new_n3867, new_n3841);
xor_3  g01572(new_n3921, new_n3885, n7670);
not_3  g01573(new_n3922, new_n3921);
nand_4 g01574(new_n3923, new_n3922, new_n3920);
not_3  g01575(new_n3924, new_n3920);
nor_4  g01576(new_n3925_1, new_n3921, new_n3924);
nor_4  g01577(new_n3926, new_n3922, new_n3920);
nor_4  g01578(new_n3927, new_n3926, new_n3925_1);
xor_3  g01579(new_n3928, new_n3882, n9598);
not_3  g01580(new_n3929, new_n3928);
not_3  g01581(new_n3930, new_n3866);
nor_4  g01582(new_n3931, new_n3865, new_n3845);
nor_4  g01583(new_n3932_1, new_n3931, new_n3930);
nor_4  g01584(new_n3933, new_n3932_1, new_n3929);
not_3  g01585(new_n3934_1, new_n3933);
not_3  g01586(new_n3935, new_n3932_1);
nor_4  g01587(new_n3936, new_n3935, new_n3928);
nor_4  g01588(new_n3937, new_n3936, new_n3933);
xor_3  g01589(new_n3938, new_n3881, n22290);
xnor_3 g01590(new_n3939, new_n3863, new_n3849);
not_3  g01591(new_n3940, new_n3939);
nor_4  g01592(new_n3941, new_n3940, new_n3938);
not_3  g01593(new_n3942, new_n3941);
not_3  g01594(new_n3943, n11273);
xor_3  g01595(new_n3944, new_n3878, new_n3943);
nor_4  g01596(new_n3945_1, new_n3853, new_n3851);
xnor_3 g01597(new_n3946, new_n3945_1, new_n3861);
not_3  g01598(new_n3947, new_n3946);
nor_4  g01599(new_n3948, new_n3947, new_n3944);
not_3  g01600(new_n3949, new_n3948);
not_3  g01601(new_n3950, new_n3944);
nor_4  g01602(new_n3951, new_n3946, new_n3950);
nor_4  g01603(new_n3952_1, new_n3951, new_n3948);
xor_3  g01604(new_n3953, n25565, n21993);
not_3  g01605(new_n3954, new_n3953);
nor_4  g01606(new_n3955, new_n3857, new_n3855);
xnor_3 g01607(new_n3956, new_n3955, new_n3859);
nand_4 g01608(new_n3957, new_n3956, new_n3954);
xor_3  g01609(new_n3958, n9246, new_n3858);
not_3  g01610(new_n3959_1, new_n3958);
nand_4 g01611(new_n3960, new_n3959_1, n21993);
not_3  g01612(new_n3961, new_n3956);
nor_4  g01613(new_n3962_1, new_n3961, new_n3953);
nor_4  g01614(new_n3963, new_n3956, new_n3954);
nor_4  g01615(new_n3964, new_n3963, new_n3962_1);
nand_4 g01616(new_n3965, new_n3964, new_n3960);
nand_4 g01617(new_n3966, new_n3965, new_n3957);
nand_4 g01618(new_n3967, new_n3966, new_n3952_1);
nand_4 g01619(new_n3968, new_n3967, new_n3949);
not_3  g01620(new_n3969, new_n3938);
nor_4  g01621(new_n3970, new_n3939, new_n3969);
nor_4  g01622(new_n3971_1, new_n3970, new_n3941);
nand_4 g01623(new_n3972, new_n3971_1, new_n3968);
nand_4 g01624(new_n3973, new_n3972, new_n3942);
nand_4 g01625(new_n3974, new_n3973, new_n3937);
nand_4 g01626(new_n3975, new_n3974, new_n3934_1);
nand_4 g01627(new_n3976, new_n3975, new_n3927);
nand_4 g01628(new_n3977, new_n3976, new_n3923);
nand_4 g01629(new_n3978, new_n3977, new_n3919);
nand_4 g01630(new_n3979, new_n3978, new_n3916);
nand_4 g01631(new_n3980, new_n3979, new_n3910);
nand_4 g01632(new_n3981, new_n3980, new_n3907);
nor_4  g01633(new_n3982, new_n3981, new_n3902);
nor_4  g01634(new_n3983_1, new_n3982, new_n3900);
xnor_3 g01635(new_n3984_1, new_n3983_1, new_n3895);
xnor_3 g01636(new_n3985, new_n3984_1, new_n3824);
xnor_3 g01637(new_n3986, new_n3819, new_n3752);
not_3  g01638(new_n3987, new_n3981);
xnor_3 g01639(new_n3988, new_n3987, new_n3902);
nor_4  g01640(new_n3989, new_n3988, new_n3986);
not_3  g01641(new_n3990, new_n3989);
not_3  g01642(new_n3991, new_n3986);
not_3  g01643(new_n3992, new_n3988);
nor_4  g01644(new_n3993, new_n3992, new_n3991);
nor_4  g01645(new_n3994, new_n3993, new_n3989);
not_3  g01646(new_n3995, new_n3758_1);
xnor_3 g01647(new_n3996, new_n3817, new_n3995);
xnor_3 g01648(new_n3997, new_n3979, new_n3910);
not_3  g01649(new_n3998, new_n3997);
nand_4 g01650(new_n3999, new_n3998, new_n3996);
xnor_3 g01651(new_n4000_1, new_n3997, new_n3996);
xnor_3 g01652(new_n4001, new_n3815, new_n3766);
xnor_3 g01653(new_n4002, new_n3977, new_n3919);
nor_4  g01654(new_n4003, new_n4002, new_n4001);
not_3  g01655(new_n4004, new_n4003);
not_3  g01656(new_n4005, new_n4001);
not_3  g01657(new_n4006, new_n4002);
nor_4  g01658(new_n4007, new_n4006, new_n4005);
nor_4  g01659(new_n4008, new_n4007, new_n4003);
xnor_3 g01660(new_n4009, new_n3813, new_n3775);
not_3  g01661(new_n4010_1, new_n4009);
not_3  g01662(new_n4011, new_n3927);
xnor_3 g01663(new_n4012, new_n3975, new_n4011);
nand_4 g01664(new_n4013, new_n4012, new_n4010_1);
xnor_3 g01665(new_n4014_1, new_n4012, new_n4009);
not_3  g01666(new_n4015, new_n3812);
nor_4  g01667(new_n4016, new_n3811, new_n3782);
nor_4  g01668(new_n4017, new_n4016, new_n4015);
not_3  g01669(new_n4018, new_n4017);
xnor_3 g01670(new_n4019, new_n3973, new_n3937);
nor_4  g01671(new_n4020, new_n4019, new_n4018);
not_3  g01672(new_n4021, new_n4020);
not_3  g01673(new_n4022, new_n4019);
nor_4  g01674(new_n4023, new_n4022, new_n4017);
nor_4  g01675(new_n4024, new_n4023, new_n4020);
xnor_3 g01676(new_n4025, new_n3809, new_n3789);
xnor_3 g01677(new_n4026, new_n3971_1, new_n3968);
nor_4  g01678(new_n4027, new_n4026, new_n4025);
not_3  g01679(new_n4028, new_n4027);
not_3  g01680(new_n4029, new_n4025);
not_3  g01681(new_n4030, new_n4026);
nor_4  g01682(new_n4031, new_n4030, new_n4029);
nor_4  g01683(new_n4032, new_n4031, new_n4027);
xnor_3 g01684(new_n4033, new_n3807, new_n3796);
not_3  g01685(new_n4034, new_n3952_1);
xnor_3 g01686(new_n4035, new_n3966, new_n4034);
nand_4 g01687(new_n4036, new_n4035, new_n4033);
not_3  g01688(new_n4037, new_n4033);
xnor_3 g01689(new_n4038, new_n4035, new_n4037);
xnor_3 g01690(new_n4039, new_n3964, new_n3960);
xnor_3 g01691(new_n4040, new_n3805, new_n3802);
not_3  g01692(new_n4041, new_n4040);
nor_4  g01693(new_n4042, new_n4041, new_n4039);
not_3  g01694(new_n4043, new_n4042);
not_3  g01695(new_n4044, new_n3802);
nor_4  g01696(new_n4045, new_n3801, n18578);
nor_4  g01697(new_n4046, new_n4045, new_n4044);
not_3  g01698(new_n4047, new_n4046);
not_3  g01699(new_n4048, new_n3960);
nor_4  g01700(new_n4049, new_n3959_1, n21993);
nor_4  g01701(new_n4050, new_n4049, new_n4048);
not_3  g01702(new_n4051, new_n4050);
nor_4  g01703(new_n4052, new_n4051, new_n4047);
not_3  g01704(new_n4053, new_n4052);
not_3  g01705(new_n4054, new_n4039);
nor_4  g01706(new_n4055, new_n4040, new_n4054);
nor_4  g01707(new_n4056, new_n4055, new_n4042);
nand_4 g01708(new_n4057, new_n4056, new_n4053);
nand_4 g01709(new_n4058, new_n4057, new_n4043);
nand_4 g01710(new_n4059, new_n4058, new_n4038);
nand_4 g01711(new_n4060, new_n4059, new_n4036);
nand_4 g01712(new_n4061, new_n4060, new_n4032);
nand_4 g01713(new_n4062, new_n4061, new_n4028);
nand_4 g01714(new_n4063, new_n4062, new_n4024);
nand_4 g01715(new_n4064, new_n4063, new_n4021);
nand_4 g01716(new_n4065, new_n4064, new_n4014_1);
nand_4 g01717(new_n4066, new_n4065, new_n4013);
nand_4 g01718(new_n4067, new_n4066, new_n4008);
nand_4 g01719(new_n4068, new_n4067, new_n4004);
nand_4 g01720(new_n4069, new_n4068, new_n4000_1);
nand_4 g01721(new_n4070, new_n4069, new_n3999);
nand_4 g01722(new_n4071_1, new_n4070, new_n3994);
nand_4 g01723(new_n4072, new_n4071_1, new_n3990);
xnor_3 g01724(n235, new_n4072, new_n3985);
not_3  g01725(new_n4074, n2113);
not_3  g01726(new_n4075, n6369);
not_3  g01727(new_n4076, n15967);
nor_4  g01728(new_n4077, n25435, n13319);
nand_4 g01729(new_n4078, new_n4077, new_n4076);
nor_4  g01730(new_n4079, new_n4078, n25797);
nand_4 g01731(new_n4080, new_n4079, new_n4075);
nor_4  g01732(new_n4081, new_n4080, n21134);
xor_3  g01733(new_n4082, new_n4081, new_n4074);
not_3  g01734(new_n4083, new_n4082);
xor_3  g01735(new_n4084, new_n4083, n19327);
xor_3  g01736(new_n4085_1, new_n4080, n21134);
nor_4  g01737(new_n4086, new_n4085_1, n22597);
not_3  g01738(new_n4087, new_n4085_1);
xor_3  g01739(new_n4088_1, new_n4087, n22597);
not_3  g01740(new_n4089_1, new_n4080);
nor_4  g01741(new_n4090, new_n4079, new_n4075);
nor_4  g01742(new_n4091, new_n4090, new_n4089_1);
nor_4  g01743(new_n4092, new_n4091, n26107);
not_3  g01744(new_n4093, n26107);
not_3  g01745(new_n4094, new_n4091);
nor_4  g01746(new_n4095, new_n4094, new_n4093);
nor_4  g01747(new_n4096, new_n4095, new_n4092);
nand_4 g01748(new_n4097, new_n4078, n25797);
not_3  g01749(new_n4098, new_n4097);
nor_4  g01750(new_n4099, new_n4098, new_n4079);
nor_4  g01751(new_n4100_1, new_n4099, n342);
not_3  g01752(new_n4101, new_n4100_1);
not_3  g01753(new_n4102, new_n4078);
nor_4  g01754(new_n4103_1, new_n4077, new_n4076);
nor_4  g01755(new_n4104, new_n4103_1, new_n4102);
nor_4  g01756(new_n4105, new_n4104, n26553);
not_3  g01757(new_n4106, new_n4105);
not_3  g01758(new_n4107, n26553);
not_3  g01759(new_n4108, new_n4104);
nor_4  g01760(new_n4109, new_n4108, new_n4107);
nor_4  g01761(new_n4110, new_n4109, new_n4105);
xnor_3 g01762(new_n4111, n25435, n13319);
not_3  g01763(new_n4112, new_n4111);
nor_4  g01764(new_n4113, new_n4112, n4964);
not_3  g01765(new_n4114, new_n4113);
nand_4 g01766(new_n4115, n25435, n7876);
not_3  g01767(new_n4116, n4964);
nor_4  g01768(new_n4117, new_n4111, new_n4116);
nor_4  g01769(new_n4118, new_n4117, new_n4113);
nand_4 g01770(new_n4119_1, new_n4118, new_n4115);
nand_4 g01771(new_n4120, new_n4119_1, new_n4114);
nand_4 g01772(new_n4121, new_n4120, new_n4110);
nand_4 g01773(new_n4122, new_n4121, new_n4106);
not_3  g01774(new_n4123_1, n342);
not_3  g01775(new_n4124, new_n4099);
nor_4  g01776(new_n4125, new_n4124, new_n4123_1);
nor_4  g01777(new_n4126, new_n4125, new_n4100_1);
nand_4 g01778(new_n4127, new_n4126, new_n4122);
nand_4 g01779(new_n4128, new_n4127, new_n4101);
nand_4 g01780(new_n4129, new_n4128, new_n4096);
not_3  g01781(new_n4130, new_n4129);
nor_4  g01782(new_n4131, new_n4130, new_n4092);
nor_4  g01783(new_n4132, new_n4131, new_n4088_1);
nor_4  g01784(new_n4133, new_n4132, new_n4086);
xnor_3 g01785(new_n4134_1, new_n4133, new_n4084);
xnor_3 g01786(new_n4135, new_n4134_1, n25749);
not_3  g01787(new_n4136, n3161);
not_3  g01788(new_n4137, new_n4131);
xnor_3 g01789(new_n4138, new_n4137, new_n4088_1);
nor_4  g01790(new_n4139, new_n4138, new_n4136);
xnor_3 g01791(new_n4140, new_n4138, new_n4136);
not_3  g01792(new_n4141, n9003);
xnor_3 g01793(new_n4142, new_n4128, new_n4096);
not_3  g01794(new_n4143, new_n4142);
nor_4  g01795(new_n4144, new_n4143, new_n4141);
not_3  g01796(new_n4145, new_n4144);
nor_4  g01797(new_n4146_1, new_n4142, n9003);
nor_4  g01798(new_n4147, new_n4146_1, new_n4144);
not_3  g01799(new_n4148, n4957);
xnor_3 g01800(new_n4149, new_n4126, new_n4122);
not_3  g01801(new_n4150_1, new_n4149);
nor_4  g01802(new_n4151_1, new_n4150_1, new_n4148);
not_3  g01803(new_n4152_1, new_n4151_1);
nor_4  g01804(new_n4153_1, new_n4149, n4957);
nor_4  g01805(new_n4154, new_n4153_1, new_n4151_1);
not_3  g01806(new_n4155, n7524);
xnor_3 g01807(new_n4156, new_n4120, new_n4110);
not_3  g01808(new_n4157, new_n4156);
nor_4  g01809(new_n4158, new_n4157, new_n4155);
not_3  g01810(new_n4159, new_n4158);
nor_4  g01811(new_n4160, new_n4156, n7524);
nor_4  g01812(new_n4161, new_n4160, new_n4158);
not_3  g01813(new_n4162, n15743);
xnor_3 g01814(new_n4163, new_n4118, new_n4115);
not_3  g01815(new_n4164, new_n4163);
nor_4  g01816(new_n4165_1, new_n4164, new_n4162);
not_3  g01817(new_n4166, new_n4165_1);
not_3  g01818(new_n4167, n20658);
not_3  g01819(new_n4168, n7876);
xor_3  g01820(new_n4169, n25435, new_n4168);
nor_4  g01821(new_n4170, new_n4169, new_n4167);
nor_4  g01822(new_n4171, new_n4163, n15743);
nor_4  g01823(new_n4172_1, new_n4171, new_n4165_1);
nand_4 g01824(new_n4173_1, new_n4172_1, new_n4170);
nand_4 g01825(new_n4174, new_n4173_1, new_n4166);
nand_4 g01826(new_n4175, new_n4174, new_n4161);
nand_4 g01827(new_n4176_1, new_n4175, new_n4159);
nand_4 g01828(new_n4177, new_n4176_1, new_n4154);
nand_4 g01829(new_n4178, new_n4177, new_n4152_1);
nand_4 g01830(new_n4179, new_n4178, new_n4147);
nand_4 g01831(new_n4180, new_n4179, new_n4145);
not_3  g01832(new_n4181, new_n4180);
nor_4  g01833(new_n4182, new_n4181, new_n4140);
nor_4  g01834(new_n4183, new_n4182, new_n4139);
xnor_3 g01835(new_n4184, new_n4183, new_n4135);
not_3  g01836(new_n4185, n22332);
xor_3  g01837(new_n4186_1, n26510, new_n4185);
not_3  g01838(new_n4187, n23068);
nand_4 g01839(new_n4188, new_n4187, n18907);
xor_3  g01840(new_n4189, n23068, new_n2443);
not_3  g01841(new_n4190, n2731);
nor_4  g01842(new_n4191, n19514, new_n4190);
not_3  g01843(new_n4192, new_n4191);
xor_3  g01844(new_n4193, n19514, new_n4190);
not_3  g01845(new_n4194, n19911);
nor_4  g01846(new_n4195, new_n4194, n10053);
not_3  g01847(new_n4196, new_n4195);
not_3  g01848(new_n4197, n10053);
xor_3  g01849(new_n4198, n19911, new_n4197);
not_3  g01850(new_n4199, n8399);
nor_4  g01851(new_n4200, n13708, new_n4199);
not_3  g01852(new_n4201, n13708);
nor_4  g01853(new_n4202, new_n4201, n8399);
not_3  g01854(new_n4203, n9507);
nor_4  g01855(new_n4204_1, n18409, new_n4203);
not_3  g01856(new_n4205_1, n18409);
nor_4  g01857(new_n4206, new_n4205_1, n9507);
nand_4 g01858(new_n4207, n26979, new_n2389);
nor_4  g01859(new_n4208, new_n4207, new_n4206);
nor_4  g01860(new_n4209, new_n4208, new_n4204_1);
nor_4  g01861(new_n4210, new_n4209, new_n4202);
nor_4  g01862(new_n4211, new_n4210, new_n4200);
nand_4 g01863(new_n4212, new_n4211, new_n4198);
nand_4 g01864(new_n4213, new_n4212, new_n4196);
nand_4 g01865(new_n4214, new_n4213, new_n4193);
nand_4 g01866(new_n4215_1, new_n4214, new_n4192);
nand_4 g01867(new_n4216, new_n4215_1, new_n4189);
nand_4 g01868(new_n4217, new_n4216, new_n4188);
xnor_3 g01869(new_n4218, new_n4217, new_n4186_1);
not_3  g01870(new_n4219, n4325);
not_3  g01871(new_n4220, n19618);
nor_4  g01872(new_n4221_1, n22043, n12121);
nand_4 g01873(new_n4222, new_n4221_1, new_n4220);
nor_4  g01874(new_n4223, new_n4222, n1204);
not_3  g01875(new_n4224_1, new_n4223);
nor_4  g01876(new_n4225, new_n4224_1, n626);
not_3  g01877(new_n4226, new_n4225);
nor_4  g01878(new_n4227, new_n4226, n5337);
xor_3  g01879(new_n4228, new_n4227, new_n4219);
xnor_3 g01880(new_n4229, new_n4228, new_n4218);
xnor_3 g01881(new_n4230, new_n4215_1, new_n4189);
not_3  g01882(new_n4231_1, n5337);
xor_3  g01883(new_n4232, new_n4225, new_n4231_1);
not_3  g01884(new_n4233, new_n4232);
nand_4 g01885(new_n4234, new_n4233, new_n4230);
xnor_3 g01886(new_n4235, new_n4232, new_n4230);
not_3  g01887(new_n4236, new_n4193);
xnor_3 g01888(new_n4237, new_n4213, new_n4236);
not_3  g01889(new_n4238, n626);
xor_3  g01890(new_n4239, new_n4223, new_n4238);
nor_4  g01891(new_n4240, new_n4239, new_n4237);
not_3  g01892(new_n4241, new_n4240);
not_3  g01893(new_n4242, new_n4237);
not_3  g01894(new_n4243, new_n4239);
nor_4  g01895(new_n4244, new_n4243, new_n4242);
nor_4  g01896(new_n4245, new_n4244, new_n4240);
not_3  g01897(new_n4246, n1204);
xor_3  g01898(new_n4247, new_n4222, new_n4246);
not_3  g01899(new_n4248, new_n4247);
not_3  g01900(new_n4249, new_n4211);
xnor_3 g01901(new_n4250, new_n4249, new_n4198);
nor_4  g01902(new_n4251, new_n4250, new_n4248);
not_3  g01903(new_n4252, new_n4251);
not_3  g01904(new_n4253, new_n4250);
nor_4  g01905(new_n4254, new_n4253, new_n4247);
nor_4  g01906(new_n4255, new_n4254, new_n4251);
xor_3  g01907(new_n4256_1, new_n4221_1, n19618);
nor_4  g01908(new_n4257, new_n4202, new_n4200);
not_3  g01909(new_n4258, new_n4257);
xnor_3 g01910(new_n4259, new_n4258, new_n4209);
not_3  g01911(new_n4260, new_n4259);
nand_4 g01912(new_n4261, new_n4260, new_n4256_1);
xnor_3 g01913(new_n4262, new_n4259, new_n4256_1);
xor_3  g01914(new_n4263, n22043, n12121);
not_3  g01915(new_n4264, new_n4263);
nor_4  g01916(new_n4265, new_n4206, new_n4204_1);
xnor_3 g01917(new_n4266_1, new_n4265, new_n4207);
nor_4  g01918(new_n4267, new_n4266_1, new_n4264);
xor_3  g01919(new_n4268, n26979, n5704);
nand_4 g01920(new_n4269, new_n4268, n12121);
not_3  g01921(new_n4270, new_n4266_1);
xnor_3 g01922(new_n4271, new_n4270, new_n4263);
nor_4  g01923(new_n4272_1, new_n4271, new_n4269);
nor_4  g01924(new_n4273, new_n4272_1, new_n4267);
nand_4 g01925(new_n4274, new_n4273, new_n4262);
nand_4 g01926(new_n4275, new_n4274, new_n4261);
nand_4 g01927(new_n4276, new_n4275, new_n4255);
nand_4 g01928(new_n4277, new_n4276, new_n4252);
nand_4 g01929(new_n4278, new_n4277, new_n4245);
nand_4 g01930(new_n4279, new_n4278, new_n4241);
nand_4 g01931(new_n4280, new_n4279, new_n4235);
nand_4 g01932(new_n4281, new_n4280, new_n4234);
xnor_3 g01933(new_n4282, new_n4281, new_n4229);
not_3  g01934(new_n4283, new_n4282);
xnor_3 g01935(new_n4284, new_n4283, new_n4184);
xnor_3 g01936(new_n4285, new_n4279, new_n4235);
not_3  g01937(new_n4286, new_n4140);
nor_4  g01938(new_n4287, new_n4180, new_n4286);
nor_4  g01939(new_n4288, new_n4287, new_n4182);
nor_4  g01940(new_n4289, new_n4288, new_n4285);
not_3  g01941(new_n4290, new_n4289);
not_3  g01942(new_n4291, new_n4285);
xnor_3 g01943(new_n4292, new_n4288, new_n4291);
xnor_3 g01944(new_n4293, new_n4277, new_n4245);
not_3  g01945(new_n4294, new_n4293);
xnor_3 g01946(new_n4295, new_n4178, new_n4147);
nand_4 g01947(new_n4296, new_n4295, new_n4294);
xnor_3 g01948(new_n4297, new_n4295, new_n4293);
xnor_3 g01949(new_n4298, new_n4275, new_n4255);
not_3  g01950(new_n4299, new_n4298);
xnor_3 g01951(new_n4300, new_n4176_1, new_n4154);
nand_4 g01952(new_n4301, new_n4300, new_n4299);
xnor_3 g01953(new_n4302, new_n4300, new_n4298);
not_3  g01954(new_n4303, new_n4267);
not_3  g01955(new_n4304, new_n4272_1);
nand_4 g01956(new_n4305, new_n4304, new_n4303);
xnor_3 g01957(new_n4306_1, new_n4305, new_n4262);
xnor_3 g01958(new_n4307, new_n4174, new_n4161);
nand_4 g01959(new_n4308, new_n4307, new_n4306_1);
not_3  g01960(new_n4309, new_n4306_1);
xnor_3 g01961(new_n4310, new_n4307, new_n4309);
xnor_3 g01962(new_n4311, new_n4271, new_n4269);
xnor_3 g01963(new_n4312, new_n4172_1, new_n4170);
nand_4 g01964(new_n4313, new_n4312, new_n4311);
not_3  g01965(new_n4314, new_n4169);
xor_3  g01966(new_n4315, new_n4314, n20658);
not_3  g01967(new_n4316, new_n4269);
nor_4  g01968(new_n4317, new_n4268, n12121);
nor_4  g01969(new_n4318, new_n4317, new_n4316);
nand_4 g01970(new_n4319_1, new_n4318, new_n4315);
not_3  g01971(new_n4320, new_n4313);
nor_4  g01972(new_n4321, new_n4312, new_n4311);
nor_4  g01973(new_n4322, new_n4321, new_n4320);
nand_4 g01974(new_n4323, new_n4322, new_n4319_1);
nand_4 g01975(new_n4324, new_n4323, new_n4313);
nand_4 g01976(new_n4325_1, new_n4324, new_n4310);
nand_4 g01977(new_n4326_1, new_n4325_1, new_n4308);
nand_4 g01978(new_n4327, new_n4326_1, new_n4302);
nand_4 g01979(new_n4328, new_n4327, new_n4301);
nand_4 g01980(new_n4329, new_n4328, new_n4297);
nand_4 g01981(new_n4330, new_n4329, new_n4296);
nand_4 g01982(new_n4331, new_n4330, new_n4292);
nand_4 g01983(new_n4332, new_n4331, new_n4290);
xor_3  g01984(n242, new_n4332, new_n4284);
not_3  g01985(new_n4334, n13677);
not_3  g01986(new_n4335, n11011);
not_3  g01987(new_n4336, n11223);
not_3  g01988(new_n4337, n26572);
nor_4  g01989(new_n4338, n21398, n11667);
nand_4 g01990(new_n4339, new_n4338, new_n4337);
nor_4  g01991(new_n4340_1, new_n4339, n5115);
nand_4 g01992(new_n4341, new_n4340_1, new_n4336);
nor_4  g01993(new_n4342, new_n4341, n19477);
nand_4 g01994(new_n4343, new_n4341, n19477);
not_3  g01995(new_n4344, new_n4343);
nor_4  g01996(new_n4345, new_n4344, new_n4342);
not_3  g01997(new_n4346, new_n4345);
nor_4  g01998(new_n4347, new_n4346, new_n4335);
nor_4  g01999(new_n4348, new_n4345, n11011);
nor_4  g02000(new_n4349, new_n4348, new_n4347);
not_3  g02001(new_n4350, new_n4341);
nor_4  g02002(new_n4351, new_n4340_1, new_n4336);
nor_4  g02003(new_n4352, new_n4351, new_n4350);
nor_4  g02004(new_n4353, new_n4352, n16029);
not_3  g02005(new_n4354, new_n4353);
not_3  g02006(new_n4355, n16029);
not_3  g02007(new_n4356, new_n4352);
nor_4  g02008(new_n4357, new_n4356, new_n4355);
nor_4  g02009(new_n4358, new_n4357, new_n4353);
not_3  g02010(new_n4359, n16476);
nand_4 g02011(new_n4360, new_n4339, n5115);
not_3  g02012(new_n4361, new_n4360);
nor_4  g02013(new_n4362, new_n4361, new_n4340_1);
not_3  g02014(new_n4363, new_n4362);
nor_4  g02015(new_n4364, new_n4363, new_n4359);
xnor_3 g02016(new_n4365, new_n4362, n16476);
not_3  g02017(new_n4366, new_n4339);
nor_4  g02018(new_n4367, new_n4338, new_n4337);
nor_4  g02019(new_n4368, new_n4367, new_n4366);
nor_4  g02020(new_n4369, new_n4368, n11615);
not_3  g02021(new_n4370, new_n4369);
not_3  g02022(new_n4371, n11615);
not_3  g02023(new_n4372, new_n4368);
nor_4  g02024(new_n4373, new_n4372, new_n4371);
nor_4  g02025(new_n4374_1, new_n4373, new_n4369);
not_3  g02026(new_n4375, n22433);
xnor_3 g02027(new_n4376_1, n21398, n11667);
nand_4 g02028(new_n4377, new_n4376_1, new_n4375);
nand_4 g02029(new_n4378, n21398, n14090);
xnor_3 g02030(new_n4379, new_n4376_1, n22433);
nand_4 g02031(new_n4380, new_n4379, new_n4378);
nand_4 g02032(new_n4381, new_n4380, new_n4377);
nand_4 g02033(new_n4382, new_n4381, new_n4374_1);
nand_4 g02034(new_n4383, new_n4382, new_n4370);
nor_4  g02035(new_n4384, new_n4383, new_n4365);
nor_4  g02036(new_n4385, new_n4384, new_n4364);
nand_4 g02037(new_n4386, new_n4385, new_n4358);
nand_4 g02038(new_n4387, new_n4386, new_n4354);
xnor_3 g02039(new_n4388, new_n4387, new_n4349);
not_3  g02040(new_n4389, new_n4388);
nor_4  g02041(new_n4390, new_n4389, new_n4334);
nor_4  g02042(new_n4391, new_n4388, n13677);
nor_4  g02043(new_n4392, new_n4391, new_n4390);
xnor_3 g02044(new_n4393, new_n4385, new_n4358);
nor_4  g02045(new_n4394, new_n4393, n18926);
not_3  g02046(new_n4395, new_n4365);
xnor_3 g02047(new_n4396, new_n4383, new_n4395);
nand_4 g02048(new_n4397, new_n4396, n5451);
not_3  g02049(new_n4398, new_n4397);
nor_4  g02050(new_n4399, new_n4396, n5451);
nor_4  g02051(new_n4400, new_n4399, new_n4398);
not_3  g02052(new_n4401_1, n5330);
xnor_3 g02053(new_n4402, new_n4381, new_n4374_1);
not_3  g02054(new_n4403, new_n4402);
nor_4  g02055(new_n4404, new_n4403, new_n4401_1);
not_3  g02056(new_n4405, new_n4404);
xnor_3 g02057(new_n4406, new_n4402, n5330);
not_3  g02058(new_n4407, new_n4406);
not_3  g02059(new_n4408, n7657);
xnor_3 g02060(new_n4409_1, new_n4379, new_n4378);
not_3  g02061(new_n4410, new_n4409_1);
nor_4  g02062(new_n4411, new_n4410, new_n4408);
not_3  g02063(new_n4412, new_n4411);
nor_4  g02064(new_n4413, new_n4409_1, n7657);
nor_4  g02065(new_n4414, new_n4413, new_n4411);
nand_4 g02066(new_n4415, new_n4414, new_n2607);
nand_4 g02067(new_n4416, new_n4415, new_n4412);
nand_4 g02068(new_n4417, new_n4416, new_n4407);
nand_4 g02069(new_n4418, new_n4417, new_n4405);
nand_4 g02070(new_n4419, new_n4418, new_n4400);
nand_4 g02071(new_n4420, new_n4419, new_n4397);
xnor_3 g02072(new_n4421, new_n4393, n18926);
nor_4  g02073(new_n4422, new_n4421, new_n4420);
nor_4  g02074(new_n4423, new_n4422, new_n4394);
not_3  g02075(new_n4424_1, new_n4423);
xnor_3 g02076(new_n4425, new_n4424_1, new_n4392);
not_3  g02077(new_n4426_1, n12398);
nor_4  g02078(new_n4427, n21687, n6729);
not_3  g02079(new_n4428, new_n4427);
nor_4  g02080(new_n4429, new_n4428, n8285);
not_3  g02081(new_n4430, new_n4429);
nor_4  g02082(new_n4431, new_n4430, n20169);
not_3  g02083(new_n4432_1, new_n4431);
nor_4  g02084(new_n4433, new_n4432_1, n19789);
xor_3  g02085(new_n4434, new_n4433, new_n4426_1);
not_3  g02086(new_n4435, new_n4434);
not_3  g02087(new_n4436, n15424);
not_3  g02088(new_n4437, n9323);
nor_4  g02089(new_n4438, n19922, n10792);
nand_4 g02090(new_n4439, new_n4438, new_n4437);
nor_4  g02091(new_n4440, new_n4439, n1949);
nand_4 g02092(new_n4441_1, new_n4440, new_n4436);
nor_4  g02093(new_n4442, new_n4441_1, n25694);
nand_4 g02094(new_n4443, new_n4441_1, n25694);
not_3  g02095(new_n4444, new_n4443);
nor_4  g02096(new_n4445, new_n4444, new_n4442);
xor_3  g02097(new_n4446, new_n4445, n20151);
not_3  g02098(new_n4447, n7693);
xnor_3 g02099(new_n4448, new_n4440, new_n4436);
nor_4  g02100(new_n4449, new_n4448, new_n4447);
not_3  g02101(new_n4450, new_n4449);
not_3  g02102(new_n4451_1, n10405);
nand_4 g02103(new_n4452, new_n4439, n1949);
not_3  g02104(new_n4453, new_n4452);
nor_4  g02105(new_n4454, new_n4453, new_n4440);
not_3  g02106(new_n4455, new_n4454);
nor_4  g02107(new_n4456, new_n4455, new_n4451_1);
nor_4  g02108(new_n4457, new_n4454, n10405);
nor_4  g02109(new_n4458, new_n4457, new_n4456);
not_3  g02110(new_n4459, new_n4458);
not_3  g02111(new_n4460, n10792);
not_3  g02112(new_n4461, n19922);
nand_4 g02113(new_n4462, new_n4461, new_n4460);
nor_4  g02114(new_n4463, new_n4462, n9323);
nor_4  g02115(new_n4464, new_n4438, new_n4437);
nor_4  g02116(new_n4465, new_n4464, new_n4463);
nor_4  g02117(new_n4466, new_n4465, n11302);
not_3  g02118(new_n4467, new_n4466);
xnor_3 g02119(new_n4468, new_n4465, n11302);
not_3  g02120(new_n4469, new_n4468);
nand_4 g02121(new_n4470, n19922, n10792);
nand_4 g02122(new_n4471, new_n4470, new_n4462);
not_3  g02123(new_n4472, new_n4471);
nor_4  g02124(new_n4473, new_n4472, n17090);
not_3  g02125(new_n4474, new_n4473);
nand_4 g02126(new_n4475, n19922, n6773);
not_3  g02127(new_n4476_1, new_n4475);
not_3  g02128(new_n4477, n17090);
xnor_3 g02129(new_n4478_1, new_n4471, new_n4477);
nor_4  g02130(new_n4479, new_n4478_1, new_n4476_1);
not_3  g02131(new_n4480, new_n4479);
nand_4 g02132(new_n4481, new_n4480, new_n4474);
nand_4 g02133(new_n4482, new_n4481, new_n4469);
nand_4 g02134(new_n4483, new_n4482, new_n4467);
nor_4  g02135(new_n4484, new_n4483, new_n4459);
nor_4  g02136(new_n4485, new_n4484, new_n4456);
not_3  g02137(new_n4486, new_n4485);
xor_3  g02138(new_n4487, new_n4448, new_n4447);
nand_4 g02139(new_n4488, new_n4487, new_n4486);
nand_4 g02140(new_n4489, new_n4488, new_n4450);
xnor_3 g02141(new_n4490, new_n4489, new_n4446);
nor_4  g02142(new_n4491, new_n4490, new_n4435);
not_3  g02143(new_n4492, new_n4490);
nor_4  g02144(new_n4493, new_n4492, new_n4434);
nor_4  g02145(new_n4494, new_n4493, new_n4491);
xor_3  g02146(new_n4495, new_n4431, n19789);
xor_3  g02147(new_n4496, new_n4448, n7693);
xnor_3 g02148(new_n4497, new_n4496, new_n4485);
nor_4  g02149(new_n4498, new_n4497, new_n4495);
not_3  g02150(new_n4499, new_n4498);
not_3  g02151(new_n4500, new_n4495);
nor_4  g02152(new_n4501, new_n4496, new_n4485);
nor_4  g02153(new_n4502, new_n4487, new_n4486);
nor_4  g02154(new_n4503, new_n4502, new_n4501);
nor_4  g02155(new_n4504, new_n4503, new_n4500);
nor_4  g02156(new_n4505, new_n4504, new_n4498);
xnor_3 g02157(new_n4506, new_n4483, new_n4458);
not_3  g02158(new_n4507, n20169);
xor_3  g02159(new_n4508, new_n4429, new_n4507);
nor_4  g02160(new_n4509, new_n4508, new_n4506);
not_3  g02161(new_n4510, new_n4506);
xnor_3 g02162(new_n4511, new_n4508, new_n4510);
not_3  g02163(new_n4512, new_n4511);
xnor_3 g02164(new_n4513, new_n4481, new_n4469);
not_3  g02165(new_n4514_1, new_n4513);
xor_3  g02166(new_n4515, new_n4427, n8285);
nor_4  g02167(new_n4516, new_n4515, new_n4514_1);
not_3  g02168(new_n4517, new_n4516);
not_3  g02169(new_n4518, new_n4515);
nor_4  g02170(new_n4519, new_n4518, new_n4513);
nor_4  g02171(new_n4520, new_n4519, new_n4516);
nand_4 g02172(new_n4521, n21687, n6729);
not_3  g02173(new_n4522, new_n4521);
nor_4  g02174(new_n4523, new_n4522, new_n4427);
not_3  g02175(new_n4524, new_n4523);
xnor_3 g02176(new_n4525, new_n4478_1, new_n4476_1);
not_3  g02177(new_n4526, new_n4525);
nor_4  g02178(new_n4527, new_n4526, new_n4524);
not_3  g02179(new_n4528, new_n4527);
nor_4  g02180(new_n4529_1, new_n2603, new_n2601);
not_3  g02181(new_n4530, new_n4529_1);
xnor_3 g02182(new_n4531, new_n4525, new_n4523);
nor_4  g02183(new_n4532, new_n4531, new_n4530);
not_3  g02184(new_n4533, new_n4532);
nand_4 g02185(new_n4534, new_n4533, new_n4528);
nand_4 g02186(new_n4535, new_n4534, new_n4520);
nand_4 g02187(new_n4536, new_n4535, new_n4517);
nor_4  g02188(new_n4537, new_n4536, new_n4512);
nor_4  g02189(new_n4538, new_n4537, new_n4509);
nand_4 g02190(new_n4539, new_n4538, new_n4505);
nand_4 g02191(new_n4540, new_n4539, new_n4499);
xnor_3 g02192(new_n4541, new_n4540, new_n4494);
xnor_3 g02193(new_n4542, new_n4541, new_n4425);
xnor_3 g02194(new_n4543, new_n4497, new_n4495);
not_3  g02195(new_n4544, new_n4538);
xnor_3 g02196(new_n4545, new_n4544, new_n4543);
xnor_3 g02197(new_n4546, new_n4421, new_n4420);
not_3  g02198(new_n4547, new_n4546);
nand_4 g02199(new_n4548, new_n4547, new_n4545);
xnor_3 g02200(new_n4549, new_n4546, new_n4545);
not_3  g02201(new_n4550, new_n4520);
nor_4  g02202(new_n4551, new_n4532, new_n4527);
nor_4  g02203(new_n4552_1, new_n4551, new_n4550);
nor_4  g02204(new_n4553, new_n4552_1, new_n4516);
nor_4  g02205(new_n4554, new_n4553, new_n4511);
nor_4  g02206(new_n4555, new_n4554, new_n4537);
not_3  g02207(new_n4556, new_n4419);
nor_4  g02208(new_n4557, new_n4418, new_n4400);
nor_4  g02209(new_n4558, new_n4557, new_n4556);
not_3  g02210(new_n4559, new_n4558);
nand_4 g02211(new_n4560, new_n4559, new_n4555);
xnor_3 g02212(new_n4561, new_n4558, new_n4555);
xnor_3 g02213(new_n4562, new_n4416, new_n4406);
not_3  g02214(new_n4563, new_n4562);
xnor_3 g02215(new_n4564, new_n4534, new_n4520);
nand_4 g02216(new_n4565, new_n4564, new_n4563);
xnor_3 g02217(new_n4566, new_n4564, new_n4562);
not_3  g02218(new_n4567, new_n4531);
nor_4  g02219(new_n4568, new_n4567, new_n4529_1);
nor_4  g02220(new_n4569, new_n4568, new_n4532);
not_3  g02221(new_n4570, new_n4414);
xnor_3 g02222(new_n4571, new_n4570, new_n2606);
not_3  g02223(new_n4572, new_n4571);
nor_4  g02224(new_n4573, new_n4572, new_n4569);
not_3  g02225(new_n4574, new_n4573);
not_3  g02226(new_n4575, new_n2604);
not_3  g02227(new_n4576, new_n2609);
nor_4  g02228(new_n4577, new_n4576, new_n4575);
not_3  g02229(new_n4578, new_n4577);
not_3  g02230(new_n4579, new_n4569);
nor_4  g02231(new_n4580, new_n4571, new_n4579);
nor_4  g02232(new_n4581, new_n4580, new_n4573);
nand_4 g02233(new_n4582, new_n4581, new_n4578);
nand_4 g02234(new_n4583, new_n4582, new_n4574);
nand_4 g02235(new_n4584, new_n4583, new_n4566);
nand_4 g02236(new_n4585, new_n4584, new_n4565);
nand_4 g02237(new_n4586, new_n4585, new_n4561);
nand_4 g02238(new_n4587, new_n4586, new_n4560);
nand_4 g02239(new_n4588_1, new_n4587, new_n4549);
nand_4 g02240(new_n4589, new_n4588_1, new_n4548);
xnor_3 g02241(n243, new_n4589, new_n4542);
xor_3  g02242(new_n4591, n24786, n11302);
nor_4  g02243(new_n4592, n27120, n17090);
not_3  g02244(new_n4593, new_n4592);
nand_4 g02245(new_n4594, n23065, n6773);
nand_4 g02246(new_n4595_1, n27120, n17090);
not_3  g02247(new_n4596, new_n4595_1);
nor_4  g02248(new_n4597, new_n4596, new_n4592);
nand_4 g02249(new_n4598, new_n4597, new_n4594);
nand_4 g02250(new_n4599, new_n4598, new_n4593);
nor_4  g02251(new_n4600, new_n4599, new_n4591);
nand_4 g02252(new_n4601, new_n4599, new_n4591);
not_3  g02253(new_n4602, new_n4601);
nor_4  g02254(new_n4603, new_n4602, new_n4600);
xor_3  g02255(new_n4604, n20036, n1689);
not_3  g02256(new_n4605, n22274);
nor_4  g02257(new_n4606, new_n4605, n11192);
not_3  g02258(new_n4607, n11192);
nor_4  g02259(new_n4608, n22274, new_n4607);
not_3  g02260(new_n4609, n9380);
nand_4 g02261(new_n4610, n24129, new_n4609);
nor_4  g02262(new_n4611, new_n4610, new_n4608);
nor_4  g02263(new_n4612, new_n4611, new_n4606);
xnor_3 g02264(new_n4613, new_n4612, new_n4604);
not_3  g02265(new_n4614, new_n4613);
xnor_3 g02266(new_n4615, new_n4614, new_n4603);
not_3  g02267(new_n4616, new_n4594);
xnor_3 g02268(new_n4617, n27120, n17090);
xor_3  g02269(new_n4618, new_n4617, new_n4616);
not_3  g02270(new_n4619, new_n4610);
nor_4  g02271(new_n4620, new_n4608, new_n4606);
xnor_3 g02272(new_n4621, new_n4620, new_n4619);
not_3  g02273(new_n4622, new_n4621);
nor_4  g02274(new_n4623, new_n4622, new_n4618);
not_3  g02275(new_n4624_1, new_n4623);
xor_3  g02276(new_n4625, n23065, n6773);
xor_3  g02277(new_n4626, n24129, n9380);
nand_4 g02278(new_n4627, new_n4626, new_n4625);
not_3  g02279(new_n4628, new_n4627);
xor_3  g02280(new_n4629, new_n4617, new_n4594);
nor_4  g02281(new_n4630, new_n4621, new_n4629);
nor_4  g02282(new_n4631, new_n4630, new_n4623);
nand_4 g02283(new_n4632, new_n4631, new_n4628);
nand_4 g02284(new_n4633, new_n4632, new_n4624_1);
nor_4  g02285(new_n4634, new_n4633, new_n4615);
not_3  g02286(new_n4635, new_n4615);
xnor_3 g02287(new_n4636, new_n4621, new_n4629);
nor_4  g02288(new_n4637, new_n4636, new_n4627);
nor_4  g02289(new_n4638, new_n4637, new_n4623);
nor_4  g02290(new_n4639, new_n4638, new_n4635);
nor_4  g02291(new_n4640, new_n4639, new_n4634);
xor_3  g02292(new_n4641, n5330, n919);
nor_4  g02293(new_n4642, n25316, n7657);
not_3  g02294(new_n4643, new_n4642);
nand_4 g02295(new_n4644, n25926, n20385);
xor_3  g02296(new_n4645, n25316, n7657);
nand_4 g02297(new_n4646_1, new_n4645, new_n4644);
nand_4 g02298(new_n4647, new_n4646_1, new_n4643);
nor_4  g02299(new_n4648, new_n4647, new_n4641);
nand_4 g02300(new_n4649, new_n4647, new_n4641);
not_3  g02301(new_n4650, new_n4649);
nor_4  g02302(new_n4651, new_n4650, new_n4648);
xnor_3 g02303(new_n4652, new_n4651, new_n4640);
not_3  g02304(new_n4653, new_n4652);
xnor_3 g02305(new_n4654, new_n4636, new_n4627);
xnor_3 g02306(new_n4655, new_n4645, new_n4644);
nand_4 g02307(new_n4656, new_n4655, new_n4654);
xor_3  g02308(new_n4657, n25926, n20385);
not_3  g02309(new_n4658, new_n4657);
nor_4  g02310(new_n4659, new_n4626, new_n4625);
nor_4  g02311(new_n4660, new_n4659, new_n4628);
nor_4  g02312(new_n4661, new_n4660, new_n4658);
not_3  g02313(new_n4662, new_n4656);
nor_4  g02314(new_n4663, new_n4655, new_n4654);
nor_4  g02315(new_n4664, new_n4663, new_n4662);
nand_4 g02316(new_n4665_1, new_n4664, new_n4661);
nand_4 g02317(new_n4666, new_n4665_1, new_n4656);
xor_3  g02318(n248, new_n4666, new_n4653);
not_3  g02319(new_n4668, n19905);
not_3  g02320(new_n4669, n14684);
nor_4  g02321(new_n4670, n24732, n6631);
nand_4 g02322(new_n4671, new_n4670, new_n4669);
nor_4  g02323(new_n4672, new_n4671, n17035);
xor_3  g02324(new_n4673, new_n4672, new_n4668);
xnor_3 g02325(new_n4674_1, new_n4673, new_n4075);
not_3  g02326(new_n4675, new_n4674_1);
not_3  g02327(new_n4676, n25797);
not_3  g02328(new_n4677, new_n4671);
xor_3  g02329(new_n4678, new_n4677, n17035);
nor_4  g02330(new_n4679, new_n4678, new_n4676);
not_3  g02331(new_n4680, n17035);
xor_3  g02332(new_n4681, new_n4677, new_n4680);
xnor_3 g02333(new_n4682, new_n4681, n25797);
xor_3  g02334(new_n4683, new_n4670, n14684);
nand_4 g02335(new_n4684, new_n4683, new_n4076);
xor_3  g02336(new_n4685, new_n4670, new_n4669);
xnor_3 g02337(new_n4686, new_n4685, new_n4076);
not_3  g02338(new_n4687, n13319);
not_3  g02339(new_n4688, n6631);
xor_3  g02340(new_n4689, n24732, new_n4688);
nand_4 g02341(new_n4690, new_n4689, new_n4687);
nand_4 g02342(new_n4691, n25435, n24732);
xnor_3 g02343(new_n4692, new_n4689, n13319);
nand_4 g02344(new_n4693_1, new_n4692, new_n4691);
nand_4 g02345(new_n4694, new_n4693_1, new_n4690);
nand_4 g02346(new_n4695, new_n4694, new_n4686);
nand_4 g02347(new_n4696, new_n4695, new_n4684);
nor_4  g02348(new_n4697, new_n4696, new_n4682);
nor_4  g02349(new_n4698, new_n4697, new_n4679);
xnor_3 g02350(new_n4699, new_n4698, new_n4675);
not_3  g02351(new_n4700, n19514);
nor_4  g02352(new_n4701, n14148, n1152);
nand_4 g02353(new_n4702, new_n4701, new_n3005);
nor_4  g02354(new_n4703, new_n4702, n18558);
nand_4 g02355(new_n4704, new_n4703, new_n3000);
not_3  g02356(new_n4705, new_n4704);
nor_4  g02357(new_n4706, new_n4703, new_n3000);
nor_4  g02358(new_n4707, new_n4706, new_n4705);
not_3  g02359(new_n4708, new_n4707);
nor_4  g02360(new_n4709, new_n4708, new_n4700);
nor_4  g02361(new_n4710, new_n4707, n19514);
nor_4  g02362(new_n4711, new_n4710, new_n4709);
nand_4 g02363(new_n4712, new_n4702, n18558);
not_3  g02364(new_n4713, new_n4712);
nor_4  g02365(new_n4714, new_n4713, new_n4703);
not_3  g02366(new_n4715, new_n4714);
nor_4  g02367(new_n4716, new_n4715, new_n4197);
not_3  g02368(new_n4717, new_n4716);
nor_4  g02369(new_n4718, new_n4714, n10053);
nor_4  g02370(new_n4719, new_n4718, new_n4716);
not_3  g02371(new_n4720, new_n4702);
nor_4  g02372(new_n4721, new_n4701, new_n3005);
nor_4  g02373(new_n4722_1, new_n4721, new_n4720);
not_3  g02374(new_n4723, new_n4722_1);
nor_4  g02375(new_n4724, new_n4723, new_n4199);
not_3  g02376(new_n4725, new_n4724);
nor_4  g02377(new_n4726, new_n4722_1, n8399);
nor_4  g02378(new_n4727, new_n4726, new_n4724);
nand_4 g02379(new_n4728, n14148, n1152);
not_3  g02380(new_n4729, new_n4728);
nor_4  g02381(new_n4730, new_n4729, new_n4701);
not_3  g02382(new_n4731_1, new_n4730);
nor_4  g02383(new_n4732, new_n4731_1, new_n4203);
not_3  g02384(new_n4733, new_n4732);
nand_4 g02385(new_n4734, n26979, n1152);
not_3  g02386(new_n4735, new_n4734);
xnor_3 g02387(new_n4736, new_n4730, new_n4203);
nand_4 g02388(new_n4737, new_n4736, new_n4735);
nand_4 g02389(new_n4738, new_n4737, new_n4733);
nand_4 g02390(new_n4739, new_n4738, new_n4727);
nand_4 g02391(new_n4740, new_n4739, new_n4725);
nand_4 g02392(new_n4741, new_n4740, new_n4719);
nand_4 g02393(new_n4742, new_n4741, new_n4717);
xnor_3 g02394(new_n4743, new_n4742, new_n4711);
not_3  g02395(new_n4744, n13668);
not_3  g02396(new_n4745_1, n26748);
nor_4  g02397(new_n4746, n10057, n8920);
nand_4 g02398(new_n4747_1, new_n4746, new_n4745_1);
nor_4  g02399(new_n4748, new_n4747_1, n21276);
xor_3  g02400(new_n4749, new_n4748, new_n4744);
xnor_3 g02401(new_n4750, new_n4749, new_n4238);
nand_4 g02402(new_n4751, new_n4747_1, n21276);
not_3  g02403(new_n4752, new_n4751);
nor_4  g02404(new_n4753, new_n4752, new_n4748);
nand_4 g02405(new_n4754, new_n4753, n1204);
xnor_3 g02406(new_n4755, new_n4753, new_n4246);
not_3  g02407(new_n4756, new_n4747_1);
nor_4  g02408(new_n4757, new_n4746, new_n4745_1);
nor_4  g02409(new_n4758, new_n4757, new_n4756);
not_3  g02410(new_n4759, new_n4758);
nor_4  g02411(new_n4760, new_n4759, new_n4220);
not_3  g02412(new_n4761, new_n4760);
nor_4  g02413(new_n4762, new_n4758, n19618);
nor_4  g02414(new_n4763, new_n4762, new_n4760);
not_3  g02415(new_n4764, new_n4746);
nand_4 g02416(new_n4765, n10057, n8920);
nand_4 g02417(new_n4766_1, new_n4765, new_n4764);
not_3  g02418(new_n4767, new_n4766_1);
nor_4  g02419(new_n4768, new_n4767, n22043);
nand_4 g02420(new_n4769, n12121, n8920);
not_3  g02421(new_n4770_1, new_n4769);
xnor_3 g02422(new_n4771, new_n4766_1, n22043);
not_3  g02423(new_n4772, new_n4771);
nor_4  g02424(new_n4773, new_n4772, new_n4770_1);
nor_4  g02425(new_n4774, new_n4773, new_n4768);
nand_4 g02426(new_n4775, new_n4774, new_n4763);
nand_4 g02427(new_n4776, new_n4775, new_n4761);
nand_4 g02428(new_n4777_1, new_n4776, new_n4755);
nand_4 g02429(new_n4778, new_n4777_1, new_n4754);
xnor_3 g02430(new_n4779, new_n4778, new_n4750);
nor_4  g02431(new_n4780, new_n4779, new_n4743);
not_3  g02432(new_n4781, new_n4743);
xnor_3 g02433(new_n4782, new_n4749, n626);
xnor_3 g02434(new_n4783, new_n4778, new_n4782);
nor_4  g02435(new_n4784, new_n4783, new_n4781);
nor_4  g02436(new_n4785_1, new_n4784, new_n4780);
xnor_3 g02437(new_n4786, new_n4740, new_n4719);
not_3  g02438(new_n4787, new_n4755);
xnor_3 g02439(new_n4788, new_n4776, new_n4787);
not_3  g02440(new_n4789, new_n4788);
nor_4  g02441(new_n4790, new_n4789, new_n4786);
not_3  g02442(new_n4791, new_n4790);
not_3  g02443(new_n4792, new_n4786);
nor_4  g02444(new_n4793, new_n4788, new_n4792);
nor_4  g02445(new_n4794, new_n4793, new_n4790);
xnor_3 g02446(new_n4795, new_n4774, new_n4763);
not_3  g02447(new_n4796, new_n4795);
xnor_3 g02448(new_n4797, new_n4736, new_n4735);
xnor_3 g02449(new_n4798, new_n4771, new_n4769);
not_3  g02450(new_n4799, new_n4798);
nor_4  g02451(new_n4800, new_n4799, new_n4797);
not_3  g02452(new_n4801, new_n4800);
xnor_3 g02453(new_n4802, n12121, n8920);
xnor_3 g02454(new_n4803, n26979, n1152);
nor_4  g02455(new_n4804_1, new_n4803, new_n4802);
not_3  g02456(new_n4805, new_n4797);
nor_4  g02457(new_n4806, new_n4798, new_n4805);
nor_4  g02458(new_n4807, new_n4806, new_n4800);
nand_4 g02459(new_n4808, new_n4807, new_n4804_1);
nand_4 g02460(new_n4809, new_n4808, new_n4801);
nand_4 g02461(new_n4810_1, new_n4809, new_n4796);
xnor_3 g02462(new_n4811, new_n4738, new_n4727);
not_3  g02463(new_n4812_1, new_n4811);
xnor_3 g02464(new_n4813, new_n4809, new_n4795);
nand_4 g02465(new_n4814_1, new_n4813, new_n4812_1);
nand_4 g02466(new_n4815, new_n4814_1, new_n4810_1);
nand_4 g02467(new_n4816, new_n4815, new_n4794);
nand_4 g02468(new_n4817, new_n4816, new_n4791);
xnor_3 g02469(new_n4818, new_n4817, new_n4785_1);
nor_4  g02470(new_n4819, new_n4818, new_n4699);
nand_4 g02471(new_n4820, new_n4818, new_n4699);
not_3  g02472(new_n4821, new_n4820);
nor_4  g02473(new_n4822, new_n4821, new_n4819);
xnor_3 g02474(new_n4823, new_n4696, new_n4682);
xnor_3 g02475(new_n4824, new_n4815, new_n4794);
nor_4  g02476(new_n4825, new_n4824, new_n4823);
xnor_3 g02477(new_n4826, new_n4824, new_n4823);
xnor_3 g02478(new_n4827, new_n4813, new_n4812_1);
xnor_3 g02479(new_n4828, new_n4694, new_n4686);
not_3  g02480(new_n4829, new_n4828);
nor_4  g02481(new_n4830, new_n4829, new_n4827);
xnor_3 g02482(new_n4831, new_n4829, new_n4827);
xnor_3 g02483(new_n4832, new_n4807, new_n4804_1);
not_3  g02484(new_n4833, new_n4832);
nor_4  g02485(new_n4834, new_n4833, new_n4692);
not_3  g02486(new_n4835, new_n4834);
not_3  g02487(new_n4836, new_n4692);
xor_3  g02488(new_n4837, new_n4836, new_n4691);
nand_4 g02489(new_n4838, new_n4837, new_n4833);
xor_3  g02490(new_n4839, n25435, n24732);
not_3  g02491(new_n4840, new_n4839);
not_3  g02492(new_n4841, new_n4803);
xor_3  g02493(new_n4842, new_n4841, new_n4802);
nor_4  g02494(new_n4843, new_n4842, new_n4840);
not_3  g02495(new_n4844, new_n4843);
nand_4 g02496(new_n4845, new_n4844, new_n4838);
nand_4 g02497(new_n4846, new_n4845, new_n4835);
nor_4  g02498(new_n4847, new_n4846, new_n4831);
nor_4  g02499(new_n4848, new_n4847, new_n4830);
nor_4  g02500(new_n4849, new_n4848, new_n4826);
nor_4  g02501(new_n4850_1, new_n4849, new_n4825);
not_3  g02502(new_n4851, new_n4850_1);
xor_3  g02503(n266, new_n4851, new_n4822);
not_3  g02504(new_n4853, n21839);
nor_4  g02505(new_n4854, n22270, new_n4853);
xor_3  g02506(new_n4855, n22270, new_n4853);
not_3  g02507(new_n4856, new_n4855);
not_3  g02508(new_n4857, n27089);
nor_4  g02509(new_n4858_1, new_n4857, n8806);
xor_3  g02510(new_n4859, new_n4857, n8806);
not_3  g02511(new_n4860, n2479);
nand_4 g02512(new_n4861, n11841, new_n4860);
xor_3  g02513(new_n4862, n11841, new_n4860);
nand_4 g02514(new_n4863, n10710, new_n2780);
xor_3  g02515(new_n4864, n10710, new_n2780);
not_3  g02516(new_n4865, n6596);
nand_4 g02517(new_n4866, n20929, new_n4865);
xor_3  g02518(new_n4867, n20929, new_n4865);
not_3  g02519(new_n4868, n8006);
nor_4  g02520(new_n4869, n15289, new_n4868);
not_3  g02521(new_n4870, new_n4869);
xor_3  g02522(new_n4871, n15289, new_n4868);
not_3  g02523(new_n4872, n25074);
nor_4  g02524(new_n4873, new_n4872, n6556);
not_3  g02525(new_n4874, new_n4873);
not_3  g02526(new_n4875, n6556);
xor_3  g02527(new_n4876, n25074, new_n4875);
not_3  g02528(new_n4877, n22871);
nor_4  g02529(new_n4878, new_n4877, n16396);
not_3  g02530(new_n4879, n16396);
nor_4  g02531(new_n4880, n22871, new_n4879);
not_3  g02532(new_n4881, n14275);
nor_4  g02533(new_n4882, new_n4881, n9399);
not_3  g02534(new_n4883, n9399);
nor_4  g02535(new_n4884, n14275, new_n4883);
not_3  g02536(new_n4885, n2088);
nand_4 g02537(new_n4886, n25023, new_n4885);
nor_4  g02538(new_n4887, new_n4886, new_n4884);
nor_4  g02539(new_n4888, new_n4887, new_n4882);
nor_4  g02540(new_n4889, new_n4888, new_n4880);
nor_4  g02541(new_n4890, new_n4889, new_n4878);
nand_4 g02542(new_n4891_1, new_n4890, new_n4876);
nand_4 g02543(new_n4892, new_n4891_1, new_n4874);
nand_4 g02544(new_n4893, new_n4892, new_n4871);
nand_4 g02545(new_n4894, new_n4893, new_n4870);
nand_4 g02546(new_n4895, new_n4894, new_n4867);
nand_4 g02547(new_n4896, new_n4895, new_n4866);
nand_4 g02548(new_n4897, new_n4896, new_n4864);
nand_4 g02549(new_n4898, new_n4897, new_n4863);
nand_4 g02550(new_n4899, new_n4898, new_n4862);
nand_4 g02551(new_n4900, new_n4899, new_n4861);
nand_4 g02552(new_n4901, new_n4900, new_n4859);
not_3  g02553(new_n4902, new_n4901);
nor_4  g02554(new_n4903, new_n4902, new_n4858_1);
nor_4  g02555(new_n4904, new_n4903, new_n4856);
nor_4  g02556(new_n4905, new_n4904, new_n4854);
not_3  g02557(new_n4906, new_n4905);
not_3  g02558(new_n4907, n23272);
xor_3  g02559(new_n4908, new_n4903, new_n4856);
not_3  g02560(new_n4909, new_n4908);
nand_4 g02561(new_n4910, new_n4909, new_n4907);
xnor_3 g02562(new_n4911, new_n4908, new_n4907);
xnor_3 g02563(new_n4912, new_n4900, new_n4859);
not_3  g02564(new_n4913_1, new_n4912);
nor_4  g02565(new_n4914, new_n4913_1, n11481);
not_3  g02566(new_n4915, new_n4914);
xor_3  g02567(new_n4916, new_n4913_1, n11481);
xnor_3 g02568(new_n4917, new_n4898, new_n4862);
not_3  g02569(new_n4918, new_n4917);
nor_4  g02570(new_n4919, new_n4918, n16439);
not_3  g02571(new_n4920, new_n4919);
xor_3  g02572(new_n4921, new_n4918, n16439);
not_3  g02573(new_n4922, n15241);
xnor_3 g02574(new_n4923, new_n4896, new_n4864);
nand_4 g02575(new_n4924, new_n4923, new_n4922);
xnor_3 g02576(new_n4925_1, new_n4923, n15241);
xnor_3 g02577(new_n4926, new_n4894, new_n4867);
not_3  g02578(new_n4927, new_n4926);
nor_4  g02579(new_n4928, new_n4927, n7678);
not_3  g02580(new_n4929, new_n4928);
xor_3  g02581(new_n4930, new_n4927, n7678);
not_3  g02582(new_n4931, new_n4871);
xnor_3 g02583(new_n4932, new_n4892, new_n4931);
nor_4  g02584(new_n4933, new_n4932, n3785);
not_3  g02585(new_n4934, new_n4933);
not_3  g02586(new_n4935, n3785);
not_3  g02587(new_n4936, new_n4932);
nor_4  g02588(new_n4937, new_n4936, new_n4935);
nor_4  g02589(new_n4938, new_n4937, new_n4933);
not_3  g02590(new_n4939_1, new_n4890);
xnor_3 g02591(new_n4940, new_n4939_1, new_n4876);
nor_4  g02592(new_n4941, new_n4940, n20250);
not_3  g02593(new_n4942, new_n4941);
not_3  g02594(new_n4943, n20250);
not_3  g02595(new_n4944, new_n4940);
nor_4  g02596(new_n4945, new_n4944, new_n4943);
nor_4  g02597(new_n4946, new_n4945, new_n4941);
not_3  g02598(new_n4947_1, n5822);
nor_4  g02599(new_n4948, new_n4880, new_n4878);
xnor_3 g02600(new_n4949, new_n4948, new_n4888);
nor_4  g02601(new_n4950, new_n4949, new_n4947_1);
not_3  g02602(new_n4951, new_n4949);
nor_4  g02603(new_n4952_1, new_n4951, n5822);
nor_4  g02604(new_n4953, new_n4884, new_n4882);
xnor_3 g02605(new_n4954, new_n4953, new_n4886);
not_3  g02606(new_n4955, new_n4954);
nor_4  g02607(new_n4956, new_n4955, n26443);
not_3  g02608(new_n4957_1, n1681);
xor_3  g02609(new_n4958, n25023, n2088);
not_3  g02610(new_n4959, new_n4958);
nor_4  g02611(new_n4960, new_n4959, new_n4957_1);
not_3  g02612(new_n4961, n26443);
nor_4  g02613(new_n4962, new_n4954, new_n4961);
nor_4  g02614(new_n4963, new_n4962, new_n4956);
not_3  g02615(new_n4964_1, new_n4963);
nor_4  g02616(new_n4965, new_n4964_1, new_n4960);
nor_4  g02617(new_n4966_1, new_n4965, new_n4956);
not_3  g02618(new_n4967_1, new_n4966_1);
nor_4  g02619(new_n4968, new_n4967_1, new_n4952_1);
nor_4  g02620(new_n4969, new_n4968, new_n4950);
nand_4 g02621(new_n4970, new_n4969, new_n4946);
nand_4 g02622(new_n4971, new_n4970, new_n4942);
nand_4 g02623(new_n4972_1, new_n4971, new_n4938);
nand_4 g02624(new_n4973, new_n4972_1, new_n4934);
nand_4 g02625(new_n4974, new_n4973, new_n4930);
nand_4 g02626(new_n4975, new_n4974, new_n4929);
nand_4 g02627(new_n4976, new_n4975, new_n4925_1);
nand_4 g02628(new_n4977, new_n4976, new_n4924);
nand_4 g02629(new_n4978, new_n4977, new_n4921);
nand_4 g02630(new_n4979, new_n4978, new_n4920);
nand_4 g02631(new_n4980, new_n4979, new_n4916);
nand_4 g02632(new_n4981, new_n4980, new_n4915);
nand_4 g02633(new_n4982, new_n4981, new_n4911);
nand_4 g02634(new_n4983, new_n4982, new_n4910);
nor_4  g02635(new_n4984, new_n4983, new_n4906);
not_3  g02636(new_n4985, n18105);
not_3  g02637(new_n4986, n6785);
nor_4  g02638(new_n4987, n24032, n22843);
nand_4 g02639(new_n4988, new_n4987, new_n4986);
nor_4  g02640(new_n4989, new_n4988, n24879);
not_3  g02641(new_n4990, new_n4989);
nor_4  g02642(new_n4991, new_n4990, n268);
not_3  g02643(new_n4992, new_n4991);
nor_4  g02644(new_n4993, new_n4992, n12587);
not_3  g02645(new_n4994, new_n4993);
nor_4  g02646(new_n4995, new_n4994, n25381);
not_3  g02647(new_n4996, new_n4995);
nor_4  g02648(new_n4997, new_n4996, n16376);
not_3  g02649(new_n4998, new_n4997);
nor_4  g02650(new_n4999, new_n4998, n24196);
xor_3  g02651(new_n5000, new_n4999, new_n4985);
not_3  g02652(new_n5001, new_n5000);
nand_4 g02653(new_n5002, new_n4342, new_n2619_1);
nor_4  g02654(new_n5003, new_n5002, n25168);
not_3  g02655(new_n5004, new_n5003);
xor_3  g02656(new_n5005, new_n5004, n1999);
nor_4  g02657(new_n5006, new_n5005, n25475);
not_3  g02658(new_n5007, n25475);
not_3  g02659(new_n5008, new_n5005);
xor_3  g02660(new_n5009, new_n5008, new_n5007);
not_3  g02661(new_n5010, new_n5009);
xor_3  g02662(new_n5011_1, new_n5002, n25168);
nor_4  g02663(new_n5012, new_n5011_1, n23849);
not_3  g02664(new_n5013, n23849);
not_3  g02665(new_n5014, new_n5011_1);
xor_3  g02666(new_n5015, new_n5014, new_n5013);
not_3  g02667(new_n5016, new_n5015);
xor_3  g02668(new_n5017, new_n4342, new_n2619_1);
nor_4  g02669(new_n5018, new_n5017, n12446);
not_3  g02670(new_n5019, new_n4348);
nand_4 g02671(new_n5020_1, new_n4387, new_n4349);
nand_4 g02672(new_n5021, new_n5020_1, new_n5019);
not_3  g02673(new_n5022, n12446);
xnor_3 g02674(new_n5023, new_n5017, new_n5022);
nand_4 g02675(new_n5024_1, new_n5023, new_n5021);
not_3  g02676(new_n5025_1, new_n5024_1);
nor_4  g02677(new_n5026_1, new_n5025_1, new_n5018);
nor_4  g02678(new_n5027, new_n5026_1, new_n5016);
nor_4  g02679(new_n5028, new_n5027, new_n5012);
nor_4  g02680(new_n5029, new_n5028, new_n5010);
nor_4  g02681(new_n5030, new_n5029, new_n5006);
nor_4  g02682(new_n5031_1, new_n5004, n1999);
xor_3  g02683(new_n5032, new_n5031_1, n9396);
not_3  g02684(new_n5033, new_n5032);
nor_4  g02685(new_n5034, new_n5033, n18880);
not_3  g02686(new_n5035, n18880);
nor_4  g02687(new_n5036, new_n5032, new_n5035);
nor_4  g02688(new_n5037, new_n5036, new_n5034);
xnor_3 g02689(new_n5038, new_n5037, new_n5030);
nor_4  g02690(new_n5039, new_n5038, new_n5001);
not_3  g02691(new_n5040, new_n4999);
nor_4  g02692(new_n5041, new_n5040, n18105);
not_3  g02693(new_n5042, new_n5041);
not_3  g02694(new_n5043, new_n5038);
nor_4  g02695(new_n5044, new_n5043, new_n5000);
nor_4  g02696(new_n5045, new_n5044, new_n5039);
not_3  g02697(new_n5046_1, n24196);
xor_3  g02698(new_n5047, new_n4997, new_n5046_1);
xnor_3 g02699(new_n5048, new_n5028, new_n5010);
nor_4  g02700(new_n5049, new_n5048, new_n5047);
not_3  g02701(new_n5050, new_n5047);
xnor_3 g02702(new_n5051, new_n5028, new_n5009);
nor_4  g02703(new_n5052, new_n5051, new_n5050);
nor_4  g02704(new_n5053, new_n5052, new_n5049);
not_3  g02705(new_n5054, new_n5053);
not_3  g02706(new_n5055, n16376);
xor_3  g02707(new_n5056, new_n4995, new_n5055);
xnor_3 g02708(new_n5057, new_n5026_1, new_n5016);
nor_4  g02709(new_n5058, new_n5057, new_n5056);
xnor_3 g02710(new_n5059, new_n5057, new_n5056);
not_3  g02711(new_n5060_1, n25381);
xor_3  g02712(new_n5061, new_n4993, new_n5060_1);
xnor_3 g02713(new_n5062_1, new_n5023, new_n5021);
nor_4  g02714(new_n5063, new_n5062_1, new_n5061);
not_3  g02715(new_n5064_1, new_n5063);
not_3  g02716(new_n5065, new_n5061);
nor_4  g02717(new_n5066, new_n5023, new_n5021);
nor_4  g02718(new_n5067, new_n5066, new_n5025_1);
nor_4  g02719(new_n5068, new_n5067, new_n5065);
nor_4  g02720(new_n5069, new_n5068, new_n5063);
not_3  g02721(new_n5070, n12587);
xor_3  g02722(new_n5071, new_n4991, new_n5070);
nor_4  g02723(new_n5072, new_n5071, new_n4388);
not_3  g02724(new_n5073, new_n5072);
not_3  g02725(new_n5074, new_n5071);
nor_4  g02726(new_n5075, new_n5074, new_n4389);
nor_4  g02727(new_n5076, new_n5075, new_n5072);
not_3  g02728(new_n5077_1, n268);
xor_3  g02729(new_n5078, new_n4989, new_n5077_1);
nor_4  g02730(new_n5079, new_n5078, new_n4393);
not_3  g02731(new_n5080, new_n5079);
not_3  g02732(new_n5081, new_n4396);
not_3  g02733(new_n5082_1, n24879);
xor_3  g02734(new_n5083, new_n4988, new_n5082_1);
nand_4 g02735(new_n5084, new_n5083, new_n5081);
xnor_3 g02736(new_n5085, new_n5083, new_n4396);
xor_3  g02737(new_n5086, new_n4987, n6785);
nor_4  g02738(new_n5087, new_n5086, new_n4403);
xnor_3 g02739(new_n5088, new_n5086, new_n4403);
not_3  g02740(new_n5089, n22843);
xor_3  g02741(new_n5090, n24032, new_n5089);
nand_4 g02742(new_n5091, new_n5090, new_n4410);
nand_4 g02743(new_n5092, new_n2605, n22843);
not_3  g02744(new_n5093, new_n5091);
nor_4  g02745(new_n5094, new_n5090, new_n4410);
nor_4  g02746(new_n5095, new_n5094, new_n5093);
nand_4 g02747(new_n5096, new_n5095, new_n5092);
nand_4 g02748(new_n5097, new_n5096, new_n5091);
nor_4  g02749(new_n5098_1, new_n5097, new_n5088);
nor_4  g02750(new_n5099, new_n5098_1, new_n5087);
nand_4 g02751(new_n5100, new_n5099, new_n5085);
nand_4 g02752(new_n5101_1, new_n5100, new_n5084);
not_3  g02753(new_n5102, new_n4393);
not_3  g02754(new_n5103, new_n5078);
nor_4  g02755(new_n5104, new_n5103, new_n5102);
nor_4  g02756(new_n5105, new_n5104, new_n5079);
nand_4 g02757(new_n5106, new_n5105, new_n5101_1);
nand_4 g02758(new_n5107, new_n5106, new_n5080);
nand_4 g02759(new_n5108, new_n5107, new_n5076);
nand_4 g02760(new_n5109, new_n5108, new_n5073);
nand_4 g02761(new_n5110, new_n5109, new_n5069);
nand_4 g02762(new_n5111, new_n5110, new_n5064_1);
not_3  g02763(new_n5112, new_n5111);
nor_4  g02764(new_n5113, new_n5112, new_n5059);
nor_4  g02765(new_n5114, new_n5113, new_n5058);
nor_4  g02766(new_n5115_1, new_n5114, new_n5054);
nor_4  g02767(new_n5116, new_n5115_1, new_n5049);
nand_4 g02768(new_n5117, new_n5116, new_n5045);
nand_4 g02769(new_n5118, new_n5117, new_n5042);
nor_4  g02770(new_n5119, new_n5118, new_n5039);
not_3  g02771(new_n5120_1, new_n5119);
not_3  g02772(new_n5121, new_n5031_1);
nor_4  g02773(new_n5122, new_n5121, n9396);
nor_4  g02774(new_n5123, new_n5036, new_n5030);
nor_4  g02775(new_n5124, new_n5123, new_n5034);
nor_4  g02776(new_n5125, new_n5124, new_n5122);
nor_4  g02777(new_n5126, new_n5125, new_n5120_1);
not_3  g02778(new_n5127, new_n5126);
nor_4  g02779(new_n5128_1, new_n5127, new_n4984);
not_3  g02780(new_n5129, new_n4984);
nor_4  g02781(new_n5130, new_n5126, new_n5129);
nor_4  g02782(new_n5131_1, new_n5130, new_n5128_1);
xnor_3 g02783(new_n5132, new_n4983, new_n4905);
not_3  g02784(new_n5133, new_n5125);
xnor_3 g02785(new_n5134, new_n5133, new_n5119);
nor_4  g02786(new_n5135, new_n5134, new_n5132);
not_3  g02787(new_n5136, new_n5132);
xnor_3 g02788(new_n5137, new_n5125, new_n5119);
xnor_3 g02789(new_n5138, new_n5137, new_n5136);
xnor_3 g02790(new_n5139, new_n5116, new_n5045);
not_3  g02791(new_n5140_1, new_n5139);
xnor_3 g02792(new_n5141, new_n4981, new_n4911);
nor_4  g02793(new_n5142, new_n5141, new_n5140_1);
not_3  g02794(new_n5143, new_n5141);
xnor_3 g02795(new_n5144, new_n5143, new_n5139);
xnor_3 g02796(new_n5145, new_n5114, new_n5054);
xnor_3 g02797(new_n5146, new_n4979, new_n4916);
nor_4  g02798(new_n5147, new_n5146, new_n5145);
not_3  g02799(new_n5148, new_n5146);
xnor_3 g02800(new_n5149, new_n5148, new_n5145);
not_3  g02801(new_n5150, new_n5149);
not_3  g02802(new_n5151, new_n5059);
nor_4  g02803(new_n5152, new_n5111, new_n5151);
nor_4  g02804(new_n5153, new_n5152, new_n5113);
not_3  g02805(new_n5154, new_n5153);
xnor_3 g02806(new_n5155, new_n4977, new_n4921);
nor_4  g02807(new_n5156, new_n5155, new_n5154);
xnor_3 g02808(new_n5157, new_n5155, new_n5153);
xnor_3 g02809(new_n5158_1, new_n5109, new_n5069);
not_3  g02810(new_n5159, new_n5158_1);
not_3  g02811(new_n5160, new_n4925_1);
xnor_3 g02812(new_n5161, new_n4975, new_n5160);
nand_4 g02813(new_n5162, new_n5161, new_n5159);
xnor_3 g02814(new_n5163, new_n5161, new_n5158_1);
xnor_3 g02815(new_n5164, new_n5107, new_n5076);
xnor_3 g02816(new_n5165, new_n4973, new_n4930);
nor_4  g02817(new_n5166, new_n5165, new_n5164);
not_3  g02818(new_n5167, new_n5166);
not_3  g02819(new_n5168_1, new_n5076);
xnor_3 g02820(new_n5169, new_n5107, new_n5168_1);
not_3  g02821(new_n5170, new_n5165);
nor_4  g02822(new_n5171, new_n5170, new_n5169);
nor_4  g02823(new_n5172, new_n5171, new_n5166);
xnor_3 g02824(new_n5173, new_n4971, new_n4938);
not_3  g02825(new_n5174, new_n5173);
not_3  g02826(new_n5175, new_n5105);
xnor_3 g02827(new_n5176, new_n5175, new_n5101_1);
nand_4 g02828(new_n5177, new_n5176, new_n5174);
xnor_3 g02829(new_n5178, new_n5176, new_n5173);
xnor_3 g02830(new_n5179, new_n5099, new_n5085);
not_3  g02831(new_n5180, new_n5179);
not_3  g02832(new_n5181, new_n4969);
xnor_3 g02833(new_n5182, new_n5181, new_n4946);
nand_4 g02834(new_n5183, new_n5182, new_n5180);
xnor_3 g02835(new_n5184_1, new_n5182, new_n5179);
xnor_3 g02836(new_n5185, new_n5097, new_n5088);
nor_4  g02837(new_n5186, new_n4952_1, new_n4950);
xnor_3 g02838(new_n5187, new_n5186, new_n4966_1);
nor_4  g02839(new_n5188, new_n5187, new_n5185);
xnor_3 g02840(new_n5189, new_n4964_1, new_n4960);
xnor_3 g02841(new_n5190, new_n5095, new_n5092);
nor_4  g02842(new_n5191, new_n5190, new_n5189);
not_3  g02843(new_n5192, new_n5191);
not_3  g02844(new_n5193, new_n5092);
nor_4  g02845(new_n5194, new_n2605, n22843);
nor_4  g02846(new_n5195, new_n5194, new_n5193);
not_3  g02847(new_n5196, new_n5195);
nor_4  g02848(new_n5197, new_n4958, n1681);
nor_4  g02849(new_n5198, new_n5197, new_n4960);
not_3  g02850(new_n5199, new_n5198);
nor_4  g02851(new_n5200, new_n5199, new_n5196);
not_3  g02852(new_n5201, new_n5200);
not_3  g02853(new_n5202, new_n5189);
not_3  g02854(new_n5203, new_n5190);
nor_4  g02855(new_n5204, new_n5203, new_n5202);
nor_4  g02856(new_n5205, new_n5204, new_n5191);
nand_4 g02857(new_n5206, new_n5205, new_n5201);
nand_4 g02858(new_n5207, new_n5206, new_n5192);
xnor_3 g02859(new_n5208, new_n5187, new_n5185);
nor_4  g02860(new_n5209, new_n5208, new_n5207);
nor_4  g02861(new_n5210, new_n5209, new_n5188);
nand_4 g02862(new_n5211_1, new_n5210, new_n5184_1);
nand_4 g02863(new_n5212, new_n5211_1, new_n5183);
nand_4 g02864(new_n5213_1, new_n5212, new_n5178);
nand_4 g02865(new_n5214, new_n5213_1, new_n5177);
nand_4 g02866(new_n5215, new_n5214, new_n5172);
nand_4 g02867(new_n5216, new_n5215, new_n5167);
nand_4 g02868(new_n5217, new_n5216, new_n5163);
nand_4 g02869(new_n5218, new_n5217, new_n5162);
nand_4 g02870(new_n5219, new_n5218, new_n5157);
not_3  g02871(new_n5220, new_n5219);
nor_4  g02872(new_n5221, new_n5220, new_n5156);
nor_4  g02873(new_n5222, new_n5221, new_n5150);
nor_4  g02874(new_n5223, new_n5222, new_n5147);
nor_4  g02875(new_n5224, new_n5223, new_n5144);
nor_4  g02876(new_n5225, new_n5224, new_n5142);
nor_4  g02877(new_n5226_1, new_n5225, new_n5138);
nor_4  g02878(new_n5227, new_n5226_1, new_n5135);
xnor_3 g02879(n298, new_n5227, new_n5131_1);
not_3  g02880(new_n5229, n20604);
xor_3  g02881(new_n5230, n21735, new_n5229);
not_3  g02882(new_n5231, n24085);
nor_4  g02883(new_n5232, new_n5231, n16158);
not_3  g02884(new_n5233, new_n5232);
not_3  g02885(new_n5234, n16158);
xor_3  g02886(new_n5235, n24085, new_n5234);
not_3  g02887(new_n5236, n14071);
nor_4  g02888(new_n5237, new_n5236, n5752);
not_3  g02889(new_n5238, new_n5237);
xor_3  g02890(new_n5239, n14071, n5752);
not_3  g02891(new_n5240, n18171);
nor_4  g02892(new_n5241, new_n5240, n1738);
not_3  g02893(new_n5242, n1738);
nor_4  g02894(new_n5243, n18171, new_n5242);
not_3  g02895(new_n5244, n25073);
nor_4  g02896(new_n5245, new_n5244, n12152);
not_3  g02897(new_n5246, n12152);
nor_4  g02898(new_n5247, n25073, new_n5246);
not_3  g02899(new_n5248, n19107);
nand_4 g02900(new_n5249, n22309, new_n5248);
nor_4  g02901(new_n5250, new_n5249, new_n5247);
nor_4  g02902(new_n5251, new_n5250, new_n5245);
nor_4  g02903(new_n5252, new_n5251, new_n5243);
nor_4  g02904(new_n5253, new_n5252, new_n5241);
not_3  g02905(new_n5254, new_n5253);
nor_4  g02906(new_n5255_1, new_n5254, new_n5239);
not_3  g02907(new_n5256_1, new_n5255_1);
nand_4 g02908(new_n5257, new_n5256_1, new_n5238);
nand_4 g02909(new_n5258, new_n5257, new_n5235);
nand_4 g02910(new_n5259, new_n5258, new_n5233);
xor_3  g02911(new_n5260, new_n5259, new_n5230);
xor_3  g02912(new_n5261, new_n3693, n1525);
not_3  g02913(new_n5262, n16988);
nor_4  g02914(new_n5263, new_n5262, n14510);
not_3  g02915(new_n5264, new_n5263);
xor_3  g02916(new_n5265_1, n16988, new_n3700);
not_3  g02917(new_n5266, n21779);
nor_4  g02918(new_n5267, new_n5266, n13263);
not_3  g02919(new_n5268, new_n5267);
xor_3  g02920(new_n5269, n21779, new_n3725_1);
nor_4  g02921(new_n5270, new_n3712, n5376);
not_3  g02922(new_n5271, n5376);
nor_4  g02923(new_n5272, n20455, new_n5271);
nor_4  g02924(new_n5273_1, n5128, new_n3716);
not_3  g02925(new_n5274_1, n5128);
nor_4  g02926(new_n5275, new_n5274_1, n1639);
not_3  g02927(new_n5276, n23120);
nand_4 g02928(new_n5277, new_n5276, n16968);
nor_4  g02929(new_n5278, new_n5277, new_n5275);
nor_4  g02930(new_n5279, new_n5278, new_n5273_1);
nor_4  g02931(new_n5280, new_n5279, new_n5272);
nor_4  g02932(new_n5281, new_n5280, new_n5270);
nand_4 g02933(new_n5282, new_n5281, new_n5269);
nand_4 g02934(new_n5283, new_n5282, new_n5268);
nand_4 g02935(new_n5284, new_n5283, new_n5265_1);
nand_4 g02936(new_n5285, new_n5284, new_n5264);
xnor_3 g02937(new_n5286, new_n5285, new_n5261);
not_3  g02938(new_n5287, n4272);
xor_3  g02939(new_n5288, n12626, new_n5287);
not_3  g02940(new_n5289, n24319);
nor_4  g02941(new_n5290, new_n5289, n6971);
not_3  g02942(new_n5291, new_n5290);
not_3  g02943(new_n5292, n6971);
xor_3  g02944(new_n5293, n24319, new_n5292);
not_3  g02945(new_n5294, n7460);
nor_4  g02946(new_n5295, n22068, new_n5294);
not_3  g02947(new_n5296, new_n5295);
xor_3  g02948(new_n5297, n22068, new_n5294);
not_3  g02949(new_n5298, n9460);
nor_4  g02950(new_n5299, new_n5298, n196);
not_3  g02951(new_n5300_1, n196);
nor_4  g02952(new_n5301, n9460, new_n5300_1);
not_3  g02953(new_n5302_1, n14954);
nor_4  g02954(new_n5303, new_n5302_1, n11749);
not_3  g02955(new_n5304, n11749);
nor_4  g02956(new_n5305, n14954, new_n5304);
not_3  g02957(new_n5306, n13424);
nand_4 g02958(new_n5307, n23831, new_n5306);
nor_4  g02959(new_n5308, new_n5307, new_n5305);
nor_4  g02960(new_n5309, new_n5308, new_n5303);
nor_4  g02961(new_n5310, new_n5309, new_n5301);
nor_4  g02962(new_n5311, new_n5310, new_n5299);
nand_4 g02963(new_n5312, new_n5311, new_n5297);
nand_4 g02964(new_n5313, new_n5312, new_n5296);
nand_4 g02965(new_n5314, new_n5313, new_n5293);
nand_4 g02966(new_n5315, new_n5314, new_n5291);
not_3  g02967(new_n5316, new_n5315);
xnor_3 g02968(new_n5317, new_n5316, new_n5288);
not_3  g02969(new_n5318, new_n5317);
nor_4  g02970(new_n5319, new_n5318, new_n5286);
not_3  g02971(new_n5320, new_n5286);
nor_4  g02972(new_n5321, new_n5317, new_n5320);
nor_4  g02973(new_n5322, new_n5321, new_n5319);
xnor_3 g02974(new_n5323, new_n5283, new_n5265_1);
xnor_3 g02975(new_n5324, new_n5313, new_n5293);
nor_4  g02976(new_n5325_1, new_n5324, new_n5323);
not_3  g02977(new_n5326, new_n5325_1);
not_3  g02978(new_n5327, new_n5323);
not_3  g02979(new_n5328, new_n5324);
nor_4  g02980(new_n5329, new_n5328, new_n5327);
nor_4  g02981(new_n5330_1, new_n5329, new_n5325_1);
not_3  g02982(new_n5331, new_n5281);
xnor_3 g02983(new_n5332, new_n5331, new_n5269);
xor_3  g02984(new_n5333, n22068, n7460);
not_3  g02985(new_n5334, new_n5311);
xnor_3 g02986(new_n5335, new_n5334, new_n5333);
not_3  g02987(new_n5336, new_n5335);
nor_4  g02988(new_n5337_1, new_n5336, new_n5332);
xnor_3 g02989(new_n5338, new_n5336, new_n5332);
nor_4  g02990(new_n5339, new_n5272, new_n5270);
not_3  g02991(new_n5340, new_n5339);
xnor_3 g02992(new_n5341, new_n5340, new_n5279);
nor_4  g02993(new_n5342, new_n5301, new_n5299);
xnor_3 g02994(new_n5343, new_n5342, new_n5309);
not_3  g02995(new_n5344, new_n5343);
nor_4  g02996(new_n5345, new_n5344, new_n5341);
not_3  g02997(new_n5346, new_n5341);
nor_4  g02998(new_n5347, new_n5343, new_n5346);
nor_4  g02999(new_n5348, new_n5347, new_n5345);
not_3  g03000(new_n5349, new_n5348);
nor_4  g03001(new_n5350, new_n5275, new_n5273_1);
xnor_3 g03002(new_n5351_1, new_n5350, new_n5277);
nor_4  g03003(new_n5352, new_n5305, new_n5303);
xnor_3 g03004(new_n5353_1, new_n5352, new_n5307);
nor_4  g03005(new_n5354, new_n5353_1, new_n5351_1);
not_3  g03006(new_n5355, new_n5354);
not_3  g03007(new_n5356, n16968);
xor_3  g03008(new_n5357, n23120, new_n5356);
xor_3  g03009(new_n5358, n23831, new_n5306);
nor_4  g03010(new_n5359, new_n5358, new_n5357);
not_3  g03011(new_n5360, new_n5351_1);
not_3  g03012(new_n5361, new_n5353_1);
nor_4  g03013(new_n5362, new_n5361, new_n5360);
nor_4  g03014(new_n5363, new_n5362, new_n5354);
nand_4 g03015(new_n5364, new_n5363, new_n5359);
nand_4 g03016(new_n5365, new_n5364, new_n5355);
nor_4  g03017(new_n5366, new_n5365, new_n5349);
nor_4  g03018(new_n5367, new_n5366, new_n5345);
nor_4  g03019(new_n5368, new_n5367, new_n5338);
nor_4  g03020(new_n5369, new_n5368, new_n5337_1);
nand_4 g03021(new_n5370, new_n5369, new_n5330_1);
nand_4 g03022(new_n5371, new_n5370, new_n5326);
xnor_3 g03023(new_n5372, new_n5371, new_n5322);
not_3  g03024(new_n5373, new_n5372);
xnor_3 g03025(new_n5374, new_n5373, new_n5260);
xor_3  g03026(new_n5375, new_n5257, new_n5235);
not_3  g03027(new_n5376_1, new_n5330_1);
xnor_3 g03028(new_n5377, new_n5369, new_n5376_1);
nor_4  g03029(new_n5378, new_n5377, new_n5375);
not_3  g03030(new_n5379, new_n5378);
not_3  g03031(new_n5380, new_n5375);
xnor_3 g03032(new_n5381, new_n5369, new_n5330_1);
nor_4  g03033(new_n5382, new_n5381, new_n5380);
nor_4  g03034(new_n5383, new_n5382, new_n5378);
xnor_3 g03035(new_n5384, new_n5367, new_n5338);
xor_3  g03036(new_n5385, new_n5254, new_n5239);
nor_4  g03037(new_n5386_1, new_n5385, new_n5384);
not_3  g03038(new_n5387, new_n5386_1);
xnor_3 g03039(new_n5388, new_n5365, new_n5348);
not_3  g03040(new_n5389, new_n5388);
nor_4  g03041(new_n5390, new_n5243, new_n5241);
xor_3  g03042(new_n5391, new_n5390, new_n5251);
nor_4  g03043(new_n5392, new_n5391, new_n5389);
xnor_3 g03044(new_n5393, new_n5391, new_n5389);
xor_3  g03045(new_n5394, n22309, new_n5248);
xor_3  g03046(new_n5395, n23120, n16968);
xor_3  g03047(new_n5396, n23831, n13424);
xnor_3 g03048(new_n5397, new_n5396, new_n5395);
nor_4  g03049(new_n5398, new_n5397, new_n5394);
nor_4  g03050(new_n5399_1, new_n5247, new_n5245);
xor_3  g03051(new_n5400_1, new_n5399_1, new_n5249);
nor_4  g03052(new_n5401, new_n5400_1, new_n5398);
not_3  g03053(new_n5402, new_n5363);
xnor_3 g03054(new_n5403_1, new_n5402, new_n5359);
xnor_3 g03055(new_n5404, new_n5400_1, new_n5398);
nor_4  g03056(new_n5405, new_n5404, new_n5403_1);
nor_4  g03057(new_n5406, new_n5405, new_n5401);
nor_4  g03058(new_n5407, new_n5406, new_n5393);
nor_4  g03059(new_n5408, new_n5407, new_n5392);
not_3  g03060(new_n5409, new_n5408);
not_3  g03061(new_n5410, new_n5384);
xnor_3 g03062(new_n5411, new_n5385, new_n5410);
nand_4 g03063(new_n5412, new_n5411, new_n5409);
nand_4 g03064(new_n5413, new_n5412, new_n5387);
nand_4 g03065(new_n5414, new_n5413, new_n5383);
nand_4 g03066(new_n5415, new_n5414, new_n5379);
xor_3  g03067(n317, new_n5415, new_n5374);
nor_4  g03068(new_n5417, n9934, n3506);
xor_3  g03069(new_n5418, n9934, n3506);
not_3  g03070(new_n5419, new_n5418);
nor_4  g03071(new_n5420, n18496, n14899);
xor_3  g03072(new_n5421, n18496, n14899);
not_3  g03073(new_n5422, new_n5421);
nor_4  g03074(new_n5423, n26224, n18444);
xor_3  g03075(new_n5424, n26224, n18444);
not_3  g03076(new_n5425, new_n5424);
not_3  g03077(new_n5426, n19327);
nand_4 g03078(new_n5427, new_n3834, new_n5426);
xor_3  g03079(new_n5428, n24638, n19327);
nor_4  g03080(new_n5429, n22597, n21674);
not_3  g03081(new_n5430_1, new_n5429);
xor_3  g03082(new_n5431, n22597, n21674);
nor_4  g03083(new_n5432, n26107, n17251);
not_3  g03084(new_n5433, new_n5432);
xor_3  g03085(new_n5434, n26107, n17251);
nor_4  g03086(new_n5435, n14790, n342);
not_3  g03087(new_n5436, new_n5435);
xor_3  g03088(new_n5437, n14790, n342);
nor_4  g03089(new_n5438_1, n26553, n10096);
not_3  g03090(new_n5439_1, new_n5438_1);
xor_3  g03091(new_n5440, n26553, n10096);
nand_4 g03092(new_n5441, new_n3854, new_n4116);
nand_4 g03093(new_n5442, n9246, n7876);
xor_3  g03094(new_n5443_1, n16994, n4964);
nand_4 g03095(new_n5444, new_n5443_1, new_n5442);
nand_4 g03096(new_n5445, new_n5444, new_n5441);
nand_4 g03097(new_n5446, new_n5445, new_n5440);
nand_4 g03098(new_n5447, new_n5446, new_n5439_1);
nand_4 g03099(new_n5448, new_n5447, new_n5437);
nand_4 g03100(new_n5449, new_n5448, new_n5436);
nand_4 g03101(new_n5450, new_n5449, new_n5434);
nand_4 g03102(new_n5451_1, new_n5450, new_n5433);
nand_4 g03103(new_n5452, new_n5451_1, new_n5431);
nand_4 g03104(new_n5453, new_n5452, new_n5430_1);
nand_4 g03105(new_n5454, new_n5453, new_n5428);
nand_4 g03106(new_n5455, new_n5454, new_n5427);
not_3  g03107(new_n5456, new_n5455);
nor_4  g03108(new_n5457, new_n5456, new_n5425);
nor_4  g03109(new_n5458, new_n5457, new_n5423);
nor_4  g03110(new_n5459, new_n5458, new_n5422);
nor_4  g03111(new_n5460, new_n5459, new_n5420);
nor_4  g03112(new_n5461, new_n5460, new_n5419);
nor_4  g03113(new_n5462, new_n5461, new_n5417);
not_3  g03114(new_n5463, new_n5462);
xor_3  g03115(new_n5464, n9554, n2979);
nor_4  g03116(new_n5465, n26408, n647);
xor_3  g03117(new_n5466, n26408, n647);
not_3  g03118(new_n5467, new_n5466);
nor_4  g03119(new_n5468, n20409, n18227);
xor_3  g03120(new_n5469, n20409, n18227);
not_3  g03121(new_n5470, new_n5469);
not_3  g03122(new_n5471, n7377);
not_3  g03123(new_n5472_1, n25749);
nand_4 g03124(new_n5473, new_n5472_1, new_n5471);
xor_3  g03125(new_n5474, n25749, n7377);
nor_4  g03126(new_n5475, n11630, n3161);
not_3  g03127(new_n5476, new_n5475);
xor_3  g03128(new_n5477, n11630, n3161);
nor_4  g03129(new_n5478, n13453, n9003);
not_3  g03130(new_n5479, new_n5478);
xor_3  g03131(new_n5480, n13453, n9003);
nor_4  g03132(new_n5481, n7421, n4957);
not_3  g03133(new_n5482, new_n5481);
nand_4 g03134(new_n5483, n7421, n4957);
not_3  g03135(new_n5484, new_n5483);
nor_4  g03136(new_n5485_1, new_n5484, new_n5481);
nor_4  g03137(new_n5486, n19680, n7524);
not_3  g03138(new_n5487, new_n5486);
nand_4 g03139(new_n5488, n19680, n7524);
not_3  g03140(new_n5489, new_n5488);
nor_4  g03141(new_n5490, new_n5489, new_n5486);
nor_4  g03142(new_n5491, n15743, n2809);
not_3  g03143(new_n5492, new_n5491);
nand_4 g03144(new_n5493, n20658, n15508);
nand_4 g03145(new_n5494, n15743, n2809);
not_3  g03146(new_n5495, new_n5494);
nor_4  g03147(new_n5496, new_n5495, new_n5491);
nand_4 g03148(new_n5497, new_n5496, new_n5493);
nand_4 g03149(new_n5498, new_n5497, new_n5492);
nand_4 g03150(new_n5499, new_n5498, new_n5490);
nand_4 g03151(new_n5500, new_n5499, new_n5487);
nand_4 g03152(new_n5501, new_n5500, new_n5485_1);
nand_4 g03153(new_n5502, new_n5501, new_n5482);
nand_4 g03154(new_n5503, new_n5502, new_n5480);
nand_4 g03155(new_n5504, new_n5503, new_n5479);
nand_4 g03156(new_n5505, new_n5504, new_n5477);
nand_4 g03157(new_n5506, new_n5505, new_n5476);
nand_4 g03158(new_n5507, new_n5506, new_n5474);
nand_4 g03159(new_n5508, new_n5507, new_n5473);
not_3  g03160(new_n5509, new_n5508);
nor_4  g03161(new_n5510, new_n5509, new_n5470);
nor_4  g03162(new_n5511, new_n5510, new_n5468);
nor_4  g03163(new_n5512, new_n5511, new_n5467);
nor_4  g03164(new_n5513, new_n5512, new_n5465);
not_3  g03165(new_n5514, new_n5513);
nor_4  g03166(new_n5515, new_n5514, new_n5464);
not_3  g03167(new_n5516, new_n5464);
nor_4  g03168(new_n5517_1, new_n5513, new_n5516);
nor_4  g03169(new_n5518, new_n5517_1, new_n5515);
not_3  g03170(new_n5519, new_n5518);
nand_4 g03171(new_n5520, new_n5519, n9259);
xnor_3 g03172(new_n5521_1, new_n5518, n9259);
xnor_3 g03173(new_n5522, new_n5511, new_n5467);
nand_4 g03174(new_n5523, new_n5522, n21489);
not_3  g03175(new_n5524_1, new_n5523);
nor_4  g03176(new_n5525, new_n5522, n21489);
nor_4  g03177(new_n5526, new_n5525, new_n5524_1);
xnor_3 g03178(new_n5527, new_n5508, new_n5469);
nor_4  g03179(new_n5528, new_n5527, n20213);
not_3  g03180(new_n5529, n20213);
xnor_3 g03181(new_n5530, new_n5527, new_n5529);
xnor_3 g03182(new_n5531, new_n5506, new_n5474);
not_3  g03183(new_n5532_1, new_n5531);
nand_4 g03184(new_n5533, new_n5532_1, new_n3913);
xnor_3 g03185(new_n5534, new_n5531, new_n3913);
not_3  g03186(new_n5535, n7670);
xnor_3 g03187(new_n5536, new_n5504, new_n5477);
not_3  g03188(new_n5537, new_n5536);
nand_4 g03189(new_n5538, new_n5537, new_n5535);
xnor_3 g03190(new_n5539, new_n5536, new_n5535);
not_3  g03191(new_n5540, n9598);
xnor_3 g03192(new_n5541, new_n5502, new_n5480);
not_3  g03193(new_n5542, new_n5541);
nand_4 g03194(new_n5543, new_n5542, new_n5540);
xnor_3 g03195(new_n5544, new_n5541, new_n5540);
not_3  g03196(new_n5545, n22290);
not_3  g03197(new_n5546, new_n5485_1);
xnor_3 g03198(new_n5547, new_n5500, new_n5546);
nand_4 g03199(new_n5548, new_n5547, new_n5545);
xnor_3 g03200(new_n5549, new_n5547, n22290);
not_3  g03201(new_n5550, new_n5493);
xnor_3 g03202(new_n5551, n15743, n2809);
nor_4  g03203(new_n5552, new_n5551, new_n5550);
nor_4  g03204(new_n5553, new_n5552, new_n5491);
xnor_3 g03205(new_n5554, new_n5553, new_n5490);
nand_4 g03206(new_n5555, new_n5554, new_n3943);
xnor_3 g03207(new_n5556, new_n5551, new_n5550);
nor_4  g03208(new_n5557, new_n5556, n25565);
not_3  g03209(new_n5558, new_n5557);
not_3  g03210(new_n5559, n21993);
xnor_3 g03211(new_n5560, n20658, n15508);
nor_4  g03212(new_n5561, new_n5560, new_n5559);
not_3  g03213(new_n5562, new_n5561);
not_3  g03214(new_n5563, n25565);
xnor_3 g03215(new_n5564_1, new_n5551, new_n5493);
nor_4  g03216(new_n5565, new_n5564_1, new_n5563);
nor_4  g03217(new_n5566, new_n5565, new_n5557);
nand_4 g03218(new_n5567, new_n5566, new_n5562);
nand_4 g03219(new_n5568, new_n5567, new_n5558);
not_3  g03220(new_n5569, new_n5555);
nor_4  g03221(new_n5570, new_n5554, new_n3943);
nor_4  g03222(new_n5571, new_n5570, new_n5569);
nand_4 g03223(new_n5572, new_n5571, new_n5568);
nand_4 g03224(new_n5573, new_n5572, new_n5555);
nand_4 g03225(new_n5574, new_n5573, new_n5549);
nand_4 g03226(new_n5575, new_n5574, new_n5548);
nand_4 g03227(new_n5576, new_n5575, new_n5544);
nand_4 g03228(new_n5577, new_n5576, new_n5543);
nand_4 g03229(new_n5578, new_n5577, new_n5539);
nand_4 g03230(new_n5579_1, new_n5578, new_n5538);
nand_4 g03231(new_n5580, new_n5579_1, new_n5534);
nand_4 g03232(new_n5581, new_n5580, new_n5533);
nand_4 g03233(new_n5582, new_n5581, new_n5530);
not_3  g03234(new_n5583, new_n5582);
nor_4  g03235(new_n5584, new_n5583, new_n5528);
nand_4 g03236(new_n5585, new_n5584, new_n5526);
nand_4 g03237(new_n5586, new_n5585, new_n5523);
nand_4 g03238(new_n5587, new_n5586, new_n5521_1);
nand_4 g03239(new_n5588, new_n5587, new_n5520);
nor_4  g03240(new_n5589, n9554, n2979);
nor_4  g03241(new_n5590, new_n5517_1, new_n5589);
nor_4  g03242(new_n5591, new_n5590, new_n5588);
nand_4 g03243(new_n5592, new_n5590, new_n5588);
not_3  g03244(new_n5593_1, new_n5592);
nor_4  g03245(new_n5594, new_n5593_1, new_n5591);
not_3  g03246(new_n5595, new_n5594);
xnor_3 g03247(new_n5596, new_n5586, new_n5521_1);
nor_4  g03248(new_n5597, new_n5596, n3740);
xnor_3 g03249(new_n5598, new_n5596, n3740);
xnor_3 g03250(new_n5599, new_n5584, new_n5526);
nor_4  g03251(new_n5600, new_n5599, n2858);
xnor_3 g03252(new_n5601, new_n5599, n2858);
not_3  g03253(new_n5602, n2659);
xnor_3 g03254(new_n5603_1, new_n5581, new_n5530);
nand_4 g03255(new_n5604, new_n5603_1, new_n5602);
xnor_3 g03256(new_n5605_1, new_n5603_1, n2659);
not_3  g03257(new_n5606, n24327);
xnor_3 g03258(new_n5607, new_n5579_1, new_n5534);
nand_4 g03259(new_n5608, new_n5607, new_n5606);
xnor_3 g03260(new_n5609_1, new_n5607, n24327);
not_3  g03261(new_n5610, n22198);
xnor_3 g03262(new_n5611, new_n5577, new_n5539);
nand_4 g03263(new_n5612, new_n5611, new_n5610);
xnor_3 g03264(new_n5613, new_n5611, n22198);
xnor_3 g03265(new_n5614, new_n5575, new_n5544);
not_3  g03266(new_n5615, new_n5614);
nor_4  g03267(new_n5616, new_n5615, n20826);
not_3  g03268(new_n5617, new_n5616);
not_3  g03269(new_n5618, n7305);
xnor_3 g03270(new_n5619, new_n5573, new_n5549);
nand_4 g03271(new_n5620, new_n5619, new_n5618);
xnor_3 g03272(new_n5621, new_n5571, new_n5568);
not_3  g03273(new_n5622, new_n5621);
nor_4  g03274(new_n5623, new_n5622, n25872);
not_3  g03275(new_n5624, new_n5623);
not_3  g03276(new_n5625, n25872);
nor_4  g03277(new_n5626, new_n5621, new_n5625);
nor_4  g03278(new_n5627, new_n5626, new_n5623);
not_3  g03279(new_n5628, n20259);
xnor_3 g03280(new_n5629, new_n5566, new_n5562);
nor_4  g03281(new_n5630, new_n5629, new_n5628);
xor_3  g03282(new_n5631, new_n5560, n21993);
nor_4  g03283(new_n5632, new_n5631, n3925);
xnor_3 g03284(new_n5633, new_n5629, new_n5628);
nor_4  g03285(new_n5634_1, new_n5633, new_n5632);
nor_4  g03286(new_n5635, new_n5634_1, new_n5630);
nand_4 g03287(new_n5636, new_n5635, new_n5627);
nand_4 g03288(new_n5637, new_n5636, new_n5624);
xnor_3 g03289(new_n5638, new_n5619, n7305);
nand_4 g03290(new_n5639, new_n5638, new_n5637);
nand_4 g03291(new_n5640, new_n5639, new_n5620);
not_3  g03292(new_n5641, n20826);
nor_4  g03293(new_n5642, new_n5614, new_n5641);
nor_4  g03294(new_n5643_1, new_n5642, new_n5616);
nand_4 g03295(new_n5644, new_n5643_1, new_n5640);
nand_4 g03296(new_n5645, new_n5644, new_n5617);
nand_4 g03297(new_n5646, new_n5645, new_n5613);
nand_4 g03298(new_n5647, new_n5646, new_n5612);
nand_4 g03299(new_n5648, new_n5647, new_n5609_1);
nand_4 g03300(new_n5649, new_n5648, new_n5608);
nand_4 g03301(new_n5650, new_n5649, new_n5605_1);
nand_4 g03302(new_n5651, new_n5650, new_n5604);
not_3  g03303(new_n5652, new_n5651);
nor_4  g03304(new_n5653, new_n5652, new_n5601);
nor_4  g03305(new_n5654, new_n5653, new_n5600);
nor_4  g03306(new_n5655, new_n5654, new_n5598);
nor_4  g03307(new_n5656, new_n5655, new_n5597);
xnor_3 g03308(new_n5657, new_n5656, new_n5595);
xnor_3 g03309(new_n5658, new_n5657, new_n5463);
xor_3  g03310(new_n5659, new_n5460, new_n5419);
not_3  g03311(new_n5660, new_n5659);
xnor_3 g03312(new_n5661, new_n5654, new_n5598);
nor_4  g03313(new_n5662, new_n5661, new_n5660);
not_3  g03314(new_n5663, new_n5662);
xnor_3 g03315(new_n5664, new_n5661, new_n5659);
xor_3  g03316(new_n5665, new_n5458, new_n5422);
not_3  g03317(new_n5666, new_n5665);
not_3  g03318(new_n5667, new_n5601);
xnor_3 g03319(new_n5668, new_n5651, new_n5667);
nor_4  g03320(new_n5669, new_n5668, new_n5666);
not_3  g03321(new_n5670, new_n5669);
xnor_3 g03322(new_n5671, new_n5668, new_n5665);
xor_3  g03323(new_n5672, new_n5456, new_n5425);
not_3  g03324(new_n5673, new_n5605_1);
xnor_3 g03325(new_n5674, new_n5649, new_n5673);
nand_4 g03326(new_n5675, new_n5674, new_n5672);
not_3  g03327(new_n5676, new_n5672);
xnor_3 g03328(new_n5677, new_n5674, new_n5676);
not_3  g03329(new_n5678, new_n5453);
xor_3  g03330(new_n5679, new_n5678, new_n5428);
not_3  g03331(new_n5680_1, new_n5679);
not_3  g03332(new_n5681, new_n5609_1);
xnor_3 g03333(new_n5682, new_n5647, new_n5681);
nand_4 g03334(new_n5683, new_n5682, new_n5680_1);
xnor_3 g03335(new_n5684, new_n5682, new_n5679);
not_3  g03336(new_n5685, new_n5451_1);
xor_3  g03337(new_n5686, new_n5685, new_n5431);
not_3  g03338(new_n5687_1, new_n5686);
not_3  g03339(new_n5688, new_n5613);
xnor_3 g03340(new_n5689, new_n5645, new_n5688);
nand_4 g03341(new_n5690, new_n5689, new_n5687_1);
xnor_3 g03342(new_n5691, new_n5689, new_n5686);
not_3  g03343(new_n5692, new_n5449);
xor_3  g03344(new_n5693, new_n5692, new_n5434);
not_3  g03345(new_n5694, new_n5693);
not_3  g03346(new_n5695, new_n5643_1);
xnor_3 g03347(new_n5696_1, new_n5695, new_n5640);
nand_4 g03348(new_n5697, new_n5696_1, new_n5694);
xnor_3 g03349(new_n5698, new_n5696_1, new_n5693);
not_3  g03350(new_n5699, new_n5448);
nor_4  g03351(new_n5700_1, new_n5447, new_n5437);
nor_4  g03352(new_n5701, new_n5700_1, new_n5699);
not_3  g03353(new_n5702, new_n5638);
xnor_3 g03354(new_n5703, new_n5702, new_n5637);
nand_4 g03355(new_n5704_1, new_n5703, new_n5701);
not_3  g03356(new_n5705, new_n5704_1);
nor_4  g03357(new_n5706, new_n5703, new_n5701);
nor_4  g03358(new_n5707, new_n5706, new_n5705);
not_3  g03359(new_n5708, new_n5627);
xnor_3 g03360(new_n5709, new_n5635, new_n5708);
not_3  g03361(new_n5710, new_n5440);
not_3  g03362(new_n5711, new_n5445);
xor_3  g03363(new_n5712, new_n5711, new_n5710);
nand_4 g03364(new_n5713, new_n5712, new_n5709);
not_3  g03365(new_n5714, new_n5713);
nor_4  g03366(new_n5715, new_n5712, new_n5709);
nor_4  g03367(new_n5716, new_n5715, new_n5714);
not_3  g03368(new_n5717, n3925);
xnor_3 g03369(new_n5718, new_n5631, new_n5717);
xor_3  g03370(new_n5719, n9246, n7876);
not_3  g03371(new_n5720, new_n5719);
nor_4  g03372(new_n5721, new_n5720, new_n5718);
nand_4 g03373(new_n5722, new_n5721, new_n5443_1);
not_3  g03374(new_n5723, new_n5722);
xnor_3 g03375(new_n5724, new_n5633, new_n5632);
not_3  g03376(new_n5725, new_n5721);
not_3  g03377(new_n5726, new_n5443_1);
xor_3  g03378(new_n5727, new_n5726, new_n5442);
not_3  g03379(new_n5728, new_n5727);
nand_4 g03380(new_n5729, new_n5728, new_n5725);
nand_4 g03381(new_n5730, new_n5729, new_n5722);
nor_4  g03382(new_n5731, new_n5730, new_n5724);
nor_4  g03383(new_n5732_1, new_n5731, new_n5723);
nand_4 g03384(new_n5733, new_n5732_1, new_n5716);
nand_4 g03385(new_n5734, new_n5733, new_n5713);
nand_4 g03386(new_n5735, new_n5734, new_n5707);
nand_4 g03387(new_n5736, new_n5735, new_n5704_1);
nand_4 g03388(new_n5737, new_n5736, new_n5698);
nand_4 g03389(new_n5738, new_n5737, new_n5697);
nand_4 g03390(new_n5739, new_n5738, new_n5691);
nand_4 g03391(new_n5740, new_n5739, new_n5690);
nand_4 g03392(new_n5741, new_n5740, new_n5684);
nand_4 g03393(new_n5742_1, new_n5741, new_n5683);
nand_4 g03394(new_n5743, new_n5742_1, new_n5677);
nand_4 g03395(new_n5744, new_n5743, new_n5675);
nand_4 g03396(new_n5745, new_n5744, new_n5671);
nand_4 g03397(new_n5746, new_n5745, new_n5670);
nand_4 g03398(new_n5747, new_n5746, new_n5664);
nand_4 g03399(new_n5748, new_n5747, new_n5663);
nor_4  g03400(new_n5749, new_n5748, new_n5658);
nor_4  g03401(new_n5750, new_n5657, new_n5463);
not_3  g03402(new_n5751, new_n5657);
nor_4  g03403(new_n5752_1, new_n5751, new_n5462);
nor_4  g03404(new_n5753, new_n5752_1, new_n5750);
not_3  g03405(new_n5754, new_n5748);
nor_4  g03406(new_n5755, new_n5754, new_n5753);
nor_4  g03407(n332, new_n5755, new_n5749);
not_3  g03408(new_n5757, n8381);
nor_4  g03409(new_n5758, n18295, n16223);
nand_4 g03410(new_n5759, n18295, n16223);
not_3  g03411(new_n5760, new_n5759);
nor_4  g03412(new_n5761, new_n5760, new_n5758);
nor_4  g03413(new_n5762, n19494, n6502);
nand_4 g03414(new_n5763, n15780, n2387);
not_3  g03415(new_n5764, new_n5763);
xnor_3 g03416(new_n5765_1, n19494, n6502);
nor_4  g03417(new_n5766, new_n5765_1, new_n5764);
nor_4  g03418(new_n5767, new_n5766, new_n5762);
not_3  g03419(new_n5768, new_n5767);
nor_4  g03420(new_n5769, new_n5768, new_n5761);
not_3  g03421(new_n5770, new_n5761);
nor_4  g03422(new_n5771, new_n5767, new_n5770);
nor_4  g03423(new_n5772, new_n5771, new_n5769);
not_3  g03424(new_n5773, new_n5772);
nand_4 g03425(new_n5774, new_n5773, new_n5757);
not_3  g03426(new_n5775, new_n5774);
nor_4  g03427(new_n5776_1, new_n5773, new_n5757);
nor_4  g03428(new_n5777, new_n5776_1, new_n5775);
not_3  g03429(new_n5778, n20235);
xnor_3 g03430(new_n5779, n15780, n2387);
nor_4  g03431(new_n5780, new_n5779, n12495);
nand_4 g03432(new_n5781, new_n5780, new_n5778);
not_3  g03433(new_n5782_1, new_n5781);
nor_4  g03434(new_n5783, new_n5780, new_n5778);
nor_4  g03435(new_n5784, new_n5783, new_n5782_1);
not_3  g03436(new_n5785, new_n5784);
not_3  g03437(new_n5786, new_n5765_1);
nor_4  g03438(new_n5787, new_n5786, new_n5763);
nor_4  g03439(new_n5788, new_n5787, new_n5766);
nor_4  g03440(new_n5789, new_n5788, new_n5785);
nor_4  g03441(new_n5790, new_n5789, new_n5782_1);
not_3  g03442(new_n5791, new_n5790);
xnor_3 g03443(new_n5792, new_n5791, new_n5777);
not_3  g03444(new_n5793, n16502);
nor_4  g03445(new_n5794, n21654, new_n5793);
not_3  g03446(new_n5795, n23842);
nor_4  g03447(new_n5796, n25471, new_n5795);
nor_4  g03448(new_n5797, new_n3291, n23842);
nor_4  g03449(new_n5798, new_n5797, new_n5796);
xnor_3 g03450(new_n5799, new_n5798, new_n5794);
nand_4 g03451(new_n5800, new_n5799, n23146);
not_3  g03452(new_n5801, new_n5800);
not_3  g03453(new_n5802, n17968);
not_3  g03454(new_n5803, n21654);
nor_4  g03455(new_n5804, new_n5803, n16502);
nor_4  g03456(new_n5805, new_n5804, new_n5794);
nor_4  g03457(new_n5806, new_n5805, new_n5802);
not_3  g03458(new_n5807, new_n5806);
not_3  g03459(new_n5808, n23146);
nor_4  g03460(new_n5809, new_n5799, new_n5808);
not_3  g03461(new_n5810, new_n5794);
xnor_3 g03462(new_n5811, new_n5798, new_n5810);
nor_4  g03463(new_n5812, new_n5811, n23146);
nor_4  g03464(new_n5813, new_n5812, new_n5809);
nor_4  g03465(new_n5814, new_n5813, new_n5807);
nor_4  g03466(new_n5815, new_n5814, new_n5801);
not_3  g03467(new_n5816, n15053);
nor_4  g03468(new_n5817, new_n5816, n3828);
not_3  g03469(new_n5818, n3828);
nor_4  g03470(new_n5819, n15053, new_n5818);
nor_4  g03471(new_n5820, new_n5819, new_n5817);
not_3  g03472(new_n5821, new_n5820);
not_3  g03473(new_n5822_1, new_n5797);
nand_4 g03474(new_n5823, new_n5798, new_n5794);
nand_4 g03475(new_n5824, new_n5823, new_n5822_1);
not_3  g03476(new_n5825, new_n5824);
nor_4  g03477(new_n5826, new_n5825, new_n5821);
nor_4  g03478(new_n5827, new_n5824, new_n5820);
nor_4  g03479(new_n5828, new_n5827, new_n5826);
nor_4  g03480(new_n5829, new_n5828, n11184);
not_3  g03481(new_n5830, n11184);
xnor_3 g03482(new_n5831, new_n5824, new_n5820);
nor_4  g03483(new_n5832, new_n5831, new_n5830);
nor_4  g03484(new_n5833_1, new_n5832, new_n5829);
xnor_3 g03485(new_n5834_1, new_n5833_1, new_n5815);
not_3  g03486(new_n5835, new_n5834_1);
nor_4  g03487(new_n5836, new_n5835, new_n5792);
not_3  g03488(new_n5837, new_n5792);
nor_4  g03489(new_n5838, new_n5834_1, new_n5837);
nor_4  g03490(new_n5839, new_n5838, new_n5836);
not_3  g03491(new_n5840_1, new_n5839);
not_3  g03492(new_n5841_1, new_n5813);
nor_4  g03493(new_n5842_1, new_n5841_1, new_n5806);
nor_4  g03494(new_n5843, new_n5842_1, new_n5814);
not_3  g03495(new_n5844, new_n5843);
not_3  g03496(new_n5845, new_n5788);
nor_4  g03497(new_n5846, new_n5845, new_n5784);
nor_4  g03498(new_n5847, new_n5846, new_n5789);
nand_4 g03499(new_n5848, new_n5847, new_n5844);
xor_3  g03500(new_n5849, new_n5779, n12495);
not_3  g03501(new_n5850_1, new_n5849);
xor_3  g03502(new_n5851, new_n5805, new_n5802);
nand_4 g03503(new_n5852, new_n5851, new_n5850_1);
not_3  g03504(new_n5853, new_n5848);
nor_4  g03505(new_n5854, new_n5847, new_n5844);
nor_4  g03506(new_n5855, new_n5854, new_n5853);
nand_4 g03507(new_n5856, new_n5855, new_n5852);
nand_4 g03508(new_n5857, new_n5856, new_n5848);
xor_3  g03509(n357, new_n5857, new_n5840_1);
nand_4 g03510(new_n5859, n22309, n9251);
not_3  g03511(new_n5860, new_n5859);
nor_4  g03512(new_n5861, n22309, n9251);
nor_4  g03513(new_n5862, new_n5861, new_n5860);
nor_4  g03514(new_n5863, n25073, n20138);
not_3  g03515(new_n5864, new_n5863);
nand_4 g03516(new_n5865, n25073, n20138);
nand_4 g03517(new_n5866, new_n5865, new_n5864);
xnor_3 g03518(new_n5867, new_n5866, new_n5860);
nor_4  g03519(new_n5868, new_n5867, new_n5862);
not_3  g03520(new_n5869, new_n5868);
nor_4  g03521(new_n5870, n18171, n6385);
nand_4 g03522(new_n5871, n18171, n6385);
not_3  g03523(new_n5872, new_n5871);
nor_4  g03524(new_n5873, new_n5872, new_n5870);
nor_4  g03525(new_n5874, new_n5866, new_n5860);
nor_4  g03526(new_n5875, new_n5874, new_n5863);
not_3  g03527(new_n5876, new_n5875);
nor_4  g03528(new_n5877, new_n5876, new_n5873);
not_3  g03529(new_n5878, new_n5873);
nor_4  g03530(new_n5879, new_n5875, new_n5878);
nor_4  g03531(new_n5880, new_n5879, new_n5877);
not_3  g03532(new_n5881, new_n5880);
nor_4  g03533(new_n5882_1, new_n5881, new_n5869);
not_3  g03534(new_n5883, new_n5882_1);
xor_3  g03535(new_n5884, n5752, n3136);
nor_4  g03536(new_n5885, new_n5879, new_n5870);
not_3  g03537(new_n5886, new_n5885);
xnor_3 g03538(new_n5887, new_n5886, new_n5884);
nor_4  g03539(new_n5888, new_n5887, new_n5883);
not_3  g03540(new_n5889, new_n5888);
xor_3  g03541(new_n5890, n16158, n9557);
nor_4  g03542(new_n5891, n5752, n3136);
not_3  g03543(new_n5892, new_n5891);
nand_4 g03544(new_n5893, new_n5886, new_n5884);
nand_4 g03545(new_n5894, new_n5893, new_n5892);
xnor_3 g03546(new_n5895, new_n5894, new_n5890);
nor_4  g03547(new_n5896, new_n5895, new_n5889);
xor_3  g03548(new_n5897, n25643, n20604);
nor_4  g03549(new_n5898, n16158, n9557);
not_3  g03550(new_n5899, new_n5898);
nand_4 g03551(new_n5900, new_n5894, new_n5890);
nand_4 g03552(new_n5901, new_n5900, new_n5899);
nor_4  g03553(new_n5902, new_n5901, new_n5897);
nand_4 g03554(new_n5903_1, new_n5901, new_n5897);
not_3  g03555(new_n5904_1, new_n5903_1);
nor_4  g03556(new_n5905, new_n5904_1, new_n5902);
xnor_3 g03557(new_n5906, new_n5905, new_n5896);
xnor_3 g03558(new_n5907, new_n5906, new_n3410);
xnor_3 g03559(new_n5908, new_n5895, new_n5889);
nand_4 g03560(new_n5909, new_n5908, new_n3414);
xnor_3 g03561(new_n5910, new_n5908, new_n3413);
xnor_3 g03562(new_n5911_1, new_n5887, new_n5883);
nand_4 g03563(new_n5912, new_n5911_1, new_n3421);
xnor_3 g03564(new_n5913, new_n5911_1, new_n3420);
xnor_3 g03565(new_n5914, new_n5880, new_n5868);
not_3  g03566(new_n5915, new_n5914);
nor_4  g03567(new_n5916, new_n5915, new_n3427);
not_3  g03568(new_n5917, new_n5916);
not_3  g03569(new_n5918, new_n5862);
nor_4  g03570(new_n5919, new_n5918, new_n3435);
nor_4  g03571(new_n5920, new_n5919, new_n3443);
not_3  g03572(new_n5921, new_n5874);
nor_4  g03573(new_n5922, new_n5921, new_n5861);
nor_4  g03574(new_n5923, new_n5922, new_n5868);
not_3  g03575(new_n5924, new_n5919);
nor_4  g03576(new_n5925, new_n5924, new_n3441);
nor_4  g03577(new_n5926, new_n5925, new_n5920);
not_3  g03578(new_n5927, new_n5926);
nor_4  g03579(new_n5928, new_n5927, new_n5923);
nor_4  g03580(new_n5929, new_n5928, new_n5920);
not_3  g03581(new_n5930, new_n5929);
nor_4  g03582(new_n5931, new_n5914, new_n3428);
nor_4  g03583(new_n5932, new_n5931, new_n5916);
nand_4 g03584(new_n5933, new_n5932, new_n5930);
nand_4 g03585(new_n5934, new_n5933, new_n5917);
nand_4 g03586(new_n5935, new_n5934, new_n5913);
nand_4 g03587(new_n5936_1, new_n5935, new_n5912);
nand_4 g03588(new_n5937, new_n5936_1, new_n5910);
nand_4 g03589(new_n5938, new_n5937, new_n5909);
xnor_3 g03590(new_n5939, new_n5938, new_n5907);
xor_3  g03591(new_n5940, n5255, new_n3693);
not_3  g03592(new_n5941, n21649);
nor_4  g03593(new_n5942, new_n5941, n14510);
not_3  g03594(new_n5943_1, new_n5942);
xor_3  g03595(new_n5944, n21649, new_n3700);
not_3  g03596(new_n5945, n18274);
nor_4  g03597(new_n5946, new_n5945, n13263);
xor_3  g03598(new_n5947, n18274, n13263);
nor_4  g03599(new_n5948, new_n3712, n3828);
nor_4  g03600(new_n5949, n20455, new_n5818);
nor_4  g03601(new_n5950, n23842, new_n3716);
nor_4  g03602(new_n5951, new_n5795, n1639);
nor_4  g03603(new_n5952, n21654, new_n5356);
not_3  g03604(new_n5953, new_n5952);
nor_4  g03605(new_n5954, new_n5953, new_n5951);
nor_4  g03606(new_n5955, new_n5954, new_n5950);
nor_4  g03607(new_n5956, new_n5955, new_n5949);
nor_4  g03608(new_n5957, new_n5956, new_n5948);
not_3  g03609(new_n5958, new_n5957);
nor_4  g03610(new_n5959, new_n5958, new_n5947);
nor_4  g03611(new_n5960, new_n5959, new_n5946);
not_3  g03612(new_n5961, new_n5960);
nand_4 g03613(new_n5962, new_n5961, new_n5944);
nand_4 g03614(new_n5963, new_n5962, new_n5943_1);
xor_3  g03615(new_n5964_1, new_n5963, new_n5940);
xnor_3 g03616(new_n5965, new_n5964_1, new_n5939);
xor_3  g03617(new_n5966, new_n5961, new_n5944);
xnor_3 g03618(new_n5967, new_n5936_1, new_n5910);
nor_4  g03619(new_n5968, new_n5967, new_n5966);
not_3  g03620(new_n5969, new_n5968);
xnor_3 g03621(new_n5970, new_n5967, new_n5966);
not_3  g03622(new_n5971, new_n5970);
xnor_3 g03623(new_n5972, new_n5934, new_n5913);
xor_3  g03624(new_n5973, new_n5958, new_n5947);
nor_4  g03625(new_n5974, new_n5973, new_n5972);
not_3  g03626(new_n5975, new_n5974);
xnor_3 g03627(new_n5976, new_n5973, new_n5972);
xnor_3 g03628(new_n5977, new_n5932, new_n5930);
nor_4  g03629(new_n5978, new_n5949, new_n5948);
xor_3  g03630(new_n5979, new_n5978, new_n5955);
nor_4  g03631(new_n5980_1, new_n5979, new_n5977);
not_3  g03632(new_n5981, new_n5977);
xnor_3 g03633(new_n5982, new_n5979, new_n5981);
not_3  g03634(new_n5983, new_n5982);
xor_3  g03635(new_n5984, n21654, new_n5356);
xor_3  g03636(new_n5985, new_n5862, new_n3508);
not_3  g03637(new_n5986, new_n5985);
nor_4  g03638(new_n5987, new_n5986, new_n5984);
nor_4  g03639(new_n5988, new_n5951, new_n5950);
xor_3  g03640(new_n5989, new_n5988, new_n5953);
nor_4  g03641(new_n5990, new_n5989, new_n5987);
not_3  g03642(new_n5991, new_n5923);
nor_4  g03643(new_n5992, new_n5926, new_n5991);
nor_4  g03644(new_n5993, new_n5992, new_n5928);
not_3  g03645(new_n5994, new_n5993);
xnor_3 g03646(new_n5995, new_n5989, new_n5987);
nor_4  g03647(new_n5996, new_n5995, new_n5994);
nor_4  g03648(new_n5997, new_n5996, new_n5990);
nor_4  g03649(new_n5998, new_n5997, new_n5983);
nor_4  g03650(new_n5999, new_n5998, new_n5980_1);
nor_4  g03651(new_n6000, new_n5999, new_n5976);
not_3  g03652(new_n6001, new_n6000);
nand_4 g03653(new_n6002, new_n6001, new_n5975);
nand_4 g03654(new_n6003, new_n6002, new_n5971);
nand_4 g03655(new_n6004, new_n6003, new_n5969);
xor_3  g03656(n422, new_n6004, new_n5965);
not_3  g03657(new_n6006, n21471);
not_3  g03658(new_n6007, n14603);
nor_4  g03659(new_n6008, n23333, n20794);
nand_4 g03660(new_n6009, new_n6008, new_n6007);
nor_4  g03661(new_n6010, new_n6009, n18737);
nand_4 g03662(new_n6011, new_n6010, new_n6006);
nor_4  g03663(new_n6012_1, new_n6011, n25738);
nand_4 g03664(new_n6013, new_n6012_1, new_n3274);
nor_4  g03665(new_n6014, new_n6013, n3228);
not_3  g03666(new_n6015, new_n6014);
xor_3  g03667(new_n6016, new_n6015, n337);
xor_3  g03668(new_n6017, new_n6016, n6485);
not_3  g03669(new_n6018, new_n6017);
xor_3  g03670(new_n6019, new_n6013, n3228);
nor_4  g03671(new_n6020, new_n6019, n26036);
xor_3  g03672(new_n6021, new_n6019, new_n3394);
xor_3  g03673(new_n6022_1, new_n6012_1, new_n3274);
nor_4  g03674(new_n6023, new_n6022_1, n19770);
not_3  g03675(new_n6024, new_n6022_1);
xor_3  g03676(new_n6025, new_n6024, new_n3401);
not_3  g03677(new_n6026, new_n6025);
xor_3  g03678(new_n6027, new_n6011, n25738);
nor_4  g03679(new_n6028, new_n6027, n8782);
not_3  g03680(new_n6029, new_n6027);
xor_3  g03681(new_n6030, new_n6029, new_n3409);
not_3  g03682(new_n6031_1, new_n6030);
xor_3  g03683(new_n6032, new_n6010, new_n6006);
nor_4  g03684(new_n6033, new_n6032, n8678);
not_3  g03685(new_n6034, new_n6032);
xor_3  g03686(new_n6035, new_n6034, new_n3417);
xor_3  g03687(new_n6036, new_n6009, n18737);
not_3  g03688(new_n6037, new_n6036);
nand_4 g03689(new_n6038, new_n6037, new_n3424);
xor_3  g03690(new_n6039, new_n6008, new_n6007);
not_3  g03691(new_n6040, new_n6039);
nand_4 g03692(new_n6041, new_n6040, new_n3431);
xor_3  g03693(new_n6042, new_n6040, new_n3431);
xor_3  g03694(new_n6043, n23333, new_n3290);
nand_4 g03695(new_n6044_1, new_n6043, new_n3434);
nand_4 g03696(new_n6045, n23333, n11424);
xnor_3 g03697(new_n6046_1, new_n6043, n25336);
nand_4 g03698(new_n6047, new_n6046_1, new_n6045);
nand_4 g03699(new_n6048, new_n6047, new_n6044_1);
nand_4 g03700(new_n6049, new_n6048, new_n6042);
nand_4 g03701(new_n6050, new_n6049, new_n6041);
xor_3  g03702(new_n6051, new_n6037, new_n3424);
nand_4 g03703(new_n6052, new_n6051, new_n6050);
nand_4 g03704(new_n6053, new_n6052, new_n6038);
nand_4 g03705(new_n6054, new_n6053, new_n6035);
not_3  g03706(new_n6055, new_n6054);
nor_4  g03707(new_n6056, new_n6055, new_n6033);
nor_4  g03708(new_n6057, new_n6056, new_n6031_1);
nor_4  g03709(new_n6058, new_n6057, new_n6028);
nor_4  g03710(new_n6059, new_n6058, new_n6026);
nor_4  g03711(new_n6060, new_n6059, new_n6023);
nor_4  g03712(new_n6061, new_n6060, new_n6021);
nor_4  g03713(new_n6062, new_n6061, new_n6020);
xnor_3 g03714(new_n6063, new_n6062, new_n6018);
xor_3  g03715(new_n6064, n22379, n9967);
nor_4  g03716(new_n6065, n20946, n1662);
not_3  g03717(new_n6066, new_n6065);
xor_3  g03718(new_n6067, n20946, n1662);
nand_4 g03719(new_n6068, new_n2989, new_n3475);
xor_3  g03720(new_n6069, n12875, n7751);
nor_4  g03721(new_n6070, n26823, n2035);
not_3  g03722(new_n6071, new_n6070);
xor_3  g03723(new_n6072, n26823, n2035);
nor_4  g03724(new_n6073, n5213, n4812);
not_3  g03725(new_n6074, new_n6073);
xor_3  g03726(new_n6075, n5213, n4812);
nor_4  g03727(new_n6076, n24278, n4665);
not_3  g03728(new_n6077, new_n6076);
xor_3  g03729(new_n6078, n24278, n4665);
nor_4  g03730(new_n6079, n24618, n19005);
not_3  g03731(new_n6080, new_n6079);
nand_4 g03732(new_n6081, n24618, n19005);
not_3  g03733(new_n6082, new_n6081);
nor_4  g03734(new_n6083, new_n6082, new_n6079);
nor_4  g03735(new_n6084_1, n4326, n3952);
not_3  g03736(new_n6085, new_n6084_1);
nand_4 g03737(new_n6086, n12315, n5438);
nand_4 g03738(new_n6087, n4326, n3952);
not_3  g03739(new_n6088, new_n6087);
nor_4  g03740(new_n6089, new_n6088, new_n6084_1);
nand_4 g03741(new_n6090, new_n6089, new_n6086);
nand_4 g03742(new_n6091, new_n6090, new_n6085);
nand_4 g03743(new_n6092, new_n6091, new_n6083);
nand_4 g03744(new_n6093, new_n6092, new_n6080);
nand_4 g03745(new_n6094, new_n6093, new_n6078);
nand_4 g03746(new_n6095, new_n6094, new_n6077);
nand_4 g03747(new_n6096, new_n6095, new_n6075);
nand_4 g03748(new_n6097, new_n6096, new_n6074);
nand_4 g03749(new_n6098, new_n6097, new_n6072);
nand_4 g03750(new_n6099, new_n6098, new_n6071);
nand_4 g03751(new_n6100, new_n6099, new_n6069);
nand_4 g03752(new_n6101, new_n6100, new_n6068);
nand_4 g03753(new_n6102, new_n6101, new_n6067);
nand_4 g03754(new_n6103, new_n6102, new_n6066);
nor_4  g03755(new_n6104_1, new_n6103, new_n6064);
not_3  g03756(new_n6105_1, new_n6064);
not_3  g03757(new_n6106, new_n6067);
not_3  g03758(new_n6107, new_n6101);
nor_4  g03759(new_n6108, new_n6107, new_n6106);
nor_4  g03760(new_n6109, new_n6108, new_n6065);
nor_4  g03761(new_n6110, new_n6109, new_n6105_1);
nor_4  g03762(new_n6111, new_n6110, new_n6104_1);
not_3  g03763(new_n6112, new_n6111);
xor_3  g03764(new_n6113, n10763, n5696);
nor_4  g03765(new_n6114, n13367, n7437);
xor_3  g03766(new_n6115, n13367, n7437);
not_3  g03767(new_n6116, new_n6115);
not_3  g03768(new_n6117, n932);
nand_4 g03769(new_n6118, new_n3037, new_n6117);
xor_3  g03770(new_n6119, n20700, n932);
nor_4  g03771(new_n6120, n7099, n6691);
not_3  g03772(new_n6121, new_n6120);
xor_3  g03773(new_n6122, n7099, n6691);
nor_4  g03774(new_n6123, n12811, n3260);
not_3  g03775(new_n6124, new_n6123);
xor_3  g03776(new_n6125, n12811, n3260);
nor_4  g03777(new_n6126, n20489, n1118);
not_3  g03778(new_n6127, new_n6126);
xor_3  g03779(new_n6128, n20489, n1118);
nor_4  g03780(new_n6129, n25974, n2355);
not_3  g03781(new_n6130, new_n6129);
nand_4 g03782(new_n6131, n25974, n2355);
not_3  g03783(new_n6132, new_n6131);
nor_4  g03784(new_n6133, new_n6132, new_n6129);
nor_4  g03785(new_n6134, n11121, n1630);
not_3  g03786(new_n6135, new_n6134);
nand_4 g03787(new_n6136, n16217, n1451);
nand_4 g03788(new_n6137, n11121, n1630);
not_3  g03789(new_n6138, new_n6137);
nor_4  g03790(new_n6139, new_n6138, new_n6134);
nand_4 g03791(new_n6140, new_n6139, new_n6136);
nand_4 g03792(new_n6141, new_n6140, new_n6135);
nand_4 g03793(new_n6142, new_n6141, new_n6133);
nand_4 g03794(new_n6143, new_n6142, new_n6130);
nand_4 g03795(new_n6144, new_n6143, new_n6128);
nand_4 g03796(new_n6145, new_n6144, new_n6127);
nand_4 g03797(new_n6146, new_n6145, new_n6125);
nand_4 g03798(new_n6147, new_n6146, new_n6124);
nand_4 g03799(new_n6148, new_n6147, new_n6122);
nand_4 g03800(new_n6149, new_n6148, new_n6121);
nand_4 g03801(new_n6150, new_n6149, new_n6119);
nand_4 g03802(new_n6151, new_n6150, new_n6118);
not_3  g03803(new_n6152, new_n6151);
nor_4  g03804(new_n6153, new_n6152, new_n6116);
nor_4  g03805(new_n6154, new_n6153, new_n6114);
xor_3  g03806(new_n6155, new_n6154, new_n6113);
xnor_3 g03807(new_n6156, new_n6155, new_n6112);
xor_3  g03808(new_n6157, new_n6152, new_n6115);
xnor_3 g03809(new_n6158, new_n6101, new_n6067);
not_3  g03810(new_n6159, new_n6158);
nand_4 g03811(new_n6160_1, new_n6159, new_n6157);
xor_3  g03812(new_n6161, new_n6152, new_n6116);
nor_4  g03813(new_n6162, new_n6158, new_n6161);
nor_4  g03814(new_n6163, new_n6159, new_n6157);
nor_4  g03815(new_n6164, new_n6163, new_n6162);
xnor_3 g03816(new_n6165, new_n6149, new_n6119);
not_3  g03817(new_n6166, new_n6069);
xnor_3 g03818(new_n6167, new_n6099, new_n6166);
nor_4  g03819(new_n6168, new_n6167, new_n6165);
xnor_3 g03820(new_n6169, new_n6167, new_n6165);
xnor_3 g03821(new_n6170, new_n6147, new_n6122);
not_3  g03822(new_n6171_1, new_n6072);
xnor_3 g03823(new_n6172, new_n6097, new_n6171_1);
nor_4  g03824(new_n6173, new_n6172, new_n6170);
not_3  g03825(new_n6174, new_n6144);
nor_4  g03826(new_n6175, new_n6143, new_n6128);
nor_4  g03827(new_n6176, new_n6175, new_n6174);
not_3  g03828(new_n6177, new_n6094);
nor_4  g03829(new_n6178, new_n6093, new_n6078);
nor_4  g03830(new_n6179, new_n6178, new_n6177);
not_3  g03831(new_n6180, new_n6179);
nand_4 g03832(new_n6181, new_n6180, new_n6176);
not_3  g03833(new_n6182, new_n6181);
xnor_3 g03834(new_n6183_1, new_n6179, new_n6176);
not_3  g03835(new_n6184, new_n6183_1);
not_3  g03836(new_n6185, new_n6142);
nor_4  g03837(new_n6186, new_n6141, new_n6133);
nor_4  g03838(new_n6187, new_n6186, new_n6185);
not_3  g03839(new_n6188, new_n6187);
not_3  g03840(new_n6189_1, new_n6092);
nor_4  g03841(new_n6190, new_n6091, new_n6083);
nor_4  g03842(new_n6191, new_n6190, new_n6189_1);
nor_4  g03843(new_n6192, new_n6191, new_n6188);
not_3  g03844(new_n6193, new_n6192);
not_3  g03845(new_n6194, new_n6090);
nor_4  g03846(new_n6195, new_n6089, new_n6086);
nor_4  g03847(new_n6196, new_n6195, new_n6194);
not_3  g03848(new_n6197, new_n6140);
nor_4  g03849(new_n6198, new_n6139, new_n6136);
nor_4  g03850(new_n6199, new_n6198, new_n6197);
not_3  g03851(new_n6200, new_n6199);
nor_4  g03852(new_n6201, new_n6200, new_n6196);
not_3  g03853(new_n6202, new_n6201);
xnor_3 g03854(new_n6203, n12315, n5438);
xor_3  g03855(new_n6204_1, n16217, n1451);
nor_4  g03856(new_n6205, new_n6204_1, new_n6203);
not_3  g03857(new_n6206, new_n6196);
nor_4  g03858(new_n6207, new_n6199, new_n6206);
nor_4  g03859(new_n6208, new_n6207, new_n6201);
nand_4 g03860(new_n6209, new_n6208, new_n6205);
nand_4 g03861(new_n6210, new_n6209, new_n6202);
not_3  g03862(new_n6211, new_n6191);
nor_4  g03863(new_n6212, new_n6211, new_n6187);
nor_4  g03864(new_n6213, new_n6212, new_n6192);
nand_4 g03865(new_n6214, new_n6213, new_n6210);
nand_4 g03866(new_n6215, new_n6214, new_n6193);
not_3  g03867(new_n6216, new_n6215);
nor_4  g03868(new_n6217, new_n6216, new_n6184);
nor_4  g03869(new_n6218_1, new_n6217, new_n6182);
not_3  g03870(new_n6219, new_n6146);
nor_4  g03871(new_n6220, new_n6145, new_n6125);
nor_4  g03872(new_n6221, new_n6220, new_n6219);
not_3  g03873(new_n6222, new_n6221);
nand_4 g03874(new_n6223_1, new_n6222, new_n6218_1);
nand_4 g03875(new_n6224, new_n6215, new_n6183_1);
nand_4 g03876(new_n6225, new_n6224, new_n6181);
xnor_3 g03877(new_n6226, new_n6222, new_n6225);
xnor_3 g03878(new_n6227, new_n6095, new_n6075);
not_3  g03879(new_n6228, new_n6227);
nand_4 g03880(new_n6229, new_n6228, new_n6226);
nand_4 g03881(new_n6230, new_n6229, new_n6223_1);
xnor_3 g03882(new_n6231, new_n6172, new_n6170);
nor_4  g03883(new_n6232, new_n6231, new_n6230);
nor_4  g03884(new_n6233_1, new_n6232, new_n6173);
nor_4  g03885(new_n6234, new_n6233_1, new_n6169);
nor_4  g03886(new_n6235, new_n6234, new_n6168);
nand_4 g03887(new_n6236, new_n6235, new_n6164);
nand_4 g03888(new_n6237, new_n6236, new_n6160_1);
xnor_3 g03889(new_n6238, new_n6237, new_n6156);
xnor_3 g03890(new_n6239, new_n6238, new_n6063);
xnor_3 g03891(new_n6240, new_n6060, new_n6021);
xnor_3 g03892(new_n6241, new_n6158, new_n6161);
xnor_3 g03893(new_n6242, new_n6235, new_n6241);
nor_4  g03894(new_n6243, new_n6242, new_n6240);
xnor_3 g03895(new_n6244, new_n6242, new_n6240);
xnor_3 g03896(new_n6245_1, new_n6058, new_n6025);
not_3  g03897(new_n6246, new_n6245_1);
not_3  g03898(new_n6247, new_n6169);
not_3  g03899(new_n6248_1, new_n6173);
not_3  g03900(new_n6249, new_n6230);
not_3  g03901(new_n6250, new_n6231);
nand_4 g03902(new_n6251, new_n6250, new_n6249);
nand_4 g03903(new_n6252, new_n6251, new_n6248_1);
xnor_3 g03904(new_n6253, new_n6252, new_n6247);
nor_4  g03905(new_n6254, new_n6253, new_n6246);
xnor_3 g03906(new_n6255, new_n6253, new_n6246);
not_3  g03907(new_n6256_1, new_n6033);
nand_4 g03908(new_n6257, new_n6054, new_n6256_1);
xnor_3 g03909(new_n6258, new_n6257, new_n6030);
xnor_3 g03910(new_n6259, new_n6231, new_n6230);
nor_4  g03911(new_n6260, new_n6259, new_n6258);
xnor_3 g03912(new_n6261, new_n6259, new_n6258);
not_3  g03913(new_n6262, new_n6035);
xnor_3 g03914(new_n6263, new_n6053, new_n6262);
xnor_3 g03915(new_n6264, new_n6221, new_n6225);
xnor_3 g03916(new_n6265, new_n6227, new_n6264);
nand_4 g03917(new_n6266, new_n6265, new_n6263);
not_3  g03918(new_n6267, new_n6266);
xnor_3 g03919(new_n6268, new_n6265, new_n6263);
nor_4  g03920(new_n6269, new_n6215, new_n6183_1);
nor_4  g03921(new_n6270, new_n6269, new_n6217);
not_3  g03922(new_n6271_1, new_n6270);
xnor_3 g03923(new_n6272, new_n6051, new_n6050);
nor_4  g03924(new_n6273, new_n6272, new_n6271_1);
xnor_3 g03925(new_n6274, new_n6272, new_n6271_1);
not_3  g03926(new_n6275, new_n6042);
xnor_3 g03927(new_n6276_1, new_n6048, new_n6275);
not_3  g03928(new_n6277, new_n6214);
nor_4  g03929(new_n6278, new_n6213, new_n6210);
nor_4  g03930(new_n6279, new_n6278, new_n6277);
nor_4  g03931(new_n6280, new_n6279, new_n6276_1);
not_3  g03932(new_n6281, new_n6280);
xnor_3 g03933(new_n6282, new_n6048, new_n6042);
not_3  g03934(new_n6283, new_n6279);
nor_4  g03935(new_n6284, new_n6283, new_n6282);
nor_4  g03936(new_n6285, new_n6284, new_n6280);
not_3  g03937(new_n6286, new_n6209);
nor_4  g03938(new_n6287, new_n6208, new_n6205);
nor_4  g03939(new_n6288, new_n6287, new_n6286);
not_3  g03940(new_n6289, new_n6288);
nor_4  g03941(new_n6290, new_n6289, new_n6046_1);
not_3  g03942(new_n6291, new_n6046_1);
xor_3  g03943(new_n6292, new_n6291, new_n6045);
not_3  g03944(new_n6293, new_n6292);
nor_4  g03945(new_n6294, new_n6293, new_n6288);
xor_3  g03946(new_n6295, n23333, n11424);
not_3  g03947(new_n6296, new_n6295);
not_3  g03948(new_n6297, new_n6204_1);
xor_3  g03949(new_n6298, new_n6297, new_n6203);
not_3  g03950(new_n6299, new_n6298);
nor_4  g03951(new_n6300, new_n6299, new_n6296);
nor_4  g03952(new_n6301, new_n6300, new_n6294);
nor_4  g03953(new_n6302, new_n6301, new_n6290);
nand_4 g03954(new_n6303, new_n6302, new_n6285);
nand_4 g03955(new_n6304, new_n6303, new_n6281);
nor_4  g03956(new_n6305, new_n6304, new_n6274);
nor_4  g03957(new_n6306, new_n6305, new_n6273);
nor_4  g03958(new_n6307, new_n6306, new_n6268);
nor_4  g03959(new_n6308_1, new_n6307, new_n6267);
nor_4  g03960(new_n6309, new_n6308_1, new_n6261);
nor_4  g03961(new_n6310, new_n6309, new_n6260);
nor_4  g03962(new_n6311_1, new_n6310, new_n6255);
nor_4  g03963(new_n6312, new_n6311_1, new_n6254);
nor_4  g03964(new_n6313, new_n6312, new_n6244);
nor_4  g03965(new_n6314, new_n6313, new_n6243);
nand_4 g03966(new_n6315, new_n6314, new_n6239);
not_3  g03967(new_n6316, new_n6315);
nor_4  g03968(new_n6317, new_n6314, new_n6239);
nor_4  g03969(n431, new_n6317, new_n6316);
not_3  g03970(new_n6319, n23895);
nor_4  g03971(new_n6320, new_n6319, n8614);
not_3  g03972(new_n6321, n8614);
xor_3  g03973(new_n6322, n23895, new_n6321);
not_3  g03974(new_n6323_1, new_n6322);
not_3  g03975(new_n6324, n17351);
nor_4  g03976(new_n6325, new_n6324, n15182);
not_3  g03977(new_n6326, n15182);
xor_3  g03978(new_n6327, n17351, new_n6326);
not_3  g03979(new_n6328, n27037);
nand_4 g03980(new_n6329, new_n6328, n11736);
not_3  g03981(new_n6330_1, n11736);
xor_3  g03982(new_n6331, n27037, new_n6330_1);
not_3  g03983(new_n6332, n8964);
nand_4 g03984(new_n6333, n23200, new_n6332);
xor_3  g03985(new_n6334, n23200, new_n6332);
not_3  g03986(new_n6335, n17959);
nor_4  g03987(new_n6336, n20151, new_n6335);
not_3  g03988(new_n6337, new_n6336);
xor_3  g03989(new_n6338, n20151, new_n6335);
not_3  g03990(new_n6339_1, n7566);
nor_4  g03991(new_n6340, n7693, new_n6339_1);
xor_3  g03992(new_n6341, n7693, new_n6339_1);
not_3  g03993(new_n6342, new_n6341);
not_3  g03994(new_n6343, n7731);
nor_4  g03995(new_n6344, n10405, new_n6343);
xor_3  g03996(new_n6345, n10405, n7731);
not_3  g03997(new_n6346, n11302);
nor_4  g03998(new_n6347, n12341, new_n6346);
not_3  g03999(new_n6348, n12341);
nor_4  g04000(new_n6349, new_n6348, n11302);
nor_4  g04001(new_n6350, n20986, new_n4477);
not_3  g04002(new_n6351, n20986);
nor_4  g04003(new_n6352, new_n6351, n17090);
not_3  g04004(new_n6353, n6773);
nor_4  g04005(new_n6354_1, n12384, new_n6353);
not_3  g04006(new_n6355, new_n6354_1);
nor_4  g04007(new_n6356_1, new_n6355, new_n6352);
nor_4  g04008(new_n6357, new_n6356_1, new_n6350);
nor_4  g04009(new_n6358, new_n6357, new_n6349);
nor_4  g04010(new_n6359, new_n6358, new_n6347);
not_3  g04011(new_n6360, new_n6359);
nor_4  g04012(new_n6361, new_n6360, new_n6345);
nor_4  g04013(new_n6362, new_n6361, new_n6344);
nor_4  g04014(new_n6363, new_n6362, new_n6342);
nor_4  g04015(new_n6364, new_n6363, new_n6340);
not_3  g04016(new_n6365, new_n6364);
nand_4 g04017(new_n6366, new_n6365, new_n6338);
nand_4 g04018(new_n6367, new_n6366, new_n6337);
nand_4 g04019(new_n6368, new_n6367, new_n6334);
nand_4 g04020(new_n6369_1, new_n6368, new_n6333);
nand_4 g04021(new_n6370, new_n6369_1, new_n6331);
nand_4 g04022(new_n6371, new_n6370, new_n6329);
nand_4 g04023(new_n6372, new_n6371, new_n6327);
not_3  g04024(new_n6373, new_n6372);
nor_4  g04025(new_n6374, new_n6373, new_n6325);
nor_4  g04026(new_n6375_1, new_n6374, new_n6323_1);
nor_4  g04027(new_n6376, new_n6375_1, new_n6320);
not_3  g04028(new_n6377, n13494);
nor_4  g04029(new_n6378, n18880, new_n6377);
xor_3  g04030(new_n6379_1, n18880, new_n6377);
not_3  g04031(new_n6380, new_n6379_1);
not_3  g04032(new_n6381_1, n25345);
nor_4  g04033(new_n6382, n25475, new_n6381_1);
xor_3  g04034(new_n6383_1, n25475, new_n6381_1);
nand_4 g04035(new_n6384, new_n5013, n9655);
not_3  g04036(new_n6385_1, n9655);
xor_3  g04037(new_n6386, n23849, new_n6385_1);
nand_4 g04038(new_n6387, n13490, new_n5022);
xor_3  g04039(new_n6388, n13490, new_n5022);
nand_4 g04040(new_n6389, n22660, new_n4335);
xor_3  g04041(new_n6390, n22660, new_n4335);
not_3  g04042(new_n6391, n1777);
nor_4  g04043(new_n6392, n16029, new_n6391);
not_3  g04044(new_n6393, new_n6392);
xor_3  g04045(new_n6394, n16029, new_n6391);
not_3  g04046(new_n6395, n8745);
nor_4  g04047(new_n6396, n16476, new_n6395);
not_3  g04048(new_n6397_1, new_n6396);
xor_3  g04049(new_n6398, n16476, new_n6395);
nor_4  g04050(new_n6399, n15636, new_n4371);
not_3  g04051(new_n6400, new_n6399);
not_3  g04052(new_n6401, n15636);
nor_4  g04053(new_n6402, new_n6401, n11615);
not_3  g04054(new_n6403, new_n6402);
nor_4  g04055(new_n6404, new_n4375, n20077);
not_3  g04056(new_n6405, new_n6404);
not_3  g04057(new_n6406, n20077);
nor_4  g04058(new_n6407_1, n22433, new_n6406);
not_3  g04059(new_n6408, new_n6407_1);
not_3  g04060(new_n6409, n14090);
nor_4  g04061(new_n6410, new_n6409, n6794);
nand_4 g04062(new_n6411, new_n6410, new_n6408);
nand_4 g04063(new_n6412, new_n6411, new_n6405);
nand_4 g04064(new_n6413, new_n6412, new_n6403);
nand_4 g04065(new_n6414, new_n6413, new_n6400);
not_3  g04066(new_n6415, new_n6414);
nand_4 g04067(new_n6416, new_n6415, new_n6398);
nand_4 g04068(new_n6417, new_n6416, new_n6397_1);
nand_4 g04069(new_n6418, new_n6417, new_n6394);
nand_4 g04070(new_n6419, new_n6418, new_n6393);
nand_4 g04071(new_n6420, new_n6419, new_n6390);
nand_4 g04072(new_n6421, new_n6420, new_n6389);
nand_4 g04073(new_n6422, new_n6421, new_n6388);
nand_4 g04074(new_n6423, new_n6422, new_n6387);
nand_4 g04075(new_n6424, new_n6423, new_n6386);
nand_4 g04076(new_n6425, new_n6424, new_n6384);
nand_4 g04077(new_n6426, new_n6425, new_n6383_1);
not_3  g04078(new_n6427_1, new_n6426);
nor_4  g04079(new_n6428, new_n6427_1, new_n6382);
nor_4  g04080(new_n6429, new_n6428, new_n6380);
nor_4  g04081(new_n6430, new_n6429, new_n6378);
not_3  g04082(new_n6431_1, new_n6430);
xnor_3 g04083(new_n6432, new_n6428, new_n6379_1);
not_3  g04084(new_n6433, n26797);
not_3  g04085(new_n6434, n22554);
not_3  g04086(new_n6435, n3909);
not_3  g04087(new_n6436, n2146);
nor_4  g04088(new_n6437_1, n22173, n583);
nand_4 g04089(new_n6438, new_n6437_1, new_n6436);
nor_4  g04090(new_n6439, new_n6438, n23974);
nand_4 g04091(new_n6440, new_n6439, new_n6435);
nor_4  g04092(new_n6441, new_n6440, n20429);
nand_4 g04093(new_n6442, new_n6441, new_n6434);
nor_4  g04094(new_n6443, new_n6442, n23913);
xor_3  g04095(new_n6444, new_n6443, new_n6433);
nor_4  g04096(new_n6445, new_n6444, n10201);
not_3  g04097(new_n6446, new_n6444);
xor_3  g04098(new_n6447, new_n6446, n10201);
xor_3  g04099(new_n6448, new_n6442, n23913);
nor_4  g04100(new_n6449, new_n6448, n10593);
not_3  g04101(new_n6450, new_n6448);
xor_3  g04102(new_n6451, new_n6450, n10593);
xor_3  g04103(new_n6452, new_n6441, new_n6434);
nor_4  g04104(new_n6453, new_n6452, n18290);
not_3  g04105(new_n6454, new_n6452);
xor_3  g04106(new_n6455, new_n6454, n18290);
nand_4 g04107(new_n6456_1, new_n6440, n20429);
not_3  g04108(new_n6457_1, new_n6456_1);
nor_4  g04109(new_n6458, new_n6457_1, new_n6441);
nor_4  g04110(new_n6459, new_n6458, n11580);
xnor_3 g04111(new_n6460, new_n6458, n11580);
xnor_3 g04112(new_n6461, new_n6439, n3909);
nor_4  g04113(new_n6462, new_n6461, n15884);
not_3  g04114(new_n6463, n15884);
not_3  g04115(new_n6464, new_n6461);
nor_4  g04116(new_n6465_1, new_n6464, new_n6463);
nor_4  g04117(new_n6466, new_n6465_1, new_n6462);
nand_4 g04118(new_n6467, new_n6438, n23974);
not_3  g04119(new_n6468, new_n6467);
nor_4  g04120(new_n6469, new_n6468, new_n6439);
nor_4  g04121(new_n6470_1, new_n6469, n6356);
not_3  g04122(new_n6471, new_n6470_1);
xnor_3 g04123(new_n6472, new_n6437_1, n2146);
nor_4  g04124(new_n6473, new_n6472, n27104);
not_3  g04125(new_n6474, new_n6473);
not_3  g04126(new_n6475, n27104);
not_3  g04127(new_n6476_1, new_n6472);
nor_4  g04128(new_n6477, new_n6476_1, new_n6475);
nor_4  g04129(new_n6478, new_n6477, new_n6473);
not_3  g04130(new_n6479, n27188);
xnor_3 g04131(new_n6480, n22173, n583);
nand_4 g04132(new_n6481, new_n6480, new_n6479);
nand_4 g04133(new_n6482, n6611, n583);
xnor_3 g04134(new_n6483, new_n6480, n27188);
nand_4 g04135(new_n6484, new_n6483, new_n6482);
nand_4 g04136(new_n6485_1, new_n6484, new_n6481);
nand_4 g04137(new_n6486, new_n6485_1, new_n6478);
nand_4 g04138(new_n6487, new_n6486, new_n6474);
not_3  g04139(new_n6488, n6356);
not_3  g04140(new_n6489, new_n6469);
nor_4  g04141(new_n6490, new_n6489, new_n6488);
nor_4  g04142(new_n6491, new_n6490, new_n6470_1);
nand_4 g04143(new_n6492, new_n6491, new_n6487);
nand_4 g04144(new_n6493, new_n6492, new_n6471);
nand_4 g04145(new_n6494, new_n6493, new_n6466);
not_3  g04146(new_n6495, new_n6494);
nor_4  g04147(new_n6496, new_n6495, new_n6462);
nor_4  g04148(new_n6497, new_n6496, new_n6460);
nor_4  g04149(new_n6498, new_n6497, new_n6459);
nor_4  g04150(new_n6499, new_n6498, new_n6455);
nor_4  g04151(new_n6500, new_n6499, new_n6453);
nor_4  g04152(new_n6501, new_n6500, new_n6451);
nor_4  g04153(new_n6502_1, new_n6501, new_n6449);
nor_4  g04154(new_n6503, new_n6502_1, new_n6447);
nor_4  g04155(new_n6504, new_n6503, new_n6445);
not_3  g04156(new_n6505, n12702);
nand_4 g04157(new_n6506_1, new_n6443, new_n6433);
not_3  g04158(new_n6507, new_n6506_1);
xor_3  g04159(new_n6508, new_n6507, new_n6505);
nor_4  g04160(new_n6509, new_n6508, n12650);
not_3  g04161(new_n6510, n12650);
not_3  g04162(new_n6511, new_n6508);
nor_4  g04163(new_n6512, new_n6511, new_n6510);
nor_4  g04164(new_n6513_1, new_n6512, new_n6509);
xnor_3 g04165(new_n6514_1, new_n6513_1, new_n6504);
not_3  g04166(new_n6515, new_n6514_1);
nor_4  g04167(new_n6516, new_n6515, new_n6432);
xnor_3 g04168(new_n6517, new_n6428, new_n6380);
xnor_3 g04169(new_n6518, new_n6514_1, new_n6517);
xnor_3 g04170(new_n6519, new_n6425, new_n6383_1);
not_3  g04171(new_n6520, new_n6519);
xnor_3 g04172(new_n6521, new_n6502_1, new_n6447);
nor_4  g04173(new_n6522, new_n6521, new_n6520);
xnor_3 g04174(new_n6523, new_n6521, new_n6520);
xnor_3 g04175(new_n6524, new_n6423, new_n6386);
not_3  g04176(new_n6525, new_n6500);
xnor_3 g04177(new_n6526, new_n6525, new_n6451);
nand_4 g04178(new_n6527, new_n6526, new_n6524);
not_3  g04179(new_n6528, new_n6386);
xnor_3 g04180(new_n6529, new_n6423, new_n6528);
xnor_3 g04181(new_n6530, new_n6526, new_n6529);
xnor_3 g04182(new_n6531, new_n6421, new_n6388);
not_3  g04183(new_n6532, new_n6498);
xnor_3 g04184(new_n6533, new_n6532, new_n6455);
nand_4 g04185(new_n6534, new_n6533, new_n6531);
not_3  g04186(new_n6535, new_n6531);
xnor_3 g04187(new_n6536, new_n6533, new_n6535);
xnor_3 g04188(new_n6537, new_n6419, new_n6390);
not_3  g04189(new_n6538, new_n6460);
not_3  g04190(new_n6539, new_n6496);
nor_4  g04191(new_n6540, new_n6539, new_n6538);
nor_4  g04192(new_n6541, new_n6540, new_n6497);
nand_4 g04193(new_n6542_1, new_n6541, new_n6537);
not_3  g04194(new_n6543, new_n6390);
xnor_3 g04195(new_n6544, new_n6419, new_n6543);
xnor_3 g04196(new_n6545, new_n6541, new_n6544);
xnor_3 g04197(new_n6546, new_n6417, new_n6394);
not_3  g04198(new_n6547, new_n6546);
xnor_3 g04199(new_n6548, new_n6493, new_n6466);
nor_4  g04200(new_n6549, new_n6548, new_n6547);
not_3  g04201(new_n6550, new_n6549);
not_3  g04202(new_n6551, new_n6548);
nor_4  g04203(new_n6552, new_n6551, new_n6546);
nor_4  g04204(new_n6553, new_n6552, new_n6549);
xor_3  g04205(new_n6554, n16476, n8745);
xnor_3 g04206(new_n6555, new_n6414, new_n6554);
xnor_3 g04207(new_n6556_1, new_n6491, new_n6487);
not_3  g04208(new_n6557, new_n6556_1);
nand_4 g04209(new_n6558_1, new_n6557, new_n6555);
not_3  g04210(new_n6559, new_n6558_1);
nor_4  g04211(new_n6560_1, new_n6557, new_n6555);
nor_4  g04212(new_n6561, new_n6560_1, new_n6559);
xnor_3 g04213(new_n6562, new_n6485_1, new_n6478);
not_3  g04214(new_n6563, new_n6562);
nor_4  g04215(new_n6564, new_n6402, new_n6399);
xnor_3 g04216(new_n6565, new_n6564, new_n6412);
not_3  g04217(new_n6566, new_n6565);
nor_4  g04218(new_n6567_1, new_n6566, new_n6563);
xnor_3 g04219(new_n6568, new_n6565, new_n6562);
xnor_3 g04220(new_n6569, new_n6483, new_n6482);
not_3  g04221(new_n6570, new_n6569);
nor_4  g04222(new_n6571, new_n6407_1, new_n6404);
xnor_3 g04223(new_n6572, new_n6571, new_n6410);
not_3  g04224(new_n6573, new_n6572);
nor_4  g04225(new_n6574, new_n6573, new_n6570);
not_3  g04226(new_n6575, n6794);
nor_4  g04227(new_n6576_1, n14090, new_n6575);
nor_4  g04228(new_n6577, new_n6576_1, new_n6410);
not_3  g04229(new_n6578, new_n6577);
xor_3  g04230(new_n6579, n6611, n583);
nand_4 g04231(new_n6580, new_n6579, new_n6578);
xnor_3 g04232(new_n6581, new_n6572, new_n6569);
nor_4  g04233(new_n6582, new_n6581, new_n6580);
nor_4  g04234(new_n6583, new_n6582, new_n6574);
nor_4  g04235(new_n6584, new_n6583, new_n6568);
nor_4  g04236(new_n6585, new_n6584, new_n6567_1);
nand_4 g04237(new_n6586, new_n6585, new_n6561);
nand_4 g04238(new_n6587_1, new_n6586, new_n6558_1);
nand_4 g04239(new_n6588, new_n6587_1, new_n6553);
nand_4 g04240(new_n6589, new_n6588, new_n6550);
nand_4 g04241(new_n6590_1, new_n6589, new_n6545);
nand_4 g04242(new_n6591, new_n6590_1, new_n6542_1);
nand_4 g04243(new_n6592, new_n6591, new_n6536);
nand_4 g04244(new_n6593, new_n6592, new_n6534);
nand_4 g04245(new_n6594, new_n6593, new_n6530);
nand_4 g04246(new_n6595, new_n6594, new_n6527);
not_3  g04247(new_n6596_1, new_n6595);
nor_4  g04248(new_n6597, new_n6596_1, new_n6523);
nor_4  g04249(new_n6598, new_n6597, new_n6522);
nor_4  g04250(new_n6599, new_n6598, new_n6518);
nor_4  g04251(new_n6600, new_n6599, new_n6516);
nor_4  g04252(new_n6601, new_n6506_1, n12702);
not_3  g04253(new_n6602, new_n6601);
not_3  g04254(new_n6603, new_n6504);
nor_4  g04255(new_n6604, new_n6509, new_n6603);
nor_4  g04256(new_n6605, new_n6604, new_n6512);
nand_4 g04257(new_n6606, new_n6605, new_n6602);
nand_4 g04258(new_n6607, new_n6606, new_n6600);
nor_4  g04259(new_n6608, new_n6607, new_n6431_1);
not_3  g04260(new_n6609, new_n6516);
not_3  g04261(new_n6610, new_n6518);
not_3  g04262(new_n6611_1, new_n6522);
not_3  g04263(new_n6612_1, new_n6523);
nand_4 g04264(new_n6613, new_n6595, new_n6612_1);
nand_4 g04265(new_n6614, new_n6613, new_n6611_1);
nand_4 g04266(new_n6615, new_n6614, new_n6610);
nand_4 g04267(new_n6616, new_n6615, new_n6609);
not_3  g04268(new_n6617, new_n6606);
nand_4 g04269(new_n6618, new_n6617, new_n6616);
nor_4  g04270(new_n6619, new_n6618, new_n6430);
nor_4  g04271(new_n6620, new_n6619, new_n6608);
nor_4  g04272(new_n6621, new_n6620, new_n6376);
not_3  g04273(new_n6622, new_n6376);
not_3  g04274(new_n6623, new_n6620);
nor_4  g04275(new_n6624, new_n6623, new_n6622);
nor_4  g04276(new_n6625, new_n6624, new_n6621);
nand_4 g04277(new_n6626, new_n6618, new_n6607);
xnor_3 g04278(new_n6627, new_n6626, new_n6430);
nor_4  g04279(new_n6628_1, new_n6627, new_n6622);
not_3  g04280(new_n6629, new_n6628_1);
xnor_3 g04281(new_n6630_1, new_n6626, new_n6431_1);
nor_4  g04282(new_n6631_1, new_n6630_1, new_n6376);
not_3  g04283(new_n6632, new_n6631_1);
xor_3  g04284(new_n6633, new_n6374, new_n6323_1);
xnor_3 g04285(new_n6634_1, new_n6598, new_n6518);
nor_4  g04286(new_n6635, new_n6634_1, new_n6633);
xnor_3 g04287(new_n6636, new_n6634_1, new_n6633);
xor_3  g04288(new_n6637, new_n6371, new_n6327);
xnor_3 g04289(new_n6638, new_n6595, new_n6612_1);
nor_4  g04290(new_n6639, new_n6638, new_n6637);
not_3  g04291(new_n6640, new_n6637);
not_3  g04292(new_n6641, new_n6638);
nor_4  g04293(new_n6642, new_n6641, new_n6640);
nor_4  g04294(new_n6643, new_n6642, new_n6639);
not_3  g04295(new_n6644, new_n6643);
xor_3  g04296(new_n6645, new_n6369_1, new_n6331);
xnor_3 g04297(new_n6646, new_n6593, new_n6530);
nor_4  g04298(new_n6647, new_n6646, new_n6645);
not_3  g04299(new_n6648, new_n6645);
not_3  g04300(new_n6649, new_n6646);
nor_4  g04301(new_n6650, new_n6649, new_n6648);
nor_4  g04302(new_n6651, new_n6650, new_n6647);
xor_3  g04303(new_n6652_1, new_n6367, new_n6334);
not_3  g04304(new_n6653, new_n6652_1);
not_3  g04305(new_n6654, new_n6536);
xnor_3 g04306(new_n6655_1, new_n6591, new_n6654);
nand_4 g04307(new_n6656, new_n6655_1, new_n6653);
xnor_3 g04308(new_n6657, new_n6655_1, new_n6652_1);
xor_3  g04309(new_n6658, new_n6365, new_n6338);
not_3  g04310(new_n6659_1, new_n6658);
not_3  g04311(new_n6660, new_n6545);
xnor_3 g04312(new_n6661, new_n6589, new_n6660);
nand_4 g04313(new_n6662, new_n6661, new_n6659_1);
xnor_3 g04314(new_n6663, new_n6661, new_n6658);
xor_3  g04315(new_n6664, new_n6362, new_n6342);
not_3  g04316(new_n6665, new_n6664);
not_3  g04317(new_n6666, new_n6587_1);
xnor_3 g04318(new_n6667, new_n6666, new_n6553);
nand_4 g04319(new_n6668, new_n6667, new_n6665);
xnor_3 g04320(new_n6669_1, new_n6667, new_n6664);
not_3  g04321(new_n6670, new_n6586);
nor_4  g04322(new_n6671_1, new_n6585, new_n6561);
nor_4  g04323(new_n6672, new_n6671_1, new_n6670);
xor_3  g04324(new_n6673_1, new_n6360, new_n6345);
not_3  g04325(new_n6674_1, new_n6673_1);
nand_4 g04326(new_n6675, new_n6674_1, new_n6672);
xnor_3 g04327(new_n6676, new_n6673_1, new_n6672);
not_3  g04328(new_n6677, new_n6568);
not_3  g04329(new_n6678, new_n6583);
nor_4  g04330(new_n6679, new_n6678, new_n6677);
nor_4  g04331(new_n6680, new_n6679, new_n6584);
not_3  g04332(new_n6681, new_n6680);
not_3  g04333(new_n6682, new_n6357);
nor_4  g04334(new_n6683, new_n6349, new_n6347);
xor_3  g04335(new_n6684_1, new_n6683, new_n6682);
nand_4 g04336(new_n6685, new_n6684_1, new_n6681);
xnor_3 g04337(new_n6686, new_n6684_1, new_n6680);
xnor_3 g04338(new_n6687, new_n6579, new_n6578);
xor_3  g04339(new_n6688, n12384, new_n6353);
nor_4  g04340(new_n6689, new_n6688, new_n6687);
nor_4  g04341(new_n6690, new_n6352, new_n6350);
xor_3  g04342(new_n6691_1, new_n6690, new_n6354_1);
not_3  g04343(new_n6692, new_n6691_1);
nor_4  g04344(new_n6693, new_n6692, new_n6689);
not_3  g04345(new_n6694, new_n6693);
not_3  g04346(new_n6695, new_n6580);
xor_3  g04347(new_n6696, new_n6581, new_n6695);
not_3  g04348(new_n6697, new_n6689);
nor_4  g04349(new_n6698, new_n6691_1, new_n6697);
nor_4  g04350(new_n6699, new_n6698, new_n6693);
nand_4 g04351(new_n6700, new_n6699, new_n6696);
nand_4 g04352(new_n6701, new_n6700, new_n6694);
nand_4 g04353(new_n6702, new_n6701, new_n6686);
nand_4 g04354(new_n6703, new_n6702, new_n6685);
nand_4 g04355(new_n6704, new_n6703, new_n6676);
nand_4 g04356(new_n6705, new_n6704, new_n6675);
nand_4 g04357(new_n6706_1, new_n6705, new_n6669_1);
nand_4 g04358(new_n6707_1, new_n6706_1, new_n6668);
nand_4 g04359(new_n6708, new_n6707_1, new_n6663);
nand_4 g04360(new_n6709, new_n6708, new_n6662);
nand_4 g04361(new_n6710, new_n6709, new_n6657);
nand_4 g04362(new_n6711, new_n6710, new_n6656);
nand_4 g04363(new_n6712, new_n6711, new_n6651);
not_3  g04364(new_n6713, new_n6712);
nor_4  g04365(new_n6714, new_n6713, new_n6647);
nor_4  g04366(new_n6715, new_n6714, new_n6644);
nor_4  g04367(new_n6716, new_n6715, new_n6639);
nor_4  g04368(new_n6717, new_n6716, new_n6636);
nor_4  g04369(new_n6718, new_n6717, new_n6635);
nand_4 g04370(new_n6719, new_n6718, new_n6632);
nand_4 g04371(new_n6720, new_n6719, new_n6629);
xnor_3 g04372(n457, new_n6720, new_n6625);
not_3  g04373(new_n6722, n24323);
nor_4  g04374(new_n6723, new_n6722, n1681);
nor_4  g04375(new_n6724, n24323, new_n4957_1);
nor_4  g04376(new_n6725, new_n6724, new_n6723);
nand_4 g04377(new_n6726, n13781, n2088);
not_3  g04378(new_n6727, new_n6726);
nor_4  g04379(new_n6728, n13781, n2088);
nor_4  g04380(new_n6729_1, new_n6728, new_n6727);
not_3  g04381(new_n6730, new_n6729_1);
xor_3  g04382(new_n6731, new_n6730, new_n6725);
nand_4 g04383(new_n6732, new_n6731, new_n6578);
not_3  g04384(new_n6733, new_n6732);
xor_3  g04385(new_n6734, new_n6733, new_n6573);
nor_4  g04386(new_n6735, new_n6730, new_n6725);
not_3  g04387(new_n6736_1, new_n6735);
not_3  g04388(new_n6737, n25877);
nor_4  g04389(new_n6738, n26443, new_n6737);
nor_4  g04390(new_n6739, new_n4961, n25877);
nor_4  g04391(new_n6740, new_n6739, new_n6738);
xnor_3 g04392(new_n6741, new_n6740, new_n6724);
not_3  g04393(new_n6742, new_n6741);
nor_4  g04394(new_n6743, new_n6742, new_n6736_1);
nor_4  g04395(new_n6744, new_n6741, new_n6735);
nor_4  g04396(new_n6745, new_n6744, new_n6743);
nor_4  g04397(new_n6746, n9399, n2088);
nand_4 g04398(new_n6747, n9399, n2088);
not_3  g04399(new_n6748, new_n6747);
nor_4  g04400(new_n6749, new_n6748, new_n6746);
not_3  g04401(new_n6750, new_n6749);
nor_4  g04402(new_n6751, new_n6727, n11486);
nand_4 g04403(new_n6752, n13781, n11486);
nor_4  g04404(new_n6753, new_n6752, new_n4885);
nor_4  g04405(new_n6754, new_n6753, new_n6751);
nor_4  g04406(new_n6755, new_n6754, new_n6750);
nand_4 g04407(new_n6756, new_n6754, new_n6750);
not_3  g04408(new_n6757, new_n6756);
nor_4  g04409(new_n6758, new_n6757, new_n6755);
not_3  g04410(new_n6759, new_n6758);
nand_4 g04411(new_n6760, new_n6759, new_n6745);
not_3  g04412(new_n6761, new_n6760);
nor_4  g04413(new_n6762, new_n6759, new_n6745);
nor_4  g04414(new_n6763, new_n6762, new_n6761);
not_3  g04415(new_n6764, new_n6763);
xor_3  g04416(n463, new_n6764, new_n6734);
xor_3  g04417(new_n6766, n12121, n6775);
nor_4  g04418(new_n6767, new_n6766, n8920);
not_3  g04419(new_n6768, n8920);
not_3  g04420(new_n6769, new_n6766);
nor_4  g04421(new_n6770, new_n6769, new_n6768);
nor_4  g04422(new_n6771, new_n6770, new_n6767);
not_3  g04423(new_n6772, n5438);
xor_3  g04424(new_n6773_1, new_n3235_1, new_n6772);
xor_3  g04425(n491, new_n6773_1, new_n6771);
not_3  g04426(new_n6775_1, new_n6676);
xor_3  g04427(n496, new_n6703, new_n6775_1);
xnor_3 g04428(new_n6777, n25926, n12384);
xor_3  g04429(new_n6778, new_n6777, new_n6353);
not_3  g04430(new_n6779, new_n6778);
not_3  g04431(new_n6780, n16167);
xor_3  g04432(new_n6781, new_n6577, new_n6780);
not_3  g04433(new_n6782, new_n6781);
nor_4  g04434(new_n6783, new_n6782, new_n6779);
nor_4  g04435(new_n6784, new_n6577, new_n6780);
nor_4  g04436(new_n6785_1, new_n6572, n18745);
not_3  g04437(new_n6786, n18745);
nor_4  g04438(new_n6787, new_n6573, new_n6786);
nor_4  g04439(new_n6788, new_n6787, new_n6785_1);
not_3  g04440(new_n6789, new_n6788);
nor_4  g04441(new_n6790_1, new_n6789, new_n6784);
not_3  g04442(new_n6791_1, new_n6784);
nor_4  g04443(new_n6792, new_n6788, new_n6791_1);
nor_4  g04444(new_n6793, new_n6792, new_n6790_1);
not_3  g04445(new_n6794_1, new_n6793);
nand_4 g04446(new_n6795, n25926, n12384);
not_3  g04447(new_n6796, new_n6795);
xnor_3 g04448(new_n6797, n25926, n7657);
xnor_3 g04449(new_n6798, new_n6797, new_n6351);
not_3  g04450(new_n6799, new_n6798);
nor_4  g04451(new_n6800, new_n6799, new_n6796);
nor_4  g04452(new_n6801, new_n6798, new_n6795);
nor_4  g04453(new_n6802_1, new_n6801, new_n6800);
nor_4  g04454(new_n6803, new_n6777, new_n6353);
not_3  g04455(new_n6804, new_n6803);
nor_4  g04456(new_n6805, new_n6804, n17090);
nor_4  g04457(new_n6806, n17090, n6773);
not_3  g04458(new_n6807, new_n6806);
nand_4 g04459(new_n6808, n17090, n6773);
not_3  g04460(new_n6809, new_n6808);
nand_4 g04461(new_n6810, new_n6809, new_n6777);
nand_4 g04462(new_n6811, new_n6810, new_n6807);
nor_4  g04463(new_n6812, new_n6811, new_n6805);
not_3  g04464(new_n6813, new_n6812);
xnor_3 g04465(new_n6814_1, new_n6813, new_n6802_1);
xnor_3 g04466(new_n6815, new_n6814_1, new_n6794_1);
not_3  g04467(new_n6816, new_n6815);
xor_3  g04468(n498, new_n6816, new_n6783);
not_3  g04469(new_n6818, new_n5554);
nor_4  g04470(new_n6819, n25872, n19618);
nand_4 g04471(new_n6820, n25872, n19618);
not_3  g04472(new_n6821, new_n6820);
nor_4  g04473(new_n6822, new_n6821, new_n6819);
nor_4  g04474(new_n6823, n22043, n20259);
not_3  g04475(new_n6824, new_n6823);
nand_4 g04476(new_n6825, n12121, n3925);
nand_4 g04477(new_n6826_1, n22043, n20259);
not_3  g04478(new_n6827, new_n6826_1);
nor_4  g04479(new_n6828, new_n6827, new_n6823);
nand_4 g04480(new_n6829, new_n6828, new_n6825);
nand_4 g04481(new_n6830, new_n6829, new_n6824);
nor_4  g04482(new_n6831, new_n6830, new_n6822);
not_3  g04483(new_n6832, new_n6822);
not_3  g04484(new_n6833, new_n6829);
nor_4  g04485(new_n6834, new_n6833, new_n6823);
nor_4  g04486(new_n6835_1, new_n6834, new_n6832);
nor_4  g04487(new_n6836, new_n6835_1, new_n6831);
xnor_3 g04488(new_n6837, new_n6836, new_n6818);
nor_4  g04489(new_n6838, new_n6828, new_n6825);
nor_4  g04490(new_n6839, new_n6838, new_n6833);
nor_4  g04491(new_n6840, new_n6839, new_n5556);
xor_3  g04492(new_n6841, n12121, n3925);
nor_4  g04493(new_n6842, new_n6841, new_n5560);
xnor_3 g04494(new_n6843, new_n6839, new_n5556);
nor_4  g04495(new_n6844, new_n6843, new_n6842);
nor_4  g04496(new_n6845, new_n6844, new_n6840);
xnor_3 g04497(new_n6846, new_n6845, new_n6837);
xnor_3 g04498(new_n6847, new_n6846, new_n4157);
xnor_3 g04499(new_n6848, new_n6843, new_n6842);
not_3  g04500(new_n6849, new_n6848);
nor_4  g04501(new_n6850, new_n6849, new_n4118);
not_3  g04502(new_n6851, new_n6850);
nand_4 g04503(new_n6852, new_n6849, new_n4163);
not_3  g04504(new_n6853_1, new_n5560);
not_3  g04505(new_n6854, new_n6841);
xor_3  g04506(new_n6855, new_n6854, new_n6853_1);
not_3  g04507(new_n6856, new_n6855);
nand_4 g04508(new_n6857, new_n6856, new_n4314);
nand_4 g04509(new_n6858, new_n6857, new_n6852);
nand_4 g04510(new_n6859, new_n6858, new_n6851);
xor_3  g04511(n521, new_n6859, new_n6847);
xor_3  g04512(n548, new_n6688, new_n6687);
xor_3  g04513(n554, new_n4848, new_n4826);
not_3  g04514(new_n6863_1, n2979);
nor_4  g04515(new_n6864, n20658, n15743);
nand_4 g04516(new_n6865, new_n6864, new_n4155);
nor_4  g04517(new_n6866, new_n6865, n4957);
nand_4 g04518(new_n6867_1, new_n6866, new_n4141);
nor_4  g04519(new_n6868, new_n6867_1, n3161);
not_3  g04520(new_n6869, new_n6868);
nor_4  g04521(new_n6870, new_n6869, n25749);
not_3  g04522(new_n6871, new_n6870);
nor_4  g04523(new_n6872, new_n6871, n20409);
not_3  g04524(new_n6873, new_n6872);
nor_4  g04525(new_n6874, new_n6873, n647);
xor_3  g04526(new_n6875, new_n6874, new_n6863_1);
not_3  g04527(new_n6876, new_n6875);
xor_3  g04528(new_n6877, n9259, n6456);
not_3  g04529(new_n6878, new_n6877);
nor_4  g04530(new_n6879, n21489, n4085);
xor_3  g04531(new_n6880, n21489, n4085);
not_3  g04532(new_n6881, new_n6880);
nor_4  g04533(new_n6882, n26725, n20213);
xor_3  g04534(new_n6883, n26725, n20213);
not_3  g04535(new_n6884, new_n6883);
not_3  g04536(new_n6885, n11980);
nand_4 g04537(new_n6886, new_n3913, new_n6885);
xor_3  g04538(new_n6887, n13912, n11980);
not_3  g04539(new_n6888, n3253);
nand_4 g04540(new_n6889, new_n5535, new_n6888);
xor_3  g04541(new_n6890, n7670, n3253);
nor_4  g04542(new_n6891, n9598, n7759);
not_3  g04543(new_n6892, new_n6891);
xor_3  g04544(new_n6893, n9598, n7759);
nor_4  g04545(new_n6894, n22290, n12562);
not_3  g04546(new_n6895, new_n6894);
xor_3  g04547(new_n6896, n22290, n12562);
nor_4  g04548(new_n6897, n11273, n7949);
not_3  g04549(new_n6898, new_n6897);
nand_4 g04550(new_n6899, n11273, n7949);
not_3  g04551(new_n6900, new_n6899);
nor_4  g04552(new_n6901, new_n6900, new_n6897);
nor_4  g04553(new_n6902, n25565, n24374);
not_3  g04554(new_n6903, new_n6902);
nand_4 g04555(new_n6904, n21993, n14575);
nand_4 g04556(new_n6905, n25565, n24374);
not_3  g04557(new_n6906, new_n6905);
nor_4  g04558(new_n6907, new_n6906, new_n6902);
nand_4 g04559(new_n6908, new_n6907, new_n6904);
nand_4 g04560(new_n6909, new_n6908, new_n6903);
nand_4 g04561(new_n6910, new_n6909, new_n6901);
nand_4 g04562(new_n6911, new_n6910, new_n6898);
nand_4 g04563(new_n6912, new_n6911, new_n6896);
nand_4 g04564(new_n6913, new_n6912, new_n6895);
nand_4 g04565(new_n6914, new_n6913, new_n6893);
nand_4 g04566(new_n6915, new_n6914, new_n6892);
nand_4 g04567(new_n6916, new_n6915, new_n6890);
nand_4 g04568(new_n6917, new_n6916, new_n6889);
nand_4 g04569(new_n6918, new_n6917, new_n6887);
nand_4 g04570(new_n6919, new_n6918, new_n6886);
not_3  g04571(new_n6920, new_n6919);
nor_4  g04572(new_n6921, new_n6920, new_n6884);
nor_4  g04573(new_n6922, new_n6921, new_n6882);
nor_4  g04574(new_n6923, new_n6922, new_n6881);
nor_4  g04575(new_n6924, new_n6923, new_n6879);
xnor_3 g04576(new_n6925, new_n6924, new_n6878);
xnor_3 g04577(new_n6926, new_n6925, new_n6876);
not_3  g04578(new_n6927, new_n6926);
xor_3  g04579(new_n6928, new_n6873, n647);
not_3  g04580(new_n6929, new_n6928);
xnor_3 g04581(new_n6930, new_n6922, new_n6881);
nor_4  g04582(new_n6931, new_n6930, new_n6929);
not_3  g04583(new_n6932, new_n6931);
not_3  g04584(new_n6933, new_n6930);
nor_4  g04585(new_n6934, new_n6933, new_n6928);
nor_4  g04586(new_n6935, new_n6934, new_n6931);
xor_3  g04587(new_n6936, new_n6871, n20409);
xnor_3 g04588(new_n6937, new_n6919, new_n6883);
not_3  g04589(new_n6938, new_n6937);
nor_4  g04590(new_n6939, new_n6938, new_n6936);
not_3  g04591(new_n6940, new_n6936);
nor_4  g04592(new_n6941, new_n6937, new_n6940);
nor_4  g04593(new_n6942, new_n6941, new_n6939);
xor_3  g04594(new_n6943, new_n6869, n25749);
not_3  g04595(new_n6944, new_n6943);
xnor_3 g04596(new_n6945, new_n6917, new_n6887);
nand_4 g04597(new_n6946, new_n6945, new_n6944);
not_3  g04598(new_n6947, new_n6945);
nor_4  g04599(new_n6948, new_n6947, new_n6943);
nor_4  g04600(new_n6949, new_n6945, new_n6944);
nor_4  g04601(new_n6950, new_n6949, new_n6948);
xor_3  g04602(new_n6951, new_n6867_1, new_n4136);
xnor_3 g04603(new_n6952, new_n6915, new_n6890);
nand_4 g04604(new_n6953, new_n6952, new_n6951);
xor_3  g04605(new_n6954, new_n6867_1, n3161);
not_3  g04606(new_n6955, new_n6952);
nor_4  g04607(new_n6956, new_n6955, new_n6954);
nor_4  g04608(new_n6957, new_n6952, new_n6951);
nor_4  g04609(new_n6958, new_n6957, new_n6956);
xnor_3 g04610(new_n6959, new_n6866, new_n4141);
xnor_3 g04611(new_n6960, new_n6913, new_n6893);
nand_4 g04612(new_n6961, new_n6960, new_n6959);
not_3  g04613(new_n6962, new_n6959);
not_3  g04614(new_n6963, new_n6960);
nor_4  g04615(new_n6964, new_n6963, new_n6962);
nor_4  g04616(new_n6965_1, new_n6960, new_n6959);
nor_4  g04617(new_n6966, new_n6965_1, new_n6964);
nand_4 g04618(new_n6967_1, new_n6865, n4957);
not_3  g04619(new_n6968, new_n6967_1);
nor_4  g04620(new_n6969, new_n6968, new_n6866);
not_3  g04621(new_n6970, new_n6969);
xnor_3 g04622(new_n6971_1, new_n6911, new_n6896);
nand_4 g04623(new_n6972, new_n6971_1, new_n6970);
not_3  g04624(new_n6973, new_n6911);
xnor_3 g04625(new_n6974, new_n6973, new_n6896);
nor_4  g04626(new_n6975_1, new_n6974, new_n6969);
nor_4  g04627(new_n6976, new_n6971_1, new_n6970);
nor_4  g04628(new_n6977, new_n6976, new_n6975_1);
not_3  g04629(new_n6978, new_n6865);
nor_4  g04630(new_n6979, new_n6864, new_n4155);
nor_4  g04631(new_n6980, new_n6979, new_n6978);
not_3  g04632(new_n6981, new_n6980);
xnor_3 g04633(new_n6982, new_n6909, new_n6901);
nor_4  g04634(new_n6983_1, new_n6982, new_n6981);
xnor_3 g04635(new_n6984, new_n6982, new_n6981);
xnor_3 g04636(new_n6985_1, n21993, n14575);
nor_4  g04637(new_n6986, new_n6985_1, n20658);
nand_4 g04638(new_n6987, new_n6986, new_n4162);
not_3  g04639(new_n6988, new_n6987);
not_3  g04640(new_n6989, new_n6904);
nand_4 g04641(new_n6990, new_n6905, new_n6903);
nor_4  g04642(new_n6991, new_n6990, new_n6989);
nor_4  g04643(new_n6992, new_n6907, new_n6904);
nor_4  g04644(new_n6993, new_n6992, new_n6991);
not_3  g04645(new_n6994, new_n6864);
nand_4 g04646(new_n6995, n20658, n15743);
nand_4 g04647(new_n6996, new_n6995, new_n6994);
nor_4  g04648(new_n6997, new_n6996, new_n6986);
not_3  g04649(new_n6998_1, new_n6997);
nand_4 g04650(new_n6999, new_n6998_1, new_n6987);
nor_4  g04651(new_n7000, new_n6999, new_n6993);
nor_4  g04652(new_n7001, new_n7000, new_n6988);
not_3  g04653(new_n7002, new_n7001);
nor_4  g04654(new_n7003, new_n7002, new_n6984);
nor_4  g04655(new_n7004, new_n7003, new_n6983_1);
nand_4 g04656(new_n7005, new_n7004, new_n6977);
nand_4 g04657(new_n7006, new_n7005, new_n6972);
nand_4 g04658(new_n7007, new_n7006, new_n6966);
nand_4 g04659(new_n7008, new_n7007, new_n6961);
nand_4 g04660(new_n7009, new_n7008, new_n6958);
nand_4 g04661(new_n7010, new_n7009, new_n6953);
nand_4 g04662(new_n7011, new_n7010, new_n6950);
nand_4 g04663(new_n7012, new_n7011, new_n6946);
nand_4 g04664(new_n7013, new_n7012, new_n6942);
not_3  g04665(new_n7014, new_n7013);
nor_4  g04666(new_n7015, new_n7014, new_n6939);
nand_4 g04667(new_n7016, new_n7015, new_n6935);
nand_4 g04668(new_n7017, new_n7016, new_n6932);
nand_4 g04669(new_n7018, new_n7017, new_n6927);
not_3  g04670(new_n7019, new_n7018);
nor_4  g04671(new_n7020, new_n7017, new_n6927);
nor_4  g04672(new_n7021, new_n7020, new_n7019);
not_3  g04673(new_n7022, n8526);
xor_3  g04674(new_n7023, n21784, n3582);
nor_4  g04675(new_n7024, n5521, n2145);
xor_3  g04676(new_n7025, n5521, n2145);
not_3  g04677(new_n7026_1, new_n7025);
nor_4  g04678(new_n7027, n11926, n5031);
xor_3  g04679(new_n7028, n11926, n5031);
not_3  g04680(new_n7029, new_n7028);
not_3  g04681(new_n7030, n11044);
nand_4 g04682(new_n7031, new_n7030, new_n4219);
xor_3  g04683(new_n7032_1, n11044, n4325);
not_3  g04684(new_n7033, n2421);
nand_4 g04685(new_n7034, new_n4231_1, new_n7033);
xor_3  g04686(new_n7035, n5337, n2421);
not_3  g04687(new_n7036, n987);
nand_4 g04688(new_n7037, new_n7036, new_n4238);
xor_3  g04689(new_n7038_1, n987, n626);
not_3  g04690(new_n7039, n20478);
nand_4 g04691(new_n7040, new_n7039, new_n4246);
xor_3  g04692(new_n7041, n20478, n1204);
nor_4  g04693(new_n7042, n26882, n19618);
not_3  g04694(new_n7043, new_n7042);
xor_3  g04695(new_n7044, n26882, n19618);
nor_4  g04696(new_n7045, n22619, n22043);
not_3  g04697(new_n7046, new_n7045);
nand_4 g04698(new_n7047, n12121, n6775);
nand_4 g04699(new_n7048, n22619, n22043);
not_3  g04700(new_n7049, new_n7048);
nor_4  g04701(new_n7050, new_n7049, new_n7045);
nand_4 g04702(new_n7051, new_n7050, new_n7047);
nand_4 g04703(new_n7052, new_n7051, new_n7046);
nand_4 g04704(new_n7053, new_n7052, new_n7044);
nand_4 g04705(new_n7054, new_n7053, new_n7043);
nand_4 g04706(new_n7055, new_n7054, new_n7041);
nand_4 g04707(new_n7056, new_n7055, new_n7040);
nand_4 g04708(new_n7057_1, new_n7056, new_n7038_1);
nand_4 g04709(new_n7058, new_n7057_1, new_n7037);
nand_4 g04710(new_n7059, new_n7058, new_n7035);
nand_4 g04711(new_n7060, new_n7059, new_n7034);
nand_4 g04712(new_n7061, new_n7060, new_n7032_1);
nand_4 g04713(new_n7062, new_n7061, new_n7031);
not_3  g04714(new_n7063, new_n7062);
nor_4  g04715(new_n7064, new_n7063, new_n7029);
nor_4  g04716(new_n7065, new_n7064, new_n7027);
nor_4  g04717(new_n7066, new_n7065, new_n7026_1);
nor_4  g04718(new_n7067, new_n7066, new_n7024);
xnor_3 g04719(new_n7068, new_n7067, new_n7023);
xnor_3 g04720(new_n7069, new_n7068, new_n7022);
not_3  g04721(new_n7070, new_n7069);
not_3  g04722(new_n7071, n2816);
xnor_3 g04723(new_n7072, new_n7065, new_n7025);
nor_4  g04724(new_n7073, new_n7072, new_n7071);
xnor_3 g04725(new_n7074, new_n7072, n2816);
not_3  g04726(new_n7075, new_n7074);
not_3  g04727(new_n7076, n20359);
xnor_3 g04728(new_n7077, new_n7062, new_n7028);
not_3  g04729(new_n7078, new_n7077);
nor_4  g04730(new_n7079_1, new_n7078, new_n7076);
xnor_3 g04731(new_n7080, new_n7077, new_n7076);
xnor_3 g04732(new_n7081, new_n7060, new_n7032_1);
nand_4 g04733(new_n7082, new_n7081, n4409);
not_3  g04734(new_n7083, n4409);
xnor_3 g04735(new_n7084, new_n7081, new_n7083);
xnor_3 g04736(new_n7085, new_n7058, new_n7035);
nand_4 g04737(new_n7086, new_n7085, n3570);
not_3  g04738(new_n7087, n3570);
xnor_3 g04739(new_n7088, new_n7085, new_n7087);
xnor_3 g04740(new_n7089, new_n7056, new_n7038_1);
nand_4 g04741(new_n7090, new_n7089, n13668);
xnor_3 g04742(new_n7091, new_n7089, new_n4744);
xnor_3 g04743(new_n7092, new_n7054, new_n7041);
nand_4 g04744(new_n7093, new_n7092, n21276);
not_3  g04745(new_n7094, new_n7093);
nor_4  g04746(new_n7095, new_n7092, n21276);
nor_4  g04747(new_n7096, new_n7095, new_n7094);
xnor_3 g04748(new_n7097, new_n7052, new_n7044);
nand_4 g04749(new_n7098, new_n7097, n26748);
not_3  g04750(new_n7099_1, new_n7051);
nor_4  g04751(new_n7100, new_n7050, new_n7047);
nor_4  g04752(new_n7101, new_n7100, new_n7099_1);
not_3  g04753(new_n7102, new_n7101);
nor_4  g04754(new_n7103, new_n7102, n10057);
not_3  g04755(new_n7104, n10057);
xnor_3 g04756(new_n7105, new_n7101, new_n7104);
nor_4  g04757(new_n7106, new_n7105, new_n6770);
nor_4  g04758(new_n7107, new_n7106, new_n7103);
not_3  g04759(new_n7108, new_n7098);
nor_4  g04760(new_n7109, new_n7097, n26748);
nor_4  g04761(new_n7110, new_n7109, new_n7108);
nand_4 g04762(new_n7111, new_n7110, new_n7107);
nand_4 g04763(new_n7112, new_n7111, new_n7098);
nand_4 g04764(new_n7113, new_n7112, new_n7096);
nand_4 g04765(new_n7114, new_n7113, new_n7093);
nand_4 g04766(new_n7115, new_n7114, new_n7091);
nand_4 g04767(new_n7116, new_n7115, new_n7090);
nand_4 g04768(new_n7117, new_n7116, new_n7088);
nand_4 g04769(new_n7118, new_n7117, new_n7086);
nand_4 g04770(new_n7119, new_n7118, new_n7084);
nand_4 g04771(new_n7120, new_n7119, new_n7082);
nand_4 g04772(new_n7121, new_n7120, new_n7080);
not_3  g04773(new_n7122, new_n7121);
nor_4  g04774(new_n7123, new_n7122, new_n7079_1);
nor_4  g04775(new_n7124, new_n7123, new_n7075);
nor_4  g04776(new_n7125, new_n7124, new_n7073);
xnor_3 g04777(new_n7126, new_n7125, new_n7070);
xnor_3 g04778(new_n7127, new_n7126, new_n7021);
xnor_3 g04779(new_n7128, new_n7123, new_n7074);
not_3  g04780(new_n7129, new_n7016);
nor_4  g04781(new_n7130, new_n7015, new_n6935);
nor_4  g04782(new_n7131, new_n7130, new_n7129);
nor_4  g04783(new_n7132, new_n7131, new_n7128);
xnor_3 g04784(new_n7133, new_n7131, new_n7128);
xnor_3 g04785(new_n7134, new_n7012, new_n6942);
not_3  g04786(new_n7135, new_n7134);
xnor_3 g04787(new_n7136, new_n7120, new_n7080);
nand_4 g04788(new_n7137, new_n7136, new_n7135);
xnor_3 g04789(new_n7138, new_n7136, new_n7134);
xnor_3 g04790(new_n7139_1, new_n7010, new_n6950);
not_3  g04791(new_n7140, new_n7139_1);
xnor_3 g04792(new_n7141, new_n7118, new_n7084);
nand_4 g04793(new_n7142, new_n7141, new_n7140);
xnor_3 g04794(new_n7143, new_n7141, new_n7139_1);
xnor_3 g04795(new_n7144, new_n7008, new_n6958);
not_3  g04796(new_n7145, new_n7088);
xnor_3 g04797(new_n7146, new_n7116, new_n7145);
nor_4  g04798(new_n7147, new_n7146, new_n7144);
not_3  g04799(new_n7148, new_n7147);
not_3  g04800(new_n7149_1, new_n7144);
xnor_3 g04801(new_n7150, new_n7116, new_n7088);
nor_4  g04802(new_n7151, new_n7150, new_n7149_1);
nor_4  g04803(new_n7152, new_n7151, new_n7147);
not_3  g04804(new_n7153, new_n6966);
xnor_3 g04805(new_n7154, new_n7006, new_n7153);
xnor_3 g04806(new_n7155, new_n7114, new_n7091);
nand_4 g04807(new_n7156, new_n7155, new_n7154);
not_3  g04808(new_n7157, new_n7155);
xnor_3 g04809(new_n7158, new_n7157, new_n7154);
not_3  g04810(new_n7159, new_n6977);
xnor_3 g04811(new_n7160, new_n7004, new_n7159);
xnor_3 g04812(new_n7161, new_n7112, new_n7096);
nand_4 g04813(new_n7162, new_n7161, new_n7160);
not_3  g04814(new_n7163, new_n7162);
nor_4  g04815(new_n7164, new_n7161, new_n7160);
nor_4  g04816(new_n7165, new_n7164, new_n7163);
and_4  g04817(new_n7166, new_n7002, new_n6984);
nor_4  g04818(new_n7167, new_n7166, new_n7003);
not_3  g04819(new_n7168, new_n7167);
xnor_3 g04820(new_n7169, new_n7110, new_n7107);
nand_4 g04821(new_n7170, new_n7169, new_n7168);
xnor_3 g04822(new_n7171, new_n7169, new_n7167);
not_3  g04823(new_n7172, new_n6770);
not_3  g04824(new_n7173, new_n7105);
nor_4  g04825(new_n7174, new_n7173, new_n7172);
nor_4  g04826(new_n7175, new_n7174, new_n7106);
xor_3  g04827(new_n7176, new_n6999, new_n6993);
nor_4  g04828(new_n7177, new_n7176, new_n7175);
xor_3  g04829(new_n7178, new_n6985_1, n20658);
not_3  g04830(new_n7179, new_n7178);
nand_4 g04831(new_n7180, new_n7179, new_n6771);
xnor_3 g04832(new_n7181, new_n7176, new_n7175);
nor_4  g04833(new_n7182, new_n7181, new_n7180);
nor_4  g04834(new_n7183, new_n7182, new_n7177);
nand_4 g04835(new_n7184, new_n7183, new_n7171);
nand_4 g04836(new_n7185, new_n7184, new_n7170);
nand_4 g04837(new_n7186, new_n7185, new_n7165);
nand_4 g04838(new_n7187, new_n7186, new_n7162);
nand_4 g04839(new_n7188, new_n7187, new_n7158);
nand_4 g04840(new_n7189, new_n7188, new_n7156);
nand_4 g04841(new_n7190_1, new_n7189, new_n7152);
nand_4 g04842(new_n7191, new_n7190_1, new_n7148);
nand_4 g04843(new_n7192, new_n7191, new_n7143);
nand_4 g04844(new_n7193, new_n7192, new_n7142);
nand_4 g04845(new_n7194, new_n7193, new_n7138);
nand_4 g04846(new_n7195, new_n7194, new_n7137);
not_3  g04847(new_n7196, new_n7195);
nor_4  g04848(new_n7197, new_n7196, new_n7133);
nor_4  g04849(new_n7198, new_n7197, new_n7132);
xnor_3 g04850(n567, new_n7198, new_n7127);
nor_4  g04851(new_n7200, n10250, n1831);
not_3  g04852(new_n7201, new_n7200);
xor_3  g04853(new_n7202, n10250, n1831);
nor_4  g04854(new_n7203, n13137, n7674);
not_3  g04855(new_n7204, new_n7203);
xor_3  g04856(new_n7205, n13137, n7674);
nor_4  g04857(new_n7206, n18452, n6397);
not_3  g04858(new_n7207, new_n7206);
xor_3  g04859(new_n7208, n18452, n6397);
not_3  g04860(new_n7209, n19196);
not_3  g04861(new_n7210, n21317);
nand_4 g04862(new_n7211, new_n7210, new_n7209);
xor_3  g04863(new_n7212, n21317, n19196);
nor_4  g04864(new_n7213, n23586, n12398);
not_3  g04865(new_n7214, new_n7213);
xor_3  g04866(new_n7215, n23586, n12398);
nor_4  g04867(new_n7216, n21226, n19789);
not_3  g04868(new_n7217, new_n7216);
xor_3  g04869(new_n7218, n21226, n19789);
nor_4  g04870(new_n7219, n20169, n4426);
not_3  g04871(new_n7220, new_n7219);
xor_3  g04872(new_n7221, n20169, n4426);
nor_4  g04873(new_n7222, n20036, n8285);
not_3  g04874(new_n7223, new_n7222);
xnor_3 g04875(new_n7224, n20036, n8285);
not_3  g04876(new_n7225, new_n7224);
nor_4  g04877(new_n7226, n11192, n6729);
not_3  g04878(new_n7227, new_n7226);
nand_4 g04879(new_n7228, n21687, n9380);
xor_3  g04880(new_n7229_1, n11192, n6729);
nand_4 g04881(new_n7230_1, new_n7229_1, new_n7228);
nand_4 g04882(new_n7231, new_n7230_1, new_n7227);
nand_4 g04883(new_n7232, new_n7231, new_n7225);
nand_4 g04884(new_n7233_1, new_n7232, new_n7223);
nand_4 g04885(new_n7234, new_n7233_1, new_n7221);
nand_4 g04886(new_n7235, new_n7234, new_n7220);
nand_4 g04887(new_n7236_1, new_n7235, new_n7218);
nand_4 g04888(new_n7237, new_n7236_1, new_n7217);
nand_4 g04889(new_n7238, new_n7237, new_n7215);
nand_4 g04890(new_n7239, new_n7238, new_n7214);
nand_4 g04891(new_n7240, new_n7239, new_n7212);
nand_4 g04892(new_n7241, new_n7240, new_n7211);
nand_4 g04893(new_n7242, new_n7241, new_n7208);
nand_4 g04894(new_n7243, new_n7242, new_n7207);
nand_4 g04895(new_n7244, new_n7243, new_n7205);
nand_4 g04896(new_n7245, new_n7244, new_n7204);
nand_4 g04897(new_n7246, new_n7245, new_n7202);
nand_4 g04898(new_n7247, new_n7246, new_n7201);
not_3  g04899(new_n7248, new_n7247);
not_3  g04900(new_n7249, n1752);
not_3  g04901(new_n7250, n13110);
nand_4 g04902(new_n7251, new_n4442, new_n7250);
not_3  g04903(new_n7252, new_n7251);
nand_4 g04904(new_n7253_1, new_n7252, new_n7249);
nor_4  g04905(new_n7254, new_n7253_1, n1288);
xor_3  g04906(new_n7255, new_n7254, n3320);
nor_4  g04907(new_n7256_1, new_n7255, new_n6321);
not_3  g04908(new_n7257, new_n7254);
nor_4  g04909(new_n7258, new_n7257, n3320);
not_3  g04910(new_n7259, new_n7258);
not_3  g04911(new_n7260, new_n7255);
nor_4  g04912(new_n7261, new_n7260, n8614);
not_3  g04913(new_n7262, new_n7261);
xor_3  g04914(new_n7263, new_n7253_1, n1288);
nor_4  g04915(new_n7264, new_n7263, n15182);
not_3  g04916(new_n7265, n1288);
xor_3  g04917(new_n7266, new_n7253_1, new_n7265);
nor_4  g04918(new_n7267, new_n7266, new_n6326);
nor_4  g04919(new_n7268_1, new_n7267, new_n7264);
not_3  g04920(new_n7269, new_n7268_1);
xor_3  g04921(new_n7270, new_n7252, new_n7249);
nor_4  g04922(new_n7271, new_n7270, n27037);
xnor_3 g04923(new_n7272, new_n7270, n27037);
xor_3  g04924(new_n7273, new_n4442, n13110);
nor_4  g04925(new_n7274, new_n7273, new_n6332);
not_3  g04926(new_n7275, new_n7274);
xor_3  g04927(new_n7276, new_n4442, new_n7250);
nor_4  g04928(new_n7277_1, new_n7276, n8964);
nor_4  g04929(new_n7278, new_n7277_1, new_n7274);
not_3  g04930(new_n7279, n20151);
not_3  g04931(new_n7280_1, new_n4445);
nor_4  g04932(new_n7281, new_n7280_1, new_n7279);
not_3  g04933(new_n7282, new_n7281);
nand_4 g04934(new_n7283, new_n4489, new_n4446);
nand_4 g04935(new_n7284, new_n7283, new_n7282);
nand_4 g04936(new_n7285, new_n7284, new_n7278);
nand_4 g04937(new_n7286, new_n7285, new_n7275);
nor_4  g04938(new_n7287, new_n7286, new_n7272);
nor_4  g04939(new_n7288, new_n7287, new_n7271);
nor_4  g04940(new_n7289, new_n7288, new_n7269);
nor_4  g04941(new_n7290, new_n7289, new_n7264);
nand_4 g04942(new_n7291, new_n7290, new_n7262);
nand_4 g04943(new_n7292, new_n7291, new_n7259);
nor_4  g04944(new_n7293, new_n7292, new_n7256_1);
nor_4  g04945(new_n7294, new_n7293, new_n7248);
not_3  g04946(new_n7295, new_n7293);
nor_4  g04947(new_n7296, new_n7295, new_n7247);
nor_4  g04948(new_n7297, new_n7296, new_n7294);
not_3  g04949(new_n7298_1, new_n7297);
not_3  g04950(new_n7299, new_n7202);
not_3  g04951(new_n7300, new_n7205);
not_3  g04952(new_n7301, new_n7208);
not_3  g04953(new_n7302, new_n7241);
nor_4  g04954(new_n7303, new_n7302, new_n7301);
nor_4  g04955(new_n7304, new_n7303, new_n7206);
nor_4  g04956(new_n7305_1, new_n7304, new_n7300);
nor_4  g04957(new_n7306, new_n7305_1, new_n7203);
xor_3  g04958(new_n7307, new_n7306, new_n7299);
not_3  g04959(new_n7308_1, new_n7307);
nor_4  g04960(new_n7309, new_n7261, new_n7256_1);
xnor_3 g04961(new_n7310, new_n7309, new_n7290);
not_3  g04962(new_n7311, new_n7310);
nor_4  g04963(new_n7312, new_n7311, new_n7308_1);
xnor_3 g04964(new_n7313_1, new_n7288, new_n7269);
xor_3  g04965(new_n7314, new_n7304, new_n7205);
nor_4  g04966(new_n7315, new_n7314, new_n7313_1);
xnor_3 g04967(new_n7316, new_n7314, new_n7313_1);
xnor_3 g04968(new_n7317, new_n7286, new_n7272);
xnor_3 g04969(new_n7318, new_n7241, new_n7208);
nor_4  g04970(new_n7319, new_n7318, new_n7317);
not_3  g04971(new_n7320, new_n7272);
not_3  g04972(new_n7321, new_n7286);
nor_4  g04973(new_n7322, new_n7321, new_n7320);
nor_4  g04974(new_n7323, new_n7322, new_n7287);
xnor_3 g04975(new_n7324, new_n7318, new_n7323);
not_3  g04976(new_n7325, new_n7212);
xnor_3 g04977(new_n7326, new_n7239, new_n7325);
xnor_3 g04978(new_n7327, new_n7284, new_n7278);
nand_4 g04979(new_n7328, new_n7327, new_n7326);
not_3  g04980(new_n7329, new_n7215);
xnor_3 g04981(new_n7330_1, new_n7237, new_n7329);
nand_4 g04982(new_n7331, new_n7330_1, new_n4490);
xnor_3 g04983(new_n7332, new_n7237, new_n7215);
xnor_3 g04984(new_n7333, new_n7332, new_n4490);
not_3  g04985(new_n7334, new_n7218);
xnor_3 g04986(new_n7335_1, new_n7235, new_n7334);
not_3  g04987(new_n7336, new_n7221);
not_3  g04988(new_n7337, new_n7228);
xnor_3 g04989(new_n7338, n11192, n6729);
nor_4  g04990(new_n7339_1, new_n7338, new_n7337);
nor_4  g04991(new_n7340, new_n7339_1, new_n7226);
nor_4  g04992(new_n7341, new_n7340, new_n7224);
nor_4  g04993(new_n7342, new_n7341, new_n7222);
xnor_3 g04994(new_n7343, new_n7342, new_n7336);
nor_4  g04995(new_n7344, new_n7343, new_n4506);
xnor_3 g04996(new_n7345, new_n7340, new_n7224);
not_3  g04997(new_n7346_1, new_n7345);
nor_4  g04998(new_n7347, new_n7346_1, new_n4514_1);
not_3  g04999(new_n7348, new_n7347);
nor_4  g05000(new_n7349_1, new_n7345, new_n4513);
nor_4  g05001(new_n7350, new_n7349_1, new_n7347);
xnor_3 g05002(new_n7351, new_n7338, new_n7228);
nor_4  g05003(new_n7352, new_n7351, new_n4526);
not_3  g05004(new_n7353, new_n7352);
xor_3  g05005(new_n7354, n21687, n9380);
not_3  g05006(new_n7355, new_n7354);
nor_4  g05007(new_n7356, new_n7355, new_n2603);
not_3  g05008(new_n7357, new_n7351);
nor_4  g05009(new_n7358, new_n7357, new_n4525);
nor_4  g05010(new_n7359, new_n7358, new_n7352);
nand_4 g05011(new_n7360, new_n7359, new_n7356);
nand_4 g05012(new_n7361, new_n7360, new_n7353);
nand_4 g05013(new_n7362, new_n7361, new_n7350);
nand_4 g05014(new_n7363_1, new_n7362, new_n7348);
xnor_3 g05015(new_n7364, new_n7343, new_n4506);
nor_4  g05016(new_n7365, new_n7364, new_n7363_1);
nor_4  g05017(new_n7366, new_n7365, new_n7344);
not_3  g05018(new_n7367, new_n7366);
nand_4 g05019(new_n7368, new_n7367, new_n7335_1);
xnor_3 g05020(new_n7369, new_n7366, new_n7335_1);
nand_4 g05021(new_n7370, new_n7369, new_n4497);
nand_4 g05022(new_n7371, new_n7370, new_n7368);
nand_4 g05023(new_n7372, new_n7371, new_n7333);
nand_4 g05024(new_n7373, new_n7372, new_n7331);
xnor_3 g05025(new_n7374, new_n7239, new_n7212);
xnor_3 g05026(new_n7375, new_n7327, new_n7374);
nand_4 g05027(new_n7376, new_n7375, new_n7373);
nand_4 g05028(new_n7377_1, new_n7376, new_n7328);
nand_4 g05029(new_n7378, new_n7377_1, new_n7324);
not_3  g05030(new_n7379, new_n7378);
nor_4  g05031(new_n7380, new_n7379, new_n7319);
nor_4  g05032(new_n7381, new_n7380, new_n7316);
nor_4  g05033(new_n7382, new_n7381, new_n7315);
xnor_3 g05034(new_n7383, new_n7310, new_n7307);
nor_4  g05035(new_n7384, new_n7383, new_n7382);
nor_4  g05036(new_n7385, new_n7384, new_n7312);
nor_4  g05037(new_n7386, new_n7385, new_n7298_1);
nor_4  g05038(new_n7387, new_n7386, new_n7294);
xnor_3 g05039(new_n7388, new_n7385, new_n7297);
not_3  g05040(new_n7389, new_n7388);
nor_4  g05041(new_n7390_1, n15766, n6105);
xor_3  g05042(new_n7391, n15766, n6105);
not_3  g05043(new_n7392, new_n7391);
not_3  g05044(new_n7393, n3795);
not_3  g05045(new_n7394, n25629);
nand_4 g05046(new_n7395, new_n7394, new_n7393);
xor_3  g05047(new_n7396, n25629, n3795);
nor_4  g05048(new_n7397, n25464, n7692);
not_3  g05049(new_n7398, new_n7397);
xor_3  g05050(new_n7399, n25464, n7692);
nor_4  g05051(new_n7400, n23039, n4590);
not_3  g05052(new_n7401, new_n7400);
xor_3  g05053(new_n7402, n23039, n4590);
nor_4  g05054(new_n7403_1, n26752, n13677);
not_3  g05055(new_n7404, new_n7403_1);
xor_3  g05056(new_n7405, n26752, n13677);
nor_4  g05057(new_n7406, n18926, n6513);
not_3  g05058(new_n7407, new_n7406);
xor_3  g05059(new_n7408_1, n18926, n6513);
nand_4 g05060(new_n7409, n5451, n3918);
not_3  g05061(new_n7410, new_n7409);
nor_4  g05062(new_n7411, n5451, n3918);
nor_4  g05063(new_n7412, n5330, n919);
not_3  g05064(new_n7413, new_n7412);
nand_4 g05065(new_n7414, new_n4649, new_n7413);
nor_4  g05066(new_n7415, new_n7414, new_n7411);
nor_4  g05067(new_n7416, new_n7415, new_n7410);
nand_4 g05068(new_n7417, new_n7416, new_n7408_1);
nand_4 g05069(new_n7418, new_n7417, new_n7407);
nand_4 g05070(new_n7419, new_n7418, new_n7405);
nand_4 g05071(new_n7420, new_n7419, new_n7404);
nand_4 g05072(new_n7421_1, new_n7420, new_n7402);
nand_4 g05073(new_n7422, new_n7421_1, new_n7401);
nand_4 g05074(new_n7423, new_n7422, new_n7399);
nand_4 g05075(new_n7424, new_n7423, new_n7398);
nand_4 g05076(new_n7425, new_n7424, new_n7396);
nand_4 g05077(new_n7426, new_n7425, new_n7395);
not_3  g05078(new_n7427, new_n7426);
nor_4  g05079(new_n7428_1, new_n7427, new_n7392);
nor_4  g05080(new_n7429, new_n7428_1, new_n7390_1);
not_3  g05081(new_n7430, new_n7429);
nor_4  g05082(new_n7431, new_n7430, new_n7389);
xnor_3 g05083(new_n7432_1, new_n7429, new_n7388);
xor_3  g05084(new_n7433, new_n7427, new_n7392);
xnor_3 g05085(new_n7434, new_n7383, new_n7382);
nor_4  g05086(new_n7435, new_n7434, new_n7433);
xnor_3 g05087(new_n7436, new_n7434, new_n7433);
xnor_3 g05088(new_n7437_1, new_n7380, new_n7316);
not_3  g05089(new_n7438, new_n7424);
xor_3  g05090(new_n7439, new_n7438, new_n7396);
not_3  g05091(new_n7440, new_n7439);
nor_4  g05092(new_n7441, new_n7440, new_n7437_1);
xnor_3 g05093(new_n7442, new_n7440, new_n7437_1);
xnor_3 g05094(new_n7443, new_n7377_1, new_n7324);
not_3  g05095(new_n7444, new_n7443);
not_3  g05096(new_n7445, new_n7422);
xor_3  g05097(new_n7446, new_n7445, new_n7399);
nand_4 g05098(new_n7447, new_n7446, new_n7444);
xnor_3 g05099(new_n7448, new_n7446, new_n7443);
not_3  g05100(new_n7449, new_n7402);
not_3  g05101(new_n7450, new_n7420);
xor_3  g05102(new_n7451, new_n7450, new_n7449);
not_3  g05103(new_n7452, new_n7451);
xnor_3 g05104(new_n7453, new_n7375, new_n7373);
not_3  g05105(new_n7454, new_n7453);
nand_4 g05106(new_n7455, new_n7454, new_n7452);
xnor_3 g05107(new_n7456, new_n7453, new_n7452);
xnor_3 g05108(new_n7457, new_n7371, new_n7333);
not_3  g05109(new_n7458, new_n7457);
not_3  g05110(new_n7459, new_n7418);
xor_3  g05111(new_n7460_1, new_n7459, new_n7405);
nand_4 g05112(new_n7461, new_n7460_1, new_n7458);
xnor_3 g05113(new_n7462, new_n7460_1, new_n7457);
xnor_3 g05114(new_n7463, new_n7369, new_n4497);
not_3  g05115(new_n7464, new_n7463);
not_3  g05116(new_n7465, new_n7416);
xor_3  g05117(new_n7466, new_n7465, new_n7408_1);
nand_4 g05118(new_n7467, new_n7466, new_n7464);
xnor_3 g05119(new_n7468, new_n7466, new_n7463);
not_3  g05120(new_n7469, new_n7363_1);
not_3  g05121(new_n7470, new_n7364);
nor_4  g05122(new_n7471, new_n7470, new_n7469);
nor_4  g05123(new_n7472, new_n7471, new_n7365);
not_3  g05124(new_n7473, new_n7414);
nor_4  g05125(new_n7474, new_n7411, new_n7410);
xor_3  g05126(new_n7475_1, new_n7474, new_n7473);
nand_4 g05127(new_n7476, new_n7475_1, new_n7472);
not_3  g05128(new_n7477_1, new_n7475_1);
xnor_3 g05129(new_n7478, new_n7477_1, new_n7472);
not_3  g05130(new_n7479, new_n7362);
nor_4  g05131(new_n7480, new_n7361, new_n7350);
nor_4  g05132(new_n7481, new_n7480, new_n7479);
nor_4  g05133(new_n7482, new_n7481, new_n4651);
not_3  g05134(new_n7483, new_n7482);
not_3  g05135(new_n7484, new_n4651);
not_3  g05136(new_n7485, new_n7481);
nor_4  g05137(new_n7486, new_n7485, new_n7484);
nor_4  g05138(new_n7487, new_n7486, new_n7482);
not_3  g05139(new_n7488, new_n4655);
xnor_3 g05140(new_n7489, new_n7359, new_n7356);
not_3  g05141(new_n7490, new_n7489);
nor_4  g05142(new_n7491, new_n7490, new_n7488);
not_3  g05143(new_n7492, new_n7491);
xor_3  g05144(new_n7493, new_n7355, new_n2603);
nor_4  g05145(new_n7494, new_n7493, new_n4658);
nor_4  g05146(new_n7495, new_n7489, new_n4655);
nor_4  g05147(new_n7496, new_n7495, new_n7491);
nand_4 g05148(new_n7497, new_n7496, new_n7494);
nand_4 g05149(new_n7498, new_n7497, new_n7492);
nand_4 g05150(new_n7499, new_n7498, new_n7487);
nand_4 g05151(new_n7500, new_n7499, new_n7483);
nand_4 g05152(new_n7501, new_n7500, new_n7478);
nand_4 g05153(new_n7502, new_n7501, new_n7476);
nand_4 g05154(new_n7503, new_n7502, new_n7468);
nand_4 g05155(new_n7504, new_n7503, new_n7467);
nand_4 g05156(new_n7505, new_n7504, new_n7462);
nand_4 g05157(new_n7506, new_n7505, new_n7461);
nand_4 g05158(new_n7507_1, new_n7506, new_n7456);
nand_4 g05159(new_n7508, new_n7507_1, new_n7455);
nand_4 g05160(new_n7509, new_n7508, new_n7448);
nand_4 g05161(new_n7510, new_n7509, new_n7447);
not_3  g05162(new_n7511, new_n7510);
nor_4  g05163(new_n7512, new_n7511, new_n7442);
nor_4  g05164(new_n7513, new_n7512, new_n7441);
nor_4  g05165(new_n7514_1, new_n7513, new_n7436);
nor_4  g05166(new_n7515, new_n7514_1, new_n7435);
nor_4  g05167(new_n7516, new_n7515, new_n7432_1);
nor_4  g05168(new_n7517, new_n7516, new_n7431);
nor_4  g05169(n588, new_n7517, new_n7387);
not_3  g05170(new_n7519, n19803);
xor_3  g05171(new_n7520, new_n7519, n18584);
nand_4 g05172(new_n7521, n12626, new_n5287);
nand_4 g05173(new_n7522, new_n5315, new_n5288);
nand_4 g05174(new_n7523, new_n7522, new_n7521);
xnor_3 g05175(new_n7524_1, new_n7523, new_n7520);
not_3  g05176(new_n7525, n7773);
xor_3  g05177(new_n7526, n16911, new_n7525);
not_3  g05178(new_n7527, n7721);
nand_4 g05179(new_n7528, new_n7527, n376);
not_3  g05180(new_n7529, n376);
xor_3  g05181(new_n7530, n7721, new_n7529);
not_3  g05182(new_n7531, n5517);
nor_4  g05183(new_n7532, n21981, new_n7531);
not_3  g05184(new_n7533, new_n7532);
xor_3  g05185(new_n7534, n21981, new_n7531);
not_3  g05186(new_n7535, n12113);
nor_4  g05187(new_n7536, n12917, new_n7535);
not_3  g05188(new_n7537, new_n7536);
xor_3  g05189(new_n7538, n12917, new_n7535);
not_3  g05190(new_n7539, n21898);
nor_4  g05191(new_n7540, new_n7539, n10614);
not_3  g05192(new_n7541, n10614);
nor_4  g05193(new_n7542, n21898, new_n7541);
not_3  g05194(new_n7543, n9926);
nor_4  g05195(new_n7544, n11266, new_n7543);
not_3  g05196(new_n7545, n11266);
nor_4  g05197(new_n7546, new_n7545, n9926);
not_3  g05198(new_n7547, n22072);
nor_4  g05199(new_n7548, new_n7547, n2646);
not_3  g05200(new_n7549, new_n7548);
nor_4  g05201(new_n7550, new_n7549, new_n7546);
nor_4  g05202(new_n7551, new_n7550, new_n7544);
nor_4  g05203(new_n7552, new_n7551, new_n7542);
nor_4  g05204(new_n7553, new_n7552, new_n7540);
nand_4 g05205(new_n7554, new_n7553, new_n7538);
nand_4 g05206(new_n7555, new_n7554, new_n7537);
nand_4 g05207(new_n7556, new_n7555, new_n7534);
nand_4 g05208(new_n7557, new_n7556, new_n7533);
nand_4 g05209(new_n7558_1, new_n7557, new_n7530);
nand_4 g05210(new_n7559, new_n7558_1, new_n7528);
xnor_3 g05211(new_n7560, new_n7559, new_n7526);
not_3  g05212(new_n7561, n16818);
not_3  g05213(new_n7562, n14576);
not_3  g05214(new_n7563, n5605);
nor_4  g05215(new_n7564, n15652, n4939);
nand_4 g05216(new_n7565, new_n7564, new_n7563);
nor_4  g05217(new_n7566_1, new_n7565, n2985);
nand_4 g05218(new_n7567, new_n7566_1, new_n7562);
nor_4  g05219(new_n7568, new_n7567, n1269);
xor_3  g05220(new_n7569_1, new_n7568, new_n7561);
nand_4 g05221(new_n7570, new_n7569_1, n1742);
not_3  g05222(new_n7571, new_n7570);
nor_4  g05223(new_n7572_1, new_n7569_1, n1742);
nor_4  g05224(new_n7573, new_n7572_1, new_n7571);
nand_4 g05225(new_n7574, new_n7567, n1269);
not_3  g05226(new_n7575_1, new_n7574);
nor_4  g05227(new_n7576, new_n7575_1, new_n7568);
nor_4  g05228(new_n7577, new_n7576, n4858);
not_3  g05229(new_n7578, new_n7577);
not_3  g05230(new_n7579, n4858);
not_3  g05231(new_n7580, new_n7576);
nor_4  g05232(new_n7581, new_n7580, new_n7579);
not_3  g05233(new_n7582, new_n7581);
not_3  g05234(new_n7583, n8244);
xnor_3 g05235(new_n7584, new_n7566_1, new_n7562);
nor_4  g05236(new_n7585_1, new_n7584, new_n7583);
not_3  g05237(new_n7586, new_n7584);
nor_4  g05238(new_n7587, new_n7586, n8244);
nor_4  g05239(new_n7588_1, new_n7587, new_n7585_1);
not_3  g05240(new_n7589, new_n7588_1);
nand_4 g05241(new_n7590, new_n7565, n2985);
not_3  g05242(new_n7591, new_n7590);
nor_4  g05243(new_n7592, new_n7591, new_n7566_1);
nor_4  g05244(new_n7593_1, new_n7592, n9493);
not_3  g05245(new_n7594, new_n7593_1);
xnor_3 g05246(new_n7595, new_n7564, new_n7563);
not_3  g05247(new_n7596, new_n7595);
nor_4  g05248(new_n7597, new_n7596, n15167);
not_3  g05249(new_n7598_1, new_n7597);
not_3  g05250(new_n7599, n15167);
nor_4  g05251(new_n7600, new_n7595, new_n7599);
nor_4  g05252(new_n7601, new_n7600, new_n7597);
not_3  g05253(new_n7602, n21095);
xnor_3 g05254(new_n7603, n15652, n4939);
nand_4 g05255(new_n7604, new_n7603, new_n7602);
nand_4 g05256(new_n7605, n8656, n4939);
not_3  g05257(new_n7606, new_n7603);
nor_4  g05258(new_n7607_1, new_n7606, n21095);
nor_4  g05259(new_n7608, new_n7603, new_n7602);
nor_4  g05260(new_n7609, new_n7608, new_n7607_1);
nand_4 g05261(new_n7610_1, new_n7609, new_n7605);
nand_4 g05262(new_n7611, new_n7610_1, new_n7604);
nand_4 g05263(new_n7612, new_n7611, new_n7601);
nand_4 g05264(new_n7613, new_n7612, new_n7598_1);
not_3  g05265(new_n7614, n9493);
not_3  g05266(new_n7615, new_n7592);
nor_4  g05267(new_n7616_1, new_n7615, new_n7614);
nor_4  g05268(new_n7617, new_n7616_1, new_n7593_1);
nand_4 g05269(new_n7618, new_n7617, new_n7613);
nand_4 g05270(new_n7619, new_n7618, new_n7594);
nor_4  g05271(new_n7620, new_n7619, new_n7589);
nor_4  g05272(new_n7621, new_n7620, new_n7585_1);
nand_4 g05273(new_n7622, new_n7621, new_n7582);
nand_4 g05274(new_n7623, new_n7622, new_n7578);
xnor_3 g05275(new_n7624, new_n7623, new_n7573);
xnor_3 g05276(new_n7625, new_n7624, new_n7560);
xnor_3 g05277(new_n7626, new_n7557, new_n7530);
not_3  g05278(new_n7627, new_n7626);
nor_4  g05279(new_n7628, new_n7581, new_n7577);
not_3  g05280(new_n7629, new_n7628);
xnor_3 g05281(new_n7630_1, new_n7629, new_n7621);
not_3  g05282(new_n7631, new_n7630_1);
nand_4 g05283(new_n7632, new_n7631, new_n7627);
not_3  g05284(new_n7633, new_n7632);
nor_4  g05285(new_n7634, new_n7631, new_n7627);
nor_4  g05286(new_n7635, new_n7634, new_n7633);
xnor_3 g05287(new_n7636, new_n7555, new_n7534);
not_3  g05288(new_n7637, new_n7636);
nand_4 g05289(new_n7638, new_n7619, new_n7589);
not_3  g05290(new_n7639, new_n7638);
nor_4  g05291(new_n7640, new_n7639, new_n7620);
nor_4  g05292(new_n7641, new_n7640, new_n7637);
not_3  g05293(new_n7642, new_n7640);
nor_4  g05294(new_n7643_1, new_n7642, new_n7636);
nor_4  g05295(new_n7644, new_n7643_1, new_n7641);
not_3  g05296(new_n7645, new_n7644);
not_3  g05297(new_n7646, new_n7538);
xnor_3 g05298(new_n7647_1, new_n7553, new_n7646);
xnor_3 g05299(new_n7648, new_n7617, new_n7613);
nand_4 g05300(new_n7649, new_n7648, new_n7647_1);
xnor_3 g05301(new_n7650, new_n7611, new_n7601);
not_3  g05302(new_n7651, new_n7551);
nor_4  g05303(new_n7652, new_n7542, new_n7540);
xnor_3 g05304(new_n7653, new_n7652, new_n7651);
nor_4  g05305(new_n7654, new_n7653, new_n7650);
xnor_3 g05306(new_n7655, new_n7653, new_n7650);
not_3  g05307(new_n7656, new_n7605);
nor_4  g05308(new_n7657_1, n8656, n4939);
nor_4  g05309(new_n7658, new_n7657_1, new_n7656);
not_3  g05310(new_n7659, new_n7658);
not_3  g05311(new_n7660, n2646);
nor_4  g05312(new_n7661, n22072, new_n7660);
nor_4  g05313(new_n7662, new_n7661, new_n7548);
nor_4  g05314(new_n7663, new_n7662, new_n7659);
nor_4  g05315(new_n7664, new_n7546, new_n7544);
xnor_3 g05316(new_n7665, new_n7664, new_n7548);
nor_4  g05317(new_n7666, new_n7665, new_n7663);
xnor_3 g05318(new_n7667, new_n7609, new_n7605);
xnor_3 g05319(new_n7668, new_n7665, new_n7663);
nor_4  g05320(new_n7669, new_n7668, new_n7667);
nor_4  g05321(new_n7670_1, new_n7669, new_n7666);
nor_4  g05322(new_n7671, new_n7670_1, new_n7655);
nor_4  g05323(new_n7672, new_n7671, new_n7654);
not_3  g05324(new_n7673, new_n7649);
nor_4  g05325(new_n7674_1, new_n7648, new_n7647_1);
nor_4  g05326(new_n7675, new_n7674_1, new_n7673);
nand_4 g05327(new_n7676, new_n7675, new_n7672);
nand_4 g05328(new_n7677, new_n7676, new_n7649);
nor_4  g05329(new_n7678_1, new_n7677, new_n7645);
nor_4  g05330(new_n7679_1, new_n7678_1, new_n7641);
nand_4 g05331(new_n7680, new_n7679_1, new_n7635);
nand_4 g05332(new_n7681, new_n7680, new_n7632);
xnor_3 g05333(new_n7682, new_n7681, new_n7625);
xnor_3 g05334(new_n7683, new_n7682, new_n7524_1);
not_3  g05335(new_n7684, new_n7680);
nor_4  g05336(new_n7685, new_n7679_1, new_n7635);
nor_4  g05337(new_n7686_1, new_n7685, new_n7684);
nor_4  g05338(new_n7687, new_n7686_1, new_n5317);
not_3  g05339(new_n7688, new_n7687);
not_3  g05340(new_n7689, new_n7686_1);
nor_4  g05341(new_n7690, new_n7689, new_n5318);
nor_4  g05342(new_n7691, new_n7690, new_n7687);
not_3  g05343(new_n7692_1, new_n7677);
nor_4  g05344(new_n7693_1, new_n7692_1, new_n7644);
nor_4  g05345(new_n7694, new_n7693_1, new_n7678_1);
nand_4 g05346(new_n7695, new_n7694, new_n5324);
xnor_3 g05347(new_n7696, new_n7694, new_n5328);
not_3  g05348(new_n7697, new_n7676);
nor_4  g05349(new_n7698_1, new_n7675, new_n7672);
nor_4  g05350(new_n7699, new_n7698_1, new_n7697);
nor_4  g05351(new_n7700, new_n7699, new_n5336);
not_3  g05352(new_n7701, new_n7700);
not_3  g05353(new_n7702, new_n7699);
nor_4  g05354(new_n7703, new_n7702, new_n5335);
nor_4  g05355(new_n7704, new_n7703, new_n7700);
xnor_3 g05356(new_n7705, new_n7670_1, new_n7655);
nor_4  g05357(new_n7706, new_n7705, new_n5344);
not_3  g05358(new_n7707, new_n7706);
not_3  g05359(new_n7708_1, new_n7705);
nor_4  g05360(new_n7709, new_n7708_1, new_n5343);
nor_4  g05361(new_n7710, new_n7709, new_n7706);
xor_3  g05362(new_n7711, new_n7662, new_n7658);
nor_4  g05363(new_n7712, new_n7711, new_n5358);
nor_4  g05364(new_n7713, new_n7712, new_n5361);
not_3  g05365(new_n7714, new_n7713);
xor_3  g05366(new_n7715, new_n7668, new_n7667);
not_3  g05367(new_n7716, new_n7712);
xor_3  g05368(new_n7717, new_n7716, new_n5353_1);
nand_4 g05369(new_n7718, new_n7717, new_n7715);
nand_4 g05370(new_n7719, new_n7718, new_n7714);
nand_4 g05371(new_n7720, new_n7719, new_n7710);
nand_4 g05372(new_n7721_1, new_n7720, new_n7707);
nand_4 g05373(new_n7722, new_n7721_1, new_n7704);
nand_4 g05374(new_n7723, new_n7722, new_n7701);
nand_4 g05375(new_n7724, new_n7723, new_n7696);
nand_4 g05376(new_n7725, new_n7724, new_n7695);
nand_4 g05377(new_n7726, new_n7725, new_n7691);
nand_4 g05378(new_n7727, new_n7726, new_n7688);
xor_3  g05379(n597, new_n7727, new_n7683);
not_3  g05380(new_n7729, n14230);
xnor_3 g05381(new_n7730, n25926, n9646);
xor_3  g05382(new_n7731_1, new_n7730, new_n7729);
xor_3  g05383(n637, new_n7731_1, new_n6781);
not_3  g05384(new_n7733, n7421);
xor_3  g05385(new_n7734, n25797, n10611);
nor_4  g05386(new_n7735, n15967, n2783);
xnor_3 g05387(new_n7736, n15967, n2783);
nor_4  g05388(new_n7737, n15490, n13319);
nand_4 g05389(new_n7738, n25435, n18);
not_3  g05390(new_n7739, new_n7738);
xnor_3 g05391(new_n7740, n15490, n13319);
nor_4  g05392(new_n7741, new_n7740, new_n7739);
nor_4  g05393(new_n7742, new_n7741, new_n7737);
nor_4  g05394(new_n7743, new_n7742, new_n7736);
nor_4  g05395(new_n7744, new_n7743, new_n7735);
not_3  g05396(new_n7745, new_n7744);
nor_4  g05397(new_n7746, new_n7745, new_n7734);
nand_4 g05398(new_n7747, new_n7745, new_n7734);
not_3  g05399(new_n7748, new_n7747);
nor_4  g05400(new_n7749, new_n7748, new_n7746);
xnor_3 g05401(new_n7750, new_n7749, new_n7733);
not_3  g05402(new_n7751_1, n19680);
not_3  g05403(new_n7752, new_n7736);
not_3  g05404(new_n7753, new_n7742);
nor_4  g05405(new_n7754, new_n7753, new_n7752);
nor_4  g05406(new_n7755, new_n7754, new_n7743);
nor_4  g05407(new_n7756, new_n7755, new_n7751_1);
not_3  g05408(new_n7757, new_n7755);
nor_4  g05409(new_n7758, new_n7757, n19680);
nor_4  g05410(new_n7759_1, new_n7758, new_n7756);
not_3  g05411(new_n7760, new_n7759_1);
not_3  g05412(new_n7761, new_n7740);
nor_4  g05413(new_n7762, new_n7761, new_n7738);
nor_4  g05414(new_n7763, new_n7762, new_n7741);
not_3  g05415(new_n7764, new_n7763);
nor_4  g05416(new_n7765, new_n7764, n2809);
not_3  g05417(new_n7766, new_n7765);
xor_3  g05418(new_n7767, n25435, n18);
nand_4 g05419(new_n7768, new_n7767, n15508);
not_3  g05420(new_n7769_1, n2809);
nor_4  g05421(new_n7770, new_n7763, new_n7769_1);
nor_4  g05422(new_n7771, new_n7770, new_n7765);
nand_4 g05423(new_n7772, new_n7771, new_n7768);
nand_4 g05424(new_n7773_1, new_n7772, new_n7766);
nor_4  g05425(new_n7774, new_n7773_1, new_n7760);
nor_4  g05426(new_n7775, new_n7774, new_n7756);
xnor_3 g05427(new_n7776, new_n7775, new_n7750);
not_3  g05428(new_n7777, new_n7776);
xor_3  g05429(new_n7778, n18157, n11056);
nor_4  g05430(new_n7779, n15271, n12161);
not_3  g05431(new_n7780_1, new_n7779);
xor_3  g05432(new_n7781, n15271, n12161);
nor_4  g05433(new_n7782, n25877, n5026);
not_3  g05434(new_n7783, new_n7782);
nand_4 g05435(new_n7784, n24323, n8581);
xor_3  g05436(new_n7785, n25877, n5026);
nand_4 g05437(new_n7786, new_n7785, new_n7784);
nand_4 g05438(new_n7787, new_n7786, new_n7783);
nand_4 g05439(new_n7788_1, new_n7787, new_n7781);
nand_4 g05440(new_n7789, new_n7788_1, new_n7780_1);
nor_4  g05441(new_n7790, new_n7789, new_n7778);
not_3  g05442(new_n7791, new_n7778);
not_3  g05443(new_n7792, n12161);
xor_3  g05444(new_n7793, n15271, new_n7792);
not_3  g05445(new_n7794_1, new_n7784);
xnor_3 g05446(new_n7795, n25877, n5026);
nor_4  g05447(new_n7796, new_n7795, new_n7794_1);
nor_4  g05448(new_n7797, new_n7796, new_n7782);
nor_4  g05449(new_n7798, new_n7797, new_n7793);
nor_4  g05450(new_n7799, new_n7798, new_n7779);
nor_4  g05451(new_n7800, new_n7799, new_n7791);
nor_4  g05452(new_n7801, new_n7800, new_n7790);
nand_4 g05453(new_n7802, new_n7801, new_n4943);
not_3  g05454(new_n7803, new_n7802);
nor_4  g05455(new_n7804, new_n7801, new_n4943);
nor_4  g05456(new_n7805, new_n7804, new_n7803);
nor_4  g05457(new_n7806, new_n7787, new_n7781);
nor_4  g05458(new_n7807, new_n7806, new_n7798);
nand_4 g05459(new_n7808, new_n7807, new_n4947_1);
xor_3  g05460(new_n7809, new_n7795, new_n7784);
nor_4  g05461(new_n7810, new_n7809, n26443);
not_3  g05462(new_n7811_1, new_n7810);
xor_3  g05463(new_n7812, n24323, n8581);
not_3  g05464(new_n7813, new_n7812);
nor_4  g05465(new_n7814, new_n7813, new_n4957_1);
not_3  g05466(new_n7815, new_n7814);
xor_3  g05467(new_n7816, new_n7795, new_n7794_1);
nor_4  g05468(new_n7817, new_n7816, new_n4961);
nor_4  g05469(new_n7818, new_n7817, new_n7810);
nand_4 g05470(new_n7819, new_n7818, new_n7815);
nand_4 g05471(new_n7820, new_n7819, new_n7811_1);
not_3  g05472(new_n7821, new_n7807);
xor_3  g05473(new_n7822, new_n7821, n5822);
nand_4 g05474(new_n7823, new_n7822, new_n7820);
nand_4 g05475(new_n7824, new_n7823, new_n7808);
xnor_3 g05476(new_n7825, new_n7824, new_n7805);
xnor_3 g05477(new_n7826, new_n7825, new_n7777);
not_3  g05478(new_n7827, new_n7826);
not_3  g05479(new_n7828, new_n7773_1);
nor_4  g05480(new_n7829, new_n7828, new_n7759_1);
nor_4  g05481(new_n7830_1, new_n7829, new_n7774);
xnor_3 g05482(new_n7831, new_n7822, new_n7820);
not_3  g05483(new_n7832, new_n7831);
nor_4  g05484(new_n7833, new_n7832, new_n7830_1);
xnor_3 g05485(new_n7834_1, new_n7832, new_n7830_1);
xnor_3 g05486(new_n7835, new_n7771, new_n7768);
xnor_3 g05487(new_n7836, new_n7816, new_n4961);
xnor_3 g05488(new_n7837, new_n7836, new_n7814);
not_3  g05489(new_n7838, new_n7837);
nand_4 g05490(new_n7839, new_n7838, new_n7835);
not_3  g05491(new_n7840, new_n7767);
xor_3  g05492(new_n7841_1, new_n7840, n15508);
xor_3  g05493(new_n7842, new_n7813, n1681);
not_3  g05494(new_n7843, new_n7842);
nor_4  g05495(new_n7844, new_n7843, new_n7841_1);
xnor_3 g05496(new_n7845, new_n7837, new_n7835);
nand_4 g05497(new_n7846, new_n7845, new_n7844);
nand_4 g05498(new_n7847, new_n7846, new_n7839);
nor_4  g05499(new_n7848, new_n7847, new_n7834_1);
nor_4  g05500(new_n7849, new_n7848, new_n7833);
xor_3  g05501(n646, new_n7849, new_n7827);
nor_4  g05502(new_n7851, n19494, n2387);
nand_4 g05503(new_n7852, new_n7851, new_n2368);
nor_4  g05504(new_n7853, new_n7852, n26913);
xor_3  g05505(new_n7854, new_n7853, n21832);
xnor_3 g05506(new_n7855, new_n2497, new_n6339_1);
nand_4 g05507(new_n7856, new_n2503, n7731);
xnor_3 g05508(new_n7857, new_n2502, n7731);
nand_4 g05509(new_n7858, new_n2510, n12341);
xnor_3 g05510(new_n7859, new_n2507, n12341);
nor_4  g05511(new_n7860, new_n2512, n12384);
not_3  g05512(new_n7861, new_n7860);
nor_4  g05513(new_n7862, new_n7861, n20986);
xnor_3 g05514(new_n7863, new_n7860, new_n6351);
nor_4  g05515(new_n7864, new_n7863, new_n2515_1);
nor_4  g05516(new_n7865, new_n7864, new_n7862);
nand_4 g05517(new_n7866, new_n7865, new_n7859);
nand_4 g05518(new_n7867, new_n7866, new_n7858);
nand_4 g05519(new_n7868, new_n7867, new_n7857);
nand_4 g05520(new_n7869, new_n7868, new_n7856);
xnor_3 g05521(new_n7870, new_n7869, new_n7855);
xnor_3 g05522(new_n7871, new_n7870, new_n7854);
xor_3  g05523(new_n7872, new_n7852, n26913);
xnor_3 g05524(new_n7873, new_n2502, new_n6343);
xnor_3 g05525(new_n7874, new_n7867, new_n7873);
nand_4 g05526(new_n7875, new_n7874, new_n7872);
not_3  g05527(new_n7876_1, new_n7875);
xor_3  g05528(new_n7877, new_n7852, new_n2361_1);
xnor_3 g05529(new_n7878, new_n7867, new_n7857);
nand_4 g05530(new_n7879, new_n7878, new_n7877);
nand_4 g05531(new_n7880, new_n7879, new_n7875);
not_3  g05532(new_n7881, n12384);
xnor_3 g05533(new_n7882, new_n2512, new_n7881);
nor_4  g05534(new_n7883, new_n7882, new_n2571);
nand_4 g05535(new_n7884_1, new_n7883, new_n2372);
xnor_3 g05536(new_n7885, new_n7863, new_n2515_1);
xnor_3 g05537(new_n7886, new_n2512, n12384);
nand_4 g05538(new_n7887, new_n7886, n2387);
nor_4  g05539(new_n7888, new_n7887, n19494);
xnor_3 g05540(new_n7889, n19494, n2387);
not_3  g05541(new_n7890, new_n7889);
nor_4  g05542(new_n7891, new_n7890, new_n7883);
nor_4  g05543(new_n7892, new_n7891, new_n7888);
nand_4 g05544(new_n7893, new_n7892, new_n7885);
nand_4 g05545(new_n7894, new_n7893, new_n7884_1);
xnor_3 g05546(new_n7895, new_n7851, new_n2368);
not_3  g05547(new_n7896, new_n7895);
nor_4  g05548(new_n7897, new_n7896, new_n7894);
not_3  g05549(new_n7898, new_n7897);
xnor_3 g05550(new_n7899, new_n7865, new_n7859);
xnor_3 g05551(new_n7900, new_n7895, new_n7894);
nand_4 g05552(new_n7901, new_n7900, new_n7899);
nand_4 g05553(new_n7902, new_n7901, new_n7898);
nor_4  g05554(new_n7903, new_n7902, new_n7880);
nor_4  g05555(new_n7904, new_n7903, new_n7876_1);
xnor_3 g05556(new_n7905, new_n7904, new_n7871);
xnor_3 g05557(new_n7906, new_n7905, new_n3590);
not_3  g05558(new_n7907, new_n7906);
xnor_3 g05559(new_n7908, new_n7902, new_n7880);
nand_4 g05560(new_n7909, new_n7908, new_n3598);
xnor_3 g05561(new_n7910, new_n7900, new_n7899);
not_3  g05562(new_n7911, new_n7910);
nor_4  g05563(new_n7912, new_n7911, new_n3607);
xnor_3 g05564(new_n7913, new_n7910, new_n3606);
xor_3  g05565(new_n7914, new_n7882, n2387);
nor_4  g05566(new_n7915, new_n7914, new_n3613);
nor_4  g05567(new_n7916, new_n7915, new_n3617_1);
not_3  g05568(new_n7917_1, new_n7916);
not_3  g05569(new_n7918, new_n7885);
xor_3  g05570(new_n7919, new_n7892, new_n7918);
xor_3  g05571(new_n7920, new_n7882, new_n2571);
nand_4 g05572(new_n7921, new_n7920, new_n3612);
nor_4  g05573(new_n7922, new_n7921, new_n3616);
nor_4  g05574(new_n7923, new_n7922, new_n7916);
nand_4 g05575(new_n7924, new_n7923, new_n7919);
nand_4 g05576(new_n7925, new_n7924, new_n7917_1);
nor_4  g05577(new_n7926, new_n7925, new_n7913);
nor_4  g05578(new_n7927, new_n7926, new_n7912);
xnor_3 g05579(new_n7928, new_n7908, new_n3599);
nand_4 g05580(new_n7929, new_n7928, new_n7927);
nand_4 g05581(new_n7930, new_n7929, new_n7909);
xor_3  g05582(n696, new_n7930, new_n7907);
xor_3  g05583(new_n7932, n25475, n23697);
not_3  g05584(new_n7933, new_n7932);
nor_4  g05585(new_n7934, n23849, n2289);
xor_3  g05586(new_n7935, n23849, n2289);
not_3  g05587(new_n7936, new_n7935);
not_3  g05588(new_n7937_1, n1112);
nand_4 g05589(new_n7938, new_n5022, new_n7937_1);
xor_3  g05590(new_n7939, n12446, n1112);
nor_4  g05591(new_n7940, n20179, n11011);
not_3  g05592(new_n7941, new_n7940);
xor_3  g05593(new_n7942, n20179, n11011);
nor_4  g05594(new_n7943_1, n19228, n16029);
not_3  g05595(new_n7944, new_n7943_1);
xor_3  g05596(new_n7945, n19228, n16029);
nor_4  g05597(new_n7946, n16476, n15539);
not_3  g05598(new_n7947, new_n7946);
nand_4 g05599(new_n7948, n16476, n15539);
not_3  g05600(new_n7949_1, new_n7948);
nor_4  g05601(new_n7950_1, new_n7949_1, new_n7946);
nor_4  g05602(new_n7951, n11615, n8052);
not_3  g05603(new_n7952, new_n7951);
nand_4 g05604(new_n7953, n11615, n8052);
not_3  g05605(new_n7954, new_n7953);
nor_4  g05606(new_n7955, new_n7954, new_n7951);
nor_4  g05607(new_n7956, n22433, n10158);
not_3  g05608(new_n7957, new_n7956);
nand_4 g05609(new_n7958, n18962, n14090);
nand_4 g05610(new_n7959_1, n22433, n10158);
not_3  g05611(new_n7960, new_n7959_1);
nor_4  g05612(new_n7961, new_n7960, new_n7956);
nand_4 g05613(new_n7962, new_n7961, new_n7958);
nand_4 g05614(new_n7963_1, new_n7962, new_n7957);
nand_4 g05615(new_n7964, new_n7963_1, new_n7955);
nand_4 g05616(new_n7965, new_n7964, new_n7952);
nand_4 g05617(new_n7966, new_n7965, new_n7950_1);
nand_4 g05618(new_n7967, new_n7966, new_n7947);
nand_4 g05619(new_n7968_1, new_n7967, new_n7945);
nand_4 g05620(new_n7969, new_n7968_1, new_n7944);
nand_4 g05621(new_n7970, new_n7969, new_n7942);
nand_4 g05622(new_n7971, new_n7970, new_n7941);
nand_4 g05623(new_n7972, new_n7971, new_n7939);
nand_4 g05624(new_n7973, new_n7972, new_n7938);
not_3  g05625(new_n7974, new_n7973);
nor_4  g05626(new_n7975, new_n7974, new_n7936);
nor_4  g05627(new_n7976, new_n7975, new_n7934);
xnor_3 g05628(new_n7977, new_n7976, new_n7933);
not_3  g05629(new_n7978, new_n7977);
nor_4  g05630(new_n7979, new_n7978, new_n6381_1);
nor_4  g05631(new_n7980, new_n7977, n25345);
nor_4  g05632(new_n7981, new_n7980, new_n7979);
xnor_3 g05633(new_n7982, new_n7973, new_n7935);
not_3  g05634(new_n7983, new_n7982);
nor_4  g05635(new_n7984, new_n7983, new_n6385_1);
not_3  g05636(new_n7985, new_n7984);
nor_4  g05637(new_n7986, new_n7982, n9655);
nor_4  g05638(new_n7987, new_n7986, new_n7984);
not_3  g05639(new_n7988, n13490);
xnor_3 g05640(new_n7989, new_n7971, new_n7939);
not_3  g05641(new_n7990, new_n7989);
nor_4  g05642(new_n7991, new_n7990, new_n7988);
not_3  g05643(new_n7992_1, new_n7991);
nor_4  g05644(new_n7993, new_n7989, n13490);
nor_4  g05645(new_n7994, new_n7993, new_n7991);
xnor_3 g05646(new_n7995, new_n7969, new_n7942);
nand_4 g05647(new_n7996, new_n7995, n22660);
xnor_3 g05648(new_n7997, new_n7967, new_n7945);
nor_4  g05649(new_n7998, new_n7997, n1777);
xnor_3 g05650(new_n7999_1, new_n7997, new_n6391);
not_3  g05651(new_n8000, new_n7999_1);
not_3  g05652(new_n8001, new_n7950_1);
xnor_3 g05653(new_n8002, new_n7965, new_n8001);
nand_4 g05654(new_n8003, new_n8002, new_n6395);
not_3  g05655(new_n8004, new_n8003);
xnor_3 g05656(new_n8005, new_n8002, new_n6395);
not_3  g05657(new_n8006_1, new_n7958);
xnor_3 g05658(new_n8007, n22433, n10158);
nor_4  g05659(new_n8008, new_n8007, new_n8006_1);
nor_4  g05660(new_n8009, new_n8008, new_n7956);
xnor_3 g05661(new_n8010, new_n8009, new_n7955);
nor_4  g05662(new_n8011, new_n8010, new_n6401);
not_3  g05663(new_n8012, new_n8011);
xnor_3 g05664(new_n8013, new_n7963_1, new_n7955);
nor_4  g05665(new_n8014, new_n8013, n15636);
nor_4  g05666(new_n8015, new_n8014, new_n8011);
nor_4  g05667(new_n8016, n18962, n14090);
nor_4  g05668(new_n8017, new_n8016, new_n8006_1);
not_3  g05669(new_n8018, new_n8017);
nand_4 g05670(new_n8019, n20077, n6794);
nor_4  g05671(new_n8020, new_n8019, new_n8018);
not_3  g05672(new_n8021, new_n8020);
xnor_3 g05673(new_n8022, new_n8007, new_n8006_1);
nor_4  g05674(new_n8023, new_n8018, new_n6575);
nor_4  g05675(new_n8024, new_n8023, n20077);
nor_4  g05676(new_n8025, new_n8024, new_n8020);
nand_4 g05677(new_n8026, new_n8025, new_n8022);
nand_4 g05678(new_n8027_1, new_n8026, new_n8021);
nand_4 g05679(new_n8028, new_n8027_1, new_n8015);
nand_4 g05680(new_n8029, new_n8028, new_n8012);
nor_4  g05681(new_n8030, new_n8029, new_n8005);
nor_4  g05682(new_n8031_1, new_n8030, new_n8004);
nor_4  g05683(new_n8032, new_n8031_1, new_n8000);
nor_4  g05684(new_n8033, new_n8032, new_n7998);
not_3  g05685(new_n8034, new_n7996);
nor_4  g05686(new_n8035, new_n7995, n22660);
nor_4  g05687(new_n8036, new_n8035, new_n8034);
nand_4 g05688(new_n8037, new_n8036, new_n8033);
nand_4 g05689(new_n8038, new_n8037, new_n7996);
nand_4 g05690(new_n8039, new_n8038, new_n7994);
nand_4 g05691(new_n8040, new_n8039, new_n7992_1);
nand_4 g05692(new_n8041, new_n8040, new_n7987);
nand_4 g05693(new_n8042_1, new_n8041, new_n7985);
xnor_3 g05694(new_n8043, new_n8042_1, new_n7981);
xor_3  g05695(new_n8044, n21915, n15182);
not_3  g05696(new_n8045, n13775);
nand_4 g05697(new_n8046, new_n6328, new_n8045);
xor_3  g05698(new_n8047, n27037, n13775);
nor_4  g05699(new_n8048, n8964, n1293);
not_3  g05700(new_n8049, new_n8048);
xor_3  g05701(new_n8050, n8964, n1293);
nor_4  g05702(new_n8051, n20151, n19042);
not_3  g05703(new_n8052_1, new_n8051);
xor_3  g05704(new_n8053, n20151, n19042);
nor_4  g05705(new_n8054, n19472, n7693);
not_3  g05706(new_n8055, new_n8054);
xor_3  g05707(new_n8056, n19472, n7693);
nand_4 g05708(new_n8057, n25370, n10405);
not_3  g05709(new_n8058, new_n8057);
nor_4  g05710(new_n8059, n25370, n10405);
nor_4  g05711(new_n8060, n24786, n11302);
not_3  g05712(new_n8061, new_n8060);
nand_4 g05713(new_n8062, new_n4601, new_n8061);
nor_4  g05714(new_n8063, new_n8062, new_n8059);
nor_4  g05715(new_n8064, new_n8063, new_n8058);
nand_4 g05716(new_n8065, new_n8064, new_n8056);
nand_4 g05717(new_n8066, new_n8065, new_n8055);
nand_4 g05718(new_n8067_1, new_n8066, new_n8053);
nand_4 g05719(new_n8068, new_n8067_1, new_n8052_1);
nand_4 g05720(new_n8069, new_n8068, new_n8050);
nand_4 g05721(new_n8070, new_n8069, new_n8049);
nand_4 g05722(new_n8071, new_n8070, new_n8047);
nand_4 g05723(new_n8072, new_n8071, new_n8046);
xnor_3 g05724(new_n8073, new_n8072, new_n8044);
not_3  g05725(new_n8074, new_n8073);
xor_3  g05726(new_n8075, new_n8074, new_n6324);
not_3  g05727(new_n8076, new_n8070);
xnor_3 g05728(new_n8077, new_n8076, new_n8047);
not_3  g05729(new_n8078, new_n8077);
nand_4 g05730(new_n8079, new_n8078, n11736);
xor_3  g05731(new_n8080, new_n8077, new_n6330_1);
not_3  g05732(new_n8081, n23200);
not_3  g05733(new_n8082, new_n8050);
not_3  g05734(new_n8083, new_n8068);
xor_3  g05735(new_n8084, new_n8083, new_n8082);
nor_4  g05736(new_n8085, new_n8084, new_n8081);
not_3  g05737(new_n8086, new_n8085);
xor_3  g05738(new_n8087, new_n8083, new_n8050);
nor_4  g05739(new_n8088, new_n8087, n23200);
nor_4  g05740(new_n8089, new_n8088, new_n8085);
not_3  g05741(new_n8090, new_n8067_1);
nor_4  g05742(new_n8091, new_n8066, new_n8053);
nor_4  g05743(new_n8092, new_n8091, new_n8090);
nor_4  g05744(new_n8093, new_n8092, new_n6335);
not_3  g05745(new_n8094, new_n8093);
not_3  g05746(new_n8095_1, new_n8092);
nor_4  g05747(new_n8096, new_n8095_1, n17959);
nor_4  g05748(new_n8097, new_n8096, new_n8093);
not_3  g05749(new_n8098, new_n8056);
xnor_3 g05750(new_n8099, new_n8064, new_n8098);
nor_4  g05751(new_n8100, new_n8099, new_n6339_1);
not_3  g05752(new_n8101, new_n8100);
not_3  g05753(new_n8102, new_n8099);
nor_4  g05754(new_n8103_1, new_n8102, n7566);
nor_4  g05755(new_n8104, new_n8103_1, new_n8100);
nor_4  g05756(new_n8105, new_n8059, new_n8058);
xnor_3 g05757(new_n8106, new_n8105, new_n8062);
not_3  g05758(new_n8107, new_n8106);
nor_4  g05759(new_n8108, new_n8107, new_n6343);
not_3  g05760(new_n8109_1, new_n8108);
xor_3  g05761(new_n8110, new_n8107, new_n6343);
nor_4  g05762(new_n8111, new_n4603, new_n6348);
not_3  g05763(new_n8112, new_n8111);
nor_4  g05764(new_n8113, new_n4629, n20986);
nand_4 g05765(new_n8114, new_n4625, n12384);
not_3  g05766(new_n8115, new_n8114);
xnor_3 g05767(new_n8116, new_n4618, new_n6351);
nor_4  g05768(new_n8117, new_n8116, new_n8115);
nor_4  g05769(new_n8118, new_n8117, new_n8113);
not_3  g05770(new_n8119, new_n4603);
nor_4  g05771(new_n8120, new_n8119, n12341);
nor_4  g05772(new_n8121, new_n8120, new_n8111);
nand_4 g05773(new_n8122, new_n8121, new_n8118);
nand_4 g05774(new_n8123, new_n8122, new_n8112);
nand_4 g05775(new_n8124, new_n8123, new_n8110);
nand_4 g05776(new_n8125, new_n8124, new_n8109_1);
nand_4 g05777(new_n8126, new_n8125, new_n8104);
nand_4 g05778(new_n8127_1, new_n8126, new_n8101);
nand_4 g05779(new_n8128, new_n8127_1, new_n8097);
nand_4 g05780(new_n8129, new_n8128, new_n8094);
nand_4 g05781(new_n8130_1, new_n8129, new_n8089);
nand_4 g05782(new_n8131, new_n8130_1, new_n8086);
nand_4 g05783(new_n8132, new_n8131, new_n8080);
nand_4 g05784(new_n8133, new_n8132, new_n8079);
xnor_3 g05785(new_n8134, new_n8133, new_n8075);
xnor_3 g05786(new_n8135_1, new_n8134, new_n8043);
xnor_3 g05787(new_n8136, new_n8131, new_n8080);
xnor_3 g05788(new_n8137, new_n8040, new_n7987);
not_3  g05789(new_n8138, new_n8137);
nand_4 g05790(new_n8139_1, new_n8138, new_n8136);
xnor_3 g05791(new_n8140, new_n8137, new_n8136);
xnor_3 g05792(new_n8141, new_n8129, new_n8089);
xnor_3 g05793(new_n8142, new_n8038, new_n7994);
not_3  g05794(new_n8143, new_n8142);
nand_4 g05795(new_n8144, new_n8143, new_n8141);
xnor_3 g05796(new_n8145, new_n8142, new_n8141);
xnor_3 g05797(new_n8146, new_n8127_1, new_n8097);
not_3  g05798(new_n8147, new_n8036);
xnor_3 g05799(new_n8148_1, new_n8147, new_n8033);
nand_4 g05800(new_n8149_1, new_n8148_1, new_n8146);
not_3  g05801(new_n8150, new_n8148_1);
xnor_3 g05802(new_n8151, new_n8150, new_n8146);
xnor_3 g05803(new_n8152, new_n8031_1, new_n8000);
xnor_3 g05804(new_n8153, new_n8125, new_n8104);
nand_4 g05805(new_n8154, new_n8153, new_n8152);
not_3  g05806(new_n8155, new_n8152);
xnor_3 g05807(new_n8156, new_n8153, new_n8155);
not_3  g05808(new_n8157, new_n8005);
not_3  g05809(new_n8158, new_n8029);
nor_4  g05810(new_n8159_1, new_n8158, new_n8157);
nor_4  g05811(new_n8160, new_n8159_1, new_n8030);
not_3  g05812(new_n8161, new_n8160);
xnor_3 g05813(new_n8162, new_n8123, new_n8110);
nand_4 g05814(new_n8163, new_n8162, new_n8161);
xnor_3 g05815(new_n8164, new_n8162, new_n8160);
not_3  g05816(new_n8165, new_n8121);
xnor_3 g05817(new_n8166, new_n8165, new_n8118);
not_3  g05818(new_n8167, new_n8166);
xnor_3 g05819(new_n8168, new_n8027_1, new_n8015);
not_3  g05820(new_n8169, new_n8168);
nand_4 g05821(new_n8170, new_n8169, new_n8167);
xnor_3 g05822(new_n8171, new_n8169, new_n8166);
xnor_3 g05823(new_n8172, new_n8116, new_n8114);
not_3  g05824(new_n8173, new_n8026);
nor_4  g05825(new_n8174, new_n8025, new_n8022);
nor_4  g05826(new_n8175, new_n8174, new_n8173);
nand_4 g05827(new_n8176, new_n8175, new_n8172);
xor_3  g05828(new_n8177, new_n8017, n6794);
not_3  g05829(new_n8178, new_n8177);
not_3  g05830(new_n8179_1, new_n4625);
xor_3  g05831(new_n8180, new_n8179_1, new_n7881);
nor_4  g05832(new_n8181, new_n8180, new_n8178);
not_3  g05833(new_n8182, new_n8176);
nor_4  g05834(new_n8183, new_n8175, new_n8172);
nor_4  g05835(new_n8184, new_n8183, new_n8182);
nand_4 g05836(new_n8185, new_n8184, new_n8181);
nand_4 g05837(new_n8186, new_n8185, new_n8176);
nand_4 g05838(new_n8187, new_n8186, new_n8171);
nand_4 g05839(new_n8188, new_n8187, new_n8170);
nand_4 g05840(new_n8189, new_n8188, new_n8164);
nand_4 g05841(new_n8190, new_n8189, new_n8163);
nand_4 g05842(new_n8191, new_n8190, new_n8156);
nand_4 g05843(new_n8192, new_n8191, new_n8154);
nand_4 g05844(new_n8193, new_n8192, new_n8151);
nand_4 g05845(new_n8194_1, new_n8193, new_n8149_1);
nand_4 g05846(new_n8195, new_n8194_1, new_n8145);
nand_4 g05847(new_n8196, new_n8195, new_n8144);
nand_4 g05848(new_n8197, new_n8196, new_n8140);
nand_4 g05849(new_n8198, new_n8197, new_n8139_1);
xnor_3 g05850(n723, new_n8198, new_n8135_1);
not_3  g05851(new_n8200, n2272);
xor_3  g05852(new_n8201, n26986, new_n8200);
not_3  g05853(new_n8202, new_n8201);
not_3  g05854(new_n8203, n25331);
nor_4  g05855(new_n8204, new_n8203, n21287);
not_3  g05856(new_n8205, n21287);
xor_3  g05857(new_n8206, n25331, new_n8205);
not_3  g05858(new_n8207, n4256);
nand_4 g05859(new_n8208, n18483, new_n8207);
xor_3  g05860(new_n8209, n18483, new_n8207);
not_3  g05861(new_n8210, n21934);
nor_4  g05862(new_n8211, n22332, new_n8210);
not_3  g05863(new_n8212, new_n8211);
xor_3  g05864(new_n8213, n22332, new_n8210);
not_3  g05865(new_n8214, n18901);
nor_4  g05866(new_n8215_1, n18907, new_n8214);
not_3  g05867(new_n8216, new_n8215_1);
xor_3  g05868(new_n8217, n18907, new_n8214);
not_3  g05869(new_n8218, n4376);
nor_4  g05870(new_n8219, new_n8218, n2731);
xor_3  g05871(new_n8220, n4376, new_n4190);
not_3  g05872(new_n8221, new_n8220);
not_3  g05873(new_n8222, n14570);
nor_4  g05874(new_n8223, n19911, new_n8222);
xor_3  g05875(new_n8224, n19911, n14570);
nor_4  g05876(new_n8225, n23775, new_n4201);
not_3  g05877(new_n8226, n23775);
nor_4  g05878(new_n8227, new_n8226, n13708);
nor_4  g05879(new_n8228, new_n4205_1, n8259);
not_3  g05880(new_n8229, n8259);
nor_4  g05881(new_n8230, n18409, new_n8229);
not_3  g05882(new_n8231, n11479);
nand_4 g05883(new_n8232, new_n8231, n5704);
nor_4  g05884(new_n8233, new_n8232, new_n8230);
nor_4  g05885(new_n8234, new_n8233, new_n8228);
nor_4  g05886(new_n8235, new_n8234, new_n8227);
nor_4  g05887(new_n8236, new_n8235, new_n8225);
not_3  g05888(new_n8237, new_n8236);
nor_4  g05889(new_n8238, new_n8237, new_n8224);
nor_4  g05890(new_n8239, new_n8238, new_n8223);
nor_4  g05891(new_n8240, new_n8239, new_n8221);
nor_4  g05892(new_n8241, new_n8240, new_n8219);
not_3  g05893(new_n8242, new_n8241);
nand_4 g05894(new_n8243, new_n8242, new_n8217);
nand_4 g05895(new_n8244_1, new_n8243, new_n8216);
nand_4 g05896(new_n8245, new_n8244_1, new_n8213);
nand_4 g05897(new_n8246, new_n8245, new_n8212);
nand_4 g05898(new_n8247, new_n8246, new_n8209);
nand_4 g05899(new_n8248, new_n8247, new_n8208);
nand_4 g05900(new_n8249, new_n8248, new_n8206);
not_3  g05901(new_n8250, new_n8249);
nor_4  g05902(new_n8251, new_n8250, new_n8204);
xor_3  g05903(new_n8252, new_n8251, new_n8202);
xor_3  g05904(new_n8253, n1255, n468);
nor_4  g05905(new_n8254, n9512, n5400);
xor_3  g05906(new_n8255_1, n9512, n5400);
not_3  g05907(new_n8256_1, new_n8255_1);
not_3  g05908(new_n8257, n16608);
not_3  g05909(new_n8258, n23923);
nand_4 g05910(new_n8259_1, new_n8258, new_n8257);
xor_3  g05911(new_n8260, n23923, n16608);
nor_4  g05912(new_n8261, n21735, n329);
not_3  g05913(new_n8262, new_n8261);
xor_3  g05914(new_n8263, n21735, n329);
nor_4  g05915(new_n8264, n24170, n24085);
not_3  g05916(new_n8265, new_n8264);
xor_3  g05917(new_n8266, n24170, n24085);
nor_4  g05918(new_n8267_1, n14071, n2409);
not_3  g05919(new_n8268, new_n8267_1);
xor_3  g05920(new_n8269, n14071, n2409);
nor_4  g05921(new_n8270, n8869, n1738);
not_3  g05922(new_n8271, new_n8270);
xor_3  g05923(new_n8272, n8869, n1738);
not_3  g05924(new_n8273, n10372);
nand_4 g05925(new_n8274, new_n5246, new_n8273);
nand_4 g05926(new_n8275, n19107, n7428);
xor_3  g05927(new_n8276_1, n12152, n10372);
nand_4 g05928(new_n8277, new_n8276_1, new_n8275);
nand_4 g05929(new_n8278, new_n8277, new_n8274);
nand_4 g05930(new_n8279, new_n8278, new_n8272);
nand_4 g05931(new_n8280, new_n8279, new_n8271);
nand_4 g05932(new_n8281, new_n8280, new_n8269);
nand_4 g05933(new_n8282, new_n8281, new_n8268);
nand_4 g05934(new_n8283, new_n8282, new_n8266);
nand_4 g05935(new_n8284, new_n8283, new_n8265);
nand_4 g05936(new_n8285_1, new_n8284, new_n8263);
nand_4 g05937(new_n8286, new_n8285_1, new_n8262);
nand_4 g05938(new_n8287, new_n8286, new_n8260);
nand_4 g05939(new_n8288_1, new_n8287, new_n8259_1);
not_3  g05940(new_n8289, new_n8288_1);
nor_4  g05941(new_n8290, new_n8289, new_n8256_1);
nor_4  g05942(new_n8291, new_n8290, new_n8254);
xor_3  g05943(new_n8292, new_n8291, new_n8253);
xor_3  g05944(new_n8293, n14130, n12861);
not_3  g05945(new_n8294, new_n8293);
nor_4  g05946(new_n8295, n16482, n13333);
xor_3  g05947(new_n8296, n16482, n13333);
not_3  g05948(new_n8297, new_n8296);
not_3  g05949(new_n8298, n2210);
nand_4 g05950(new_n8299, new_n2349, new_n8298);
xor_3  g05951(new_n8300, n9942, n2210);
nor_4  g05952(new_n8301, n25643, n20604);
not_3  g05953(new_n8302, new_n8301);
nand_4 g05954(new_n8303, new_n5903_1, new_n8302);
nand_4 g05955(new_n8304, new_n8303, new_n8300);
nand_4 g05956(new_n8305_1, new_n8304, new_n8299);
not_3  g05957(new_n8306_1, new_n8305_1);
nor_4  g05958(new_n8307, new_n8306_1, new_n8297);
nor_4  g05959(new_n8308, new_n8307, new_n8295);
xnor_3 g05960(new_n8309_1, new_n8308, new_n8294);
not_3  g05961(new_n8310, new_n8309_1);
nor_4  g05962(new_n8311, new_n8310, new_n8292);
not_3  g05963(new_n8312, new_n8311);
not_3  g05964(new_n8313, new_n8253);
xor_3  g05965(new_n8314, new_n8291, new_n8313);
xnor_3 g05966(new_n8315, new_n8309_1, new_n8314);
not_3  g05967(new_n8316, new_n8315);
xor_3  g05968(new_n8317, new_n8289, new_n8255_1);
nor_4  g05969(new_n8318, new_n8305_1, new_n8296);
nor_4  g05970(new_n8319, new_n8318, new_n8307);
nor_4  g05971(new_n8320_1, new_n8319, new_n8317);
not_3  g05972(new_n8321_1, new_n8320_1);
not_3  g05973(new_n8322, new_n8319);
xnor_3 g05974(new_n8323, new_n8322, new_n8317);
xnor_3 g05975(new_n8324_1, new_n8303, new_n8300);
xnor_3 g05976(new_n8325, new_n8286, new_n8260);
not_3  g05977(new_n8326, new_n8325);
nand_4 g05978(new_n8327, new_n8326, new_n8324_1);
xnor_3 g05979(new_n8328, new_n8325, new_n8324_1);
not_3  g05980(new_n8329, new_n5905);
xnor_3 g05981(new_n8330, new_n8284, new_n8263);
not_3  g05982(new_n8331, new_n8330);
nand_4 g05983(new_n8332, new_n8331, new_n8329);
xnor_3 g05984(new_n8333, new_n8330, new_n8329);
not_3  g05985(new_n8334, new_n5895);
xnor_3 g05986(new_n8335, new_n8282, new_n8266);
nor_4  g05987(new_n8336, new_n8335, new_n8334);
not_3  g05988(new_n8337, new_n8336);
xnor_3 g05989(new_n8338, new_n8335, new_n5895);
not_3  g05990(new_n8339_1, new_n8269);
xnor_3 g05991(new_n8340, new_n8280, new_n8339_1);
nand_4 g05992(new_n8341, new_n8340, new_n5887);
not_3  g05993(new_n8342, new_n5887);
xnor_3 g05994(new_n8343, new_n8340, new_n8342);
not_3  g05995(new_n8344, new_n8272);
xnor_3 g05996(new_n8345, new_n8278, new_n8344);
nand_4 g05997(new_n8346, new_n8345, new_n5881);
xnor_3 g05998(new_n8347, new_n8345, new_n5880);
not_3  g05999(new_n8348, new_n5867);
xnor_3 g06000(new_n8349, n12152, n10372);
xor_3  g06001(new_n8350, new_n8349, new_n8275);
nor_4  g06002(new_n8351, new_n8350, new_n8348);
not_3  g06003(new_n8352, new_n8351);
xor_3  g06004(new_n8353, n19107, n7428);
nor_4  g06005(new_n8354, new_n8353, new_n5918);
not_3  g06006(new_n8355, new_n8275);
xor_3  g06007(new_n8356, new_n8349, new_n8355);
nor_4  g06008(new_n8357, new_n8356, new_n5867);
nor_4  g06009(new_n8358, new_n8357, new_n8351);
nand_4 g06010(new_n8359, new_n8358, new_n8354);
nand_4 g06011(new_n8360, new_n8359, new_n8352);
nand_4 g06012(new_n8361, new_n8360, new_n8347);
nand_4 g06013(new_n8362, new_n8361, new_n8346);
nand_4 g06014(new_n8363_1, new_n8362, new_n8343);
nand_4 g06015(new_n8364, new_n8363_1, new_n8341);
nand_4 g06016(new_n8365, new_n8364, new_n8338);
nand_4 g06017(new_n8366, new_n8365, new_n8337);
nand_4 g06018(new_n8367, new_n8366, new_n8333);
nand_4 g06019(new_n8368, new_n8367, new_n8332);
nand_4 g06020(new_n8369, new_n8368, new_n8328);
nand_4 g06021(new_n8370, new_n8369, new_n8327);
nand_4 g06022(new_n8371, new_n8370, new_n8323);
nand_4 g06023(new_n8372, new_n8371, new_n8321_1);
nand_4 g06024(new_n8373, new_n8372, new_n8316);
nand_4 g06025(new_n8374, new_n8373, new_n8312);
xor_3  g06026(new_n8375, n22442, n22253);
not_3  g06027(new_n8376_1, new_n8375);
nor_4  g06028(new_n8377, n1255, n468);
nor_4  g06029(new_n8378, new_n8291, new_n8313);
nor_4  g06030(new_n8379, new_n8378, new_n8377);
xor_3  g06031(new_n8380, new_n8379, new_n8376_1);
xor_3  g06032(new_n8381_1, n8856, n8305);
nor_4  g06033(new_n8382, n14130, n12861);
nor_4  g06034(new_n8383, new_n8308, new_n8294);
nor_4  g06035(new_n8384, new_n8383, new_n8382);
xnor_3 g06036(new_n8385, new_n8384, new_n8381_1);
not_3  g06037(new_n8386, new_n8385);
xnor_3 g06038(new_n8387, new_n8386, new_n8380);
not_3  g06039(new_n8388, new_n8387);
xnor_3 g06040(new_n8389, new_n8388, new_n8374);
nor_4  g06041(new_n8390, new_n8389, new_n8252);
xnor_3 g06042(new_n8391, new_n8389, new_n8252);
xor_3  g06043(new_n8392, new_n8248, new_n8206);
not_3  g06044(new_n8393, new_n8371);
nor_4  g06045(new_n8394, new_n8393, new_n8320_1);
xnor_3 g06046(new_n8395, new_n8394, new_n8315);
nor_4  g06047(new_n8396, new_n8395, new_n8392);
not_3  g06048(new_n8397, new_n8392);
xnor_3 g06049(new_n8398, new_n8394, new_n8316);
xnor_3 g06050(new_n8399_1, new_n8398, new_n8397);
xnor_3 g06051(new_n8400, new_n8246, new_n8209);
xnor_3 g06052(new_n8401, new_n8370, new_n8323);
not_3  g06053(new_n8402, new_n8401);
nand_4 g06054(new_n8403, new_n8402, new_n8400);
xnor_3 g06055(new_n8404, new_n8401, new_n8400);
not_3  g06056(new_n8405_1, new_n8213);
xor_3  g06057(new_n8406, new_n8244_1, new_n8405_1);
xnor_3 g06058(new_n8407, new_n8368, new_n8328);
not_3  g06059(new_n8408_1, new_n8407);
nand_4 g06060(new_n8409, new_n8408_1, new_n8406);
xnor_3 g06061(new_n8410, new_n8407, new_n8406);
xor_3  g06062(new_n8411, new_n8242, new_n8217);
not_3  g06063(new_n8412, new_n8411);
xnor_3 g06064(new_n8413, new_n8330, new_n5905);
xnor_3 g06065(new_n8414, new_n8366, new_n8413);
nand_4 g06066(new_n8415, new_n8414, new_n8412);
xnor_3 g06067(new_n8416, new_n8414, new_n8411);
xor_3  g06068(new_n8417_1, new_n8239, new_n8221);
not_3  g06069(new_n8418, new_n8417_1);
xnor_3 g06070(new_n8419, new_n8335, new_n8334);
xnor_3 g06071(new_n8420, new_n8364, new_n8419);
nand_4 g06072(new_n8421, new_n8420, new_n8418);
xnor_3 g06073(new_n8422, new_n8420, new_n8417_1);
xnor_3 g06074(new_n8423, new_n8340, new_n5887);
xnor_3 g06075(new_n8424, new_n8362, new_n8423);
xor_3  g06076(new_n8425, new_n8237, new_n8224);
not_3  g06077(new_n8426, new_n8425);
nand_4 g06078(new_n8427, new_n8426, new_n8424);
xnor_3 g06079(new_n8428, new_n8360, new_n8347);
not_3  g06080(new_n8429, new_n8428);
nor_4  g06081(new_n8430, new_n8227, new_n8225);
not_3  g06082(new_n8431, new_n8430);
xor_3  g06083(new_n8432_1, new_n8431, new_n8234);
nand_4 g06084(new_n8433, new_n8432_1, new_n8429);
xnor_3 g06085(new_n8434, new_n8432_1, new_n8428);
xnor_3 g06086(new_n8435, new_n8353, new_n5862);
xor_3  g06087(new_n8436, n11479, new_n2389);
nor_4  g06088(new_n8437, new_n8436, new_n8435);
nor_4  g06089(new_n8438, new_n8230, new_n8228);
xor_3  g06090(new_n8439_1, new_n8438, new_n8232);
nand_4 g06091(new_n8440, new_n8439_1, new_n8437);
not_3  g06092(new_n8441, new_n8440);
not_3  g06093(new_n8442, new_n8358);
xnor_3 g06094(new_n8443, new_n8442, new_n8354);
xnor_3 g06095(new_n8444, new_n8439_1, new_n8437);
nor_4  g06096(new_n8445, new_n8444, new_n8443);
nor_4  g06097(new_n8446, new_n8445, new_n8441);
nand_4 g06098(new_n8447, new_n8446, new_n8434);
nand_4 g06099(new_n8448, new_n8447, new_n8433);
xnor_3 g06100(new_n8449, new_n8425, new_n8424);
nand_4 g06101(new_n8450, new_n8449, new_n8448);
nand_4 g06102(new_n8451, new_n8450, new_n8427);
nand_4 g06103(new_n8452, new_n8451, new_n8422);
nand_4 g06104(new_n8453_1, new_n8452, new_n8421);
nand_4 g06105(new_n8454, new_n8453_1, new_n8416);
nand_4 g06106(new_n8455, new_n8454, new_n8415);
nand_4 g06107(new_n8456, new_n8455, new_n8410);
nand_4 g06108(new_n8457, new_n8456, new_n8409);
nand_4 g06109(new_n8458, new_n8457, new_n8404);
nand_4 g06110(new_n8459, new_n8458, new_n8403);
not_3  g06111(new_n8460, new_n8459);
nor_4  g06112(new_n8461, new_n8460, new_n8399_1);
nor_4  g06113(new_n8462, new_n8461, new_n8396);
nor_4  g06114(new_n8463, new_n8462, new_n8391);
nor_4  g06115(new_n8464, new_n8463, new_n8390);
nor_4  g06116(new_n8465, n26986, new_n8200);
nor_4  g06117(new_n8466, new_n8251, new_n8202);
nor_4  g06118(new_n8467, new_n8466, new_n8465);
not_3  g06119(new_n8468, new_n8467);
nor_4  g06120(new_n8469, n22442, n22253);
nor_4  g06121(new_n8470, new_n8379, new_n8376_1);
nor_4  g06122(new_n8471, new_n8470, new_n8469);
nor_4  g06123(new_n8472, n8856, n8305);
not_3  g06124(new_n8473, new_n8381_1);
nor_4  g06125(new_n8474, new_n8384, new_n8473);
nor_4  g06126(new_n8475, new_n8474, new_n8472);
xor_3  g06127(new_n8476, new_n8475, new_n8471);
nand_4 g06128(new_n8477, new_n8386, new_n8380);
nand_4 g06129(new_n8478, new_n8388, new_n8374);
nand_4 g06130(new_n8479, new_n8478, new_n8477);
nor_4  g06131(new_n8480_1, new_n8479, new_n8476);
not_3  g06132(new_n8481, new_n8476);
not_3  g06133(new_n8482, new_n8479);
nor_4  g06134(new_n8483, new_n8482, new_n8481);
nor_4  g06135(new_n8484, new_n8483, new_n8480_1);
nor_4  g06136(new_n8485, new_n8484, new_n8468);
xnor_3 g06137(new_n8486, new_n8479, new_n8476);
nor_4  g06138(new_n8487, new_n8486, new_n8467);
nor_4  g06139(new_n8488, new_n8487, new_n8485);
xnor_3 g06140(n735, new_n8488, new_n8464);
xor_3  g06141(new_n8490, n21138, n14230);
not_3  g06142(new_n8491, n26167);
xnor_3 g06143(new_n8492, new_n8017, n19234);
not_3  g06144(new_n8493, new_n8492);
xor_3  g06145(new_n8494, new_n8493, new_n8491);
not_3  g06146(new_n8495, new_n8494);
xor_3  g06147(n779, new_n8495, new_n8490);
nor_4  g06148(new_n8497, n17458, new_n7022);
xor_3  g06149(new_n8498, n17458, new_n7022);
not_3  g06150(new_n8499, new_n8498);
nor_4  g06151(new_n8500, new_n7071, n1222);
not_3  g06152(new_n8501, n1222);
xor_3  g06153(new_n8502, n2816, new_n8501);
not_3  g06154(new_n8503, n25240);
nand_4 g06155(new_n8504, new_n8503, n20359);
xor_3  g06156(new_n8505_1, n25240, new_n7076);
not_3  g06157(new_n8506, n10125);
nand_4 g06158(new_n8507, new_n8506, n4409);
xor_3  g06159(new_n8508, n10125, new_n7083);
not_3  g06160(new_n8509, n8067);
nand_4 g06161(new_n8510_1, new_n8509, n3570);
xor_3  g06162(new_n8511, n8067, new_n7087);
nor_4  g06163(new_n8512, n20923, new_n4744);
not_3  g06164(new_n8513, new_n8512);
xor_3  g06165(new_n8514, n20923, n13668);
not_3  g06166(new_n8515, new_n8514);
not_3  g06167(new_n8516, n21276);
nor_4  g06168(new_n8517, new_n8516, n18157);
not_3  g06169(new_n8518, new_n8517);
not_3  g06170(new_n8519_1, n18157);
nor_4  g06171(new_n8520, n21276, new_n8519_1);
nor_4  g06172(new_n8521, new_n8520, new_n8517);
nor_4  g06173(new_n8522, n26748, new_n7792);
nor_4  g06174(new_n8523, new_n4745_1, n12161);
not_3  g06175(new_n8524, n5026);
nor_4  g06176(new_n8525, n10057, new_n8524);
nor_4  g06177(new_n8526_1, new_n7104, n5026);
nand_4 g06178(new_n8527, new_n6768, n8581);
nor_4  g06179(new_n8528, new_n8527, new_n8526_1);
nor_4  g06180(new_n8529, new_n8528, new_n8525);
nor_4  g06181(new_n8530, new_n8529, new_n8523);
nor_4  g06182(new_n8531, new_n8530, new_n8522);
nand_4 g06183(new_n8532, new_n8531, new_n8521);
nand_4 g06184(new_n8533, new_n8532, new_n8518);
nand_4 g06185(new_n8534, new_n8533, new_n8515);
nand_4 g06186(new_n8535_1, new_n8534, new_n8513);
nand_4 g06187(new_n8536, new_n8535_1, new_n8511);
nand_4 g06188(new_n8537, new_n8536, new_n8510_1);
nand_4 g06189(new_n8538, new_n8537, new_n8508);
nand_4 g06190(new_n8539, new_n8538, new_n8507);
nand_4 g06191(new_n8540, new_n8539, new_n8505_1);
nand_4 g06192(new_n8541, new_n8540, new_n8504);
nand_4 g06193(new_n8542, new_n8541, new_n8502);
not_3  g06194(new_n8543, new_n8542);
nor_4  g06195(new_n8544, new_n8543, new_n8500);
nor_4  g06196(new_n8545, new_n8544, new_n8499);
nor_4  g06197(new_n8546, new_n8545, new_n8497);
not_3  g06198(new_n8547, n26986);
nor_4  g06199(new_n8548, new_n8547, n19282);
not_3  g06200(new_n8549, n19282);
xor_3  g06201(new_n8550_1, n26986, new_n8549);
not_3  g06202(new_n8551, new_n8550_1);
nor_4  g06203(new_n8552, new_n8205, n12657);
not_3  g06204(new_n8553, n12657);
xor_3  g06205(new_n8554, n21287, new_n8553);
not_3  g06206(new_n8555, n17077);
nand_4 g06207(new_n8556, new_n8555, n4256);
xor_3  g06208(new_n8557, n17077, new_n8207);
nand_4 g06209(new_n8558, new_n3081, n22332);
nand_4 g06210(new_n8559, new_n4217, new_n4186_1);
nand_4 g06211(new_n8560, new_n8559, new_n8558);
nand_4 g06212(new_n8561, new_n8560, new_n8557);
nand_4 g06213(new_n8562, new_n8561, new_n8556);
nand_4 g06214(new_n8563_1, new_n8562, new_n8554);
not_3  g06215(new_n8564, new_n8563_1);
nor_4  g06216(new_n8565, new_n8564, new_n8552);
nor_4  g06217(new_n8566, new_n8565, new_n8551);
nor_4  g06218(new_n8567, new_n8566, new_n8548);
xor_3  g06219(new_n8568, new_n8567, new_n8546);
not_3  g06220(new_n8569, new_n8544);
nor_4  g06221(new_n8570, new_n8569, new_n8498);
nor_4  g06222(new_n8571, new_n8570, new_n8545);
not_3  g06223(new_n8572, new_n8571);
xor_3  g06224(new_n8573, new_n8565, new_n8551);
not_3  g06225(new_n8574, new_n8573);
nor_4  g06226(new_n8575, new_n8574, new_n8572);
xnor_3 g06227(new_n8576, new_n8573, new_n8571);
nor_4  g06228(new_n8577, new_n8541, new_n8502);
nor_4  g06229(new_n8578, new_n8577, new_n8543);
nor_4  g06230(new_n8579, new_n8562, new_n8554);
nor_4  g06231(new_n8580, new_n8579, new_n8564);
nor_4  g06232(new_n8581_1, new_n8580, new_n8578);
not_3  g06233(new_n8582, new_n8581_1);
not_3  g06234(new_n8583, new_n8578);
not_3  g06235(new_n8584, new_n8580);
nor_4  g06236(new_n8585, new_n8584, new_n8583);
nor_4  g06237(new_n8586, new_n8585, new_n8581_1);
xnor_3 g06238(new_n8587, new_n8539, new_n8505_1);
not_3  g06239(new_n8588, new_n8587);
xnor_3 g06240(new_n8589, new_n8560, new_n8557);
not_3  g06241(new_n8590, new_n8589);
nor_4  g06242(new_n8591, new_n8590, new_n8588);
not_3  g06243(new_n8592, new_n8591);
nor_4  g06244(new_n8593, new_n8589, new_n8587);
nor_4  g06245(new_n8594_1, new_n8593, new_n8591);
not_3  g06246(new_n8595, new_n8508);
xnor_3 g06247(new_n8596, new_n8537, new_n8595);
not_3  g06248(new_n8597, new_n8596);
nand_4 g06249(new_n8598, new_n8597, new_n4218);
xnor_3 g06250(new_n8599, new_n8596, new_n4218);
xnor_3 g06251(new_n8600, new_n8535_1, new_n8511);
nand_4 g06252(new_n8601, new_n8600, new_n4230);
not_3  g06253(new_n8602, new_n8600);
xnor_3 g06254(new_n8603, new_n8602, new_n4230);
xnor_3 g06255(new_n8604, new_n8533, new_n8514);
nor_4  g06256(new_n8605, new_n8604, new_n4237);
not_3  g06257(new_n8606, new_n8605);
not_3  g06258(new_n8607, new_n8604);
nor_4  g06259(new_n8608_1, new_n8607, new_n4242);
nor_4  g06260(new_n8609, new_n8608_1, new_n8605);
xnor_3 g06261(new_n8610, new_n8531, new_n8521);
not_3  g06262(new_n8611, new_n8610);
nor_4  g06263(new_n8612, new_n8611, new_n4250);
not_3  g06264(new_n8613, new_n8612);
nor_4  g06265(new_n8614_1, new_n8610, new_n4253);
nor_4  g06266(new_n8615, new_n8614_1, new_n8612);
nor_4  g06267(new_n8616, new_n8523, new_n8522);
xnor_3 g06268(new_n8617, new_n8616, new_n8529);
not_3  g06269(new_n8618, new_n8617);
nor_4  g06270(new_n8619, new_n8618, new_n4259);
not_3  g06271(new_n8620_1, new_n8619);
nor_4  g06272(new_n8621, new_n8617, new_n4260);
nor_4  g06273(new_n8622, new_n8621, new_n8619);
nor_4  g06274(new_n8623, new_n8526_1, new_n8525);
xnor_3 g06275(new_n8624, new_n8623, new_n8527);
nor_4  g06276(new_n8625, new_n8624, new_n4266_1);
not_3  g06277(new_n8626, n8581);
xnor_3 g06278(new_n8627, n8920, new_n8626);
nand_4 g06279(new_n8628, new_n8627, new_n4268);
not_3  g06280(new_n8629, new_n8624);
nor_4  g06281(new_n8630, new_n8629, new_n4270);
nor_4  g06282(new_n8631, new_n8630, new_n8625);
not_3  g06283(new_n8632, new_n8631);
nor_4  g06284(new_n8633, new_n8632, new_n8628);
nor_4  g06285(new_n8634, new_n8633, new_n8625);
nand_4 g06286(new_n8635, new_n8634, new_n8622);
nand_4 g06287(new_n8636, new_n8635, new_n8620_1);
nand_4 g06288(new_n8637_1, new_n8636, new_n8615);
nand_4 g06289(new_n8638_1, new_n8637_1, new_n8613);
nand_4 g06290(new_n8639, new_n8638_1, new_n8609);
nand_4 g06291(new_n8640, new_n8639, new_n8606);
nand_4 g06292(new_n8641, new_n8640, new_n8603);
nand_4 g06293(new_n8642, new_n8641, new_n8601);
nand_4 g06294(new_n8643, new_n8642, new_n8599);
nand_4 g06295(new_n8644, new_n8643, new_n8598);
nand_4 g06296(new_n8645, new_n8644, new_n8594_1);
nand_4 g06297(new_n8646, new_n8645, new_n8592);
nand_4 g06298(new_n8647, new_n8646, new_n8586);
nand_4 g06299(new_n8648, new_n8647, new_n8582);
nor_4  g06300(new_n8649, new_n8648, new_n8576);
nor_4  g06301(new_n8650, new_n8649, new_n8575);
xnor_3 g06302(new_n8651, new_n8650, new_n8568);
not_3  g06303(new_n8652, new_n8651);
nor_4  g06304(new_n8653, n11898, new_n6863_1);
xor_3  g06305(new_n8654, n11898, new_n6863_1);
not_3  g06306(new_n8655, new_n8654);
not_3  g06307(new_n8656_1, n647);
nor_4  g06308(new_n8657, n19941, new_n8656_1);
xor_3  g06309(new_n8658, n19941, new_n8656_1);
not_3  g06310(new_n8659, n20409);
nor_4  g06311(new_n8660, new_n8659, n1099);
not_3  g06312(new_n8661, new_n8660);
not_3  g06313(new_n8662_1, n1099);
xor_3  g06314(new_n8663, n20409, new_n8662_1);
nor_4  g06315(new_n8664, new_n5472_1, n2113);
not_3  g06316(new_n8665, new_n8664);
xor_3  g06317(new_n8666, n25749, new_n4074);
nor_4  g06318(new_n8667, n21134, new_n4136);
not_3  g06319(new_n8668, new_n8667);
xor_3  g06320(new_n8669, n21134, new_n4136);
nor_4  g06321(new_n8670, new_n4141, n6369);
xor_3  g06322(new_n8671, n9003, new_n4075);
not_3  g06323(new_n8672, new_n8671);
nor_4  g06324(new_n8673, n25797, new_n4148);
xor_3  g06325(new_n8674, n25797, n4957);
nor_4  g06326(new_n8675, new_n4076, n7524);
nor_4  g06327(new_n8676, n15967, new_n4155);
nor_4  g06328(new_n8677, n15743, new_n4687);
nand_4 g06329(new_n8678_1, n15743, new_n4687);
not_3  g06330(new_n8679, new_n8678_1);
not_3  g06331(new_n8680, n25435);
nor_4  g06332(new_n8681, new_n8680, n20658);
not_3  g06333(new_n8682, new_n8681);
nor_4  g06334(new_n8683, new_n8682, new_n8679);
nor_4  g06335(new_n8684, new_n8683, new_n8677);
nor_4  g06336(new_n8685, new_n8684, new_n8676);
nor_4  g06337(new_n8686, new_n8685, new_n8675);
not_3  g06338(new_n8687_1, new_n8686);
nor_4  g06339(new_n8688, new_n8687_1, new_n8674);
nor_4  g06340(new_n8689, new_n8688, new_n8673);
nor_4  g06341(new_n8690, new_n8689, new_n8672);
nor_4  g06342(new_n8691, new_n8690, new_n8670);
not_3  g06343(new_n8692, new_n8691);
nand_4 g06344(new_n8693, new_n8692, new_n8669);
nand_4 g06345(new_n8694_1, new_n8693, new_n8668);
nand_4 g06346(new_n8695, new_n8694_1, new_n8666);
nand_4 g06347(new_n8696, new_n8695, new_n8665);
nand_4 g06348(new_n8697, new_n8696, new_n8663);
nand_4 g06349(new_n8698, new_n8697, new_n8661);
nand_4 g06350(new_n8699, new_n8698, new_n8658);
not_3  g06351(new_n8700, new_n8699);
nor_4  g06352(new_n8701, new_n8700, new_n8657);
nor_4  g06353(new_n8702, new_n8701, new_n8655);
nor_4  g06354(new_n8703, new_n8702, new_n8653);
not_3  g06355(new_n8704, new_n8703);
nor_4  g06356(new_n8705, new_n8704, new_n8652);
nor_4  g06357(new_n8706, new_n8703, new_n8651);
nor_4  g06358(new_n8707, new_n8706, new_n8705);
xor_3  g06359(new_n8708, new_n8701, new_n8654);
xnor_3 g06360(new_n8709, new_n8648, new_n8576);
nand_4 g06361(new_n8710, new_n8709, new_n8708);
not_3  g06362(new_n8711, new_n8709);
xnor_3 g06363(new_n8712, new_n8711, new_n8708);
xnor_3 g06364(new_n8713, new_n8698, new_n8658);
xnor_3 g06365(new_n8714, new_n8646, new_n8586);
not_3  g06366(new_n8715, new_n8714);
nand_4 g06367(new_n8716_1, new_n8715, new_n8713);
xnor_3 g06368(new_n8717, new_n8714, new_n8713);
xor_3  g06369(new_n8718, new_n8696, new_n8663);
not_3  g06370(new_n8719, new_n8645);
nor_4  g06371(new_n8720, new_n8644, new_n8594_1);
nor_4  g06372(new_n8721_1, new_n8720, new_n8719);
not_3  g06373(new_n8722, new_n8721_1);
nor_4  g06374(new_n8723, new_n8722, new_n8718);
not_3  g06375(new_n8724, new_n8723);
not_3  g06376(new_n8725, new_n8718);
nor_4  g06377(new_n8726, new_n8721_1, new_n8725);
nor_4  g06378(new_n8727, new_n8726, new_n8723);
not_3  g06379(new_n8728, new_n8666);
xor_3  g06380(new_n8729, new_n8694_1, new_n8728);
xnor_3 g06381(new_n8730, new_n8642, new_n8599);
not_3  g06382(new_n8731, new_n8730);
nand_4 g06383(new_n8732, new_n8731, new_n8729);
xnor_3 g06384(new_n8733, new_n8730, new_n8729);
xor_3  g06385(new_n8734, new_n8692, new_n8669);
not_3  g06386(new_n8735, new_n8734);
not_3  g06387(new_n8736, new_n8603);
xnor_3 g06388(new_n8737, new_n8640, new_n8736);
nand_4 g06389(new_n8738, new_n8737, new_n8735);
xnor_3 g06390(new_n8739, new_n8737, new_n8734);
xor_3  g06391(new_n8740, new_n8689, new_n8672);
not_3  g06392(new_n8741, new_n8740);
not_3  g06393(new_n8742, new_n8609);
xnor_3 g06394(new_n8743, new_n8638_1, new_n8742);
nand_4 g06395(new_n8744_1, new_n8743, new_n8741);
xnor_3 g06396(new_n8745_1, new_n8743, new_n8740);
xnor_3 g06397(new_n8746, new_n8636, new_n8615);
not_3  g06398(new_n8747, new_n8746);
xor_3  g06399(new_n8748, new_n8686, new_n8674);
nand_4 g06400(new_n8749, new_n8748, new_n8747);
not_3  g06401(new_n8750, new_n8622);
xnor_3 g06402(new_n8751, new_n8634, new_n8750);
xor_3  g06403(new_n8752, n15967, n7524);
xor_3  g06404(new_n8753, new_n8752, new_n8684);
nand_4 g06405(new_n8754, new_n8753, new_n8751);
not_3  g06406(new_n8755, new_n8753);
xnor_3 g06407(new_n8756, new_n8755, new_n8751);
xor_3  g06408(new_n8757, n25435, new_n4167);
xnor_3 g06409(new_n8758, new_n8627, new_n4268);
nor_4  g06410(new_n8759, new_n8758, new_n8757);
nor_4  g06411(new_n8760, new_n8679, new_n8677);
xor_3  g06412(new_n8761, new_n8760, new_n8681);
not_3  g06413(new_n8762, new_n8761);
nor_4  g06414(new_n8763, new_n8762, new_n8759);
not_3  g06415(new_n8764, new_n8763);
xnor_3 g06416(new_n8765, new_n8632, new_n8628);
not_3  g06417(new_n8766, new_n8759);
nor_4  g06418(new_n8767, new_n8761, new_n8766);
nor_4  g06419(new_n8768, new_n8767, new_n8763);
nand_4 g06420(new_n8769, new_n8768, new_n8765);
nand_4 g06421(new_n8770, new_n8769, new_n8764);
nand_4 g06422(new_n8771, new_n8770, new_n8756);
nand_4 g06423(new_n8772, new_n8771, new_n8754);
xnor_3 g06424(new_n8773, new_n8748, new_n8746);
nand_4 g06425(new_n8774, new_n8773, new_n8772);
nand_4 g06426(new_n8775, new_n8774, new_n8749);
nand_4 g06427(new_n8776, new_n8775, new_n8745_1);
nand_4 g06428(new_n8777, new_n8776, new_n8744_1);
nand_4 g06429(new_n8778, new_n8777, new_n8739);
nand_4 g06430(new_n8779, new_n8778, new_n8738);
nand_4 g06431(new_n8780, new_n8779, new_n8733);
nand_4 g06432(new_n8781, new_n8780, new_n8732);
nand_4 g06433(new_n8782_1, new_n8781, new_n8727);
nand_4 g06434(new_n8783, new_n8782_1, new_n8724);
nand_4 g06435(new_n8784, new_n8783, new_n8717);
nand_4 g06436(new_n8785, new_n8784, new_n8716_1);
nand_4 g06437(new_n8786, new_n8785, new_n8712);
nand_4 g06438(new_n8787, new_n8786, new_n8710);
xnor_3 g06439(n809, new_n8787, new_n8707);
not_3  g06440(new_n8789, n2978);
nor_4  g06441(new_n8790, n19282, new_n8789);
xor_3  g06442(new_n8791, n19282, new_n8789);
not_3  g06443(new_n8792, new_n8791);
not_3  g06444(new_n8793, n23697);
nor_4  g06445(new_n8794, new_n8793, n12657);
xor_3  g06446(new_n8795, n23697, new_n8553);
not_3  g06447(new_n8796, n2289);
nor_4  g06448(new_n8797, n17077, new_n8796);
not_3  g06449(new_n8798, new_n8797);
xor_3  g06450(new_n8799, n17077, new_n8796);
nor_4  g06451(new_n8800, n26510, new_n7937_1);
not_3  g06452(new_n8801, new_n8800);
xor_3  g06453(new_n8802, n26510, new_n7937_1);
not_3  g06454(new_n8803_1, n20179);
nor_4  g06455(new_n8804, n23068, new_n8803_1);
not_3  g06456(new_n8805, new_n8804);
xor_3  g06457(new_n8806_1, n23068, new_n8803_1);
not_3  g06458(new_n8807, n19228);
nor_4  g06459(new_n8808, n19514, new_n8807);
xor_3  g06460(new_n8809_1, n19514, new_n8807);
not_3  g06461(new_n8810, new_n8809_1);
not_3  g06462(new_n8811, n15539);
nor_4  g06463(new_n8812, new_n8811, n10053);
xor_3  g06464(new_n8813, n15539, n10053);
nor_4  g06465(new_n8814, new_n4199, n8052);
not_3  g06466(new_n8815, n8052);
nor_4  g06467(new_n8816, n8399, new_n8815);
nor_4  g06468(new_n8817, n10158, new_n4203);
nand_4 g06469(new_n8818, n10158, new_n4203);
not_3  g06470(new_n8819, new_n8818);
not_3  g06471(new_n8820, n26979);
nor_4  g06472(new_n8821_1, new_n8820, n18962);
not_3  g06473(new_n8822, new_n8821_1);
nor_4  g06474(new_n8823, new_n8822, new_n8819);
nor_4  g06475(new_n8824_1, new_n8823, new_n8817);
nor_4  g06476(new_n8825, new_n8824_1, new_n8816);
nor_4  g06477(new_n8826, new_n8825, new_n8814);
not_3  g06478(new_n8827_1, new_n8826);
nor_4  g06479(new_n8828, new_n8827_1, new_n8813);
nor_4  g06480(new_n8829, new_n8828, new_n8812);
nor_4  g06481(new_n8830, new_n8829, new_n8810);
nor_4  g06482(new_n8831, new_n8830, new_n8808);
not_3  g06483(new_n8832, new_n8831);
nand_4 g06484(new_n8833, new_n8832, new_n8806_1);
nand_4 g06485(new_n8834, new_n8833, new_n8805);
nand_4 g06486(new_n8835, new_n8834, new_n8802);
nand_4 g06487(new_n8836, new_n8835, new_n8801);
nand_4 g06488(new_n8837, new_n8836, new_n8799);
nand_4 g06489(new_n8838, new_n8837, new_n8798);
nand_4 g06490(new_n8839, new_n8838, new_n8795);
not_3  g06491(new_n8840, new_n8839);
nor_4  g06492(new_n8841, new_n8840, new_n8794);
nor_4  g06493(new_n8842, new_n8841, new_n8792);
nor_4  g06494(new_n8843, new_n8842, new_n8790);
not_3  g06495(new_n8844, new_n8843);
nor_4  g06496(new_n8845, n26986, n22626);
not_3  g06497(new_n8846, new_n8845);
nand_4 g06498(new_n8847, new_n2448, new_n2440_1);
xor_3  g06499(new_n8848, n4256, n1654);
not_3  g06500(new_n8849_1, n13783);
nand_4 g06501(new_n8850, new_n4185, new_n8849_1);
nand_4 g06502(new_n8851, new_n2447, new_n2441);
nand_4 g06503(new_n8852, new_n8851, new_n8850);
xnor_3 g06504(new_n8853, new_n8852, new_n8848);
nor_4  g06505(new_n8854, new_n8853, new_n8847);
xor_3  g06506(new_n8855, n21287, n14440);
nor_4  g06507(new_n8856_1, n4256, n1654);
not_3  g06508(new_n8857, new_n8848);
not_3  g06509(new_n8858, new_n8852);
nor_4  g06510(new_n8859, new_n8858, new_n8857);
nor_4  g06511(new_n8860, new_n8859, new_n8856_1);
xnor_3 g06512(new_n8861_1, new_n8860, new_n8855);
nand_4 g06513(new_n8862_1, new_n8861_1, new_n8854);
xor_3  g06514(new_n8863, n26986, n22626);
not_3  g06515(new_n8864, new_n8863);
nor_4  g06516(new_n8865, n21287, n14440);
not_3  g06517(new_n8866, new_n8855);
nor_4  g06518(new_n8867, new_n8860, new_n8866);
nor_4  g06519(new_n8868, new_n8867, new_n8865);
xnor_3 g06520(new_n8869_1, new_n8868, new_n8864);
nor_4  g06521(new_n8870, new_n8869_1, new_n8862_1);
not_3  g06522(new_n8871, new_n8870);
nor_4  g06523(new_n8872, new_n8871, new_n8846);
nor_4  g06524(new_n8873, new_n8868, new_n8864);
nor_4  g06525(new_n8874, new_n8873, new_n8845);
not_3  g06526(new_n8875, new_n8874);
nor_4  g06527(new_n8876, new_n8875, new_n8870);
nor_4  g06528(new_n8877, new_n8876, new_n8872);
not_3  g06529(new_n8878, new_n8877);
nor_4  g06530(new_n8879, n13494, n3425);
xor_3  g06531(new_n8880, n13494, n3425);
not_3  g06532(new_n8881, new_n8880);
nor_4  g06533(new_n8882, n25345, n9967);
xor_3  g06534(new_n8883, n25345, n9967);
not_3  g06535(new_n8884_1, n20946);
nand_4 g06536(new_n8885, new_n8884_1, new_n6385_1);
xor_3  g06537(new_n8886, n20946, n9655);
nor_4  g06538(new_n8887, n13490, n7751);
not_3  g06539(new_n8888, new_n8887);
nand_4 g06540(new_n8889, new_n2482, new_n2450);
nand_4 g06541(new_n8890, new_n8889, new_n8888);
nand_4 g06542(new_n8891, new_n8890, new_n8886);
nand_4 g06543(new_n8892, new_n8891, new_n8885);
nand_4 g06544(new_n8893, new_n8892, new_n8883);
not_3  g06545(new_n8894, new_n8893);
nor_4  g06546(new_n8895, new_n8894, new_n8882);
nor_4  g06547(new_n8896, new_n8895, new_n8881);
nor_4  g06548(new_n8897, new_n8896, new_n8879);
not_3  g06549(new_n8898, new_n8897);
nor_4  g06550(new_n8899, new_n8898, new_n8878);
nor_4  g06551(new_n8900, new_n8897, new_n8877);
xnor_3 g06552(new_n8901, new_n8869_1, new_n8862_1);
not_3  g06553(new_n8902, new_n8901);
xnor_3 g06554(new_n8903, new_n8895, new_n8880);
not_3  g06555(new_n8904, new_n8903);
nor_4  g06556(new_n8905, new_n8904, new_n8902);
not_3  g06557(new_n8906, new_n8905);
nor_4  g06558(new_n8907, new_n8903, new_n8901);
nor_4  g06559(new_n8908, new_n8907, new_n8905);
xnor_3 g06560(new_n8909_1, new_n8861_1, new_n8854);
nor_4  g06561(new_n8910, new_n8892, new_n8883);
nor_4  g06562(new_n8911_1, new_n8910, new_n8894);
nand_4 g06563(new_n8912, new_n8911_1, new_n8909_1);
not_3  g06564(new_n8913, new_n8912);
nor_4  g06565(new_n8914, new_n8911_1, new_n8909_1);
nor_4  g06566(new_n8915, new_n8914, new_n8913);
xnor_3 g06567(new_n8916, new_n8853, new_n8847);
xnor_3 g06568(new_n8917, new_n8890, new_n8886);
not_3  g06569(new_n8918, new_n8917);
nand_4 g06570(new_n8919, new_n8918, new_n8916);
not_3  g06571(new_n8920_1, new_n8919);
nor_4  g06572(new_n8921, new_n8918, new_n8916);
nor_4  g06573(new_n8922, new_n8921, new_n8920_1);
not_3  g06574(new_n8923, new_n2483);
nand_4 g06575(new_n8924, new_n8923, new_n2449);
nand_4 g06576(new_n8925, new_n2538, new_n2484);
nand_4 g06577(new_n8926, new_n8925, new_n8924);
nand_4 g06578(new_n8927, new_n8926, new_n8922);
nand_4 g06579(new_n8928, new_n8927, new_n8919);
nand_4 g06580(new_n8929, new_n8928, new_n8915);
nand_4 g06581(new_n8930, new_n8929, new_n8912);
nand_4 g06582(new_n8931, new_n8930, new_n8908);
nand_4 g06583(new_n8932, new_n8931, new_n8906);
nor_4  g06584(new_n8933, new_n8932, new_n8900);
nor_4  g06585(new_n8934, new_n8933, new_n8872);
not_3  g06586(new_n8935, new_n8934);
nor_4  g06587(new_n8936, new_n8935, new_n8899);
nand_4 g06588(new_n8937, new_n8936, new_n8844);
not_3  g06589(new_n8938, new_n8936);
nand_4 g06590(new_n8939, new_n8938, new_n8843);
nand_4 g06591(new_n8940, new_n8939, new_n8937);
not_3  g06592(new_n8941, new_n8932);
nor_4  g06593(new_n8942, new_n8900, new_n8899);
xnor_3 g06594(new_n8943_1, new_n8942, new_n8941);
nand_4 g06595(new_n8944, new_n8943_1, new_n8844);
xnor_3 g06596(new_n8945, new_n8943_1, new_n8843);
xor_3  g06597(new_n8946, new_n8841, new_n8792);
xnor_3 g06598(new_n8947, new_n8930, new_n8908);
nor_4  g06599(new_n8948, new_n8947, new_n8946);
not_3  g06600(new_n8949, new_n8948);
not_3  g06601(new_n8950, new_n8946);
not_3  g06602(new_n8951, new_n8908);
xnor_3 g06603(new_n8952, new_n8930, new_n8951);
nor_4  g06604(new_n8953, new_n8952, new_n8950);
nor_4  g06605(new_n8954, new_n8953, new_n8948);
xnor_3 g06606(new_n8955, new_n8838, new_n8795);
xnor_3 g06607(new_n8956, new_n8928, new_n8915);
not_3  g06608(new_n8957, new_n8956);
nand_4 g06609(new_n8958, new_n8957, new_n8955);
xnor_3 g06610(new_n8959, new_n8956, new_n8955);
not_3  g06611(new_n8960, new_n8799);
xor_3  g06612(new_n8961, new_n8836, new_n8960);
not_3  g06613(new_n8962, new_n8926);
xnor_3 g06614(new_n8963, new_n8962, new_n8922);
nand_4 g06615(new_n8964_1, new_n8963, new_n8961);
xnor_3 g06616(new_n8965, new_n8926, new_n8922);
xnor_3 g06617(new_n8966, new_n8965, new_n8961);
not_3  g06618(new_n8967, new_n8802);
xor_3  g06619(new_n8968, new_n8834, new_n8967);
nand_4 g06620(new_n8969, new_n8968, new_n2539);
xnor_3 g06621(new_n8970, new_n2538, new_n2484);
xnor_3 g06622(new_n8971_1, new_n8968, new_n8970);
xor_3  g06623(new_n8972, new_n8832, new_n8806_1);
nor_4  g06624(new_n8973, new_n8972, new_n2542);
not_3  g06625(new_n8974, new_n8973);
not_3  g06626(new_n8975, new_n8972);
nor_4  g06627(new_n8976, new_n8975, new_n2545);
nor_4  g06628(new_n8977, new_n8976, new_n8973);
xor_3  g06629(new_n8978, new_n8829, new_n8810);
nor_4  g06630(new_n8979, new_n8978, new_n2548);
not_3  g06631(new_n8980, new_n8979);
not_3  g06632(new_n8981, new_n8978);
nor_4  g06633(new_n8982_1, new_n8981, new_n2552);
nor_4  g06634(new_n8983, new_n8982_1, new_n8979);
xor_3  g06635(new_n8984, new_n8826, new_n8813);
nand_4 g06636(new_n8985, new_n8984, new_n2560_1);
not_3  g06637(new_n8986, new_n8985);
nor_4  g06638(new_n8987, new_n8984, new_n2560_1);
nor_4  g06639(new_n8988, new_n8987, new_n8986);
not_3  g06640(new_n8989, new_n8824_1);
nor_4  g06641(new_n8990, new_n8816, new_n8814);
xor_3  g06642(new_n8991, new_n8990, new_n8989);
not_3  g06643(new_n8992, new_n8991);
nor_4  g06644(new_n8993_1, new_n8992, new_n2563);
not_3  g06645(new_n8994, new_n8993_1);
nor_4  g06646(new_n8995, new_n8991, new_n2569);
nor_4  g06647(new_n8996, new_n8995, new_n8993_1);
not_3  g06648(new_n8997, n18962);
xor_3  g06649(new_n8998, n26979, new_n8997);
nor_4  g06650(new_n8999, new_n8998, new_n2574);
nor_4  g06651(new_n9000, new_n8819, new_n8817);
xor_3  g06652(new_n9001, new_n9000, new_n8821_1);
not_3  g06653(new_n9002, new_n9001);
nor_4  g06654(new_n9003_1, new_n9002, new_n8999);
not_3  g06655(new_n9004, new_n9003_1);
not_3  g06656(new_n9005, new_n2579);
not_3  g06657(new_n9006, new_n8999);
nor_4  g06658(new_n9007, new_n9001, new_n9006);
nor_4  g06659(new_n9008, new_n9007, new_n9003_1);
nand_4 g06660(new_n9009, new_n9008, new_n9005);
nand_4 g06661(new_n9010, new_n9009, new_n9004);
nand_4 g06662(new_n9011, new_n9010, new_n8996);
nand_4 g06663(new_n9012_1, new_n9011, new_n8994);
nand_4 g06664(new_n9013, new_n9012_1, new_n8988);
nand_4 g06665(new_n9014, new_n9013, new_n8985);
nand_4 g06666(new_n9015, new_n9014, new_n8983);
nand_4 g06667(new_n9016, new_n9015, new_n8980);
nand_4 g06668(new_n9017, new_n9016, new_n8977);
nand_4 g06669(new_n9018, new_n9017, new_n8974);
nand_4 g06670(new_n9019, new_n9018, new_n8971_1);
nand_4 g06671(new_n9020, new_n9019, new_n8969);
nand_4 g06672(new_n9021, new_n9020, new_n8966);
nand_4 g06673(new_n9022, new_n9021, new_n8964_1);
nand_4 g06674(new_n9023, new_n9022, new_n8959);
nand_4 g06675(new_n9024, new_n9023, new_n8958);
nand_4 g06676(new_n9025, new_n9024, new_n8954);
nand_4 g06677(new_n9026, new_n9025, new_n8949);
nand_4 g06678(new_n9027, new_n9026, new_n8945);
nand_4 g06679(new_n9028, new_n9027, new_n8944);
xnor_3 g06680(n819, new_n9028, new_n8940);
nor_4  g06681(new_n9030, n22626, new_n3662);
xor_3  g06682(new_n9031, n22626, new_n3662);
not_3  g06683(new_n9032_1, new_n9031);
not_3  g06684(new_n9033, n14130);
nor_4  g06685(new_n9034, n14440, new_n9033);
xor_3  g06686(new_n9035, n14440, new_n9033);
not_3  g06687(new_n9036, n1654);
nand_4 g06688(new_n9037, n16482, new_n9036);
xor_3  g06689(new_n9038, n16482, new_n9036);
nand_4 g06690(new_n9039, new_n8849_1, n9942);
xor_3  g06691(new_n9040, n13783, new_n2349);
nand_4 g06692(new_n9041, new_n2444_1, n25643);
xor_3  g06693(new_n9042_1, n26660, new_n2352);
nor_4  g06694(new_n9043, new_n2359, n3018);
not_3  g06695(new_n9044, new_n9043);
not_3  g06696(new_n9045, n3018);
xor_3  g06697(new_n9046_1, n9557, new_n9045);
nor_4  g06698(new_n9047_1, n3480, new_n2364);
not_3  g06699(new_n9048, new_n9047_1);
xor_3  g06700(new_n9049, n3480, new_n2364);
not_3  g06701(new_n9050, n16722);
nor_4  g06702(new_n9051, new_n9050, n6385);
nor_4  g06703(new_n9052, n16722, new_n2366);
not_3  g06704(new_n9053, n11486);
nor_4  g06705(new_n9054, n20138, new_n9053);
nor_4  g06706(new_n9055, new_n2370, n11486);
nand_4 g06707(new_n9056, n13781, new_n2374_1);
nor_4  g06708(new_n9057, new_n9056, new_n9055);
nor_4  g06709(new_n9058, new_n9057, new_n9054);
nor_4  g06710(new_n9059, new_n9058, new_n9052);
nor_4  g06711(new_n9060, new_n9059, new_n9051);
nand_4 g06712(new_n9061, new_n9060, new_n9049);
nand_4 g06713(new_n9062, new_n9061, new_n9048);
nand_4 g06714(new_n9063, new_n9062, new_n9046_1);
nand_4 g06715(new_n9064, new_n9063, new_n9044);
nand_4 g06716(new_n9065, new_n9064, new_n9042_1);
nand_4 g06717(new_n9066, new_n9065, new_n9041);
nand_4 g06718(new_n9067, new_n9066, new_n9040);
nand_4 g06719(new_n9068, new_n9067, new_n9039);
nand_4 g06720(new_n9069, new_n9068, new_n9038);
nand_4 g06721(new_n9070, new_n9069, new_n9037);
nand_4 g06722(new_n9071, new_n9070, new_n9035);
not_3  g06723(new_n9072, new_n9071);
nor_4  g06724(new_n9073, new_n9072, new_n9034);
nor_4  g06725(new_n9074, new_n9073, new_n9032_1);
nor_4  g06726(new_n9075, new_n9074, new_n9030);
not_3  g06727(new_n9076, n3582);
nor_4  g06728(new_n9077, n25120, new_n9076);
xor_3  g06729(new_n9078, n25120, new_n9076);
not_3  g06730(new_n9079, new_n9078);
not_3  g06731(new_n9080, n2145);
nor_4  g06732(new_n9081, n8363, new_n9080);
xor_3  g06733(new_n9082, n8363, new_n9080);
not_3  g06734(new_n9083, n14680);
nand_4 g06735(new_n9084, new_n9083, n5031);
not_3  g06736(new_n9085, n5031);
xor_3  g06737(new_n9086, n14680, new_n9085);
not_3  g06738(new_n9087, n17250);
nand_4 g06739(new_n9088, new_n9087, n11044);
xor_3  g06740(new_n9089, n17250, new_n7030);
not_3  g06741(new_n9090_1, n23160);
nand_4 g06742(new_n9091, new_n9090_1, n2421);
xor_3  g06743(new_n9092, n23160, new_n7033);
nor_4  g06744(new_n9093, n16524, new_n7036);
not_3  g06745(new_n9094, new_n9093);
xor_3  g06746(new_n9095, n16524, new_n7036);
nor_4  g06747(new_n9096, new_n7039, n11056);
not_3  g06748(new_n9097, new_n9096);
not_3  g06749(new_n9098, n11056);
xor_3  g06750(new_n9099, n20478, new_n9098);
not_3  g06751(new_n9100, n15271);
nor_4  g06752(new_n9101, n26882, new_n9100);
not_3  g06753(new_n9102, n26882);
nor_4  g06754(new_n9103, new_n9102, n15271);
nor_4  g06755(new_n9104_1, new_n6737, n22619);
not_3  g06756(new_n9105, n22619);
nor_4  g06757(new_n9106, n25877, new_n9105);
not_3  g06758(new_n9107, n6775);
nand_4 g06759(new_n9108, n24323, new_n9107);
nor_4  g06760(new_n9109, new_n9108, new_n9106);
nor_4  g06761(new_n9110, new_n9109, new_n9104_1);
nor_4  g06762(new_n9111, new_n9110, new_n9103);
nor_4  g06763(new_n9112, new_n9111, new_n9101);
nand_4 g06764(new_n9113, new_n9112, new_n9099);
nand_4 g06765(new_n9114, new_n9113, new_n9097);
nand_4 g06766(new_n9115, new_n9114, new_n9095);
nand_4 g06767(new_n9116, new_n9115, new_n9094);
nand_4 g06768(new_n9117, new_n9116, new_n9092);
nand_4 g06769(new_n9118, new_n9117, new_n9091);
nand_4 g06770(new_n9119, new_n9118, new_n9089);
nand_4 g06771(new_n9120, new_n9119, new_n9088);
nand_4 g06772(new_n9121, new_n9120, new_n9086);
nand_4 g06773(new_n9122, new_n9121, new_n9084);
nand_4 g06774(new_n9123, new_n9122, new_n9082);
not_3  g06775(new_n9124, new_n9123);
nor_4  g06776(new_n9125, new_n9124, new_n9081);
nor_4  g06777(new_n9126, new_n9125, new_n9079);
nor_4  g06778(new_n9127, new_n9126, new_n9077);
xor_3  g06779(new_n9128, new_n9127, new_n9075);
xor_3  g06780(new_n9129_1, new_n9125, new_n9078);
not_3  g06781(new_n9130, new_n9129_1);
and_4  g06782(new_n9131, new_n9073, new_n9032_1);
nor_4  g06783(new_n9132, new_n9131, new_n9074);
nor_4  g06784(new_n9133, new_n9132, new_n9130);
not_3  g06785(new_n9134, new_n9133);
not_3  g06786(new_n9135, new_n9132);
xnor_3 g06787(new_n9136, new_n9135, new_n9129_1);
not_3  g06788(new_n9137, new_n9136);
nor_4  g06789(new_n9138, new_n9122, new_n9082);
nor_4  g06790(new_n9139, new_n9138, new_n9124);
nor_4  g06791(new_n9140, new_n9070, new_n9035);
nor_4  g06792(new_n9141, new_n9140, new_n9072);
nor_4  g06793(new_n9142, new_n9141, new_n9139);
not_3  g06794(new_n9143, new_n9142);
not_3  g06795(new_n9144, new_n9139);
not_3  g06796(new_n9145, new_n9141);
nor_4  g06797(new_n9146_1, new_n9145, new_n9144);
nor_4  g06798(new_n9147, new_n9146_1, new_n9142);
not_3  g06799(new_n9148, new_n9086);
xnor_3 g06800(new_n9149, new_n9120, new_n9148);
not_3  g06801(new_n9150, new_n9038);
xnor_3 g06802(new_n9151, new_n9068, new_n9150);
nor_4  g06803(new_n9152, new_n9151, new_n9149);
not_3  g06804(new_n9153, new_n9152);
not_3  g06805(new_n9154, new_n9149);
xnor_3 g06806(new_n9155, new_n9068, new_n9038);
nor_4  g06807(new_n9156, new_n9155, new_n9154);
nor_4  g06808(new_n9157, new_n9156, new_n9152);
not_3  g06809(new_n9158, new_n9089);
xnor_3 g06810(new_n9159, new_n9118, new_n9158);
not_3  g06811(new_n9160, new_n9040);
xnor_3 g06812(new_n9161, new_n9066, new_n9160);
nor_4  g06813(new_n9162, new_n9161, new_n9159);
not_3  g06814(new_n9163, new_n9162);
not_3  g06815(new_n9164_1, new_n9159);
xnor_3 g06816(new_n9165, new_n9066, new_n9040);
nor_4  g06817(new_n9166_1, new_n9165, new_n9164_1);
nor_4  g06818(new_n9167, new_n9166_1, new_n9162);
not_3  g06819(new_n9168, new_n9092);
not_3  g06820(new_n9169, new_n9095);
xor_3  g06821(new_n9170, n20478, n11056);
not_3  g06822(new_n9171, new_n9112);
nor_4  g06823(new_n9172_1, new_n9171, new_n9170);
nor_4  g06824(new_n9173, new_n9172_1, new_n9096);
nor_4  g06825(new_n9174, new_n9173, new_n9169);
nor_4  g06826(new_n9175, new_n9174, new_n9093);
xnor_3 g06827(new_n9176, new_n9175, new_n9168);
not_3  g06828(new_n9177, new_n9176);
not_3  g06829(new_n9178, new_n9042_1);
xnor_3 g06830(new_n9179, new_n9064, new_n9178);
nor_4  g06831(new_n9180, new_n9179, new_n9177);
not_3  g06832(new_n9181, new_n9180);
xnor_3 g06833(new_n9182_1, new_n9064, new_n9042_1);
nor_4  g06834(new_n9183, new_n9182_1, new_n9176);
nor_4  g06835(new_n9184, new_n9183, new_n9180);
xnor_3 g06836(new_n9185, new_n9173, new_n9169);
not_3  g06837(new_n9186, new_n9185);
not_3  g06838(new_n9187, new_n9046_1);
xnor_3 g06839(new_n9188, new_n9062, new_n9187);
nor_4  g06840(new_n9189, new_n9188, new_n9186);
not_3  g06841(new_n9190, new_n9189);
xnor_3 g06842(new_n9191_1, new_n9062, new_n9046_1);
nor_4  g06843(new_n9192, new_n9191_1, new_n9185);
nor_4  g06844(new_n9193, new_n9192, new_n9189);
xnor_3 g06845(new_n9194, new_n9171, new_n9170);
not_3  g06846(new_n9195, new_n9194);
not_3  g06847(new_n9196, new_n9060);
xnor_3 g06848(new_n9197, new_n9196, new_n9049);
nor_4  g06849(new_n9198, new_n9197, new_n9195);
not_3  g06850(new_n9199, new_n9198);
xnor_3 g06851(new_n9200, new_n9060, new_n9049);
nor_4  g06852(new_n9201, new_n9200, new_n9194);
nor_4  g06853(new_n9202, new_n9201, new_n9198);
nor_4  g06854(new_n9203, new_n9103, new_n9101);
xnor_3 g06855(new_n9204, new_n9203, new_n9110);
nor_4  g06856(new_n9205, new_n9052, new_n9051);
xnor_3 g06857(new_n9206, new_n9205, new_n9058);
nand_4 g06858(new_n9207, new_n9206, new_n9204);
xnor_3 g06859(new_n9208, new_n9206, new_n9204);
not_3  g06860(new_n9209, new_n9208);
nor_4  g06861(new_n9210, new_n6722, n6775);
nor_4  g06862(new_n9211, new_n9106, new_n9104_1);
xnor_3 g06863(new_n9212, new_n9211, new_n9210);
not_3  g06864(new_n9213, new_n9212);
nor_4  g06865(new_n9214, new_n9055, new_n9054);
xnor_3 g06866(new_n9215, new_n9214, new_n9056);
nand_4 g06867(new_n9216, new_n9215, new_n9213);
nor_4  g06868(new_n9217_1, n24323, new_n9107);
nor_4  g06869(new_n9218, new_n9217_1, new_n9210);
not_3  g06870(new_n9219, new_n9056);
nor_4  g06871(new_n9220_1, n13781, new_n2374_1);
nor_4  g06872(new_n9221, new_n9220_1, new_n9219);
nor_4  g06873(new_n9222, new_n9221, new_n9218);
not_3  g06874(new_n9223, new_n9222);
not_3  g06875(new_n9224, new_n9215);
xnor_3 g06876(new_n9225, new_n9224, new_n9212);
not_3  g06877(new_n9226, new_n9225);
nand_4 g06878(new_n9227, new_n9226, new_n9223);
nand_4 g06879(new_n9228, new_n9227, new_n9216);
nand_4 g06880(new_n9229, new_n9228, new_n9209);
nand_4 g06881(new_n9230, new_n9229, new_n9207);
nand_4 g06882(new_n9231, new_n9230, new_n9202);
nand_4 g06883(new_n9232, new_n9231, new_n9199);
nand_4 g06884(new_n9233, new_n9232, new_n9193);
nand_4 g06885(new_n9234, new_n9233, new_n9190);
nand_4 g06886(new_n9235, new_n9234, new_n9184);
nand_4 g06887(new_n9236, new_n9235, new_n9181);
nand_4 g06888(new_n9237, new_n9236, new_n9167);
nand_4 g06889(new_n9238, new_n9237, new_n9163);
nand_4 g06890(new_n9239, new_n9238, new_n9157);
nand_4 g06891(new_n9240, new_n9239, new_n9153);
nand_4 g06892(new_n9241, new_n9240, new_n9147);
nand_4 g06893(new_n9242, new_n9241, new_n9143);
nand_4 g06894(new_n9243, new_n9242, new_n9137);
nand_4 g06895(new_n9244, new_n9243, new_n9134);
xnor_3 g06896(new_n9245, new_n9244, new_n9128);
not_3  g06897(new_n9246_1, n13453);
nor_4  g06898(new_n9247, n15508, n2809);
nand_4 g06899(new_n9248, new_n9247, new_n7751_1);
nor_4  g06900(new_n9249, new_n9248, n7421);
nand_4 g06901(new_n9250, new_n9249, new_n9246_1);
nor_4  g06902(new_n9251_1, new_n9250, n11630);
nand_4 g06903(new_n9252, new_n9251_1, new_n5471);
nor_4  g06904(new_n9253, new_n9252, n18227);
not_3  g06905(new_n9254, new_n9253);
nor_4  g06906(new_n9255, new_n9254, n26408);
not_3  g06907(new_n9256, new_n9255);
nor_4  g06908(new_n9257, new_n9256, n9554);
not_3  g06909(new_n9258, n9554);
xor_3  g06910(new_n9259_1, new_n9255, new_n9258);
nor_4  g06911(new_n9260, new_n9259_1, n9259);
xor_3  g06912(new_n9261_1, new_n9254, n26408);
nor_4  g06913(new_n9262, new_n9261_1, n21489);
xor_3  g06914(new_n9263, new_n9261_1, new_n3897);
xor_3  g06915(new_n9264, new_n9252, n18227);
nor_4  g06916(new_n9265, new_n9264, n20213);
xor_3  g06917(new_n9266, new_n9264, new_n5529);
xor_3  g06918(new_n9267, new_n9251_1, new_n5471);
nor_4  g06919(new_n9268, new_n9267, n13912);
not_3  g06920(new_n9269, new_n9267);
xor_3  g06921(new_n9270, new_n9269, new_n3913);
not_3  g06922(new_n9271, new_n9270);
xor_3  g06923(new_n9272, new_n9250, n11630);
nor_4  g06924(new_n9273, new_n9272, n7670);
not_3  g06925(new_n9274, new_n9272);
xor_3  g06926(new_n9275, new_n9274, new_n5535);
not_3  g06927(new_n9276, new_n9275);
xor_3  g06928(new_n9277, new_n9249, new_n9246_1);
nor_4  g06929(new_n9278, new_n9277, n9598);
not_3  g06930(new_n9279, new_n9277);
xor_3  g06931(new_n9280, new_n9279, new_n5540);
xor_3  g06932(new_n9281, new_n9248, n7421);
not_3  g06933(new_n9282, new_n9281);
nand_4 g06934(new_n9283, new_n9282, new_n5545);
xor_3  g06935(new_n9284, new_n9247, new_n7751_1);
not_3  g06936(new_n9285, new_n9284);
nand_4 g06937(new_n9286, new_n9285, new_n3943);
xor_3  g06938(new_n9287_1, new_n9285, new_n3943);
xnor_3 g06939(new_n9288, n15508, n2809);
nand_4 g06940(new_n9289, new_n9288, new_n5563);
nand_4 g06941(new_n9290, n21993, n15508);
xnor_3 g06942(new_n9291, new_n9288, n25565);
nand_4 g06943(new_n9292, new_n9291, new_n9290);
nand_4 g06944(new_n9293, new_n9292, new_n9289);
nand_4 g06945(new_n9294, new_n9293, new_n9287_1);
nand_4 g06946(new_n9295, new_n9294, new_n9286);
xor_3  g06947(new_n9296, new_n9282, new_n5545);
nand_4 g06948(new_n9297, new_n9296, new_n9295);
nand_4 g06949(new_n9298, new_n9297, new_n9283);
nand_4 g06950(new_n9299, new_n9298, new_n9280);
not_3  g06951(new_n9300, new_n9299);
nor_4  g06952(new_n9301, new_n9300, new_n9278);
nor_4  g06953(new_n9302, new_n9301, new_n9276);
nor_4  g06954(new_n9303, new_n9302, new_n9273);
nor_4  g06955(new_n9304, new_n9303, new_n9271);
nor_4  g06956(new_n9305, new_n9304, new_n9268);
nor_4  g06957(new_n9306, new_n9305, new_n9266);
nor_4  g06958(new_n9307, new_n9306, new_n9265);
nor_4  g06959(new_n9308_1, new_n9307, new_n9263);
nor_4  g06960(new_n9309, new_n9308_1, new_n9262);
and_4  g06961(new_n9310, new_n9259_1, n9259);
nor_4  g06962(new_n9311, new_n9310, new_n9309);
nor_4  g06963(new_n9312, new_n9311, new_n9260);
nor_4  g06964(new_n9313, new_n9312, new_n9257);
xnor_3 g06965(new_n9314, new_n9313, new_n9245);
not_3  g06966(new_n9315, new_n9314);
xnor_3 g06967(new_n9316, new_n9242, new_n9136);
nor_4  g06968(new_n9317, new_n9310, new_n9260);
xnor_3 g06969(new_n9318_1, new_n9317, new_n9309);
nand_4 g06970(new_n9319, new_n9318_1, new_n9316);
not_3  g06971(new_n9320, new_n9316);
xnor_3 g06972(new_n9321, new_n9318_1, new_n9320);
xnor_3 g06973(new_n9322, new_n9240, new_n9147);
not_3  g06974(new_n9323_1, new_n9322);
xnor_3 g06975(new_n9324, new_n9307, new_n9263);
not_3  g06976(new_n9325, new_n9324);
nor_4  g06977(new_n9326, new_n9325, new_n9323_1);
xnor_3 g06978(new_n9327, new_n9324, new_n9322);
xnor_3 g06979(new_n9328, new_n9238, new_n9157);
not_3  g06980(new_n9329, new_n9328);
not_3  g06981(new_n9330, new_n9305);
xnor_3 g06982(new_n9331, new_n9330, new_n9266);
nor_4  g06983(new_n9332, new_n9331, new_n9329);
xnor_3 g06984(new_n9333, new_n9331, new_n9329);
xnor_3 g06985(new_n9334, new_n9236, new_n9167);
not_3  g06986(new_n9335, new_n9334);
not_3  g06987(new_n9336, new_n9303);
nor_4  g06988(new_n9337, new_n9336, new_n9270);
nor_4  g06989(new_n9338, new_n9337, new_n9304);
nand_4 g06990(new_n9339, new_n9338, new_n9335);
not_3  g06991(new_n9340, new_n9338);
nand_4 g06992(new_n9341, new_n9340, new_n9334);
not_3  g06993(new_n9342, new_n9184);
xnor_3 g06994(new_n9343, new_n9234, new_n9342);
xnor_3 g06995(new_n9344_1, new_n9301, new_n9275);
nand_4 g06996(new_n9345, new_n9344_1, new_n9343);
not_3  g06997(new_n9346, new_n9344_1);
xnor_3 g06998(new_n9347, new_n9346, new_n9343);
xnor_3 g06999(new_n9348, new_n9298, new_n9280);
not_3  g07000(new_n9349, new_n9348);
not_3  g07001(new_n9350, new_n9193);
xnor_3 g07002(new_n9351, new_n9232, new_n9350);
nand_4 g07003(new_n9352, new_n9351, new_n9349);
xnor_3 g07004(new_n9353, new_n9351, new_n9348);
xnor_3 g07005(new_n9354, new_n9230, new_n9202);
not_3  g07006(new_n9355, new_n9354);
xnor_3 g07007(new_n9356, new_n9296, new_n9295);
not_3  g07008(new_n9357, new_n9356);
nand_4 g07009(new_n9358, new_n9357, new_n9355);
nand_4 g07010(new_n9359, new_n9356, new_n9354);
xnor_3 g07011(new_n9360, new_n9228, new_n9208);
xnor_3 g07012(new_n9361, new_n9225, new_n9222);
not_3  g07013(new_n9362, new_n9361);
and_4  g07014(new_n9363, new_n9291, new_n9290);
nor_4  g07015(new_n9364_1, new_n9291, new_n9290);
nor_4  g07016(new_n9365, new_n9364_1, new_n9363);
nand_4 g07017(new_n9366, new_n9365, new_n9362);
xor_3  g07018(new_n9367, n21993, n15508);
not_3  g07019(new_n9368, new_n9218);
xor_3  g07020(new_n9369, new_n9221, new_n9368);
not_3  g07021(new_n9370, new_n9369);
nand_4 g07022(new_n9371_1, new_n9370, new_n9367);
xnor_3 g07023(new_n9372_1, new_n9365, new_n9361);
nand_4 g07024(new_n9373, new_n9372_1, new_n9371_1);
nand_4 g07025(new_n9374, new_n9373, new_n9366);
nor_4  g07026(new_n9375, new_n9374, new_n9360);
not_3  g07027(new_n9376, new_n9287_1);
xnor_3 g07028(new_n9377, new_n9293, new_n9376);
xnor_3 g07029(new_n9378, new_n9374, new_n9360);
nor_4  g07030(new_n9379, new_n9378, new_n9377);
nor_4  g07031(new_n9380_1, new_n9379, new_n9375);
nand_4 g07032(new_n9381, new_n9380_1, new_n9359);
nand_4 g07033(new_n9382_1, new_n9381, new_n9358);
nand_4 g07034(new_n9383, new_n9382_1, new_n9353);
nand_4 g07035(new_n9384, new_n9383, new_n9352);
nand_4 g07036(new_n9385, new_n9384, new_n9347);
nand_4 g07037(new_n9386, new_n9385, new_n9345);
nand_4 g07038(new_n9387, new_n9386, new_n9341);
nand_4 g07039(new_n9388, new_n9387, new_n9339);
nor_4  g07040(new_n9389, new_n9388, new_n9333);
nor_4  g07041(new_n9390, new_n9389, new_n9332);
nor_4  g07042(new_n9391, new_n9390, new_n9327);
nor_4  g07043(new_n9392, new_n9391, new_n9326);
nand_4 g07044(new_n9393, new_n9392, new_n9321);
nand_4 g07045(new_n9394, new_n9393, new_n9319);
xnor_3 g07046(n829, new_n9394, new_n9315);
xor_3  g07047(new_n9396_1, n23272, n14826);
nor_4  g07048(new_n9397, n23493, n11481);
xor_3  g07049(new_n9398, n23493, n11481);
not_3  g07050(new_n9399_1, new_n9398);
nor_4  g07051(new_n9400, n16439, n10275);
xor_3  g07052(new_n9401, n16439, n10275);
not_3  g07053(new_n9402, new_n9401);
not_3  g07054(new_n9403_1, n15146);
nand_4 g07055(new_n9404, new_n4922, new_n9403_1);
xor_3  g07056(new_n9405, n15241, n15146);
nor_4  g07057(new_n9406, n11579, n7678);
not_3  g07058(new_n9407, new_n9406);
xor_3  g07059(new_n9408, n11579, n7678);
nor_4  g07060(new_n9409, n3785, n21);
not_3  g07061(new_n9410, new_n9409);
xor_3  g07062(new_n9411, n3785, n21);
nor_4  g07063(new_n9412, n20250, n1682);
not_3  g07064(new_n9413, new_n9412);
xor_3  g07065(new_n9414, n20250, n1682);
nor_4  g07066(new_n9415, n7963, n5822);
not_3  g07067(new_n9416, new_n9415);
xnor_3 g07068(new_n9417, n7963, n5822);
not_3  g07069(new_n9418, new_n9417);
nor_4  g07070(new_n9419_1, n26443, n10017);
not_3  g07071(new_n9420, new_n9419_1);
nand_4 g07072(new_n9421, n3618, n1681);
nand_4 g07073(new_n9422, n26443, n10017);
not_3  g07074(new_n9423_1, new_n9422);
nor_4  g07075(new_n9424, new_n9423_1, new_n9419_1);
nand_4 g07076(new_n9425, new_n9424, new_n9421);
nand_4 g07077(new_n9426, new_n9425, new_n9420);
nand_4 g07078(new_n9427, new_n9426, new_n9418);
nand_4 g07079(new_n9428, new_n9427, new_n9416);
nand_4 g07080(new_n9429, new_n9428, new_n9414);
nand_4 g07081(new_n9430_1, new_n9429, new_n9413);
nand_4 g07082(new_n9431, new_n9430_1, new_n9411);
nand_4 g07083(new_n9432, new_n9431, new_n9410);
nand_4 g07084(new_n9433, new_n9432, new_n9408);
nand_4 g07085(new_n9434, new_n9433, new_n9407);
nand_4 g07086(new_n9435_1, new_n9434, new_n9405);
nand_4 g07087(new_n9436, new_n9435_1, new_n9404);
not_3  g07088(new_n9437, new_n9436);
nor_4  g07089(new_n9438, new_n9437, new_n9402);
nor_4  g07090(new_n9439, new_n9438, new_n9400);
nor_4  g07091(new_n9440, new_n9439, new_n9399_1);
nor_4  g07092(new_n9441, new_n9440, new_n9397);
not_3  g07093(new_n9442, new_n9441);
nor_4  g07094(new_n9443, new_n9442, new_n9396_1);
not_3  g07095(new_n9444, new_n9396_1);
nor_4  g07096(new_n9445_1, new_n9441, new_n9444);
nor_4  g07097(new_n9446, new_n9445_1, new_n9443);
nor_4  g07098(new_n9447, new_n9446, n22764);
xnor_3 g07099(new_n9448, new_n9446, n22764);
not_3  g07100(new_n9449, new_n9439);
nor_4  g07101(new_n9450, new_n9449, new_n9398);
nor_4  g07102(new_n9451_1, new_n9450, new_n9440);
nor_4  g07103(new_n9452, new_n9451_1, n26264);
xnor_3 g07104(new_n9453, new_n9451_1, n26264);
xnor_3 g07105(new_n9454, new_n9436, new_n9401);
not_3  g07106(new_n9455, new_n9454);
nor_4  g07107(new_n9456, new_n9455, n7841);
not_3  g07108(new_n9457, n7841);
nor_4  g07109(new_n9458_1, new_n9454, new_n9457);
nor_4  g07110(new_n9459_1, new_n9458_1, new_n9456);
not_3  g07111(new_n9460_1, n16812);
xnor_3 g07112(new_n9461, new_n9434, new_n9405);
nand_4 g07113(new_n9462, new_n9461, new_n9460_1);
not_3  g07114(new_n9463, new_n9461);
nor_4  g07115(new_n9464, new_n9463, n16812);
nor_4  g07116(new_n9465, new_n9461, new_n9460_1);
nor_4  g07117(new_n9466, new_n9465, new_n9464);
not_3  g07118(new_n9467, n25068);
xnor_3 g07119(new_n9468, new_n9432, new_n9408);
nand_4 g07120(new_n9469, new_n9468, new_n9467);
not_3  g07121(new_n9470, new_n9468);
nor_4  g07122(new_n9471, new_n9470, n25068);
nor_4  g07123(new_n9472, new_n9468, new_n9467);
nor_4  g07124(new_n9473, new_n9472, new_n9471);
not_3  g07125(new_n9474, n2331);
xnor_3 g07126(new_n9475, new_n9430_1, new_n9411);
nand_4 g07127(new_n9476, new_n9475, new_n9474);
not_3  g07128(new_n9477, new_n9475);
nor_4  g07129(new_n9478, new_n9477, n2331);
nor_4  g07130(new_n9479, new_n9475, new_n9474);
nor_4  g07131(new_n9480, new_n9479, new_n9478);
xnor_3 g07132(new_n9481, new_n9428, new_n9414);
not_3  g07133(new_n9482, new_n9481);
nor_4  g07134(new_n9483, new_n9482, n22631);
not_3  g07135(new_n9484, new_n9483);
not_3  g07136(new_n9485, n22631);
nor_4  g07137(new_n9486, new_n9481, new_n9485);
nor_4  g07138(new_n9487, new_n9486, new_n9483);
not_3  g07139(new_n9488, n16743);
xnor_3 g07140(new_n9489, new_n9426, new_n9418);
nor_4  g07141(new_n9490, new_n9489, new_n9488);
xnor_3 g07142(new_n9491, new_n9489, new_n9488);
not_3  g07143(new_n9492, n15258);
nor_4  g07144(new_n9493_1, new_n2593, n4588);
nor_4  g07145(new_n9494, new_n9493_1, new_n9492);
nand_4 g07146(new_n9495, new_n9422, new_n9420);
xnor_3 g07147(new_n9496, new_n9495, new_n9421);
not_3  g07148(new_n9497, new_n9496);
nor_4  g07149(new_n9498, n15258, n4588);
not_3  g07150(new_n9499, new_n9498);
nor_4  g07151(new_n9500, new_n9499, new_n2593);
nor_4  g07152(new_n9501, new_n9500, new_n9494);
not_3  g07153(new_n9502, new_n9501);
nor_4  g07154(new_n9503, new_n9502, new_n9497);
nor_4  g07155(new_n9504, new_n9503, new_n9494);
nor_4  g07156(new_n9505, new_n9504, new_n9491);
nor_4  g07157(new_n9506, new_n9505, new_n9490);
nand_4 g07158(new_n9507_1, new_n9506, new_n9487);
nand_4 g07159(new_n9508_1, new_n9507_1, new_n9484);
nand_4 g07160(new_n9509, new_n9508_1, new_n9480);
nand_4 g07161(new_n9510, new_n9509, new_n9476);
nand_4 g07162(new_n9511, new_n9510, new_n9473);
nand_4 g07163(new_n9512_1, new_n9511, new_n9469);
nand_4 g07164(new_n9513, new_n9512_1, new_n9466);
nand_4 g07165(new_n9514, new_n9513, new_n9462);
nand_4 g07166(new_n9515, new_n9514, new_n9459_1);
not_3  g07167(new_n9516, new_n9515);
nor_4  g07168(new_n9517, new_n9516, new_n9456);
nor_4  g07169(new_n9518, new_n9517, new_n9453);
nor_4  g07170(new_n9519, new_n9518, new_n9452);
nor_4  g07171(new_n9520, new_n9519, new_n9448);
nor_4  g07172(new_n9521, new_n9520, new_n9447);
not_3  g07173(new_n9522, new_n9521);
nor_4  g07174(new_n9523, n23272, n14826);
nor_4  g07175(new_n9524, new_n9445_1, new_n9523);
nor_4  g07176(new_n9525, new_n9524, new_n9522);
not_3  g07177(new_n9526, new_n9525);
nor_4  g07178(new_n9527, n18105, new_n6505);
xor_3  g07179(new_n9528, n18105, new_n6505);
not_3  g07180(new_n9529, new_n9528);
nor_4  g07181(new_n9530, new_n6433, n24196);
xor_3  g07182(new_n9531, n26797, new_n5046_1);
nand_4 g07183(new_n9532, n23913, new_n5055);
xor_3  g07184(new_n9533, n23913, new_n5055);
nand_4 g07185(new_n9534, new_n5060_1, n22554);
xor_3  g07186(new_n9535, n25381, new_n6434);
nand_4 g07187(new_n9536, n20429, new_n5070);
xor_3  g07188(new_n9537, n20429, new_n5070);
nor_4  g07189(new_n9538, new_n6435, n268);
not_3  g07190(new_n9539, new_n9538);
xor_3  g07191(new_n9540, n3909, new_n5077_1);
not_3  g07192(new_n9541, n23974);
nor_4  g07193(new_n9542, n24879, new_n9541);
not_3  g07194(new_n9543, new_n9542);
xor_3  g07195(new_n9544, n24879, new_n9541);
nor_4  g07196(new_n9545, new_n4986, n2146);
nor_4  g07197(new_n9546, n6785, new_n6436);
not_3  g07198(new_n9547, n24032);
nor_4  g07199(new_n9548, new_n9547, n22173);
not_3  g07200(new_n9549, n583);
nand_4 g07201(new_n9550, n22843, new_n9549);
not_3  g07202(new_n9551, n22173);
nor_4  g07203(new_n9552_1, n24032, new_n9551);
nor_4  g07204(new_n9553, new_n9552_1, new_n9550);
nor_4  g07205(new_n9554_1, new_n9553, new_n9548);
nor_4  g07206(new_n9555, new_n9554_1, new_n9546);
nor_4  g07207(new_n9556_1, new_n9555, new_n9545);
nand_4 g07208(new_n9557_1, new_n9556_1, new_n9544);
nand_4 g07209(new_n9558_1, new_n9557_1, new_n9543);
nand_4 g07210(new_n9559, new_n9558_1, new_n9540);
nand_4 g07211(new_n9560, new_n9559, new_n9539);
nand_4 g07212(new_n9561, new_n9560, new_n9537);
nand_4 g07213(new_n9562, new_n9561, new_n9536);
nand_4 g07214(new_n9563, new_n9562, new_n9535);
nand_4 g07215(new_n9564, new_n9563, new_n9534);
nand_4 g07216(new_n9565, new_n9564, new_n9533);
nand_4 g07217(new_n9566, new_n9565, new_n9532);
nand_4 g07218(new_n9567, new_n9566, new_n9531);
not_3  g07219(new_n9568, new_n9567);
nor_4  g07220(new_n9569, new_n9568, new_n9530);
nor_4  g07221(new_n9570, new_n9569, new_n9529);
nor_4  g07222(new_n9571, new_n9570, new_n9527);
not_3  g07223(new_n9572, new_n9571);
not_3  g07224(new_n9573, n1536);
xor_3  g07225(new_n9574, new_n9569, new_n9529);
not_3  g07226(new_n9575, new_n9574);
nand_4 g07227(new_n9576, new_n9575, new_n9573);
xnor_3 g07228(new_n9577, new_n9574, new_n9573);
not_3  g07229(new_n9578, n19454);
xnor_3 g07230(new_n9579, new_n9566, new_n9531);
nand_4 g07231(new_n9580, new_n9579, new_n9578);
not_3  g07232(new_n9581, new_n9579);
xor_3  g07233(new_n9582, new_n9581, n19454);
not_3  g07234(new_n9583, n9445);
xnor_3 g07235(new_n9584, new_n9564, new_n9533);
nand_4 g07236(new_n9585, new_n9584, new_n9583);
not_3  g07237(new_n9586, new_n9584);
xor_3  g07238(new_n9587, new_n9586, n9445);
not_3  g07239(new_n9588, n1279);
xnor_3 g07240(new_n9589, new_n9562, new_n9535);
nand_4 g07241(new_n9590, new_n9589, new_n9588);
xnor_3 g07242(new_n9591, new_n9589, n1279);
not_3  g07243(new_n9592, n8324);
xnor_3 g07244(new_n9593, new_n9560, new_n9537);
nand_4 g07245(new_n9594, new_n9593, new_n9592);
xnor_3 g07246(new_n9595, new_n9593, n8324);
not_3  g07247(new_n9596, new_n9540);
xnor_3 g07248(new_n9597, new_n9558_1, new_n9596);
nor_4  g07249(new_n9598_1, new_n9597, n12546);
not_3  g07250(new_n9599, new_n9598_1);
not_3  g07251(new_n9600, n12546);
not_3  g07252(new_n9601, new_n9597);
nor_4  g07253(new_n9602, new_n9601, new_n9600);
nor_4  g07254(new_n9603, new_n9602, new_n9598_1);
xor_3  g07255(new_n9604, n24879, n23974);
xnor_3 g07256(new_n9605, new_n9556_1, new_n9604);
nor_4  g07257(new_n9606, new_n9605, n21078);
not_3  g07258(new_n9607, new_n9606);
not_3  g07259(new_n9608, n21078);
not_3  g07260(new_n9609, new_n9605);
nor_4  g07261(new_n9610, new_n9609, new_n9608);
nor_4  g07262(new_n9611, new_n9610, new_n9606);
not_3  g07263(new_n9612, n24485);
not_3  g07264(new_n9613, new_n9554_1);
nor_4  g07265(new_n9614, new_n9546, new_n9545);
xnor_3 g07266(new_n9615, new_n9614, new_n9613);
not_3  g07267(new_n9616_1, new_n9615);
nor_4  g07268(new_n9617, new_n9616_1, new_n9612);
not_3  g07269(new_n9618, new_n9617);
nor_4  g07270(new_n9619, new_n9615, n24485);
not_3  g07271(new_n9620, new_n9619);
nor_4  g07272(new_n9621, new_n9552_1, new_n9548);
xnor_3 g07273(new_n9622_1, new_n9621, new_n9550);
not_3  g07274(new_n9623, new_n9622_1);
nor_4  g07275(new_n9624, new_n9623, n2420);
nor_4  g07276(new_n9625, new_n2598, new_n2596);
not_3  g07277(new_n9626_1, n2420);
nor_4  g07278(new_n9627, new_n9622_1, new_n9626_1);
nor_4  g07279(new_n9628, new_n9627, new_n9624);
not_3  g07280(new_n9629, new_n9628);
nor_4  g07281(new_n9630, new_n9629, new_n9625);
nor_4  g07282(new_n9631, new_n9630, new_n9624);
nand_4 g07283(new_n9632, new_n9631, new_n9620);
nand_4 g07284(new_n9633_1, new_n9632, new_n9618);
not_3  g07285(new_n9634, new_n9633_1);
nand_4 g07286(new_n9635_1, new_n9634, new_n9611);
nand_4 g07287(new_n9636, new_n9635_1, new_n9607);
nand_4 g07288(new_n9637, new_n9636, new_n9603);
nand_4 g07289(new_n9638, new_n9637, new_n9599);
nand_4 g07290(new_n9639, new_n9638, new_n9595);
nand_4 g07291(new_n9640, new_n9639, new_n9594);
nand_4 g07292(new_n9641, new_n9640, new_n9591);
nand_4 g07293(new_n9642, new_n9641, new_n9590);
nand_4 g07294(new_n9643, new_n9642, new_n9587);
nand_4 g07295(new_n9644, new_n9643, new_n9585);
nand_4 g07296(new_n9645, new_n9644, new_n9582);
nand_4 g07297(new_n9646_1, new_n9645, new_n9580);
nand_4 g07298(new_n9647, new_n9646_1, new_n9577);
nand_4 g07299(new_n9648_1, new_n9647, new_n9576);
nor_4  g07300(new_n9649, new_n9648_1, new_n9572);
not_3  g07301(new_n9650, new_n9649);
not_3  g07302(new_n9651, new_n9524);
xnor_3 g07303(new_n9652, new_n9651, new_n9521);
xnor_3 g07304(new_n9653, new_n9648_1, new_n9571);
not_3  g07305(new_n9654, new_n9653);
nand_4 g07306(new_n9655_1, new_n9654, new_n9652);
xnor_3 g07307(new_n9656, new_n9653, new_n9652);
not_3  g07308(new_n9657, new_n9448);
not_3  g07309(new_n9658, new_n9519);
nor_4  g07310(new_n9659, new_n9658, new_n9657);
nor_4  g07311(new_n9660, new_n9659, new_n9520);
not_3  g07312(new_n9661, new_n9660);
xnor_3 g07313(new_n9662, new_n9646_1, new_n9577);
nor_4  g07314(new_n9663, new_n9662, new_n9661);
not_3  g07315(new_n9664, new_n9663);
xnor_3 g07316(new_n9665, new_n9662, new_n9660);
xnor_3 g07317(new_n9666, new_n9517, new_n9453);
not_3  g07318(new_n9667, new_n9666);
not_3  g07319(new_n9668, new_n9645);
nor_4  g07320(new_n9669, new_n9644, new_n9582);
nor_4  g07321(new_n9670, new_n9669, new_n9668);
nand_4 g07322(new_n9671, new_n9670, new_n9667);
xnor_3 g07323(new_n9672, new_n9670, new_n9666);
nor_4  g07324(new_n9673, new_n9514, new_n9459_1);
nor_4  g07325(new_n9674, new_n9673, new_n9516);
not_3  g07326(new_n9675, new_n9674);
xnor_3 g07327(new_n9676, new_n9642, new_n9587);
nor_4  g07328(new_n9677, new_n9676, new_n9675);
not_3  g07329(new_n9678, new_n9677);
not_3  g07330(new_n9679, new_n9676);
nor_4  g07331(new_n9680, new_n9679, new_n9674);
nor_4  g07332(new_n9681, new_n9680, new_n9677);
xnor_3 g07333(new_n9682, new_n9512_1, new_n9466);
xnor_3 g07334(new_n9683, new_n9640, new_n9591);
nor_4  g07335(new_n9684, new_n9683, new_n9682);
not_3  g07336(new_n9685, new_n9684);
not_3  g07337(new_n9686, new_n9682);
not_3  g07338(new_n9687, new_n9683);
nor_4  g07339(new_n9688, new_n9687, new_n9686);
nor_4  g07340(new_n9689_1, new_n9688, new_n9684);
xnor_3 g07341(new_n9690, new_n9510, new_n9473);
not_3  g07342(new_n9691, new_n9690);
not_3  g07343(new_n9692, new_n9595);
xnor_3 g07344(new_n9693, new_n9638, new_n9692);
nand_4 g07345(new_n9694, new_n9693, new_n9691);
xnor_3 g07346(new_n9695_1, new_n9693, new_n9690);
not_3  g07347(new_n9696, new_n9480);
xnor_3 g07348(new_n9697, new_n9508_1, new_n9696);
xnor_3 g07349(new_n9698, new_n9636, new_n9603);
not_3  g07350(new_n9699_1, new_n9698);
nand_4 g07351(new_n9700, new_n9699_1, new_n9697);
xnor_3 g07352(new_n9701, new_n9698, new_n9697);
xnor_3 g07353(new_n9702, new_n9506, new_n9487);
not_3  g07354(new_n9703, new_n9702);
xnor_3 g07355(new_n9704, new_n9633_1, new_n9611);
nand_4 g07356(new_n9705, new_n9704, new_n9703);
not_3  g07357(new_n9706, new_n9705);
nor_4  g07358(new_n9707, new_n9704, new_n9703);
nor_4  g07359(new_n9708, new_n9707, new_n9706);
xnor_3 g07360(new_n9709, new_n9504, new_n9491);
not_3  g07361(new_n9710, new_n9709);
not_3  g07362(new_n9711, new_n9631);
nor_4  g07363(new_n9712, new_n9619, new_n9617);
xnor_3 g07364(new_n9713, new_n9712, new_n9711);
nor_4  g07365(new_n9714, new_n9713, new_n9710);
not_3  g07366(new_n9715, new_n9714);
not_3  g07367(new_n9716, new_n9713);
nor_4  g07368(new_n9717, new_n9716, new_n9709);
nor_4  g07369(new_n9718, new_n9717, new_n9714);
not_3  g07370(new_n9719, new_n9625);
nor_4  g07371(new_n9720, new_n9628, new_n9719);
nor_4  g07372(new_n9721, new_n9720, new_n9630);
xor_3  g07373(new_n9722, new_n9502, new_n9496);
nor_4  g07374(new_n9723, new_n9722, new_n9721);
nand_4 g07375(new_n9724, new_n2599, new_n2595);
xnor_3 g07376(new_n9725, new_n9722, new_n9721);
nor_4  g07377(new_n9726_1, new_n9725, new_n9724);
nor_4  g07378(new_n9727, new_n9726_1, new_n9723);
nand_4 g07379(new_n9728, new_n9727, new_n9718);
nand_4 g07380(new_n9729, new_n9728, new_n9715);
nand_4 g07381(new_n9730, new_n9729, new_n9708);
nand_4 g07382(new_n9731, new_n9730, new_n9705);
nand_4 g07383(new_n9732, new_n9731, new_n9701);
nand_4 g07384(new_n9733, new_n9732, new_n9700);
nand_4 g07385(new_n9734, new_n9733, new_n9695_1);
nand_4 g07386(new_n9735, new_n9734, new_n9694);
nand_4 g07387(new_n9736, new_n9735, new_n9689_1);
nand_4 g07388(new_n9737, new_n9736, new_n9685);
nand_4 g07389(new_n9738, new_n9737, new_n9681);
nand_4 g07390(new_n9739, new_n9738, new_n9678);
nand_4 g07391(new_n9740, new_n9739, new_n9672);
nand_4 g07392(new_n9741, new_n9740, new_n9671);
nand_4 g07393(new_n9742, new_n9741, new_n9665);
nand_4 g07394(new_n9743, new_n9742, new_n9664);
nand_4 g07395(new_n9744, new_n9743, new_n9656);
nand_4 g07396(new_n9745, new_n9744, new_n9655_1);
xnor_3 g07397(new_n9746, new_n9745, new_n9650);
nand_4 g07398(new_n9747, new_n9746, new_n9526);
xnor_3 g07399(new_n9748, new_n9745, new_n9649);
nand_4 g07400(new_n9749, new_n9748, new_n9525);
nand_4 g07401(n849, new_n9749, new_n9747);
xor_3  g07402(n858, new_n2580, new_n9005);
not_3  g07403(new_n9752, n22442);
not_3  g07404(new_n9753_1, n3506);
not_3  g07405(new_n9754, n17251);
nor_4  g07406(new_n9755, n16994, n9246);
nand_4 g07407(new_n9756, new_n9755, new_n3850_1);
nor_4  g07408(new_n9757, new_n9756, n14790);
nand_4 g07409(new_n9758, new_n9757, new_n9754);
nor_4  g07410(new_n9759, new_n9758, n21674);
nand_4 g07411(new_n9760, new_n9759, new_n3834);
nor_4  g07412(new_n9761_1, new_n9760, n18444);
not_3  g07413(new_n9762, new_n9761_1);
nor_4  g07414(new_n9763_1, new_n9762, n14899);
xor_3  g07415(new_n9764, new_n9763_1, new_n9753_1);
nor_4  g07416(new_n9765, new_n9764, n1314);
not_3  g07417(new_n9766, n1314);
not_3  g07418(new_n9767_1, new_n9764);
nor_4  g07419(new_n9768, new_n9767_1, new_n9766);
nor_4  g07420(new_n9769, new_n9768, new_n9765);
not_3  g07421(new_n9770, n3306);
xor_3  g07422(new_n9771_1, new_n9762, n14899);
not_3  g07423(new_n9772, new_n9771_1);
nor_4  g07424(new_n9773, new_n9772, new_n9770);
not_3  g07425(new_n9774, new_n9773);
nor_4  g07426(new_n9775, new_n9771_1, n3306);
not_3  g07427(new_n9776, new_n9775);
xor_3  g07428(new_n9777, new_n9760, n18444);
nor_4  g07429(new_n9778_1, new_n9777, n22335);
xnor_3 g07430(new_n9779, new_n9777, n22335);
xor_3  g07431(new_n9780, new_n9759, new_n3834);
nor_4  g07432(new_n9781, new_n9780, n24048);
xnor_3 g07433(new_n9782, new_n9780, n24048);
nand_4 g07434(new_n9783_1, new_n9758, n21674);
not_3  g07435(new_n9784, new_n9783_1);
nor_4  g07436(new_n9785, new_n9784, new_n9759);
nor_4  g07437(new_n9786, new_n9785, n1525);
xnor_3 g07438(new_n9787, new_n9785, n1525);
xnor_3 g07439(new_n9788, new_n9757, n17251);
nor_4  g07440(new_n9789, new_n9788, n16988);
not_3  g07441(new_n9790, new_n9788);
nor_4  g07442(new_n9791, new_n9790, new_n5262);
nor_4  g07443(new_n9792, new_n9791, new_n9789);
nand_4 g07444(new_n9793, new_n9756, n14790);
not_3  g07445(new_n9794, new_n9793);
nor_4  g07446(new_n9795, new_n9794, new_n9757);
nor_4  g07447(new_n9796, new_n9795, n21779);
not_3  g07448(new_n9797, new_n9796);
xnor_3 g07449(new_n9798, new_n9755, n10096);
nor_4  g07450(new_n9799, new_n9798, n5376);
not_3  g07451(new_n9800, new_n9799);
not_3  g07452(new_n9801, new_n9798);
nor_4  g07453(new_n9802, new_n9801, new_n5271);
nor_4  g07454(new_n9803_1, new_n9802, new_n9799);
xnor_3 g07455(new_n9804, n16994, n9246);
nand_4 g07456(new_n9805, new_n9804, new_n5274_1);
nand_4 g07457(new_n9806, n23120, n9246);
not_3  g07458(new_n9807, new_n9805);
nor_4  g07459(new_n9808, new_n9804, new_n5274_1);
nor_4  g07460(new_n9809, new_n9808, new_n9807);
nand_4 g07461(new_n9810, new_n9809, new_n9806);
nand_4 g07462(new_n9811, new_n9810, new_n9805);
nand_4 g07463(new_n9812, new_n9811, new_n9803_1);
nand_4 g07464(new_n9813, new_n9812, new_n9800);
not_3  g07465(new_n9814, new_n9795);
nor_4  g07466(new_n9815, new_n9814, new_n5266);
nor_4  g07467(new_n9816, new_n9815, new_n9796);
nand_4 g07468(new_n9817, new_n9816, new_n9813);
nand_4 g07469(new_n9818, new_n9817, new_n9797);
nand_4 g07470(new_n9819, new_n9818, new_n9792);
not_3  g07471(new_n9820, new_n9819);
nor_4  g07472(new_n9821, new_n9820, new_n9789);
nor_4  g07473(new_n9822, new_n9821, new_n9787);
nor_4  g07474(new_n9823, new_n9822, new_n9786);
nor_4  g07475(new_n9824, new_n9823, new_n9782);
nor_4  g07476(new_n9825, new_n9824, new_n9781);
nor_4  g07477(new_n9826, new_n9825, new_n9779);
nor_4  g07478(new_n9827, new_n9826, new_n9778_1);
nand_4 g07479(new_n9828, new_n9827, new_n9776);
nand_4 g07480(new_n9829, new_n9828, new_n9774);
xnor_3 g07481(new_n9830, new_n9829, new_n9769);
not_3  g07482(new_n9831, new_n9830);
nand_4 g07483(new_n9832_1, new_n9831, new_n9752);
xnor_3 g07484(new_n9833_1, new_n9830, new_n9752);
not_3  g07485(new_n9834, n468);
nor_4  g07486(new_n9835, new_n9775, new_n9773);
xnor_3 g07487(new_n9836, new_n9835, new_n9827);
not_3  g07488(new_n9837, new_n9836);
nor_4  g07489(new_n9838_1, new_n9837, new_n9834);
xnor_3 g07490(new_n9839, new_n9836, n468);
not_3  g07491(new_n9840, n5400);
xnor_3 g07492(new_n9841, new_n9825, new_n9779);
nand_4 g07493(new_n9842, new_n9841, new_n9840);
not_3  g07494(new_n9843, n24048);
xnor_3 g07495(new_n9844, new_n9780, new_n9843);
xnor_3 g07496(new_n9845, new_n9823, new_n9844);
not_3  g07497(new_n9846, new_n9845);
nor_4  g07498(new_n9847, new_n9846, new_n8258);
xnor_3 g07499(new_n9848, new_n9845, n23923);
not_3  g07500(new_n9849, n329);
not_3  g07501(new_n9850, new_n9787);
not_3  g07502(new_n9851, new_n9821);
nor_4  g07503(new_n9852, new_n9851, new_n9850);
nor_4  g07504(new_n9853, new_n9852, new_n9822);
not_3  g07505(new_n9854, new_n9853);
nor_4  g07506(new_n9855, new_n9854, new_n9849);
nor_4  g07507(new_n9856, new_n9853, n329);
not_3  g07508(new_n9857, n24170);
not_3  g07509(new_n9858, n2409);
xnor_3 g07510(new_n9859, new_n9816, new_n9813);
nand_4 g07511(new_n9860, new_n9859, new_n9858);
not_3  g07512(new_n9861, new_n9860);
nor_4  g07513(new_n9862, new_n9859, new_n9858);
nor_4  g07514(new_n9863, new_n9862, new_n9861);
not_3  g07515(new_n9864, n8869);
xnor_3 g07516(new_n9865, new_n9811, new_n9803_1);
nand_4 g07517(new_n9866, new_n9865, new_n9864);
xnor_3 g07518(new_n9867_1, new_n9809, new_n9806);
nand_4 g07519(new_n9868, new_n9867_1, new_n8273);
not_3  g07520(new_n9869, n7428);
xnor_3 g07521(new_n9870, n23120, n9246);
not_3  g07522(new_n9871, new_n9870);
nor_4  g07523(new_n9872_1, new_n9871, new_n9869);
not_3  g07524(new_n9873, new_n9872_1);
not_3  g07525(new_n9874, new_n9868);
nor_4  g07526(new_n9875, new_n9867_1, new_n8273);
nor_4  g07527(new_n9876, new_n9875, new_n9874);
nand_4 g07528(new_n9877, new_n9876, new_n9873);
nand_4 g07529(new_n9878, new_n9877, new_n9868);
not_3  g07530(new_n9879, new_n9866);
nor_4  g07531(new_n9880, new_n9865, new_n9864);
nor_4  g07532(new_n9881, new_n9880, new_n9879);
nand_4 g07533(new_n9882, new_n9881, new_n9878);
nand_4 g07534(new_n9883, new_n9882, new_n9866);
nand_4 g07535(new_n9884, new_n9883, new_n9863);
nand_4 g07536(new_n9885, new_n9884, new_n9860);
nor_4  g07537(new_n9886, new_n9885, new_n9857);
nand_4 g07538(new_n9887, new_n9885, new_n9857);
nor_4  g07539(new_n9888, new_n9818, new_n9792);
nor_4  g07540(new_n9889, new_n9888, new_n9820);
nand_4 g07541(new_n9890_1, new_n9889, new_n9887);
not_3  g07542(new_n9891, new_n9890_1);
nor_4  g07543(new_n9892, new_n9891, new_n9886);
nor_4  g07544(new_n9893, new_n9892, new_n9856);
nor_4  g07545(new_n9894, new_n9893, new_n9855);
nor_4  g07546(new_n9895, new_n9894, new_n9848);
nor_4  g07547(new_n9896, new_n9895, new_n9847);
not_3  g07548(new_n9897, new_n9842);
nor_4  g07549(new_n9898, new_n9841, new_n9840);
nor_4  g07550(new_n9899, new_n9898, new_n9897);
nand_4 g07551(new_n9900, new_n9899, new_n9896);
nand_4 g07552(new_n9901, new_n9900, new_n9842);
nor_4  g07553(new_n9902, new_n9901, new_n9839);
nor_4  g07554(new_n9903, new_n9902, new_n9838_1);
nand_4 g07555(new_n9904, new_n9903, new_n9833_1);
nand_4 g07556(new_n9905, new_n9904, new_n9832_1);
not_3  g07557(new_n9906, new_n9763_1);
nor_4  g07558(new_n9907, new_n9906, n3506);
not_3  g07559(new_n9908, new_n9768);
not_3  g07560(new_n9909, new_n9765);
nand_4 g07561(new_n9910, new_n9829, new_n9909);
nand_4 g07562(new_n9911, new_n9910, new_n9908);
nor_4  g07563(new_n9912, new_n9911, new_n9907);
not_3  g07564(new_n9913, new_n9912);
xnor_3 g07565(new_n9914, new_n9913, new_n9905);
not_3  g07566(new_n9915, new_n3746);
nor_4  g07567(new_n9916, new_n3822, new_n9915);
nor_4  g07568(new_n9917_1, new_n9916, new_n3745);
not_3  g07569(new_n9918, new_n3671);
nor_4  g07570(new_n9919_1, new_n9918, n8856);
not_3  g07571(new_n9920, new_n3741);
nor_4  g07572(new_n9921, new_n9920, new_n3675);
nor_4  g07573(new_n9922, new_n9921, new_n9919_1);
not_3  g07574(new_n9923, new_n9922);
nor_4  g07575(new_n9924, new_n9923, new_n3674);
xnor_3 g07576(new_n9925, new_n9924, new_n9917_1);
nor_4  g07577(new_n9926_1, new_n9925, new_n9914);
nand_4 g07578(new_n9927, new_n9925, new_n9914);
not_3  g07579(new_n9928, new_n9927);
nor_4  g07580(new_n9929, new_n9928, new_n9926_1);
not_3  g07581(new_n9930, new_n9833_1);
xnor_3 g07582(new_n9931, new_n9903, new_n9930);
nor_4  g07583(new_n9932, new_n9931, new_n3824);
xnor_3 g07584(new_n9933, new_n9931, new_n3823);
not_3  g07585(new_n9934_1, new_n9839);
xnor_3 g07586(new_n9935, new_n9901, new_n9934_1);
nand_4 g07587(new_n9936, new_n9935, new_n3991);
xnor_3 g07588(new_n9937, new_n9935, new_n3986);
not_3  g07589(new_n9938_1, new_n9896);
xnor_3 g07590(new_n9939, new_n9899, new_n9938_1);
not_3  g07591(new_n9940, new_n9939);
nand_4 g07592(new_n9941, new_n9940, new_n3996);
xnor_3 g07593(new_n9942_1, new_n9939, new_n3996);
not_3  g07594(new_n9943, new_n9894);
xnor_3 g07595(new_n9944, new_n9943, new_n9848);
nand_4 g07596(new_n9945, new_n9944, new_n4005);
nor_4  g07597(new_n9946_1, new_n9856, new_n9855);
xnor_3 g07598(new_n9947, new_n9946_1, new_n9892);
nand_4 g07599(new_n9948, new_n9947, new_n4010_1);
xnor_3 g07600(new_n9949, new_n9947, new_n4009);
not_3  g07601(new_n9950, new_n9887);
nor_4  g07602(new_n9951, new_n9950, new_n9886);
xnor_3 g07603(new_n9952, new_n9951, new_n9889);
not_3  g07604(new_n9953, new_n9952);
nor_4  g07605(new_n9954, new_n9953, new_n4017);
nor_4  g07606(new_n9955, new_n9952, new_n4018);
xnor_3 g07607(new_n9956, new_n9883, new_n9863);
not_3  g07608(new_n9957, new_n9956);
nor_4  g07609(new_n9958, new_n9957, new_n4025);
not_3  g07610(new_n9959, new_n9958);
nor_4  g07611(new_n9960, new_n9956, new_n4029);
nor_4  g07612(new_n9961, new_n9960, new_n9958);
xnor_3 g07613(new_n9962, new_n9881, new_n9878);
nand_4 g07614(new_n9963, new_n9962, new_n4033);
not_3  g07615(new_n9964, new_n9877);
nor_4  g07616(new_n9965, new_n9876, new_n9873);
nor_4  g07617(new_n9966, new_n9965, new_n9964);
nor_4  g07618(new_n9967_1, new_n9966, new_n4041);
not_3  g07619(new_n9968_1, new_n9967_1);
xor_3  g07620(new_n9969, new_n9870, n7428);
not_3  g07621(new_n9970, new_n9969);
nand_4 g07622(new_n9971, new_n9970, new_n4046);
not_3  g07623(new_n9972, new_n9966);
nor_4  g07624(new_n9973, new_n9972, new_n4040);
nor_4  g07625(new_n9974, new_n9973, new_n9967_1);
nand_4 g07626(new_n9975, new_n9974, new_n9971);
nand_4 g07627(new_n9976, new_n9975, new_n9968_1);
not_3  g07628(new_n9977, new_n9963);
nor_4  g07629(new_n9978, new_n9962, new_n4033);
nor_4  g07630(new_n9979, new_n9978, new_n9977);
nand_4 g07631(new_n9980, new_n9979, new_n9976);
nand_4 g07632(new_n9981, new_n9980, new_n9963);
nand_4 g07633(new_n9982, new_n9981, new_n9961);
nand_4 g07634(new_n9983, new_n9982, new_n9959);
nor_4  g07635(new_n9984, new_n9983, new_n9955);
nor_4  g07636(new_n9985, new_n9984, new_n9954);
nand_4 g07637(new_n9986, new_n9985, new_n9949);
nand_4 g07638(new_n9987, new_n9986, new_n9948);
xnor_3 g07639(new_n9988, new_n9944, new_n4001);
nand_4 g07640(new_n9989, new_n9988, new_n9987);
nand_4 g07641(new_n9990, new_n9989, new_n9945);
nand_4 g07642(new_n9991, new_n9990, new_n9942_1);
nand_4 g07643(new_n9992, new_n9991, new_n9941);
nand_4 g07644(new_n9993, new_n9992, new_n9937);
nand_4 g07645(new_n9994, new_n9993, new_n9936);
nand_4 g07646(new_n9995, new_n9994, new_n9933);
not_3  g07647(new_n9996, new_n9995);
nor_4  g07648(new_n9997, new_n9996, new_n9932);
not_3  g07649(new_n9998, new_n9997);
xnor_3 g07650(n873, new_n9998, new_n9929);
not_3  g07651(new_n10000, new_n5967);
xor_3  g07652(new_n10001, n4812, new_n4190);
not_3  g07653(new_n10002, n24278);
nor_4  g07654(new_n10003, new_n10002, n19911);
xor_3  g07655(new_n10004, n24278, n19911);
nor_4  g07656(new_n10005, n24618, new_n4201);
nor_4  g07657(new_n10006, new_n3314, n13708);
nor_4  g07658(new_n10007, new_n4205_1, n3952);
nand_4 g07659(new_n10008, new_n4205_1, n3952);
nor_4  g07660(new_n10009_1, n12315, new_n2389);
nand_4 g07661(new_n10010_1, new_n10009_1, new_n10008);
not_3  g07662(new_n10011, new_n10010_1);
nor_4  g07663(new_n10012, new_n10011, new_n10007);
nor_4  g07664(new_n10013, new_n10012, new_n10006);
nor_4  g07665(new_n10014, new_n10013, new_n10005);
not_3  g07666(new_n10015, new_n10014);
nor_4  g07667(new_n10016, new_n10015, new_n10004);
nor_4  g07668(new_n10017_1, new_n10016, new_n10003);
xor_3  g07669(new_n10018_1, new_n10017_1, new_n10001);
xnor_3 g07670(new_n10019_1, new_n10018_1, new_n10000);
not_3  g07671(new_n10020, new_n5972);
xor_3  g07672(new_n10021_1, new_n10014, new_n10004);
nand_4 g07673(new_n10022, new_n10021_1, new_n10020);
not_3  g07674(new_n10023, new_n10012);
not_3  g07675(new_n10024, new_n10005);
not_3  g07676(new_n10025, new_n10006);
nand_4 g07677(new_n10026, new_n10025, new_n10024);
xor_3  g07678(new_n10027, new_n10026, new_n10023);
not_3  g07679(new_n10028, new_n10027);
nor_4  g07680(new_n10029, new_n10028, new_n5981);
xnor_3 g07681(new_n10030, new_n10027, new_n5977);
xor_3  g07682(new_n10031, n12315, new_n2389);
not_3  g07683(new_n10032, new_n10031);
nand_4 g07684(new_n10033, new_n10032, new_n5985);
nor_4  g07685(new_n10034, new_n10033, new_n5993);
xnor_3 g07686(new_n10035, new_n10033, new_n5993);
not_3  g07687(new_n10036, new_n10008);
nor_4  g07688(new_n10037, new_n10036, new_n10007);
xor_3  g07689(new_n10038, new_n10037, new_n10009_1);
nor_4  g07690(new_n10039, new_n10038, new_n10035);
nor_4  g07691(new_n10040, new_n10039, new_n10034);
nor_4  g07692(new_n10041, new_n10040, new_n10030);
nor_4  g07693(new_n10042, new_n10041, new_n10029);
not_3  g07694(new_n10043, new_n10022);
nor_4  g07695(new_n10044, new_n10021_1, new_n10020);
nor_4  g07696(new_n10045, new_n10044, new_n10043);
nand_4 g07697(new_n10046, new_n10045, new_n10042);
nand_4 g07698(new_n10047, new_n10046, new_n10022);
xor_3  g07699(n879, new_n10047, new_n10019_1);
xor_3  g07700(new_n10049, new_n9482, new_n8519_1);
not_3  g07701(new_n10050, new_n9489);
nand_4 g07702(new_n10051, new_n10050, new_n7792);
nor_4  g07703(new_n10052, new_n9496, new_n8524);
nor_4  g07704(new_n10053_1, new_n2593, new_n8626);
not_3  g07705(new_n10054, new_n10053_1);
xnor_3 g07706(new_n10055_1, new_n9496, new_n8524);
nor_4  g07707(new_n10056, new_n10055_1, new_n10054);
nor_4  g07708(new_n10057_1, new_n10056, new_n10052);
xnor_3 g07709(new_n10058, new_n9489, n12161);
not_3  g07710(new_n10059, new_n10058);
nand_4 g07711(new_n10060, new_n10059, new_n10057_1);
and_4  g07712(new_n10061, new_n10060, new_n10051);
xnor_3 g07713(new_n10062, new_n10061, new_n10049);
xnor_3 g07714(new_n10063, new_n10058, new_n10057_1);
nor_4  g07715(new_n10064, new_n7755, new_n4669);
nor_4  g07716(new_n10065, new_n7757, n14684);
nor_4  g07717(new_n10066, new_n10065, new_n10064);
nor_4  g07718(new_n10067, new_n7764, n6631);
not_3  g07719(new_n10068, new_n10067);
nand_4 g07720(new_n10069, new_n7767, n24732);
xnor_3 g07721(new_n10070, new_n7763, new_n4688);
not_3  g07722(new_n10071, new_n10070);
nand_4 g07723(new_n10072, new_n10071, new_n10069);
nand_4 g07724(new_n10073, new_n10072, new_n10068);
xnor_3 g07725(new_n10074, new_n10073, new_n10066);
nand_4 g07726(new_n10075, new_n10074, new_n10063);
not_3  g07727(new_n10076, new_n10075);
nor_4  g07728(new_n10077, new_n10074, new_n10063);
nor_4  g07729(new_n10078, new_n10077, new_n10076);
xnor_3 g07730(new_n10079, new_n10071, new_n10069);
xnor_3 g07731(new_n10080, new_n10055_1, new_n10053_1);
not_3  g07732(new_n10081, new_n10080);
nand_4 g07733(new_n10082, new_n10081, new_n10079);
xor_3  g07734(new_n10083, new_n7840, n24732);
xor_3  g07735(new_n10084, new_n2593, new_n8626);
nor_4  g07736(new_n10085, new_n10084, new_n10083);
not_3  g07737(new_n10086, new_n10082);
nor_4  g07738(new_n10087, new_n10081, new_n10079);
nor_4  g07739(new_n10088, new_n10087, new_n10086);
nand_4 g07740(new_n10089, new_n10088, new_n10085);
nand_4 g07741(new_n10090, new_n10089, new_n10082);
nand_4 g07742(new_n10091, new_n10090, new_n10078);
nand_4 g07743(new_n10092, new_n10091, new_n10075);
xnor_3 g07744(new_n10093, new_n10092, new_n10062);
nor_4  g07745(new_n10094, new_n7749, new_n4680);
not_3  g07746(new_n10095, new_n7749);
nor_4  g07747(new_n10096_1, new_n10095, n17035);
nor_4  g07748(new_n10097, new_n10096_1, new_n10094);
nand_4 g07749(new_n10098, new_n10073, new_n10066);
not_3  g07750(new_n10099, new_n10098);
nor_4  g07751(new_n10100, new_n10099, new_n10065);
nand_4 g07752(new_n10101_1, new_n10100, new_n10097);
not_3  g07753(new_n10102, new_n10101_1);
nor_4  g07754(new_n10103, new_n10100, new_n10097);
nor_4  g07755(new_n10104, new_n10103, new_n10102);
xor_3  g07756(n887, new_n10104, new_n10093);
xnor_3 g07757(new_n10106, new_n7081, new_n5606);
not_3  g07758(new_n10107, new_n10106);
nand_4 g07759(new_n10108, new_n7085, n22198);
xnor_3 g07760(new_n10109, new_n7085, new_n5610);
nand_4 g07761(new_n10110, new_n7089, n20826);
xnor_3 g07762(new_n10111_1, new_n7089, new_n5641);
nand_4 g07763(new_n10112, new_n7092, n7305);
not_3  g07764(new_n10113, new_n10112);
nor_4  g07765(new_n10114, new_n7092, n7305);
nor_4  g07766(new_n10115, new_n10114, new_n10113);
nand_4 g07767(new_n10116, new_n7097, n25872);
nor_4  g07768(new_n10117_1, new_n7102, n20259);
nor_4  g07769(new_n10118, new_n6769, new_n5717);
nor_4  g07770(new_n10119, new_n7101, new_n5628);
nor_4  g07771(new_n10120, new_n10119, new_n10117_1);
not_3  g07772(new_n10121, new_n10120);
nor_4  g07773(new_n10122, new_n10121, new_n10118);
nor_4  g07774(new_n10123, new_n10122, new_n10117_1);
not_3  g07775(new_n10124, new_n10116);
nor_4  g07776(new_n10125_1, new_n7097, n25872);
nor_4  g07777(new_n10126, new_n10125_1, new_n10124);
nand_4 g07778(new_n10127, new_n10126, new_n10123);
nand_4 g07779(new_n10128, new_n10127, new_n10116);
nand_4 g07780(new_n10129, new_n10128, new_n10115);
nand_4 g07781(new_n10130, new_n10129, new_n10112);
nand_4 g07782(new_n10131, new_n10130, new_n10111_1);
nand_4 g07783(new_n10132, new_n10131, new_n10110);
nand_4 g07784(new_n10133, new_n10132, new_n10109);
nand_4 g07785(new_n10134, new_n10133, new_n10108);
xnor_3 g07786(new_n10135, new_n10134, new_n10107);
not_3  g07787(new_n10136, new_n10135);
not_3  g07788(new_n10137, n25119);
xor_3  g07789(new_n10138, new_n3128, new_n10137);
not_3  g07790(new_n10139, n1163);
nor_4  g07791(new_n10140, new_n3133, new_n10139);
nor_4  g07792(new_n10141, new_n3137, n18537);
not_3  g07793(new_n10142, new_n10141);
not_3  g07794(new_n10143, n18537);
xor_3  g07795(new_n10144, new_n3138, new_n10143);
not_3  g07796(new_n10145, new_n3143);
nor_4  g07797(new_n10146, new_n10145, n7057);
not_3  g07798(new_n10147, new_n10146);
not_3  g07799(new_n10148, n7057);
nor_4  g07800(new_n10149, new_n3143, new_n10148);
nor_4  g07801(new_n10150, new_n10149, new_n10146);
nor_4  g07802(new_n10151, new_n3152, new_n5757);
xnor_3 g07803(new_n10152, new_n3152, new_n5757);
nand_4 g07804(new_n10153, new_n3165, n12495);
nand_4 g07805(new_n10154, new_n10153, new_n5778);
not_3  g07806(new_n10155, new_n10153);
xor_3  g07807(new_n10156, new_n10155, n20235);
nand_4 g07808(new_n10157, new_n10156, new_n3169);
nand_4 g07809(new_n10158_1, new_n10157, new_n10154);
nor_4  g07810(new_n10159, new_n10158_1, new_n10152);
nor_4  g07811(new_n10160, new_n10159, new_n10151);
nand_4 g07812(new_n10161, new_n10160, new_n10150);
nand_4 g07813(new_n10162, new_n10161, new_n10147);
nand_4 g07814(new_n10163, new_n10162, new_n10144);
nand_4 g07815(new_n10164, new_n10163, new_n10142);
xor_3  g07816(new_n10165_1, new_n3133, n1163);
nor_4  g07817(new_n10166, new_n10165_1, new_n10164);
nor_4  g07818(new_n10167, new_n10166, new_n10140);
nand_4 g07819(new_n10168, new_n10167, new_n10138);
not_3  g07820(new_n10169, new_n10168);
nor_4  g07821(new_n10170, new_n10167, new_n10138);
nor_4  g07822(new_n10171, new_n10170, new_n10169);
xnor_3 g07823(new_n10172, new_n10171, new_n10136);
xnor_3 g07824(new_n10173, new_n10132, new_n10109);
not_3  g07825(new_n10174, new_n10173);
xnor_3 g07826(new_n10175, new_n10165_1, new_n10164);
nand_4 g07827(new_n10176, new_n10175, new_n10174);
xnor_3 g07828(new_n10177, new_n10175, new_n10173);
not_3  g07829(new_n10178, new_n10163);
nor_4  g07830(new_n10179, new_n10162, new_n10144);
nor_4  g07831(new_n10180, new_n10179, new_n10178);
xnor_3 g07832(new_n10181, new_n10130, new_n10111_1);
not_3  g07833(new_n10182, new_n10181);
nand_4 g07834(new_n10183, new_n10182, new_n10180);
xnor_3 g07835(new_n10184, new_n10181, new_n10180);
not_3  g07836(new_n10185, new_n10161);
nor_4  g07837(new_n10186, new_n10160, new_n10150);
nor_4  g07838(new_n10187, new_n10186, new_n10185);
xnor_3 g07839(new_n10188, new_n10128, new_n10115);
not_3  g07840(new_n10189, new_n10188);
nand_4 g07841(new_n10190, new_n10189, new_n10187);
not_3  g07842(new_n10191, new_n10190);
nor_4  g07843(new_n10192, new_n10189, new_n10187);
nor_4  g07844(new_n10193, new_n10192, new_n10191);
not_3  g07845(new_n10194, new_n10152);
xnor_3 g07846(new_n10195, new_n10158_1, new_n10194);
xnor_3 g07847(new_n10196, new_n10126, new_n10123);
nor_4  g07848(new_n10197, new_n10196, new_n10195);
not_3  g07849(new_n10198, new_n10197);
not_3  g07850(new_n10199, new_n10195);
not_3  g07851(new_n10200, new_n10196);
nor_4  g07852(new_n10201_1, new_n10200, new_n10199);
nor_4  g07853(new_n10202, new_n10201_1, new_n10197);
xnor_3 g07854(new_n10203, new_n10121, new_n10118);
xnor_3 g07855(new_n10204, new_n10156, new_n3159);
nand_4 g07856(new_n10205, new_n10204, new_n10203);
nor_4  g07857(new_n10206, new_n6766, n3925);
nor_4  g07858(new_n10207, new_n10206, new_n10118);
not_3  g07859(new_n10208, new_n10207);
not_3  g07860(new_n10209, n12495);
xor_3  g07861(new_n10210, new_n3235_1, new_n10209);
nor_4  g07862(new_n10211, new_n10210, new_n10208);
not_3  g07863(new_n10212, new_n10205);
nor_4  g07864(new_n10213, new_n10204, new_n10203);
nor_4  g07865(new_n10214, new_n10213, new_n10212);
nand_4 g07866(new_n10215, new_n10214, new_n10211);
nand_4 g07867(new_n10216, new_n10215, new_n10205);
nand_4 g07868(new_n10217, new_n10216, new_n10202);
nand_4 g07869(new_n10218, new_n10217, new_n10198);
nand_4 g07870(new_n10219, new_n10218, new_n10193);
nand_4 g07871(new_n10220, new_n10219, new_n10190);
nand_4 g07872(new_n10221, new_n10220, new_n10184);
nand_4 g07873(new_n10222, new_n10221, new_n10183);
nand_4 g07874(new_n10223, new_n10222, new_n10177);
nand_4 g07875(new_n10224, new_n10223, new_n10176);
xnor_3 g07876(n904, new_n10224, new_n10172);
nor_4  g07877(new_n10226, n18962, n10158);
nand_4 g07878(new_n10227, new_n10226, new_n8815);
nor_4  g07879(new_n10228, new_n10227, n15539);
nand_4 g07880(new_n10229, new_n10228, new_n8807);
not_3  g07881(new_n10230, new_n10229);
nor_4  g07882(new_n10231, new_n10228, new_n8807);
nor_4  g07883(new_n10232, new_n10231, new_n10230);
xnor_3 g07884(new_n10233, new_n10232, n21471);
not_3  g07885(new_n10234, n18737);
nand_4 g07886(new_n10235, new_n10227, n15539);
not_3  g07887(new_n10236_1, new_n10235);
nor_4  g07888(new_n10237, new_n10236_1, new_n10228);
not_3  g07889(new_n10238, new_n10237);
nor_4  g07890(new_n10239_1, new_n10238, new_n10234);
not_3  g07891(new_n10240, new_n10239_1);
nor_4  g07892(new_n10241, new_n10237, n18737);
nor_4  g07893(new_n10242, new_n10241, new_n10239_1);
not_3  g07894(new_n10243, new_n10227);
nor_4  g07895(new_n10244_1, new_n10226, new_n8815);
nor_4  g07896(new_n10245, new_n10244_1, new_n10243);
nand_4 g07897(new_n10246, new_n10245, n14603);
xnor_3 g07898(new_n10247, new_n10245, n14603);
not_3  g07899(new_n10248, new_n10247);
nand_4 g07900(new_n10249, n18962, n10158);
not_3  g07901(new_n10250_1, new_n10249);
nor_4  g07902(new_n10251, new_n10250_1, new_n10226);
nor_4  g07903(new_n10252, new_n10251, n20794);
nand_4 g07904(new_n10253, n23333, n18962);
not_3  g07905(new_n10254, new_n10253);
xnor_3 g07906(new_n10255, n18962, n10158);
xnor_3 g07907(new_n10256, new_n10255, new_n3290);
nor_4  g07908(new_n10257, new_n10256, new_n10254);
nor_4  g07909(new_n10258, new_n10257, new_n10252);
nand_4 g07910(new_n10259, new_n10258, new_n10248);
nand_4 g07911(new_n10260, new_n10259, new_n10246);
nand_4 g07912(new_n10261_1, new_n10260, new_n10242);
nand_4 g07913(new_n10262_1, new_n10261_1, new_n10240);
xnor_3 g07914(new_n10263, new_n10262_1, new_n10233);
nor_4  g07915(new_n10264, new_n10263, n19472);
not_3  g07916(new_n10265, n19472);
not_3  g07917(new_n10266, new_n10263);
nor_4  g07918(new_n10267, new_n10266, new_n10265);
nor_4  g07919(new_n10268, new_n10267, new_n10264);
xnor_3 g07920(new_n10269, new_n10260, new_n10242);
not_3  g07921(new_n10270, new_n10269);
nor_4  g07922(new_n10271, new_n10270, n25370);
not_3  g07923(new_n10272, n24786);
xnor_3 g07924(new_n10273, new_n10258, new_n10248);
nor_4  g07925(new_n10274, new_n10273, new_n10272);
not_3  g07926(new_n10275_1, new_n10274);
xnor_3 g07927(new_n10276, new_n10273, new_n10272);
not_3  g07928(new_n10277, new_n10276);
nor_4  g07929(new_n10278, n23333, n18962);
nor_4  g07930(new_n10279, new_n10278, new_n10254);
nand_4 g07931(new_n10280, new_n10279, n23065);
nor_4  g07932(new_n10281, new_n10280, new_n10256);
not_3  g07933(new_n10282, new_n10281);
not_3  g07934(new_n10283, new_n10280);
xnor_3 g07935(new_n10284, new_n10256, new_n10254);
nor_4  g07936(new_n10285, new_n10284, new_n10283);
nor_4  g07937(new_n10286, new_n10285, new_n10281);
nand_4 g07938(new_n10287_1, new_n10286, n27120);
nand_4 g07939(new_n10288, new_n10287_1, new_n10282);
nand_4 g07940(new_n10289, new_n10288, new_n10277);
nand_4 g07941(new_n10290, new_n10289, new_n10275_1);
not_3  g07942(new_n10291, n25370);
xnor_3 g07943(new_n10292, new_n10269, new_n10291);
nor_4  g07944(new_n10293, new_n10292, new_n10290);
nor_4  g07945(new_n10294, new_n10293, new_n10271);
xnor_3 g07946(new_n10295_1, new_n10294, new_n10268);
xnor_3 g07947(new_n10296, new_n10295_1, new_n7870);
not_3  g07948(new_n10297, new_n10296);
xnor_3 g07949(new_n10298, new_n10292, new_n10290);
not_3  g07950(new_n10299, new_n10298);
nand_4 g07951(new_n10300, new_n10299, new_n7878);
not_3  g07952(new_n10301, new_n10300);
xnor_3 g07953(new_n10302, new_n10298, new_n7874);
not_3  g07954(new_n10303, new_n10287_1);
nor_4  g07955(new_n10304, new_n10286, n27120);
nor_4  g07956(new_n10305, new_n10304, new_n10303);
not_3  g07957(new_n10306, new_n10305);
nor_4  g07958(new_n10307, new_n10306, new_n7918);
nor_4  g07959(new_n10308, new_n10305, new_n7885);
xor_3  g07960(new_n10309, new_n10279, n23065);
nand_4 g07961(new_n10310, new_n10309, new_n7886);
nor_4  g07962(new_n10311, new_n10310, new_n10308);
nor_4  g07963(new_n10312, new_n10311, new_n10307);
nor_4  g07964(new_n10313, new_n10312, new_n7899);
not_3  g07965(new_n10314, new_n10313);
nand_4 g07966(new_n10315, new_n10312, new_n7899);
not_3  g07967(new_n10316, new_n10288);
xnor_3 g07968(new_n10317, new_n10316, new_n10276);
not_3  g07969(new_n10318, new_n10317);
nand_4 g07970(new_n10319, new_n10318, new_n10315);
nand_4 g07971(new_n10320, new_n10319, new_n10314);
nor_4  g07972(new_n10321_1, new_n10320, new_n10302);
nor_4  g07973(new_n10322, new_n10321_1, new_n10301);
xor_3  g07974(n948, new_n10322, new_n10297);
not_3  g07975(new_n10324, n10250);
xor_3  g07976(new_n10325, n25972, new_n10324);
not_3  g07977(new_n10326_1, new_n10325);
not_3  g07978(new_n10327_1, n21915);
nor_4  g07979(new_n10328, new_n10327_1, n7674);
not_3  g07980(new_n10329, n7674);
xor_3  g07981(new_n10330_1, n21915, new_n10329);
not_3  g07982(new_n10331, n6397);
nand_4 g07983(new_n10332, n13775, new_n10331);
xor_3  g07984(new_n10333, n13775, new_n10331);
nand_4 g07985(new_n10334, new_n7209, n1293);
not_3  g07986(new_n10335, n1293);
xor_3  g07987(new_n10336, n19196, new_n10335);
not_3  g07988(new_n10337, n19042);
nor_4  g07989(new_n10338, n23586, new_n10337);
not_3  g07990(new_n10339, new_n10338);
xor_3  g07991(new_n10340_1, n23586, new_n10337);
nor_4  g07992(new_n10341, n21226, new_n10265);
xor_3  g07993(new_n10342, n21226, new_n10265);
not_3  g07994(new_n10343, new_n10342);
nor_4  g07995(new_n10344, new_n10291, n4426);
xor_3  g07996(new_n10345_1, n25370, n4426);
not_3  g07997(new_n10346, n20036);
nor_4  g07998(new_n10347, n24786, new_n10346);
nor_4  g07999(new_n10348, new_n10272, n20036);
not_3  g08000(new_n10349, new_n10348);
nor_4  g08001(new_n10350, n27120, new_n4607);
not_3  g08002(new_n10351, new_n10350);
nand_4 g08003(new_n10352, n27120, new_n4607);
nor_4  g08004(new_n10353, n23065, new_n4609);
nand_4 g08005(new_n10354, new_n10353, new_n10352);
nand_4 g08006(new_n10355, new_n10354, new_n10351);
nand_4 g08007(new_n10356_1, new_n10355, new_n10349);
not_3  g08008(new_n10357, new_n10356_1);
nor_4  g08009(new_n10358, new_n10357, new_n10347);
not_3  g08010(new_n10359, new_n10358);
nor_4  g08011(new_n10360, new_n10359, new_n10345_1);
nor_4  g08012(new_n10361, new_n10360, new_n10344);
nor_4  g08013(new_n10362, new_n10361, new_n10343);
nor_4  g08014(new_n10363, new_n10362, new_n10341);
not_3  g08015(new_n10364, new_n10363);
nand_4 g08016(new_n10365, new_n10364, new_n10340_1);
nand_4 g08017(new_n10366, new_n10365, new_n10339);
nand_4 g08018(new_n10367, new_n10366, new_n10336);
nand_4 g08019(new_n10368, new_n10367, new_n10334);
nand_4 g08020(new_n10369, new_n10368, new_n10333);
nand_4 g08021(new_n10370, new_n10369, new_n10332);
nand_4 g08022(new_n10371, new_n10370, new_n10330_1);
not_3  g08023(new_n10372_1, new_n10371);
nor_4  g08024(new_n10373, new_n10372_1, new_n10328);
xor_3  g08025(new_n10374, new_n10373, new_n10326_1);
not_3  g08026(new_n10375, new_n10374);
xor_3  g08027(new_n10376, n20040, new_n8789);
not_3  g08028(new_n10377, new_n10376);
nor_4  g08029(new_n10378, new_n8793, n19531);
not_3  g08030(new_n10379, n19531);
xor_3  g08031(new_n10380, n23697, new_n10379);
not_3  g08032(new_n10381, n18345);
nand_4 g08033(new_n10382, new_n10381, n2289);
xor_3  g08034(new_n10383, n18345, new_n8796);
nand_4 g08035(new_n10384, new_n2620, n1112);
xor_3  g08036(new_n10385_1, n13190, new_n7937_1);
not_3  g08037(new_n10386, n3460);
nand_4 g08038(new_n10387_1, n20179, new_n10386);
xor_3  g08039(new_n10388_1, n20179, new_n10386);
nor_4  g08040(new_n10389, new_n8807, n5226);
not_3  g08041(new_n10390_1, new_n10389);
not_3  g08042(new_n10391, n5226);
xor_3  g08043(new_n10392, n19228, new_n10391);
nor_4  g08044(new_n10393, n17664, new_n8811);
not_3  g08045(new_n10394, new_n10393);
xor_3  g08046(new_n10395, n17664, new_n8811);
not_3  g08047(new_n10396, n23369);
nor_4  g08048(new_n10397, new_n10396, n8052);
nor_4  g08049(new_n10398, n23369, new_n8815);
not_3  g08050(new_n10399, n1136);
nor_4  g08051(new_n10400, n10158, new_n10399);
not_3  g08052(new_n10401, n10158);
nor_4  g08053(new_n10402, new_n10401, n1136);
nand_4 g08054(new_n10403, n19234, new_n8997);
nor_4  g08055(new_n10404_1, new_n10403, new_n10402);
nor_4  g08056(new_n10405_1, new_n10404_1, new_n10400);
nor_4  g08057(new_n10406, new_n10405_1, new_n10398);
nor_4  g08058(new_n10407, new_n10406, new_n10397);
nand_4 g08059(new_n10408, new_n10407, new_n10395);
nand_4 g08060(new_n10409_1, new_n10408, new_n10394);
nand_4 g08061(new_n10410, new_n10409_1, new_n10392);
nand_4 g08062(new_n10411_1, new_n10410, new_n10390_1);
nand_4 g08063(new_n10412, new_n10411_1, new_n10388_1);
nand_4 g08064(new_n10413, new_n10412, new_n10387_1);
nand_4 g08065(new_n10414, new_n10413, new_n10385_1);
nand_4 g08066(new_n10415, new_n10414, new_n10384);
nand_4 g08067(new_n10416, new_n10415, new_n10383);
nand_4 g08068(new_n10417, new_n10416, new_n10382);
nand_4 g08069(new_n10418, new_n10417, new_n10380);
not_3  g08070(new_n10419, new_n10418);
nor_4  g08071(new_n10420_1, new_n10419, new_n10378);
xor_3  g08072(new_n10421, new_n10420_1, new_n10377);
not_3  g08073(new_n10422, new_n10421);
not_3  g08074(new_n10423, n12507);
not_3  g08075(new_n10424, n22764);
nand_4 g08076(new_n10425, new_n9498, new_n9488);
nor_4  g08077(new_n10426, new_n10425, n22631);
nand_4 g08078(new_n10427, new_n10426, new_n9474);
nor_4  g08079(new_n10428, new_n10427, n25068);
nand_4 g08080(new_n10429, new_n10428, new_n9460_1);
nor_4  g08081(new_n10430, new_n10429, n7841);
not_3  g08082(new_n10431, new_n10430);
nor_4  g08083(new_n10432_1, new_n10431, n26264);
xor_3  g08084(new_n10433, new_n10432_1, new_n10424);
not_3  g08085(new_n10434, new_n10433);
nor_4  g08086(new_n10435, new_n10434, new_n10423);
nor_4  g08087(new_n10436, new_n10433, n12507);
nor_4  g08088(new_n10437, new_n10436, new_n10435);
not_3  g08089(new_n10438, n15077);
xor_3  g08090(new_n10439, new_n10431, n26264);
not_3  g08091(new_n10440, new_n10439);
nor_4  g08092(new_n10441, new_n10440, new_n10438);
not_3  g08093(new_n10442, new_n10441);
nor_4  g08094(new_n10443, new_n10439, n15077);
not_3  g08095(new_n10444, new_n10443);
not_3  g08096(new_n10445, n3710);
xor_3  g08097(new_n10446, new_n10429, n7841);
not_3  g08098(new_n10447, new_n10446);
nor_4  g08099(new_n10448, new_n10447, new_n10445);
not_3  g08100(new_n10449, new_n10448);
nor_4  g08101(new_n10450, new_n10446, n3710);
not_3  g08102(new_n10451, new_n10450);
xor_3  g08103(new_n10452, new_n10428, new_n9460_1);
nor_4  g08104(new_n10453, new_n10452, n26318);
not_3  g08105(new_n10454, n26318);
xnor_3 g08106(new_n10455, new_n10452, new_n10454);
not_3  g08107(new_n10456, new_n10455);
xor_3  g08108(new_n10457, new_n10427, n25068);
nor_4  g08109(new_n10458, new_n10457, n26054);
xnor_3 g08110(new_n10459, new_n10457, n26054);
xor_3  g08111(new_n10460, new_n10426, new_n9474);
nor_4  g08112(new_n10461, new_n10460, n19081);
not_3  g08113(new_n10462, n19081);
xnor_3 g08114(new_n10463, new_n10460, new_n10462);
nand_4 g08115(new_n10464, new_n10425, n22631);
not_3  g08116(new_n10465, new_n10464);
nor_4  g08117(new_n10466, new_n10465, new_n10426);
nor_4  g08118(new_n10467, new_n10466, n8309);
not_3  g08119(new_n10468, new_n10467);
not_3  g08120(new_n10469, new_n10425);
nor_4  g08121(new_n10470, new_n9498, new_n9488);
nor_4  g08122(new_n10471, new_n10470, new_n10469);
nor_4  g08123(new_n10472, new_n10471, n19144);
not_3  g08124(new_n10473, new_n10472);
not_3  g08125(new_n10474, n19144);
not_3  g08126(new_n10475, new_n10471);
nor_4  g08127(new_n10476, new_n10475, new_n10474);
nor_4  g08128(new_n10477, new_n10476, new_n10472);
xnor_3 g08129(new_n10478, n15258, n4588);
not_3  g08130(new_n10479, new_n10478);
nor_4  g08131(new_n10480, new_n10479, n12593);
not_3  g08132(new_n10481, new_n10480);
nand_4 g08133(new_n10482, n13714, n4588);
not_3  g08134(new_n10483, n12593);
nor_4  g08135(new_n10484_1, new_n10478, new_n10483);
nor_4  g08136(new_n10485, new_n10484_1, new_n10480);
nand_4 g08137(new_n10486, new_n10485, new_n10482);
nand_4 g08138(new_n10487, new_n10486, new_n10481);
nand_4 g08139(new_n10488, new_n10487, new_n10477);
nand_4 g08140(new_n10489_1, new_n10488, new_n10473);
not_3  g08141(new_n10490, n8309);
not_3  g08142(new_n10491, new_n10466);
nor_4  g08143(new_n10492, new_n10491, new_n10490);
nor_4  g08144(new_n10493, new_n10492, new_n10467);
nand_4 g08145(new_n10494, new_n10493, new_n10489_1);
nand_4 g08146(new_n10495, new_n10494, new_n10468);
nand_4 g08147(new_n10496, new_n10495, new_n10463);
not_3  g08148(new_n10497, new_n10496);
nor_4  g08149(new_n10498, new_n10497, new_n10461);
nor_4  g08150(new_n10499, new_n10498, new_n10459);
nor_4  g08151(new_n10500, new_n10499, new_n10458);
nor_4  g08152(new_n10501, new_n10500, new_n10456);
nor_4  g08153(new_n10502, new_n10501, new_n10453);
nand_4 g08154(new_n10503, new_n10502, new_n10451);
nand_4 g08155(new_n10504, new_n10503, new_n10449);
nand_4 g08156(new_n10505, new_n10504, new_n10444);
nand_4 g08157(new_n10506, new_n10505, new_n10442);
xnor_3 g08158(new_n10507, new_n10506, new_n10437);
xnor_3 g08159(new_n10508, new_n10507, new_n10422);
not_3  g08160(new_n10509, new_n10508);
xnor_3 g08161(new_n10510, new_n10417, new_n10380);
nor_4  g08162(new_n10511, new_n10443, new_n10441);
xnor_3 g08163(new_n10512, new_n10511, new_n10504);
nor_4  g08164(new_n10513, new_n10512, new_n10510);
not_3  g08165(new_n10514_1, new_n10513);
xnor_3 g08166(new_n10515, new_n10512, new_n10510);
not_3  g08167(new_n10516, new_n10515);
xnor_3 g08168(new_n10517, new_n10415, new_n10383);
nand_4 g08169(new_n10518, new_n10451, new_n10449);
not_3  g08170(new_n10519, new_n10518);
xnor_3 g08171(new_n10520, new_n10519, new_n10502);
nand_4 g08172(new_n10521, new_n10520, new_n10517);
not_3  g08173(new_n10522, new_n10517);
xnor_3 g08174(new_n10523, new_n10520, new_n10522);
xnor_3 g08175(new_n10524, new_n10413, new_n10385_1);
xnor_3 g08176(new_n10525_1, new_n10500, new_n10455);
nand_4 g08177(new_n10526, new_n10525_1, new_n10524);
not_3  g08178(new_n10527, new_n10524);
xnor_3 g08179(new_n10528, new_n10525_1, new_n10527);
xnor_3 g08180(new_n10529, new_n10411_1, new_n10388_1);
not_3  g08181(new_n10530, new_n10459);
xnor_3 g08182(new_n10531, new_n10498, new_n10530);
nand_4 g08183(new_n10532, new_n10531, new_n10529);
not_3  g08184(new_n10533, new_n10529);
xnor_3 g08185(new_n10534, new_n10531, new_n10533);
xnor_3 g08186(new_n10535, new_n10409_1, new_n10392);
nor_4  g08187(new_n10536, new_n10495, new_n10463);
nor_4  g08188(new_n10537, new_n10536, new_n10497);
nand_4 g08189(new_n10538, new_n10537, new_n10535);
not_3  g08190(new_n10539, new_n10535);
xnor_3 g08191(new_n10540_1, new_n10537, new_n10539);
xnor_3 g08192(new_n10541, new_n10407, new_n10395);
not_3  g08193(new_n10542, new_n10541);
xnor_3 g08194(new_n10543, new_n10493, new_n10489_1);
nor_4  g08195(new_n10544, new_n10543, new_n10542);
not_3  g08196(new_n10545, new_n10544);
not_3  g08197(new_n10546, new_n10543);
nor_4  g08198(new_n10547, new_n10546, new_n10541);
nor_4  g08199(new_n10548, new_n10547, new_n10544);
xnor_3 g08200(new_n10549, new_n10487, new_n10477);
not_3  g08201(new_n10550, new_n10549);
nor_4  g08202(new_n10551, new_n10398, new_n10397);
xnor_3 g08203(new_n10552, new_n10551, new_n10405_1);
nor_4  g08204(new_n10553, new_n10552, new_n10550);
xnor_3 g08205(new_n10554, new_n10552, new_n10550);
xnor_3 g08206(new_n10555, new_n10485, new_n10482);
not_3  g08207(new_n10556, new_n10555);
nor_4  g08208(new_n10557, new_n10402, new_n10400);
xnor_3 g08209(new_n10558, new_n10557, new_n10403);
nor_4  g08210(new_n10559, new_n10558, new_n10556);
xor_3  g08211(new_n10560, n19234, new_n8997);
xor_3  g08212(new_n10561_1, n13714, n4588);
not_3  g08213(new_n10562, new_n10561_1);
nor_4  g08214(new_n10563, new_n10562, new_n10560);
not_3  g08215(new_n10564_1, new_n10563);
not_3  g08216(new_n10565, new_n10558);
xnor_3 g08217(new_n10566, new_n10565, new_n10555);
nor_4  g08218(new_n10567, new_n10566, new_n10564_1);
nor_4  g08219(new_n10568, new_n10567, new_n10559);
nor_4  g08220(new_n10569, new_n10568, new_n10554);
nor_4  g08221(new_n10570, new_n10569, new_n10553);
nand_4 g08222(new_n10571, new_n10570, new_n10548);
nand_4 g08223(new_n10572, new_n10571, new_n10545);
nand_4 g08224(new_n10573, new_n10572, new_n10540_1);
nand_4 g08225(new_n10574, new_n10573, new_n10538);
nand_4 g08226(new_n10575, new_n10574, new_n10534);
nand_4 g08227(new_n10576, new_n10575, new_n10532);
nand_4 g08228(new_n10577_1, new_n10576, new_n10528);
nand_4 g08229(new_n10578, new_n10577_1, new_n10526);
nand_4 g08230(new_n10579, new_n10578, new_n10523);
nand_4 g08231(new_n10580, new_n10579, new_n10521);
not_3  g08232(new_n10581, new_n10580);
nand_4 g08233(new_n10582, new_n10581, new_n10516);
nand_4 g08234(new_n10583, new_n10582, new_n10514_1);
xnor_3 g08235(new_n10584, new_n10583, new_n10509);
xnor_3 g08236(new_n10585, new_n10584, new_n10375);
not_3  g08237(new_n10586, new_n10330_1);
xor_3  g08238(new_n10587, new_n10370, new_n10586);
xnor_3 g08239(new_n10588_1, new_n10580, new_n10515);
nand_4 g08240(new_n10589, new_n10588_1, new_n10587);
xnor_3 g08241(new_n10590, new_n10588_1, new_n10587);
not_3  g08242(new_n10591, new_n10590);
xor_3  g08243(new_n10592, new_n10368, new_n10333);
xnor_3 g08244(new_n10593_1, new_n10578, new_n10523);
nor_4  g08245(new_n10594, new_n10593_1, new_n10592);
not_3  g08246(new_n10595_1, new_n10594);
not_3  g08247(new_n10596, new_n10592);
not_3  g08248(new_n10597, new_n10593_1);
nor_4  g08249(new_n10598, new_n10597, new_n10596);
nor_4  g08250(new_n10599, new_n10598, new_n10594);
xnor_3 g08251(new_n10600, new_n10366, new_n10336);
xnor_3 g08252(new_n10601, new_n10576, new_n10528);
not_3  g08253(new_n10602, new_n10601);
nand_4 g08254(new_n10603, new_n10602, new_n10600);
xnor_3 g08255(new_n10604, new_n10601, new_n10600);
xor_3  g08256(new_n10605, new_n10364, new_n10340_1);
not_3  g08257(new_n10606, new_n10605);
not_3  g08258(new_n10607, new_n10534);
xnor_3 g08259(new_n10608, new_n10574, new_n10607);
nand_4 g08260(new_n10609, new_n10608, new_n10606);
xnor_3 g08261(new_n10610, new_n10608, new_n10605);
xor_3  g08262(new_n10611_1, new_n10361, new_n10343);
not_3  g08263(new_n10612, new_n10611_1);
not_3  g08264(new_n10613, new_n10572);
xnor_3 g08265(new_n10614_1, new_n10613, new_n10540_1);
nand_4 g08266(new_n10615, new_n10614_1, new_n10612);
xnor_3 g08267(new_n10616, new_n10614_1, new_n10611_1);
not_3  g08268(new_n10617_1, new_n10571);
nor_4  g08269(new_n10618, new_n10570, new_n10548);
nor_4  g08270(new_n10619, new_n10618, new_n10617_1);
xor_3  g08271(new_n10620, new_n10359, new_n10345_1);
not_3  g08272(new_n10621, new_n10620);
nand_4 g08273(new_n10622, new_n10621, new_n10619);
xnor_3 g08274(new_n10623, new_n10620, new_n10619);
not_3  g08275(new_n10624, new_n10554);
not_3  g08276(new_n10625, new_n10568);
nor_4  g08277(new_n10626, new_n10625, new_n10624);
nor_4  g08278(new_n10627, new_n10626, new_n10569);
not_3  g08279(new_n10628_1, new_n10627);
nor_4  g08280(new_n10629, new_n10348, new_n10347);
xor_3  g08281(new_n10630, new_n10629, new_n10355);
nand_4 g08282(new_n10631, new_n10630, new_n10628_1);
xnor_3 g08283(new_n10632, new_n10630, new_n10627);
xor_3  g08284(new_n10633, n23065, new_n4609);
xor_3  g08285(new_n10634, n19234, n18962);
xnor_3 g08286(new_n10635, new_n10561_1, new_n10634);
nor_4  g08287(new_n10636, new_n10635, new_n10633);
not_3  g08288(new_n10637, new_n10352);
nor_4  g08289(new_n10638, new_n10637, new_n10350);
xor_3  g08290(new_n10639, new_n10638, new_n10353);
not_3  g08291(new_n10640, new_n10639);
nor_4  g08292(new_n10641, new_n10640, new_n10636);
not_3  g08293(new_n10642, new_n10641);
xnor_3 g08294(new_n10643, new_n10566, new_n10564_1);
not_3  g08295(new_n10644, new_n10636);
nor_4  g08296(new_n10645, new_n10639, new_n10644);
nor_4  g08297(new_n10646, new_n10645, new_n10641);
nand_4 g08298(new_n10647_1, new_n10646, new_n10643);
nand_4 g08299(new_n10648, new_n10647_1, new_n10642);
nand_4 g08300(new_n10649, new_n10648, new_n10632);
nand_4 g08301(new_n10650_1, new_n10649, new_n10631);
nand_4 g08302(new_n10651, new_n10650_1, new_n10623);
nand_4 g08303(new_n10652, new_n10651, new_n10622);
nand_4 g08304(new_n10653_1, new_n10652, new_n10616);
nand_4 g08305(new_n10654, new_n10653_1, new_n10615);
nand_4 g08306(new_n10655, new_n10654, new_n10610);
nand_4 g08307(new_n10656, new_n10655, new_n10609);
nand_4 g08308(new_n10657, new_n10656, new_n10604);
nand_4 g08309(new_n10658, new_n10657, new_n10603);
nand_4 g08310(new_n10659, new_n10658, new_n10599);
nand_4 g08311(new_n10660, new_n10659, new_n10595_1);
nand_4 g08312(new_n10661, new_n10660, new_n10591);
nand_4 g08313(new_n10662, new_n10661, new_n10589);
nor_4  g08314(new_n10663, new_n10662, new_n10585);
not_3  g08315(new_n10664, new_n10585);
not_3  g08316(new_n10665, new_n10662);
nor_4  g08317(new_n10666, new_n10665, new_n10664);
nor_4  g08318(n957, new_n10666, new_n10663);
nor_4  g08319(new_n10668, new_n10634, n20385);
not_3  g08320(new_n10669, n20385);
nor_4  g08321(new_n10670, new_n10560, new_n10669);
nor_4  g08322(new_n10671, new_n10670, new_n10668);
not_3  g08323(new_n10672, new_n10671);
xnor_3 g08324(new_n10673, n26167, n24129);
xor_3  g08325(new_n10674, new_n10673, n21138);
xor_3  g08326(n980, new_n10674, new_n10672);
nor_4  g08327(new_n10676, new_n9129_1, new_n4909);
xnor_3 g08328(new_n10677, new_n9130, new_n4908);
nor_4  g08329(new_n10678, new_n9139, new_n4913_1);
not_3  g08330(new_n10679, new_n10678);
nor_4  g08331(new_n10680, new_n9144, new_n4912);
nor_4  g08332(new_n10681, new_n10680, new_n10678);
nor_4  g08333(new_n10682, new_n9149, new_n4918);
not_3  g08334(new_n10683, new_n10682);
nor_4  g08335(new_n10684, new_n9154, new_n4917);
nor_4  g08336(new_n10685, new_n10684, new_n10682);
nand_4 g08337(new_n10686, new_n9164_1, new_n4923);
xnor_3 g08338(new_n10687, new_n9159, new_n4923);
nor_4  g08339(new_n10688, new_n9177, new_n4927);
not_3  g08340(new_n10689, new_n10688);
nor_4  g08341(new_n10690, new_n9176, new_n4926);
nor_4  g08342(new_n10691, new_n10690, new_n10688);
nor_4  g08343(new_n10692_1, new_n9186, new_n4932);
not_3  g08344(new_n10693, new_n10692_1);
nor_4  g08345(new_n10694_1, new_n9185, new_n4936);
nor_4  g08346(new_n10695, new_n10694_1, new_n10692_1);
nor_4  g08347(new_n10696, new_n9195, new_n4940);
not_3  g08348(new_n10697, new_n10696);
nor_4  g08349(new_n10698, new_n9194, new_n4944);
nor_4  g08350(new_n10699, new_n10698, new_n10696);
nand_4 g08351(new_n10700, new_n9204, new_n4949);
xnor_3 g08352(new_n10701_1, new_n9204, new_n4951);
nor_4  g08353(new_n10702, new_n9213, new_n4954);
nand_4 g08354(new_n10703, new_n9368, new_n4958);
nor_4  g08355(new_n10704, new_n9212, new_n4955);
nor_4  g08356(new_n10705, new_n10704, new_n10702);
not_3  g08357(new_n10706, new_n10705);
nor_4  g08358(new_n10707, new_n10706, new_n10703);
nor_4  g08359(new_n10708, new_n10707, new_n10702);
nand_4 g08360(new_n10709, new_n10708, new_n10701_1);
nand_4 g08361(new_n10710_1, new_n10709, new_n10700);
nand_4 g08362(new_n10711, new_n10710_1, new_n10699);
nand_4 g08363(new_n10712_1, new_n10711, new_n10697);
nand_4 g08364(new_n10713, new_n10712_1, new_n10695);
nand_4 g08365(new_n10714, new_n10713, new_n10693);
nand_4 g08366(new_n10715, new_n10714, new_n10691);
nand_4 g08367(new_n10716, new_n10715, new_n10689);
nand_4 g08368(new_n10717, new_n10716, new_n10687);
nand_4 g08369(new_n10718, new_n10717, new_n10686);
nand_4 g08370(new_n10719, new_n10718, new_n10685);
nand_4 g08371(new_n10720, new_n10719, new_n10683);
nand_4 g08372(new_n10721, new_n10720, new_n10681);
nand_4 g08373(new_n10722, new_n10721, new_n10679);
nor_4  g08374(new_n10723, new_n10722, new_n10677);
nor_4  g08375(new_n10724, new_n10723, new_n10676);
xor_3  g08376(new_n10725, new_n9127, new_n4905);
not_3  g08377(new_n10726, new_n10725);
xnor_3 g08378(new_n10727, new_n10726, new_n10724);
not_3  g08379(new_n10728, n16544);
nor_4  g08380(new_n10729, new_n10728, n12650);
xor_3  g08381(new_n10730, n16544, new_n6510);
not_3  g08382(new_n10731, new_n10730);
not_3  g08383(new_n10732, n6814);
nor_4  g08384(new_n10733, n10201, new_n10732);
xor_3  g08385(new_n10734, n10201, new_n10732);
not_3  g08386(new_n10735, n10593);
nand_4 g08387(new_n10736, n19701, new_n10735);
xor_3  g08388(new_n10737, n19701, new_n10735);
not_3  g08389(new_n10738, n18290);
nand_4 g08390(new_n10739_1, n23529, new_n10738);
xor_3  g08391(new_n10740, n23529, new_n10738);
not_3  g08392(new_n10741, n24620);
nor_4  g08393(new_n10742, new_n10741, n11580);
not_3  g08394(new_n10743, new_n10742);
not_3  g08395(new_n10744, n11580);
xor_3  g08396(new_n10745, n24620, new_n10744);
not_3  g08397(new_n10746, n5211);
nor_4  g08398(new_n10747, n15884, new_n10746);
not_3  g08399(new_n10748, new_n10747);
xor_3  g08400(new_n10749, n15884, new_n10746);
not_3  g08401(new_n10750, n12956);
nor_4  g08402(new_n10751, new_n10750, n6356);
not_3  g08403(new_n10752, new_n10751);
xor_3  g08404(new_n10753, n12956, new_n6488);
nor_4  g08405(new_n10754, new_n6475, n18295);
not_3  g08406(new_n10755, new_n10754);
not_3  g08407(new_n10756_1, n18295);
nor_4  g08408(new_n10757, n27104, new_n10756_1);
not_3  g08409(new_n10758, new_n10757);
nor_4  g08410(new_n10759, new_n6479, n6502);
not_3  g08411(new_n10760, new_n10759);
nand_4 g08412(new_n10761, new_n6479, n6502);
not_3  g08413(new_n10762, n6611);
nor_4  g08414(new_n10763_1, n15780, new_n10762);
nand_4 g08415(new_n10764, new_n10763_1, new_n10761);
nand_4 g08416(new_n10765, new_n10764, new_n10760);
nand_4 g08417(new_n10766, new_n10765, new_n10758);
nand_4 g08418(new_n10767, new_n10766, new_n10755);
not_3  g08419(new_n10768, new_n10767);
nand_4 g08420(new_n10769, new_n10768, new_n10753);
nand_4 g08421(new_n10770, new_n10769, new_n10752);
nand_4 g08422(new_n10771, new_n10770, new_n10749);
nand_4 g08423(new_n10772, new_n10771, new_n10748);
nand_4 g08424(new_n10773, new_n10772, new_n10745);
nand_4 g08425(new_n10774, new_n10773, new_n10743);
nand_4 g08426(new_n10775_1, new_n10774, new_n10740);
nand_4 g08427(new_n10776, new_n10775_1, new_n10739_1);
nand_4 g08428(new_n10777, new_n10776, new_n10737);
nand_4 g08429(new_n10778, new_n10777, new_n10736);
nand_4 g08430(new_n10779, new_n10778, new_n10734);
not_3  g08431(new_n10780_1, new_n10779);
nor_4  g08432(new_n10781, new_n10780_1, new_n10733);
nor_4  g08433(new_n10782, new_n10781, new_n10731);
nor_4  g08434(new_n10783, new_n10782, new_n10729);
not_3  g08435(new_n10784, new_n10783);
xnor_3 g08436(new_n10785, new_n10784, new_n10727);
xor_3  g08437(new_n10786, new_n10781, new_n10731);
not_3  g08438(new_n10787, new_n10722);
xnor_3 g08439(new_n10788, new_n10787, new_n10677);
nor_4  g08440(new_n10789, new_n10788, new_n10786);
xnor_3 g08441(new_n10790, new_n10788, new_n10786);
xor_3  g08442(new_n10791, new_n10778, new_n10734);
xnor_3 g08443(new_n10792_1, new_n10720, new_n10681);
nor_4  g08444(new_n10793, new_n10792_1, new_n10791);
xnor_3 g08445(new_n10794, new_n10792_1, new_n10791);
xor_3  g08446(new_n10795, new_n10776, new_n10737);
not_3  g08447(new_n10796, new_n10719);
nor_4  g08448(new_n10797, new_n10718, new_n10685);
nor_4  g08449(new_n10798, new_n10797, new_n10796);
not_3  g08450(new_n10799, new_n10798);
nor_4  g08451(new_n10800, new_n10799, new_n10795);
xnor_3 g08452(new_n10801, new_n10798, new_n10795);
xnor_3 g08453(new_n10802, new_n10774, new_n10740);
xnor_3 g08454(new_n10803, new_n10716, new_n10687);
not_3  g08455(new_n10804, new_n10803);
nand_4 g08456(new_n10805, new_n10804, new_n10802);
xnor_3 g08457(new_n10806, new_n10803, new_n10802);
xor_3  g08458(new_n10807, new_n10772, new_n10745);
not_3  g08459(new_n10808, new_n10807);
not_3  g08460(new_n10809, new_n10691);
xnor_3 g08461(new_n10810, new_n10714, new_n10809);
nand_4 g08462(new_n10811, new_n10810, new_n10808);
xnor_3 g08463(new_n10812, new_n10810, new_n10807);
xor_3  g08464(new_n10813, new_n10770, new_n10749);
not_3  g08465(new_n10814, new_n10813);
not_3  g08466(new_n10815, new_n10695);
xnor_3 g08467(new_n10816, new_n10712_1, new_n10815);
nand_4 g08468(new_n10817_1, new_n10816, new_n10814);
xnor_3 g08469(new_n10818, new_n10816, new_n10813);
xnor_3 g08470(new_n10819, new_n10710_1, new_n10699);
not_3  g08471(new_n10820, new_n10819);
xor_3  g08472(new_n10821, new_n10767, new_n10753);
nand_4 g08473(new_n10822, new_n10821, new_n10820);
not_3  g08474(new_n10823, new_n10708);
xnor_3 g08475(new_n10824, new_n10823, new_n10701_1);
not_3  g08476(new_n10825, new_n10824);
nand_4 g08477(new_n10826, new_n10758, new_n10755);
xor_3  g08478(new_n10827, new_n10826, new_n10765);
nor_4  g08479(new_n10828, new_n10827, new_n10825);
not_3  g08480(new_n10829, new_n10828);
not_3  g08481(new_n10830, new_n10827);
nor_4  g08482(new_n10831, new_n10830, new_n10824);
nor_4  g08483(new_n10832, new_n10831, new_n10828);
xor_3  g08484(new_n10833, n15780, new_n10762);
xor_3  g08485(new_n10834_1, new_n9368, new_n4959);
nor_4  g08486(new_n10835, new_n10834_1, new_n10833);
not_3  g08487(new_n10836, new_n10761);
nor_4  g08488(new_n10837, new_n10836, new_n10759);
xor_3  g08489(new_n10838, new_n10837, new_n10763_1);
not_3  g08490(new_n10839, new_n10838);
nor_4  g08491(new_n10840, new_n10839, new_n10835);
not_3  g08492(new_n10841, new_n10840);
not_3  g08493(new_n10842, new_n10703);
xor_3  g08494(new_n10843, new_n10706, new_n10842);
not_3  g08495(new_n10844, new_n10835);
nor_4  g08496(new_n10845, new_n10838, new_n10844);
nor_4  g08497(new_n10846, new_n10845, new_n10840);
nand_4 g08498(new_n10847, new_n10846, new_n10843);
nand_4 g08499(new_n10848, new_n10847, new_n10841);
nand_4 g08500(new_n10849, new_n10848, new_n10832);
nand_4 g08501(new_n10850, new_n10849, new_n10829);
xnor_3 g08502(new_n10851_1, new_n10821, new_n10819);
nand_4 g08503(new_n10852, new_n10851_1, new_n10850);
nand_4 g08504(new_n10853, new_n10852, new_n10822);
nand_4 g08505(new_n10854, new_n10853, new_n10818);
nand_4 g08506(new_n10855, new_n10854, new_n10817_1);
nand_4 g08507(new_n10856, new_n10855, new_n10812);
nand_4 g08508(new_n10857, new_n10856, new_n10811);
nand_4 g08509(new_n10858, new_n10857, new_n10806);
nand_4 g08510(new_n10859, new_n10858, new_n10805);
nand_4 g08511(new_n10860, new_n10859, new_n10801);
not_3  g08512(new_n10861, new_n10860);
nor_4  g08513(new_n10862, new_n10861, new_n10800);
nor_4  g08514(new_n10863, new_n10862, new_n10794);
nor_4  g08515(new_n10864, new_n10863, new_n10793);
nor_4  g08516(new_n10865, new_n10864, new_n10790);
nor_4  g08517(new_n10866, new_n10865, new_n10789);
xnor_3 g08518(n982, new_n10866, new_n10785);
not_3  g08519(new_n10868, n4306);
not_3  g08520(new_n10869, n1667);
nor_4  g08521(new_n10870, n26808, n7339);
nand_4 g08522(new_n10871, new_n10870, new_n10869);
nor_4  g08523(new_n10872, new_n10871, n2680);
not_3  g08524(new_n10873, new_n10872);
nor_4  g08525(new_n10874_1, new_n10873, n2547);
not_3  g08526(new_n10875, new_n10874_1);
nor_4  g08527(new_n10876, new_n10875, n2999);
not_3  g08528(new_n10877, new_n10876);
nor_4  g08529(new_n10878, new_n10877, n14702);
not_3  g08530(new_n10879, new_n10878);
nor_4  g08531(new_n10880, new_n10879, n13914);
not_3  g08532(new_n10881, new_n10880);
nor_4  g08533(new_n10882, new_n10881, n3279);
xor_3  g08534(new_n10883, new_n10882, new_n10868);
xor_3  g08535(new_n10884, n23166, new_n4985);
not_3  g08536(new_n10885, new_n10884);
not_3  g08537(new_n10886, n10577);
nor_4  g08538(new_n10887, n24196, new_n10886);
xor_3  g08539(new_n10888, n24196, new_n10886);
nand_4 g08540(new_n10889, new_n5055, n6381);
not_3  g08541(new_n10890, n6381);
xor_3  g08542(new_n10891, n16376, new_n10890);
nand_4 g08543(new_n10892, new_n5060_1, n14345);
not_3  g08544(new_n10893, n14345);
xor_3  g08545(new_n10894, n25381, new_n10893);
nand_4 g08546(new_n10895, new_n5070, n11356);
not_3  g08547(new_n10896, n11356);
xor_3  g08548(new_n10897, n12587, new_n10896);
not_3  g08549(new_n10898, n3164);
nor_4  g08550(new_n10899, new_n10898, n268);
not_3  g08551(new_n10900, new_n10899);
xor_3  g08552(new_n10901, n3164, new_n5077_1);
not_3  g08553(new_n10902, n10611);
nor_4  g08554(new_n10903, n24879, new_n10902);
not_3  g08555(new_n10904, new_n10903);
xor_3  g08556(new_n10905, n24879, new_n10902);
nor_4  g08557(new_n10906, new_n4986, n2783);
not_3  g08558(new_n10907, n2783);
nor_4  g08559(new_n10908, n6785, new_n10907);
nor_4  g08560(new_n10909, new_n9547, n15490);
not_3  g08561(new_n10910, n15490);
nor_4  g08562(new_n10911, n24032, new_n10910);
not_3  g08563(new_n10912, n18);
nand_4 g08564(new_n10913, n22843, new_n10912);
nor_4  g08565(new_n10914, new_n10913, new_n10911);
nor_4  g08566(new_n10915, new_n10914, new_n10909);
nor_4  g08567(new_n10916, new_n10915, new_n10908);
nor_4  g08568(new_n10917, new_n10916, new_n10906);
nand_4 g08569(new_n10918, new_n10917, new_n10905);
nand_4 g08570(new_n10919, new_n10918, new_n10904);
nand_4 g08571(new_n10920, new_n10919, new_n10901);
nand_4 g08572(new_n10921, new_n10920, new_n10900);
nand_4 g08573(new_n10922, new_n10921, new_n10897);
nand_4 g08574(new_n10923, new_n10922, new_n10895);
nand_4 g08575(new_n10924_1, new_n10923, new_n10894);
nand_4 g08576(new_n10925, new_n10924_1, new_n10892);
nand_4 g08577(new_n10926, new_n10925, new_n10891);
nand_4 g08578(new_n10927, new_n10926, new_n10889);
nand_4 g08579(new_n10928, new_n10927, new_n10888);
not_3  g08580(new_n10929, new_n10928);
nor_4  g08581(new_n10930, new_n10929, new_n10887);
xor_3  g08582(new_n10931, new_n10930, new_n10885);
xnor_3 g08583(new_n10932, new_n10931, new_n10883);
not_3  g08584(new_n10933, n3279);
xor_3  g08585(new_n10934, new_n10880, new_n10933);
not_3  g08586(new_n10935, new_n10934);
xnor_3 g08587(new_n10936, new_n10927, new_n10888);
nor_4  g08588(new_n10937, new_n10936, new_n10935);
not_3  g08589(new_n10938, new_n10937);
not_3  g08590(new_n10939, new_n10936);
xor_3  g08591(new_n10940, new_n10939, new_n10935);
not_3  g08592(new_n10941, new_n10940);
not_3  g08593(new_n10942, n13914);
xor_3  g08594(new_n10943_1, new_n10878, new_n10942);
xnor_3 g08595(new_n10944, new_n10925, new_n10891);
not_3  g08596(new_n10945, new_n10944);
nor_4  g08597(new_n10946, new_n10945, new_n10943_1);
not_3  g08598(new_n10947, new_n10943_1);
xor_3  g08599(new_n10948, new_n10945, new_n10947);
not_3  g08600(new_n10949, n14702);
xor_3  g08601(new_n10950, new_n10876, new_n10949);
xnor_3 g08602(new_n10951, new_n10923, new_n10894);
not_3  g08603(new_n10952, new_n10951);
nor_4  g08604(new_n10953, new_n10952, new_n10950);
not_3  g08605(new_n10954, new_n10953);
not_3  g08606(new_n10955, new_n10950);
nor_4  g08607(new_n10956, new_n10951, new_n10955);
nor_4  g08608(new_n10957, new_n10956, new_n10953);
not_3  g08609(new_n10958, n2999);
xor_3  g08610(new_n10959, new_n10874_1, new_n10958);
xnor_3 g08611(new_n10960, new_n10921, new_n10897);
not_3  g08612(new_n10961_1, new_n10960);
nor_4  g08613(new_n10962, new_n10961_1, new_n10959);
not_3  g08614(new_n10963, new_n10962);
not_3  g08615(new_n10964, n2547);
xor_3  g08616(new_n10965, new_n10872, new_n10964);
not_3  g08617(new_n10966, new_n10901);
xor_3  g08618(new_n10967, n24879, n10611);
not_3  g08619(new_n10968, new_n10917);
nor_4  g08620(new_n10969, new_n10968, new_n10967);
nor_4  g08621(new_n10970, new_n10969, new_n10903);
nor_4  g08622(new_n10971, new_n10970, new_n10966);
nor_4  g08623(new_n10972, new_n10919, new_n10901);
nor_4  g08624(new_n10973, new_n10972, new_n10971);
nor_4  g08625(new_n10974, new_n10973, new_n10965);
not_3  g08626(new_n10975, new_n10974);
not_3  g08627(new_n10976, new_n10965);
not_3  g08628(new_n10977, new_n10973);
nor_4  g08629(new_n10978, new_n10977, new_n10976);
nor_4  g08630(new_n10979, new_n10978, new_n10974);
not_3  g08631(new_n10980, n2680);
xor_3  g08632(new_n10981, new_n10871, new_n10980);
nor_4  g08633(new_n10982, new_n10917, new_n10905);
nor_4  g08634(new_n10983, new_n10982, new_n10969);
not_3  g08635(new_n10984, new_n10983);
nand_4 g08636(new_n10985, new_n10984, new_n10981);
xor_3  g08637(new_n10986, new_n10870, n1667);
nor_4  g08638(new_n10987, new_n10908, new_n10906);
not_3  g08639(new_n10988, new_n10987);
xnor_3 g08640(new_n10989, new_n10988, new_n10915);
not_3  g08641(new_n10990, new_n10989);
nand_4 g08642(new_n10991, new_n10990, new_n10986);
xnor_3 g08643(new_n10992, new_n10989, new_n10986);
xor_3  g08644(new_n10993, n26808, n7339);
not_3  g08645(new_n10994, new_n10993);
nor_4  g08646(new_n10995, new_n10911, new_n10909);
xnor_3 g08647(new_n10996, new_n10995, new_n10913);
nor_4  g08648(new_n10997, new_n10996, new_n10994);
xor_3  g08649(new_n10998, n22843, n18);
nand_4 g08650(new_n10999, new_n10998, n26808);
not_3  g08651(new_n11000, new_n10996);
xnor_3 g08652(new_n11001, new_n11000, new_n10993);
nor_4  g08653(new_n11002, new_n11001, new_n10999);
nor_4  g08654(new_n11003, new_n11002, new_n10997);
nand_4 g08655(new_n11004, new_n11003, new_n10992);
nand_4 g08656(new_n11005_1, new_n11004, new_n10991);
xnor_3 g08657(new_n11006, new_n10983, new_n10981);
nand_4 g08658(new_n11007, new_n11006, new_n11005_1);
nand_4 g08659(new_n11008, new_n11007, new_n10985);
nand_4 g08660(new_n11009, new_n11008, new_n10979);
nand_4 g08661(new_n11010, new_n11009, new_n10975);
not_3  g08662(new_n11011_1, new_n10959);
nor_4  g08663(new_n11012, new_n10960, new_n11011_1);
nor_4  g08664(new_n11013, new_n11012, new_n10962);
nand_4 g08665(new_n11014, new_n11013, new_n11010);
nand_4 g08666(new_n11015, new_n11014, new_n10963);
nand_4 g08667(new_n11016, new_n11015, new_n10957);
nand_4 g08668(new_n11017, new_n11016, new_n10954);
not_3  g08669(new_n11018, new_n11017);
nor_4  g08670(new_n11019, new_n11018, new_n10948);
nor_4  g08671(new_n11020, new_n11019, new_n10946);
nand_4 g08672(new_n11021, new_n11020, new_n10941);
nand_4 g08673(new_n11022, new_n11021, new_n10938);
xnor_3 g08674(new_n11023_1, new_n11022, new_n10932);
xnor_3 g08675(new_n11024, new_n11023_1, new_n5141);
xnor_3 g08676(new_n11025_1, new_n11020, new_n10940);
nor_4  g08677(new_n11026, new_n11025_1, new_n5146);
xnor_3 g08678(new_n11027, new_n11025_1, new_n5146);
not_3  g08679(new_n11028, new_n5155);
not_3  g08680(new_n11029, new_n10948);
nor_4  g08681(new_n11030, new_n11017, new_n11029);
nor_4  g08682(new_n11031, new_n11030, new_n11019);
nand_4 g08683(new_n11032, new_n11031, new_n11028);
xnor_3 g08684(new_n11033, new_n11031, new_n5155);
xnor_3 g08685(new_n11034, new_n11015, new_n10957);
not_3  g08686(new_n11035, new_n11034);
nand_4 g08687(new_n11036, new_n11035, new_n5161);
xnor_3 g08688(new_n11037, new_n11034, new_n5161);
not_3  g08689(new_n11038, new_n11013);
xnor_3 g08690(new_n11039, new_n11038, new_n11010);
nand_4 g08691(new_n11040, new_n11039, new_n5170);
xnor_3 g08692(new_n11041, new_n11039, new_n5165);
xnor_3 g08693(new_n11042, new_n11008, new_n10979);
nor_4  g08694(new_n11043, new_n11042, new_n5173);
not_3  g08695(new_n11044_1, new_n11043);
not_3  g08696(new_n11045, new_n11042);
nor_4  g08697(new_n11046, new_n11045, new_n5174);
nor_4  g08698(new_n11047, new_n11046, new_n11043);
xnor_3 g08699(new_n11048, new_n11006, new_n11005_1);
not_3  g08700(new_n11049, new_n11048);
nand_4 g08701(new_n11050, new_n11049, new_n5182);
xnor_3 g08702(new_n11051, new_n11048, new_n5182);
not_3  g08703(new_n11052, new_n11003);
xnor_3 g08704(new_n11053, new_n11052, new_n10992);
nor_4  g08705(new_n11054, new_n11053, new_n5187);
xnor_3 g08706(new_n11055, new_n11053, new_n5187);
xnor_3 g08707(new_n11056_1, new_n11001, new_n10999);
nor_4  g08708(new_n11057, new_n11056_1, new_n5202);
not_3  g08709(new_n11058, new_n10999);
nor_4  g08710(new_n11059, new_n10998, n26808);
nor_4  g08711(new_n11060, new_n11059, new_n11058);
nand_4 g08712(new_n11061, new_n11060, new_n5198);
xnor_3 g08713(new_n11062, new_n11056_1, new_n5202);
nor_4  g08714(new_n11063_1, new_n11062, new_n11061);
nor_4  g08715(new_n11064, new_n11063_1, new_n11057);
nor_4  g08716(new_n11065, new_n11064, new_n11055);
nor_4  g08717(new_n11066, new_n11065, new_n11054);
nand_4 g08718(new_n11067, new_n11066, new_n11051);
nand_4 g08719(new_n11068, new_n11067, new_n11050);
nand_4 g08720(new_n11069, new_n11068, new_n11047);
nand_4 g08721(new_n11070, new_n11069, new_n11044_1);
nand_4 g08722(new_n11071, new_n11070, new_n11041);
nand_4 g08723(new_n11072, new_n11071, new_n11040);
nand_4 g08724(new_n11073, new_n11072, new_n11037);
nand_4 g08725(new_n11074, new_n11073, new_n11036);
nand_4 g08726(new_n11075, new_n11074, new_n11033);
nand_4 g08727(new_n11076, new_n11075, new_n11032);
not_3  g08728(new_n11077, new_n11076);
nor_4  g08729(new_n11078_1, new_n11077, new_n11027);
nor_4  g08730(new_n11079, new_n11078_1, new_n11026);
xnor_3 g08731(n984, new_n11079, new_n11024);
xnor_3 g08732(n1005, new_n11072, new_n11037);
not_3  g08733(new_n11082, new_n3573);
xor_3  g08734(n1016, new_n3637, new_n11082);
not_3  g08735(new_n11084, new_n4561);
xor_3  g08736(n1020, new_n4585, new_n11084);
xor_3  g08737(new_n11086, n18290, n12875);
nor_4  g08738(new_n11087, n11580, n2035);
not_3  g08739(new_n11088, new_n11087);
xor_3  g08740(new_n11089, n11580, n2035);
nor_4  g08741(new_n11090, n15884, n5213);
not_3  g08742(new_n11091, new_n11090);
xor_3  g08743(new_n11092, n15884, n5213);
nor_4  g08744(new_n11093, n6356, n4665);
not_3  g08745(new_n11094_1, new_n11093);
xor_3  g08746(new_n11095, n6356, n4665);
nor_4  g08747(new_n11096, n27104, n19005);
not_3  g08748(new_n11097, new_n11096);
xor_3  g08749(new_n11098, n27104, n19005);
nand_4 g08750(new_n11099, new_n6479, new_n3011);
nand_4 g08751(new_n11100, n6611, n5438);
xor_3  g08752(new_n11101_1, n27188, n4326);
nand_4 g08753(new_n11102, new_n11101_1, new_n11100);
nand_4 g08754(new_n11103_1, new_n11102, new_n11099);
nand_4 g08755(new_n11104, new_n11103_1, new_n11098);
nand_4 g08756(new_n11105, new_n11104, new_n11097);
nand_4 g08757(new_n11106, new_n11105, new_n11095);
nand_4 g08758(new_n11107, new_n11106, new_n11094_1);
nand_4 g08759(new_n11108, new_n11107, new_n11092);
nand_4 g08760(new_n11109, new_n11108, new_n11091);
nand_4 g08761(new_n11110, new_n11109, new_n11089);
nand_4 g08762(new_n11111, new_n11110, new_n11088);
xnor_3 g08763(new_n11112, new_n11111, new_n11086);
xnor_3 g08764(new_n11113, new_n11112, new_n3038);
not_3  g08765(new_n11114, new_n11089);
xnor_3 g08766(new_n11115, new_n11109, new_n11114);
nand_4 g08767(new_n11116, new_n11115, new_n10741);
xnor_3 g08768(new_n11117, new_n11109, new_n11089);
xnor_3 g08769(new_n11118, new_n11117, new_n10741);
not_3  g08770(new_n11119, new_n11095);
not_3  g08771(new_n11120_1, new_n11098);
not_3  g08772(new_n11121_1, new_n11099);
not_3  g08773(new_n11122, new_n11100);
xnor_3 g08774(new_n11123, n27188, n4326);
nor_4  g08775(new_n11124, new_n11123, new_n11122);
nor_4  g08776(new_n11125, new_n11124, new_n11121_1);
nor_4  g08777(new_n11126, new_n11125, new_n11120_1);
nor_4  g08778(new_n11127_1, new_n11126, new_n11096);
nor_4  g08779(new_n11128, new_n11127_1, new_n11119);
nor_4  g08780(new_n11129, new_n11128, new_n11093);
xnor_3 g08781(new_n11130, new_n11129, new_n11092);
not_3  g08782(new_n11131, new_n11130);
nor_4  g08783(new_n11132_1, new_n11131, n5211);
not_3  g08784(new_n11133, new_n11132_1);
nor_4  g08785(new_n11134_1, new_n11130, new_n10746);
nor_4  g08786(new_n11135, new_n11134_1, new_n11132_1);
xnor_3 g08787(new_n11136, new_n11127_1, new_n11095);
not_3  g08788(new_n11137, new_n11136);
nor_4  g08789(new_n11138_1, new_n11137, n12956);
not_3  g08790(new_n11139, new_n11138_1);
nor_4  g08791(new_n11140, new_n11136, new_n10750);
nor_4  g08792(new_n11141, new_n11140, new_n11138_1);
xnor_3 g08793(new_n11142, new_n11125, new_n11098);
not_3  g08794(new_n11143, new_n11142);
nor_4  g08795(new_n11144, new_n11143, n18295);
not_3  g08796(new_n11145, new_n11144);
not_3  g08797(new_n11146, n6502);
xnor_3 g08798(new_n11147, new_n11123, new_n11100);
nor_4  g08799(new_n11148, new_n11147, new_n11146);
not_3  g08800(new_n11149, n15780);
xnor_3 g08801(new_n11150, n6611, n5438);
nor_4  g08802(new_n11151, new_n11150, new_n11149);
not_3  g08803(new_n11152, new_n11151);
not_3  g08804(new_n11153, new_n11147);
xor_3  g08805(new_n11154, new_n11153, new_n11146);
nor_4  g08806(new_n11155, new_n11154, new_n11152);
nor_4  g08807(new_n11156, new_n11155, new_n11148);
xor_3  g08808(new_n11157, new_n11143, n18295);
nand_4 g08809(new_n11158, new_n11157, new_n11156);
nand_4 g08810(new_n11159, new_n11158, new_n11145);
nand_4 g08811(new_n11160, new_n11159, new_n11141);
nand_4 g08812(new_n11161, new_n11160, new_n11139);
nand_4 g08813(new_n11162, new_n11161, new_n11135);
nand_4 g08814(new_n11163, new_n11162, new_n11133);
nand_4 g08815(new_n11164, new_n11163, new_n11118);
nand_4 g08816(new_n11165, new_n11164, new_n11116);
xnor_3 g08817(new_n11166, new_n11165, new_n11113);
xor_3  g08818(new_n11167, n17250, n4409);
nor_4  g08819(new_n11168, n23160, n3570);
not_3  g08820(new_n11169, new_n11168);
xor_3  g08821(new_n11170, n23160, n3570);
nor_4  g08822(new_n11171, n16524, n13668);
not_3  g08823(new_n11172, new_n11171);
xor_3  g08824(new_n11173, n16524, n13668);
nor_4  g08825(new_n11174, n21276, n11056);
not_3  g08826(new_n11175, new_n11174);
xor_3  g08827(new_n11176, n21276, n11056);
nor_4  g08828(new_n11177, n26748, n15271);
nand_4 g08829(new_n11178, n26748, n15271);
not_3  g08830(new_n11179, new_n11178);
nor_4  g08831(new_n11180, new_n11179, new_n11177);
not_3  g08832(new_n11181, new_n11180);
nor_4  g08833(new_n11182_1, n25877, n10057);
nand_4 g08834(new_n11183, n24323, n8920);
not_3  g08835(new_n11184_1, new_n11183);
xnor_3 g08836(new_n11185, n25877, n10057);
nor_4  g08837(new_n11186, new_n11185, new_n11184_1);
nor_4  g08838(new_n11187, new_n11186, new_n11182_1);
nor_4  g08839(new_n11188, new_n11187, new_n11181);
nor_4  g08840(new_n11189, new_n11188, new_n11177);
not_3  g08841(new_n11190, new_n11189);
nand_4 g08842(new_n11191, new_n11190, new_n11176);
nand_4 g08843(new_n11192_1, new_n11191, new_n11175);
nand_4 g08844(new_n11193, new_n11192_1, new_n11173);
nand_4 g08845(new_n11194, new_n11193, new_n11172);
nand_4 g08846(new_n11195, new_n11194, new_n11170);
nand_4 g08847(new_n11196, new_n11195, new_n11169);
xnor_3 g08848(new_n11197, new_n11196, new_n11167);
not_3  g08849(new_n11198, new_n11197);
nor_4  g08850(new_n11199, new_n11198, new_n7030);
nor_4  g08851(new_n11200, new_n11197, n11044);
nor_4  g08852(new_n11201_1, new_n11200, new_n11199);
xnor_3 g08853(new_n11202, new_n11194, new_n11170);
not_3  g08854(new_n11203, new_n11202);
nor_4  g08855(new_n11204, new_n11203, new_n7033);
not_3  g08856(new_n11205, new_n11204);
nor_4  g08857(new_n11206, new_n11202, n2421);
nor_4  g08858(new_n11207, new_n11206, new_n11204);
xnor_3 g08859(new_n11208, new_n11192_1, new_n11173);
not_3  g08860(new_n11209, new_n11208);
nor_4  g08861(new_n11210, new_n11209, new_n7036);
not_3  g08862(new_n11211, new_n11210);
nor_4  g08863(new_n11212, new_n11208, n987);
nor_4  g08864(new_n11213, new_n11212, new_n11210);
xnor_3 g08865(new_n11214, new_n11189, new_n11176);
not_3  g08866(new_n11215, new_n11214);
nand_4 g08867(new_n11216, new_n11215, n20478);
xnor_3 g08868(new_n11217, new_n11214, n20478);
not_3  g08869(new_n11218, new_n11187);
nor_4  g08870(new_n11219, new_n11218, new_n11180);
nor_4  g08871(new_n11220_1, new_n11219, new_n11188);
nor_4  g08872(new_n11221, new_n11220_1, new_n9102);
not_3  g08873(new_n11222, new_n11221);
not_3  g08874(new_n11223_1, new_n11185);
nor_4  g08875(new_n11224, new_n11223_1, new_n11183);
nor_4  g08876(new_n11225, new_n11224, new_n11186);
not_3  g08877(new_n11226, new_n11225);
nor_4  g08878(new_n11227, new_n11226, n22619);
xnor_3 g08879(new_n11228, n24323, n8920);
nor_4  g08880(new_n11229, new_n11228, new_n9107);
xnor_3 g08881(new_n11230, new_n11225, new_n9105);
nor_4  g08882(new_n11231, new_n11230, new_n11229);
nor_4  g08883(new_n11232, new_n11231, new_n11227);
xnor_3 g08884(new_n11233, new_n11220_1, n26882);
nand_4 g08885(new_n11234_1, new_n11233, new_n11232);
nand_4 g08886(new_n11235, new_n11234_1, new_n11222);
nand_4 g08887(new_n11236, new_n11235, new_n11217);
nand_4 g08888(new_n11237, new_n11236, new_n11216);
nand_4 g08889(new_n11238, new_n11237, new_n11213);
nand_4 g08890(new_n11239, new_n11238, new_n11211);
nand_4 g08891(new_n11240, new_n11239, new_n11207);
nand_4 g08892(new_n11241, new_n11240, new_n11205);
xnor_3 g08893(new_n11242, new_n11241, new_n11201_1);
not_3  g08894(new_n11243, new_n11242);
xnor_3 g08895(new_n11244, new_n11243, new_n11166);
xnor_3 g08896(new_n11245_1, new_n11163, new_n11118);
not_3  g08897(new_n11246, new_n11245_1);
xnor_3 g08898(new_n11247, new_n11239, new_n11207);
not_3  g08899(new_n11248, new_n11247);
nand_4 g08900(new_n11249, new_n11248, new_n11246);
xnor_3 g08901(new_n11250, new_n11248, new_n11245_1);
not_3  g08902(new_n11251, new_n11135);
xnor_3 g08903(new_n11252, new_n11161, new_n11251);
xnor_3 g08904(new_n11253, new_n11237, new_n11213);
not_3  g08905(new_n11254, new_n11253);
nand_4 g08906(new_n11255, new_n11254, new_n11252);
xnor_3 g08907(new_n11256, new_n11253, new_n11252);
not_3  g08908(new_n11257, new_n11141);
xnor_3 g08909(new_n11258, new_n11159, new_n11257);
not_3  g08910(new_n11259, new_n11236);
nor_4  g08911(new_n11260, new_n11235, new_n11217);
nor_4  g08912(new_n11261_1, new_n11260, new_n11259);
nand_4 g08913(new_n11262, new_n11261_1, new_n11258);
not_3  g08914(new_n11263, new_n11262);
nor_4  g08915(new_n11264, new_n11261_1, new_n11258);
nor_4  g08916(new_n11265, new_n11264, new_n11263);
xor_3  g08917(new_n11266_1, new_n11143, new_n10756_1);
xnor_3 g08918(new_n11267, new_n11266_1, new_n11156);
xnor_3 g08919(new_n11268, new_n11233, new_n11232);
not_3  g08920(new_n11269, new_n11268);
nand_4 g08921(new_n11270, new_n11269, new_n11267);
not_3  g08922(new_n11271, new_n11270);
nor_4  g08923(new_n11272, new_n11269, new_n11267);
nor_4  g08924(new_n11273_1, new_n11272, new_n11271);
xnor_3 g08925(new_n11274, new_n11230, new_n11229);
xnor_3 g08926(new_n11275_1, new_n11154, new_n11152);
nand_4 g08927(new_n11276, new_n11275_1, new_n11274);
xor_3  g08928(new_n11277, new_n11228, new_n9107);
not_3  g08929(new_n11278, new_n11277);
xor_3  g08930(new_n11279, new_n11150, new_n11149);
nor_4  g08931(new_n11280, new_n11279, new_n11278);
not_3  g08932(new_n11281, new_n11276);
nor_4  g08933(new_n11282, new_n11275_1, new_n11274);
nor_4  g08934(new_n11283, new_n11282, new_n11281);
nand_4 g08935(new_n11284, new_n11283, new_n11280);
nand_4 g08936(new_n11285, new_n11284, new_n11276);
nand_4 g08937(new_n11286, new_n11285, new_n11273_1);
nand_4 g08938(new_n11287, new_n11286, new_n11270);
nand_4 g08939(new_n11288, new_n11287, new_n11265);
nand_4 g08940(new_n11289, new_n11288, new_n11262);
nand_4 g08941(new_n11290_1, new_n11289, new_n11256);
nand_4 g08942(new_n11291, new_n11290_1, new_n11255);
nand_4 g08943(new_n11292, new_n11291, new_n11250);
nand_4 g08944(new_n11293, new_n11292, new_n11249);
xnor_3 g08945(n1044, new_n11293, new_n11244);
nor_4  g08946(new_n11295, n22619, n6775);
nand_4 g08947(new_n11296, new_n11295, new_n9102);
nor_4  g08948(new_n11297, new_n11296, n20478);
nand_4 g08949(new_n11298, new_n11296, n20478);
not_3  g08950(new_n11299, new_n11298);
nor_4  g08951(new_n11300, new_n11299, new_n11297);
xnor_3 g08952(new_n11301, new_n11300, new_n5618);
not_3  g08953(new_n11302_1, new_n11296);
nor_4  g08954(new_n11303, new_n11295, new_n9102);
nor_4  g08955(new_n11304, new_n11303, new_n11302_1);
nand_4 g08956(new_n11305, new_n11304, n25872);
xnor_3 g08957(new_n11306, new_n11304, new_n5625);
nand_4 g08958(new_n11307, n22619, n6775);
not_3  g08959(new_n11308, new_n11307);
nor_4  g08960(new_n11309, new_n11308, new_n11295);
nand_4 g08961(new_n11310, new_n11309, n20259);
nand_4 g08962(new_n11311, n6775, n3925);
not_3  g08963(new_n11312, new_n11311);
xnor_3 g08964(new_n11313_1, new_n11309, new_n5628);
nand_4 g08965(new_n11314, new_n11313_1, new_n11312);
nand_4 g08966(new_n11315, new_n11314, new_n11310);
nand_4 g08967(new_n11316, new_n11315, new_n11306);
nand_4 g08968(new_n11317, new_n11316, new_n11305);
xnor_3 g08969(new_n11318, new_n11317, new_n11301);
nand_4 g08970(new_n11319, new_n6746, new_n4879);
nor_4  g08971(new_n11320, new_n11319, n25074);
nand_4 g08972(new_n11321, new_n11319, n25074);
not_3  g08973(new_n11322, new_n11321);
nor_4  g08974(new_n11323, new_n11322, new_n11320);
not_3  g08975(new_n11324, new_n11323);
nor_4  g08976(new_n11325_1, new_n11324, new_n2426);
nor_4  g08977(new_n11326_1, new_n11323, n3480);
nor_4  g08978(new_n11327, new_n11326_1, new_n11325_1);
not_3  g08979(new_n11328, new_n11327);
not_3  g08980(new_n11329, new_n11319);
nor_4  g08981(new_n11330_1, new_n6746, new_n4879);
nor_4  g08982(new_n11331, new_n11330_1, new_n11329);
not_3  g08983(new_n11332, new_n11331);
nor_4  g08984(new_n11333, new_n11332, new_n9050);
not_3  g08985(new_n11334, new_n11333);
nor_4  g08986(new_n11335, new_n11331, n16722);
nor_4  g08987(new_n11336, new_n11335, new_n11333);
not_3  g08988(new_n11337, new_n6751);
nand_4 g08989(new_n11338, new_n6756, new_n11337);
not_3  g08990(new_n11339, new_n11338);
nand_4 g08991(new_n11340, new_n11339, new_n11336);
nand_4 g08992(new_n11341, new_n11340, new_n11334);
nor_4  g08993(new_n11342, new_n11341, new_n11328);
not_3  g08994(new_n11343, new_n11341);
nor_4  g08995(new_n11344, new_n11343, new_n11327);
nor_4  g08996(new_n11345, new_n11344, new_n11342);
nor_4  g08997(new_n11346, new_n11345, new_n11318);
not_3  g08998(new_n11347_1, new_n11301);
xnor_3 g08999(new_n11348_1, new_n11317, new_n11347_1);
not_3  g09000(new_n11349, new_n11345);
nor_4  g09001(new_n11350, new_n11349, new_n11348_1);
nor_4  g09002(new_n11351, new_n11350, new_n11346);
xnor_3 g09003(new_n11352_1, new_n11339, new_n11336);
xnor_3 g09004(new_n11353, new_n11315, new_n11306);
nor_4  g09005(new_n11354, new_n11353, new_n11352_1);
not_3  g09006(new_n11355, new_n11354);
not_3  g09007(new_n11356_1, new_n11352_1);
not_3  g09008(new_n11357, new_n11353);
nor_4  g09009(new_n11358, new_n11357, new_n11356_1);
nor_4  g09010(new_n11359, new_n11358, new_n11354);
xnor_3 g09011(new_n11360, new_n11313_1, new_n11312);
nor_4  g09012(new_n11361, new_n11360, new_n6758);
not_3  g09013(new_n11362, new_n11361);
xor_3  g09014(new_n11363, n6775, n3925);
not_3  g09015(new_n11364, new_n11363);
nor_4  g09016(new_n11365, new_n11364, new_n6730);
not_3  g09017(new_n11366, new_n11360);
nor_4  g09018(new_n11367, new_n11366, new_n6759);
nor_4  g09019(new_n11368, new_n11367, new_n11361);
nand_4 g09020(new_n11369, new_n11368, new_n11365);
nand_4 g09021(new_n11370, new_n11369, new_n11362);
nand_4 g09022(new_n11371, new_n11370, new_n11359);
nand_4 g09023(new_n11372, new_n11371, new_n11355);
xnor_3 g09024(new_n11373, new_n11372, new_n11351);
xor_3  g09025(new_n11374, n12956, new_n10148);
nor_4  g09026(new_n11375_1, new_n10756_1, n8381);
not_3  g09027(new_n11376, new_n11375_1);
nor_4  g09028(new_n11377, n18295, new_n5757);
not_3  g09029(new_n11378, new_n11377);
nor_4  g09030(new_n11379_1, n20235, new_n11146);
not_3  g09031(new_n11380, new_n11379_1);
nor_4  g09032(new_n11381, new_n5778, n6502);
not_3  g09033(new_n11382, new_n11381);
nor_4  g09034(new_n11383, new_n11149, n12495);
nand_4 g09035(new_n11384, new_n11383, new_n11382);
nand_4 g09036(new_n11385, new_n11384, new_n11380);
nand_4 g09037(new_n11386_1, new_n11385, new_n11378);
nand_4 g09038(new_n11387, new_n11386_1, new_n11376);
xor_3  g09039(new_n11388, new_n11387, new_n11374);
xnor_3 g09040(new_n11389, new_n11388, new_n11373);
not_3  g09041(new_n11390, new_n11359);
xnor_3 g09042(new_n11391_1, new_n11370, new_n11390);
nor_4  g09043(new_n11392, new_n11377, new_n11375_1);
xor_3  g09044(new_n11393, new_n11392, new_n11385);
not_3  g09045(new_n11394, new_n11393);
nor_4  g09046(new_n11395, new_n11394, new_n11391_1);
not_3  g09047(new_n11396, new_n11395);
not_3  g09048(new_n11397, new_n11391_1);
nor_4  g09049(new_n11398_1, new_n11393, new_n11397);
nor_4  g09050(new_n11399, new_n11398_1, new_n11395);
xor_3  g09051(new_n11400, n15780, new_n10209);
xor_3  g09052(new_n11401, new_n11364, new_n6729_1);
nor_4  g09053(new_n11402, new_n11401, new_n11400);
nor_4  g09054(new_n11403_1, new_n11381, new_n11379_1);
xor_3  g09055(new_n11404, new_n11403_1, new_n11383);
not_3  g09056(new_n11405, new_n11404);
nor_4  g09057(new_n11406, new_n11405, new_n11402);
not_3  g09058(new_n11407, new_n11406);
xnor_3 g09059(new_n11408, new_n11368, new_n11365);
not_3  g09060(new_n11409, new_n11402);
nor_4  g09061(new_n11410, new_n11404, new_n11409);
nor_4  g09062(new_n11411, new_n11410, new_n11406);
nand_4 g09063(new_n11412, new_n11411, new_n11408);
nand_4 g09064(new_n11413, new_n11412, new_n11407);
nand_4 g09065(new_n11414, new_n11413, new_n11399);
nand_4 g09066(new_n11415, new_n11414, new_n11396);
xor_3  g09067(n1060, new_n11415, new_n11389);
not_3  g09068(new_n11417, new_n3581);
xor_3  g09069(n1069, new_n3634, new_n11417);
xor_3  g09070(new_n11419_1, n9832, n3959);
nor_4  g09071(new_n11420, n11566, n1558);
not_3  g09072(new_n11421, new_n11420);
xor_3  g09073(new_n11422, n11566, n1558);
nor_4  g09074(new_n11423, n26744, n21749);
not_3  g09075(new_n11424_1, new_n11423);
xor_3  g09076(new_n11425, n26744, n21749);
nor_4  g09077(new_n11426, n26625, n7769);
not_3  g09078(new_n11427, new_n11426);
nand_4 g09079(new_n11428, n21138, n14230);
xor_3  g09080(new_n11429, n26625, n7769);
nand_4 g09081(new_n11430, new_n11429, new_n11428);
nand_4 g09082(new_n11431, new_n11430, new_n11427);
nand_4 g09083(new_n11432, new_n11431, new_n11425);
nand_4 g09084(new_n11433, new_n11432, new_n11424_1);
nand_4 g09085(new_n11434, new_n11433, new_n11422);
nand_4 g09086(new_n11435, new_n11434, new_n11421);
nor_4  g09087(new_n11436, new_n11435, new_n11419_1);
nand_4 g09088(new_n11437, new_n11435, new_n11419_1);
not_3  g09089(new_n11438, new_n11437);
nor_4  g09090(new_n11439_1, new_n11438, new_n11436);
not_3  g09091(new_n11440, new_n11439_1);
not_3  g09092(new_n11441, n19575);
not_3  g09093(new_n11442, n17095);
nor_4  g09094(new_n11443, n26167, n22591);
nand_4 g09095(new_n11444, new_n11443, new_n11442);
nor_4  g09096(new_n11445, new_n11444, n15378);
xor_3  g09097(new_n11446, new_n11445, new_n11441);
xnor_3 g09098(new_n11447, new_n7997, new_n10391);
not_3  g09099(new_n11448, new_n11447);
not_3  g09100(new_n11449, n17664);
nor_4  g09101(new_n11450, new_n8002, new_n11449);
not_3  g09102(new_n11451, new_n11450);
xnor_3 g09103(new_n11452, new_n8002, n17664);
nor_4  g09104(new_n11453, new_n8010, new_n10396);
not_3  g09105(new_n11454, new_n11453);
nor_4  g09106(new_n11455_1, new_n8013, n23369);
nor_4  g09107(new_n11456, new_n11455_1, new_n11453);
nor_4  g09108(new_n11457, new_n8022, n1136);
not_3  g09109(new_n11458, n19234);
nor_4  g09110(new_n11459, new_n8018, new_n11458);
xnor_3 g09111(new_n11460, new_n8007, new_n7958);
xnor_3 g09112(new_n11461, new_n11460, new_n10399);
nor_4  g09113(new_n11462_1, new_n11461, new_n11459);
nor_4  g09114(new_n11463, new_n11462_1, new_n11457);
nand_4 g09115(new_n11464, new_n11463, new_n11456);
nand_4 g09116(new_n11465, new_n11464, new_n11454);
nand_4 g09117(new_n11466, new_n11465, new_n11452);
nand_4 g09118(new_n11467, new_n11466, new_n11451);
not_3  g09119(new_n11468, new_n11467);
nor_4  g09120(new_n11469, new_n11468, new_n11448);
nor_4  g09121(new_n11470_1, new_n11467, new_n11447);
nor_4  g09122(new_n11471, new_n11470_1, new_n11469);
xnor_3 g09123(new_n11472_1, new_n11471, new_n11446);
not_3  g09124(new_n11473_1, new_n11472_1);
xnor_3 g09125(new_n11474, new_n8002, new_n11449);
xnor_3 g09126(new_n11475, new_n8010, new_n10396);
not_3  g09127(new_n11476, new_n11457);
not_3  g09128(new_n11477, new_n11459);
nor_4  g09129(new_n11478, new_n11460, new_n10399);
nor_4  g09130(new_n11479_1, new_n11478, new_n11457);
nand_4 g09131(new_n11480, new_n11479_1, new_n11477);
nand_4 g09132(new_n11481_1, new_n11480, new_n11476);
nor_4  g09133(new_n11482, new_n11481_1, new_n11475);
nor_4  g09134(new_n11483, new_n11482, new_n11453);
nor_4  g09135(new_n11484, new_n11483, new_n11474);
nor_4  g09136(new_n11485, new_n11465, new_n11452);
nor_4  g09137(new_n11486_1, new_n11485, new_n11484);
xor_3  g09138(new_n11487, new_n11444, n15378);
nor_4  g09139(new_n11488, new_n11487, new_n11486_1);
xnor_3 g09140(new_n11489, new_n11487, new_n11486_1);
xnor_3 g09141(new_n11490, new_n11481_1, new_n11475);
not_3  g09142(new_n11491, new_n11490);
xor_3  g09143(new_n11492, new_n11443, new_n11442);
nor_4  g09144(new_n11493, new_n11492, new_n11491);
xnor_3 g09145(new_n11494, new_n11492, new_n11491);
nor_4  g09146(new_n11495, new_n11479_1, new_n11477);
nor_4  g09147(new_n11496_1, new_n11495, new_n11462_1);
not_3  g09148(new_n11497, n22591);
nor_4  g09149(new_n11498, new_n8493, new_n8491);
xnor_3 g09150(new_n11499, new_n11498, new_n11497);
not_3  g09151(new_n11500, new_n11499);
nor_4  g09152(new_n11501, new_n11500, new_n11496_1);
nor_4  g09153(new_n11502, new_n8492, new_n8491);
not_3  g09154(new_n11503_1, new_n11502);
nor_4  g09155(new_n11504, new_n11503_1, n22591);
nor_4  g09156(new_n11505, new_n11504, new_n11501);
not_3  g09157(new_n11506_1, new_n11505);
nor_4  g09158(new_n11507, new_n11506_1, new_n11494);
nor_4  g09159(new_n11508, new_n11507, new_n11493);
nor_4  g09160(new_n11509, new_n11508, new_n11489);
nor_4  g09161(new_n11510, new_n11509, new_n11488);
not_3  g09162(new_n11511, new_n11510);
nor_4  g09163(new_n11512, new_n11511, new_n11473_1);
nor_4  g09164(new_n11513, new_n11510, new_n11472_1);
nor_4  g09165(new_n11514, new_n11513, new_n11512);
xnor_3 g09166(new_n11515_1, new_n11514, new_n11440);
xnor_3 g09167(new_n11516, new_n11508, new_n11489);
not_3  g09168(new_n11517, new_n11516);
not_3  g09169(new_n11518, new_n11422);
not_3  g09170(new_n11519, new_n11433);
xor_3  g09171(new_n11520, new_n11519, new_n11518);
not_3  g09172(new_n11521, new_n11520);
nand_4 g09173(new_n11522, new_n11521, new_n11517);
not_3  g09174(new_n11523, new_n11522);
nor_4  g09175(new_n11524, new_n11521, new_n11517);
nor_4  g09176(new_n11525, new_n11524, new_n11523);
not_3  g09177(new_n11526, new_n11494);
nor_4  g09178(new_n11527, new_n11505, new_n11526);
nor_4  g09179(new_n11528, new_n11527, new_n11507);
xnor_3 g09180(new_n11529, new_n11431, new_n11425);
nor_4  g09181(new_n11530, new_n11529, new_n11528);
xnor_3 g09182(new_n11531, new_n11529, new_n11528);
xnor_3 g09183(new_n11532, new_n11500, new_n11496_1);
not_3  g09184(new_n11533, new_n11532);
not_3  g09185(new_n11534, new_n11428);
xnor_3 g09186(new_n11535, new_n11429, new_n11534);
nor_4  g09187(new_n11536, new_n11535, new_n11533);
not_3  g09188(new_n11537, new_n11536);
not_3  g09189(new_n11538_1, new_n8490);
nor_4  g09190(new_n11539, new_n8495, new_n11538_1);
not_3  g09191(new_n11540, new_n11535);
nor_4  g09192(new_n11541, new_n11540, new_n11532);
nor_4  g09193(new_n11542, new_n11541, new_n11536);
nand_4 g09194(new_n11543, new_n11542, new_n11539);
nand_4 g09195(new_n11544, new_n11543, new_n11537);
nor_4  g09196(new_n11545, new_n11544, new_n11531);
nor_4  g09197(new_n11546, new_n11545, new_n11530);
nand_4 g09198(new_n11547, new_n11546, new_n11525);
nand_4 g09199(new_n11548_1, new_n11547, new_n11522);
xor_3  g09200(n1111, new_n11548_1, new_n11515_1);
xnor_3 g09201(new_n11550, new_n2672, new_n5007);
nor_4  g09202(new_n11551, new_n2680_1, new_n5013);
xnor_3 g09203(new_n11552, new_n2680_1, new_n5013);
nand_4 g09204(new_n11553, new_n2687, new_n5022);
nand_4 g09205(new_n11554, new_n2691, new_n4335);
not_3  g09206(new_n11555, new_n11554);
nor_4  g09207(new_n11556, new_n2691, new_n4335);
nor_4  g09208(new_n11557, new_n11556, new_n11555);
not_3  g09209(new_n11558, new_n2698);
nand_4 g09210(new_n11559, new_n11558, new_n4355);
xnor_3 g09211(new_n11560, new_n2698, new_n4355);
nor_4  g09212(new_n11561, new_n2706_1, n16476);
not_3  g09213(new_n11562, new_n11561);
nor_4  g09214(new_n11563, new_n2703_1, new_n4359);
nor_4  g09215(new_n11564_1, new_n11563, new_n11561);
nor_4  g09216(new_n11565, new_n2731_1, n11615);
not_3  g09217(new_n11566_1, new_n11565);
nor_4  g09218(new_n11567, new_n2716, n22433);
not_3  g09219(new_n11568, new_n11567);
nor_4  g09220(new_n11569, new_n2720, new_n6409);
not_3  g09221(new_n11570, new_n11569);
nor_4  g09222(new_n11571, new_n2726, new_n4375);
nor_4  g09223(new_n11572, new_n11571, new_n11567);
nand_4 g09224(new_n11573, new_n11572, new_n11570);
nand_4 g09225(new_n11574, new_n11573, new_n11568);
nor_4  g09226(new_n11575, new_n2711_1, new_n4371);
nor_4  g09227(new_n11576, new_n11575, new_n11565);
nand_4 g09228(new_n11577, new_n11576, new_n11574);
nand_4 g09229(new_n11578, new_n11577, new_n11566_1);
nand_4 g09230(new_n11579_1, new_n11578, new_n11564_1);
nand_4 g09231(new_n11580_1, new_n11579_1, new_n11562);
nand_4 g09232(new_n11581, new_n11580_1, new_n11560);
nand_4 g09233(new_n11582, new_n11581, new_n11559);
nand_4 g09234(new_n11583, new_n11582, new_n11557);
nand_4 g09235(new_n11584, new_n11583, new_n11554);
not_3  g09236(new_n11585, new_n11553);
nor_4  g09237(new_n11586, new_n2687, new_n5022);
nor_4  g09238(new_n11587, new_n11586, new_n11585);
nand_4 g09239(new_n11588, new_n11587, new_n11584);
nand_4 g09240(new_n11589, new_n11588, new_n11553);
nor_4  g09241(new_n11590, new_n11589, new_n11552);
nor_4  g09242(new_n11591_1, new_n11590, new_n11551);
xnor_3 g09243(new_n11592, new_n11591_1, new_n11550);
not_3  g09244(new_n11593, new_n11592);
nand_4 g09245(new_n11594, new_n11320, new_n4868);
nor_4  g09246(new_n11595, new_n11594, n20929);
nand_4 g09247(new_n11596, new_n11595, new_n3080);
nor_4  g09248(new_n11597, new_n11596, n11841);
not_3  g09249(new_n11598, new_n11597);
xor_3  g09250(new_n11599, new_n11598, n27089);
not_3  g09251(new_n11600, new_n11599);
xnor_3 g09252(new_n11601, new_n11600, new_n2826_1);
xor_3  g09253(new_n11602, new_n11596, n11841);
not_3  g09254(new_n11603, new_n11602);
nor_4  g09255(new_n11604, new_n11603, new_n2831);
xnor_3 g09256(new_n11605, new_n11603, new_n2831);
xor_3  g09257(new_n11606, new_n11595, new_n3080);
not_3  g09258(new_n11607_1, new_n11606);
nand_4 g09259(new_n11608, new_n11607_1, new_n2842);
xnor_3 g09260(new_n11609, new_n11606, new_n2842);
not_3  g09261(new_n11610, n20929);
xor_3  g09262(new_n11611, new_n11594, new_n11610);
nand_4 g09263(new_n11612, new_n11611, new_n2851);
xor_3  g09264(new_n11613, new_n11594, n20929);
xnor_3 g09265(new_n11614, new_n11613, new_n2851);
xor_3  g09266(new_n11615_1, new_n11320, new_n4868);
not_3  g09267(new_n11616, new_n11615_1);
nand_4 g09268(new_n11617, new_n11616, new_n2895);
nand_4 g09269(new_n11618, new_n11324, new_n2862);
not_3  g09270(new_n11619, new_n2792);
xnor_3 g09271(new_n11620, new_n2805, new_n11619);
xnor_3 g09272(new_n11621, new_n11324, new_n11620);
nor_4  g09273(new_n11622, new_n11331, new_n2869);
not_3  g09274(new_n11623, new_n11622);
nor_4  g09275(new_n11624, new_n11332, new_n2873);
nor_4  g09276(new_n11625, new_n11624, new_n11622);
nor_4  g09277(new_n11626, new_n6749, new_n2879);
nand_4 g09278(new_n11627, new_n2883, new_n4885);
xnor_3 g09279(new_n11628, new_n6749, new_n2879);
nor_4  g09280(new_n11629, new_n11628, new_n11627);
nor_4  g09281(new_n11630_1, new_n11629, new_n11626);
not_3  g09282(new_n11631, new_n11630_1);
nand_4 g09283(new_n11632, new_n11631, new_n11625);
nand_4 g09284(new_n11633, new_n11632, new_n11623);
nand_4 g09285(new_n11634, new_n11633, new_n11621);
nand_4 g09286(new_n11635, new_n11634, new_n11618);
xnor_3 g09287(new_n11636, new_n11615_1, new_n2895);
nand_4 g09288(new_n11637, new_n11636, new_n11635);
nand_4 g09289(new_n11638, new_n11637, new_n11617);
nand_4 g09290(new_n11639, new_n11638, new_n11614);
nand_4 g09291(new_n11640, new_n11639, new_n11612);
nand_4 g09292(new_n11641, new_n11640, new_n11609);
nand_4 g09293(new_n11642, new_n11641, new_n11608);
nor_4  g09294(new_n11643, new_n11642, new_n11605);
nor_4  g09295(new_n11644, new_n11643, new_n11604);
xnor_3 g09296(new_n11645, new_n11644, new_n11601);
xnor_3 g09297(new_n11646, new_n11645, new_n11593);
xnor_3 g09298(new_n11647_1, new_n11589, new_n11552);
not_3  g09299(new_n11648, new_n11647_1);
not_3  g09300(new_n11649, new_n11642);
xnor_3 g09301(new_n11650, new_n11649, new_n11605);
nand_4 g09302(new_n11651, new_n11650, new_n11648);
xnor_3 g09303(new_n11652, new_n11650, new_n11647_1);
xnor_3 g09304(new_n11653, new_n11587, new_n11584);
xnor_3 g09305(new_n11654, new_n11640, new_n11609);
nor_4  g09306(new_n11655, new_n11654, new_n11653);
xnor_3 g09307(new_n11656, new_n11654, new_n11653);
not_3  g09308(new_n11657, new_n11582);
xnor_3 g09309(new_n11658, new_n11657, new_n11557);
not_3  g09310(new_n11659, new_n11658);
xnor_3 g09311(new_n11660, new_n11638, new_n11614);
nand_4 g09312(new_n11661, new_n11660, new_n11659);
xnor_3 g09313(new_n11662, new_n11660, new_n11658);
xnor_3 g09314(new_n11663, new_n11580_1, new_n11560);
not_3  g09315(new_n11664, new_n11635);
xnor_3 g09316(new_n11665, new_n11636, new_n11664);
not_3  g09317(new_n11666, new_n11665);
nand_4 g09318(new_n11667_1, new_n11666, new_n11663);
xnor_3 g09319(new_n11668, new_n11665, new_n11663);
xnor_3 g09320(new_n11669, new_n11633, new_n11621);
xnor_3 g09321(new_n11670, new_n11578, new_n11564_1);
nand_4 g09322(new_n11671, new_n11670, new_n11669);
xnor_3 g09323(new_n11672, new_n2716, n22433);
nor_4  g09324(new_n11673, new_n11672, new_n11569);
nor_4  g09325(new_n11674_1, new_n11673, new_n11567);
xnor_3 g09326(new_n11675, new_n2711_1, new_n4371);
nor_4  g09327(new_n11676, new_n11675, new_n11674_1);
nor_4  g09328(new_n11677, new_n11676, new_n11565);
xnor_3 g09329(new_n11678, new_n11677, new_n11564_1);
xnor_3 g09330(new_n11679, new_n11678, new_n11669);
xnor_3 g09331(new_n11680, new_n11631, new_n11625);
xnor_3 g09332(new_n11681, new_n11675, new_n11674_1);
nand_4 g09333(new_n11682_1, new_n11681, new_n11680);
not_3  g09334(new_n11683, new_n11681);
xnor_3 g09335(new_n11684, new_n11683, new_n11680);
xnor_3 g09336(new_n11685, new_n11628, new_n11627);
nor_4  g09337(new_n11686, new_n11572, new_n11570);
nor_4  g09338(new_n11687, new_n11686, new_n11673);
not_3  g09339(new_n11688, new_n11687);
nor_4  g09340(new_n11689, new_n11688, new_n11685);
xnor_3 g09341(new_n11690, new_n2720, n14090);
not_3  g09342(new_n11691, new_n11690);
not_3  g09343(new_n11692, new_n11627);
nor_4  g09344(new_n11693, new_n2883, new_n4885);
nor_4  g09345(new_n11694, new_n11693, new_n11692);
nor_4  g09346(new_n11695, new_n11694, new_n11691);
xnor_3 g09347(new_n11696, new_n11688, new_n11685);
nor_4  g09348(new_n11697, new_n11696, new_n11695);
nor_4  g09349(new_n11698, new_n11697, new_n11689);
nand_4 g09350(new_n11699, new_n11698, new_n11684);
nand_4 g09351(new_n11700, new_n11699, new_n11682_1);
nand_4 g09352(new_n11701, new_n11700, new_n11679);
nand_4 g09353(new_n11702, new_n11701, new_n11671);
nand_4 g09354(new_n11703, new_n11702, new_n11668);
nand_4 g09355(new_n11704, new_n11703, new_n11667_1);
nand_4 g09356(new_n11705, new_n11704, new_n11662);
nand_4 g09357(new_n11706, new_n11705, new_n11661);
nor_4  g09358(new_n11707, new_n11706, new_n11656);
nor_4  g09359(new_n11708, new_n11707, new_n11655);
nand_4 g09360(new_n11709, new_n11708, new_n11652);
nand_4 g09361(new_n11710_1, new_n11709, new_n11651);
xnor_3 g09362(n1119, new_n11710_1, new_n11646);
nand_4 g09363(new_n11712_1, new_n9359, new_n9358);
xor_3  g09364(n1120, new_n11712_1, new_n9380_1);
xnor_3 g09365(new_n11714, n9246, n3925);
not_3  g09366(new_n11715, new_n11714);
xor_3  g09367(new_n11716, new_n11715, new_n9221);
xor_3  g09368(new_n11717, n12495, new_n9869);
xor_3  g09369(n1196, new_n11717, new_n11716);
not_3  g09370(new_n11719, new_n9360);
xor_3  g09371(new_n11720, n16223, n15636);
nor_4  g09372(new_n11721, new_n6406, n19494);
nor_4  g09373(new_n11722, n20077, new_n2372);
nor_4  g09374(new_n11723, new_n6575, n2387);
not_3  g09375(new_n11724_1, new_n11723);
nor_4  g09376(new_n11725, new_n11724_1, new_n11722);
nor_4  g09377(new_n11726, new_n11725, new_n11721);
xor_3  g09378(new_n11727, new_n11726, new_n11720);
xnor_3 g09379(new_n11728, new_n11727, new_n11719);
xor_3  g09380(new_n11729, n6794, new_n2571);
nor_4  g09381(new_n11730, new_n11729, new_n9369);
nor_4  g09382(new_n11731, new_n11722, new_n11721);
xor_3  g09383(new_n11732, new_n11731, new_n11723);
not_3  g09384(new_n11733, new_n11732);
nor_4  g09385(new_n11734, new_n11733, new_n11730);
not_3  g09386(new_n11735, new_n11734);
not_3  g09387(new_n11736_1, new_n11730);
nor_4  g09388(new_n11737, new_n11732, new_n11736_1);
nor_4  g09389(new_n11738, new_n11737, new_n11734);
nand_4 g09390(new_n11739, new_n11738, new_n9362);
nand_4 g09391(new_n11740, new_n11739, new_n11735);
not_3  g09392(new_n11741_1, new_n11740);
xor_3  g09393(n1237, new_n11741_1, new_n11728);
not_3  g09394(new_n11743, new_n6635);
not_3  g09395(new_n11744, new_n6633);
not_3  g09396(new_n11745, new_n6634_1);
nor_4  g09397(new_n11746, new_n11745, new_n11744);
nor_4  g09398(new_n11747, new_n11746, new_n6635);
not_3  g09399(new_n11748, new_n6639);
not_3  g09400(new_n11749_1, new_n6647);
nand_4 g09401(new_n11750, new_n6712, new_n11749_1);
nand_4 g09402(new_n11751, new_n11750, new_n6643);
nand_4 g09403(new_n11752, new_n11751, new_n11748);
nand_4 g09404(new_n11753, new_n11752, new_n11747);
nand_4 g09405(new_n11754, new_n11753, new_n11743);
nor_4  g09406(new_n11755, new_n6631_1, new_n6628_1);
xnor_3 g09407(n1239, new_n11755, new_n11754);
xor_3  g09408(new_n11757, n22764, n1536);
not_3  g09409(new_n11758, new_n11757);
nor_4  g09410(new_n11759, n26264, n19454);
xor_3  g09411(new_n11760, n26264, n19454);
not_3  g09412(new_n11761, new_n11760);
nor_4  g09413(new_n11762, n9445, n7841);
xor_3  g09414(new_n11763, n9445, n7841);
not_3  g09415(new_n11764, new_n11763);
nand_4 g09416(new_n11765, new_n9460_1, new_n9588);
xor_3  g09417(new_n11766, n16812, n1279);
nor_4  g09418(new_n11767, n25068, n8324);
not_3  g09419(new_n11768, new_n11767);
xor_3  g09420(new_n11769, n25068, n8324);
nor_4  g09421(new_n11770_1, n12546, n2331);
not_3  g09422(new_n11771_1, new_n11770_1);
xor_3  g09423(new_n11772, n12546, n2331);
nor_4  g09424(new_n11773, n22631, n21078);
not_3  g09425(new_n11774, new_n11773);
xor_3  g09426(new_n11775_1, n22631, n21078);
nor_4  g09427(new_n11776, n24485, n16743);
not_3  g09428(new_n11777, new_n11776);
xor_3  g09429(new_n11778, n24485, n16743);
nand_4 g09430(new_n11779, new_n9492, new_n9626_1);
nand_4 g09431(new_n11780, n22201, n4588);
xor_3  g09432(new_n11781, n15258, n2420);
nand_4 g09433(new_n11782, new_n11781, new_n11780);
nand_4 g09434(new_n11783, new_n11782, new_n11779);
nand_4 g09435(new_n11784, new_n11783, new_n11778);
nand_4 g09436(new_n11785, new_n11784, new_n11777);
nand_4 g09437(new_n11786, new_n11785, new_n11775_1);
nand_4 g09438(new_n11787, new_n11786, new_n11774);
nand_4 g09439(new_n11788, new_n11787, new_n11772);
nand_4 g09440(new_n11789, new_n11788, new_n11771_1);
nand_4 g09441(new_n11790, new_n11789, new_n11769);
nand_4 g09442(new_n11791, new_n11790, new_n11768);
nand_4 g09443(new_n11792, new_n11791, new_n11766);
nand_4 g09444(new_n11793, new_n11792, new_n11765);
not_3  g09445(new_n11794, new_n11793);
nor_4  g09446(new_n11795, new_n11794, new_n11764);
nor_4  g09447(new_n11796, new_n11795, new_n11762);
nor_4  g09448(new_n11797, new_n11796, new_n11761);
nor_4  g09449(new_n11798, new_n11797, new_n11759);
xor_3  g09450(new_n11799, new_n11798, new_n11758);
not_3  g09451(new_n11800, new_n11799);
nor_4  g09452(new_n11801, new_n11800, n2416);
not_3  g09453(new_n11802, n2416);
xnor_3 g09454(new_n11803, new_n11799, new_n11802);
xor_3  g09455(new_n11804, new_n11796, new_n11760);
nor_4  g09456(new_n11805, new_n11804, n21905);
not_3  g09457(new_n11806, n21905);
xor_3  g09458(new_n11807, new_n11796, new_n11761);
nor_4  g09459(new_n11808, new_n11807, new_n11806);
nor_4  g09460(new_n11809, new_n11808, new_n11805);
not_3  g09461(new_n11810, new_n11809);
xor_3  g09462(new_n11811, new_n11794, new_n11763);
nor_4  g09463(new_n11812, new_n11811, n22918);
not_3  g09464(new_n11813, n22918);
xnor_3 g09465(new_n11814, new_n11811, new_n11813);
not_3  g09466(new_n11815, n25923);
xnor_3 g09467(new_n11816, new_n11791, new_n11766);
not_3  g09468(new_n11817, new_n11816);
nand_4 g09469(new_n11818_1, new_n11817, new_n11815);
xnor_3 g09470(new_n11819, new_n11816, new_n11815);
not_3  g09471(new_n11820, n6790);
xnor_3 g09472(new_n11821, new_n11789, new_n11769);
not_3  g09473(new_n11822, new_n11821);
nand_4 g09474(new_n11823, new_n11822, new_n11820);
xnor_3 g09475(new_n11824, new_n11821, new_n11820);
xnor_3 g09476(new_n11825, new_n11787, new_n11772);
nor_4  g09477(new_n11826, new_n11825, n22879);
not_3  g09478(new_n11827, new_n11826);
not_3  g09479(new_n11828, n22879);
xnor_3 g09480(new_n11829, new_n11825, new_n11828);
not_3  g09481(new_n11830, n2117);
not_3  g09482(new_n11831, new_n11775_1);
xnor_3 g09483(new_n11832, new_n11785, new_n11831);
nand_4 g09484(new_n11833, new_n11832, new_n11830);
xnor_3 g09485(new_n11834, new_n11832, n2117);
xnor_3 g09486(new_n11835, new_n11783, new_n11778);
nor_4  g09487(new_n11836, new_n11835, n5882);
not_3  g09488(new_n11837_1, new_n11836);
xnor_3 g09489(new_n11838, n15258, n2420);
xor_3  g09490(new_n11839, new_n11838, new_n11780);
nor_4  g09491(new_n11840, new_n11839, n11775);
not_3  g09492(new_n11841_1, new_n11840);
not_3  g09493(new_n11842_1, n27134);
xor_3  g09494(new_n11843_1, n22201, n4588);
not_3  g09495(new_n11844, new_n11843_1);
nor_4  g09496(new_n11845, new_n11844, new_n11842_1);
not_3  g09497(new_n11846, new_n11845);
not_3  g09498(new_n11847, n11775);
not_3  g09499(new_n11848, new_n11780);
xor_3  g09500(new_n11849, new_n11838, new_n11848);
xnor_3 g09501(new_n11850, new_n11849, new_n11847);
not_3  g09502(new_n11851, new_n11850);
nand_4 g09503(new_n11852, new_n11851, new_n11846);
nand_4 g09504(new_n11853, new_n11852, new_n11841_1);
not_3  g09505(new_n11854, n5882);
not_3  g09506(new_n11855, new_n11778);
xnor_3 g09507(new_n11856, new_n11783, new_n11855);
nor_4  g09508(new_n11857, new_n11856, new_n11854);
nor_4  g09509(new_n11858, new_n11857, new_n11836);
nand_4 g09510(new_n11859, new_n11858, new_n11853);
nand_4 g09511(new_n11860, new_n11859, new_n11837_1);
nand_4 g09512(new_n11861, new_n11860, new_n11834);
nand_4 g09513(new_n11862, new_n11861, new_n11833);
nand_4 g09514(new_n11863, new_n11862, new_n11829);
nand_4 g09515(new_n11864, new_n11863, new_n11827);
nand_4 g09516(new_n11865, new_n11864, new_n11824);
nand_4 g09517(new_n11866, new_n11865, new_n11823);
nand_4 g09518(new_n11867, new_n11866, new_n11819);
nand_4 g09519(new_n11868, new_n11867, new_n11818_1);
nand_4 g09520(new_n11869, new_n11868, new_n11814);
not_3  g09521(new_n11870, new_n11869);
nor_4  g09522(new_n11871, new_n11870, new_n11812);
nor_4  g09523(new_n11872, new_n11871, new_n11810);
nor_4  g09524(new_n11873, new_n11872, new_n11805);
nor_4  g09525(new_n11874, new_n11873, new_n11803);
nor_4  g09526(new_n11875, new_n11874, new_n11801);
nor_4  g09527(new_n11876, n22764, n1536);
nor_4  g09528(new_n11877, new_n11798, new_n11758);
nor_4  g09529(new_n11878, new_n11877, new_n11876);
nand_4 g09530(new_n11879, new_n11878, new_n11875);
nor_4  g09531(new_n11880, n23493, n8405);
nor_4  g09532(new_n11881, n22359, n10275);
not_3  g09533(new_n11882, n5532);
nand_4 g09534(new_n11883, new_n9403_1, new_n11882);
not_3  g09535(new_n11884, n3962);
not_3  g09536(new_n11885, n11579);
nand_4 g09537(new_n11886, new_n11885, new_n11884);
not_3  g09538(new_n11887, n21);
not_3  g09539(new_n11888, n23513);
nand_4 g09540(new_n11889, new_n11888, new_n11887);
xor_3  g09541(new_n11890, n23513, n21);
not_3  g09542(new_n11891, n1682);
not_3  g09543(new_n11892, n6427);
nand_4 g09544(new_n11893, new_n11892, new_n11891);
nand_4 g09545(new_n11894, n6427, n1682);
not_3  g09546(new_n11895, n6590);
not_3  g09547(new_n11896, n7963);
nand_4 g09548(new_n11897, new_n11896, new_n11895);
not_3  g09549(new_n11898_1, n10017);
not_3  g09550(new_n11899, n20349);
nand_4 g09551(new_n11900, new_n11899, new_n11898_1);
nand_4 g09552(new_n11901, n15936, n3618);
nand_4 g09553(new_n11902, n20349, n10017);
nand_4 g09554(new_n11903, new_n11902, new_n11901);
nand_4 g09555(new_n11904, new_n11903, new_n11900);
nand_4 g09556(new_n11905_1, n7963, n6590);
nand_4 g09557(new_n11906, new_n11905_1, new_n11904);
nand_4 g09558(new_n11907, new_n11906, new_n11897);
nand_4 g09559(new_n11908, new_n11907, new_n11894);
nand_4 g09560(new_n11909, new_n11908, new_n11893);
nand_4 g09561(new_n11910, new_n11909, new_n11890);
nand_4 g09562(new_n11911, new_n11910, new_n11889);
xor_3  g09563(new_n11912, n11579, n3962);
nand_4 g09564(new_n11913, new_n11912, new_n11911);
nand_4 g09565(new_n11914, new_n11913, new_n11886);
xor_3  g09566(new_n11915, n15146, new_n11882);
not_3  g09567(new_n11916, new_n11915);
nand_4 g09568(new_n11917, new_n11916, new_n11914);
nand_4 g09569(new_n11918, new_n11917, new_n11883);
not_3  g09570(new_n11919, n10275);
xor_3  g09571(new_n11920, n22359, new_n11919);
not_3  g09572(new_n11921, new_n11920);
nand_4 g09573(new_n11922, new_n11921, new_n11918);
not_3  g09574(new_n11923, new_n11922);
nor_4  g09575(new_n11924, new_n11923, new_n11881);
not_3  g09576(new_n11925, n23493);
xor_3  g09577(new_n11926_1, new_n11925, n8405);
nor_4  g09578(new_n11927, new_n11926_1, new_n11924);
nor_4  g09579(new_n11928, new_n11927, new_n11880);
not_3  g09580(new_n11929, n14826);
xor_3  g09581(new_n11930, new_n11929, n13549);
not_3  g09582(new_n11931, new_n11930);
xor_3  g09583(new_n11932, new_n11931, new_n11928);
nor_4  g09584(new_n11933, new_n11932, n18105);
not_3  g09585(new_n11934, new_n11933);
not_3  g09586(new_n11935, new_n11932);
nor_4  g09587(new_n11936, new_n11935, new_n4985);
nor_4  g09588(new_n11937, new_n11936, new_n11933);
not_3  g09589(new_n11938, new_n11926_1);
xor_3  g09590(new_n11939, new_n11938, new_n11924);
nor_4  g09591(new_n11940, new_n11939, n24196);
xnor_3 g09592(new_n11941, new_n11939, n24196);
xnor_3 g09593(new_n11942, new_n11921, new_n11918);
nor_4  g09594(new_n11943, new_n11942, n16376);
not_3  g09595(new_n11944, new_n11942);
xor_3  g09596(new_n11945, new_n11944, new_n5055);
not_3  g09597(new_n11946, new_n11945);
xnor_3 g09598(new_n11947, new_n11915, new_n11914);
not_3  g09599(new_n11948, new_n11947);
nor_4  g09600(new_n11949, new_n11948, n25381);
xor_3  g09601(new_n11950, new_n11948, n25381);
not_3  g09602(new_n11951, new_n11950);
xnor_3 g09603(new_n11952, new_n11912, new_n11911);
nor_4  g09604(new_n11953, new_n11952, n12587);
not_3  g09605(new_n11954, new_n11952);
xor_3  g09606(new_n11955, new_n11954, new_n5070);
not_3  g09607(new_n11956, new_n11955);
xor_3  g09608(new_n11957, n23513, new_n11887);
xnor_3 g09609(new_n11958, new_n11909, new_n11957);
nand_4 g09610(new_n11959, new_n11958, new_n5077_1);
xnor_3 g09611(new_n11960, new_n11958, n268);
nand_4 g09612(new_n11961, new_n11894, new_n11893);
xor_3  g09613(new_n11962, new_n11961, new_n11907);
not_3  g09614(new_n11963, new_n11962);
nand_4 g09615(new_n11964, new_n11963, new_n5082_1);
xnor_3 g09616(new_n11965_1, new_n11962, new_n5082_1);
nor_4  g09617(new_n11966, new_n11896, n6590);
nor_4  g09618(new_n11967, n7963, new_n11895);
nor_4  g09619(new_n11968, new_n11967, new_n11966);
not_3  g09620(new_n11969, new_n11968);
xor_3  g09621(new_n11970, new_n11969, new_n11904);
nand_4 g09622(new_n11971, new_n11970, new_n4986);
not_3  g09623(new_n11972, new_n11901);
nor_4  g09624(new_n11973, n20349, new_n11898_1);
nor_4  g09625(new_n11974, new_n11899, n10017);
nor_4  g09626(new_n11975, new_n11974, new_n11973);
xnor_3 g09627(new_n11976, new_n11975, new_n11972);
nor_4  g09628(new_n11977, new_n11976, n24032);
not_3  g09629(new_n11978, new_n11977);
not_3  g09630(new_n11979, n15936);
nor_4  g09631(new_n11980_1, new_n11979, n3618);
not_3  g09632(new_n11981, n3618);
nor_4  g09633(new_n11982, n15936, new_n11981);
nor_4  g09634(new_n11983, new_n11982, new_n11980_1);
nor_4  g09635(new_n11984, new_n11983, new_n5089);
not_3  g09636(new_n11985, new_n11984);
not_3  g09637(new_n11986, new_n11976);
nor_4  g09638(new_n11987, new_n11986, new_n9547);
nor_4  g09639(new_n11988, new_n11987, new_n11977);
nand_4 g09640(new_n11989, new_n11988, new_n11985);
nand_4 g09641(new_n11990, new_n11989, new_n11978);
xnor_3 g09642(new_n11991, new_n11970, n6785);
nand_4 g09643(new_n11992, new_n11991, new_n11990);
nand_4 g09644(new_n11993, new_n11992, new_n11971);
nand_4 g09645(new_n11994, new_n11993, new_n11965_1);
nand_4 g09646(new_n11995, new_n11994, new_n11964);
nand_4 g09647(new_n11996, new_n11995, new_n11960);
nand_4 g09648(new_n11997, new_n11996, new_n11959);
not_3  g09649(new_n11998, new_n11997);
nor_4  g09650(new_n11999, new_n11998, new_n11956);
nor_4  g09651(new_n12000_1, new_n11999, new_n11953);
nor_4  g09652(new_n12001, new_n12000_1, new_n11951);
nor_4  g09653(new_n12002, new_n12001, new_n11949);
nor_4  g09654(new_n12003_1, new_n12002, new_n11946);
nor_4  g09655(new_n12004, new_n12003_1, new_n11943);
nor_4  g09656(new_n12005, new_n12004, new_n11941);
nor_4  g09657(new_n12006, new_n12005, new_n11940);
not_3  g09658(new_n12007, new_n12006);
nand_4 g09659(new_n12008, new_n12007, new_n11937);
nand_4 g09660(new_n12009, new_n12008, new_n11934);
nor_4  g09661(new_n12010, new_n11930, new_n11928);
nor_4  g09662(new_n12011_1, n14826, n13549);
nor_4  g09663(new_n12012, new_n12011_1, new_n12010);
not_3  g09664(new_n12013, new_n12012);
nor_4  g09665(new_n12014, new_n12013, new_n12009);
not_3  g09666(new_n12015, new_n12014);
xnor_3 g09667(new_n12016, new_n12015, new_n11879);
xnor_3 g09668(new_n12017, new_n11878, new_n11875);
xnor_3 g09669(new_n12018, new_n12012, new_n12009);
nand_4 g09670(new_n12019, new_n12018, new_n12017);
xnor_3 g09671(new_n12020, new_n12013, new_n12009);
xnor_3 g09672(new_n12021, new_n12020, new_n12017);
not_3  g09673(new_n12022, new_n11803);
xnor_3 g09674(new_n12023, new_n11873, new_n12022);
xnor_3 g09675(new_n12024, new_n12006, new_n11937);
not_3  g09676(new_n12025, new_n12024);
nand_4 g09677(new_n12026, new_n12025, new_n12023);
xnor_3 g09678(new_n12027, new_n12024, new_n12023);
xnor_3 g09679(new_n12028, new_n11871, new_n11809);
xnor_3 g09680(new_n12029, new_n12004, new_n11941);
nand_4 g09681(new_n12030, new_n12029, new_n12028);
not_3  g09682(new_n12031, new_n12029);
xnor_3 g09683(new_n12032, new_n12031, new_n12028);
xnor_3 g09684(new_n12033, new_n11868, new_n11814);
not_3  g09685(new_n12034, new_n12033);
xnor_3 g09686(new_n12035, new_n12002, new_n11946);
nand_4 g09687(new_n12036, new_n12035, new_n12034);
xnor_3 g09688(new_n12037, new_n12035, new_n12033);
xnor_3 g09689(new_n12038, new_n11866, new_n11819);
not_3  g09690(new_n12039, new_n12038);
xnor_3 g09691(new_n12040, new_n12000_1, new_n11951);
nand_4 g09692(new_n12041, new_n12040, new_n12039);
xnor_3 g09693(new_n12042, new_n12040, new_n12038);
xnor_3 g09694(new_n12043, new_n11864, new_n11824);
not_3  g09695(new_n12044, new_n12043);
xnor_3 g09696(new_n12045, new_n11997, new_n11955);
nand_4 g09697(new_n12046, new_n12045, new_n12044);
xnor_3 g09698(new_n12047, new_n12045, new_n12043);
not_3  g09699(new_n12048, new_n11829);
xnor_3 g09700(new_n12049, new_n11862, new_n12048);
xnor_3 g09701(new_n12050, new_n11995, new_n11960);
nand_4 g09702(new_n12051, new_n12050, new_n12049);
not_3  g09703(new_n12052, new_n11960);
xnor_3 g09704(new_n12053, new_n11995, new_n12052);
xnor_3 g09705(new_n12054, new_n12053, new_n12049);
xnor_3 g09706(new_n12055, new_n11860, new_n11834);
not_3  g09707(new_n12056, new_n12055);
xnor_3 g09708(new_n12057, new_n11993, new_n11965_1);
nand_4 g09709(new_n12058, new_n12057, new_n12056);
xnor_3 g09710(new_n12059, new_n12057, new_n12055);
xnor_3 g09711(new_n12060, new_n11858, new_n11853);
not_3  g09712(new_n12061, new_n12060);
xnor_3 g09713(new_n12062, new_n11991, new_n11990);
nand_4 g09714(new_n12063, new_n12062, new_n12061);
xnor_3 g09715(new_n12064, new_n12062, new_n12060);
xor_3  g09716(new_n12065, new_n11851, new_n11845);
not_3  g09717(new_n12066, new_n12065);
xnor_3 g09718(new_n12067, new_n11988, new_n11985);
nand_4 g09719(new_n12068, new_n12067, new_n12066);
nor_4  g09720(new_n12069, new_n11843_1, n27134);
nor_4  g09721(new_n12070, new_n12069, new_n11845);
xor_3  g09722(new_n12071, new_n11983, n22843);
nor_4  g09723(new_n12072_1, new_n12071, new_n12070);
xnor_3 g09724(new_n12073, new_n12067, new_n12065);
nand_4 g09725(new_n12074, new_n12073, new_n12072_1);
nand_4 g09726(new_n12075, new_n12074, new_n12068);
nand_4 g09727(new_n12076, new_n12075, new_n12064);
nand_4 g09728(new_n12077, new_n12076, new_n12063);
nand_4 g09729(new_n12078, new_n12077, new_n12059);
nand_4 g09730(new_n12079, new_n12078, new_n12058);
nand_4 g09731(new_n12080, new_n12079, new_n12054);
nand_4 g09732(new_n12081, new_n12080, new_n12051);
nand_4 g09733(new_n12082, new_n12081, new_n12047);
nand_4 g09734(new_n12083, new_n12082, new_n12046);
nand_4 g09735(new_n12084, new_n12083, new_n12042);
nand_4 g09736(new_n12085, new_n12084, new_n12041);
nand_4 g09737(new_n12086, new_n12085, new_n12037);
nand_4 g09738(new_n12087, new_n12086, new_n12036);
nand_4 g09739(new_n12088, new_n12087, new_n12032);
nand_4 g09740(new_n12089, new_n12088, new_n12030);
nand_4 g09741(new_n12090, new_n12089, new_n12027);
nand_4 g09742(new_n12091, new_n12090, new_n12026);
nand_4 g09743(new_n12092, new_n12091, new_n12021);
nand_4 g09744(new_n12093, new_n12092, new_n12019);
xnor_3 g09745(n1302, new_n12093, new_n12016);
nor_4  g09746(new_n12095, n13951, new_n10423);
xor_3  g09747(new_n12096, n13951, new_n10423);
not_3  g09748(new_n12097, new_n12096);
nor_4  g09749(new_n12098, n22793, new_n10438);
xor_3  g09750(new_n12099, n22793, new_n10438);
nand_4 g09751(new_n12100, new_n2758, n3710);
xor_3  g09752(new_n12101, n8439, new_n10445);
nor_4  g09753(new_n12102, new_n10454, n25523);
not_3  g09754(new_n12103, new_n12102);
not_3  g09755(new_n12104, n25523);
xor_3  g09756(new_n12105, n26318, new_n12104);
not_3  g09757(new_n12106, n26054);
nor_4  g09758(new_n12107, new_n12106, n5579);
not_3  g09759(new_n12108, new_n12107);
xor_3  g09760(new_n12109, n26054, new_n2759);
nor_4  g09761(new_n12110, n23430, new_n10462);
xor_3  g09762(new_n12111, n23430, new_n10462);
not_3  g09763(new_n12112, new_n12111);
nor_4  g09764(new_n12113_1, n10411, new_n10490);
xor_3  g09765(new_n12114, n10411, n8309);
nor_4  g09766(new_n12115, n19144, new_n2760);
nor_4  g09767(new_n12116, new_n10474, n16971);
not_3  g09768(new_n12117, n11503);
nor_4  g09769(new_n12118, n12593, new_n12117);
nor_4  g09770(new_n12119, new_n10483, n11503);
nor_4  g09771(new_n12120, new_n2882, n13714);
not_3  g09772(new_n12121_1, new_n12120);
nor_4  g09773(new_n12122, new_n12121_1, new_n12119);
nor_4  g09774(new_n12123, new_n12122, new_n12118);
nor_4  g09775(new_n12124, new_n12123, new_n12116);
nor_4  g09776(new_n12125, new_n12124, new_n12115);
not_3  g09777(new_n12126, new_n12125);
nor_4  g09778(new_n12127, new_n12126, new_n12114);
nor_4  g09779(new_n12128, new_n12127, new_n12113_1);
nor_4  g09780(new_n12129, new_n12128, new_n12112);
nor_4  g09781(new_n12130, new_n12129, new_n12110);
not_3  g09782(new_n12131_1, new_n12130);
nand_4 g09783(new_n12132, new_n12131_1, new_n12109);
nand_4 g09784(new_n12133, new_n12132, new_n12108);
nand_4 g09785(new_n12134, new_n12133, new_n12105);
nand_4 g09786(new_n12135, new_n12134, new_n12103);
nand_4 g09787(new_n12136, new_n12135, new_n12101);
nand_4 g09788(new_n12137, new_n12136, new_n12100);
nand_4 g09789(new_n12138, new_n12137, new_n12099);
not_3  g09790(new_n12139, new_n12138);
nor_4  g09791(new_n12140, new_n12139, new_n12098);
nor_4  g09792(new_n12141, new_n12140, new_n12097);
nor_4  g09793(new_n12142, new_n12141, new_n12095);
nor_4  g09794(new_n12143, n12650, n11220);
xor_3  g09795(new_n12144, n12650, n11220);
not_3  g09796(new_n12145, new_n12144);
nor_4  g09797(new_n12146_1, n22379, n10201);
xor_3  g09798(new_n12147, n22379, n10201);
not_3  g09799(new_n12148, new_n12147);
nor_4  g09800(new_n12149, n10593, n1662);
xor_3  g09801(new_n12150, n10593, n1662);
not_3  g09802(new_n12151, new_n12150);
nand_4 g09803(new_n12152_1, new_n10738, new_n2989);
nand_4 g09804(new_n12153_1, new_n11111, new_n11086);
nand_4 g09805(new_n12154, new_n12153_1, new_n12152_1);
not_3  g09806(new_n12155, new_n12154);
nor_4  g09807(new_n12156, new_n12155, new_n12151);
nor_4  g09808(new_n12157_1, new_n12156, new_n12149);
nor_4  g09809(new_n12158_1, new_n12157_1, new_n12148);
nor_4  g09810(new_n12159, new_n12158_1, new_n12146_1);
nor_4  g09811(new_n12160, new_n12159, new_n12145);
nor_4  g09812(new_n12161_1, new_n12160, new_n12143);
nor_4  g09813(new_n12162, n22270, n2944);
nor_4  g09814(new_n12163, new_n2818, new_n2773);
nor_4  g09815(new_n12164, new_n12163, new_n12162);
xor_3  g09816(new_n12165, new_n12164, new_n12161_1);
xor_3  g09817(new_n12166, new_n12159, new_n12145);
nor_4  g09818(new_n12167, new_n12166, new_n2819);
not_3  g09819(new_n12168, new_n12167);
not_3  g09820(new_n12169, new_n2826_1);
xor_3  g09821(new_n12170, new_n12157_1, new_n12148);
nand_4 g09822(new_n12171, new_n12170, new_n12169);
xor_3  g09823(new_n12172, new_n12157_1, new_n12147);
nor_4  g09824(new_n12173, new_n12172, new_n2826_1);
nor_4  g09825(new_n12174, new_n12170, new_n12169);
nor_4  g09826(new_n12175, new_n12174, new_n12173);
xor_3  g09827(new_n12176, new_n12155, new_n12150);
nor_4  g09828(new_n12177, new_n12176, new_n2832);
not_3  g09829(new_n12178, new_n12177);
xor_3  g09830(new_n12179_1, new_n12155, new_n12151);
nor_4  g09831(new_n12180, new_n12179_1, new_n2831);
nor_4  g09832(new_n12181, new_n12180, new_n12177);
nor_4  g09833(new_n12182, new_n11112, new_n2838);
not_3  g09834(new_n12183, new_n12182);
nor_4  g09835(new_n12184, new_n11117, new_n2847);
not_3  g09836(new_n12185, new_n12184);
nor_4  g09837(new_n12186, new_n11115, new_n2851);
nor_4  g09838(new_n12187, new_n12186, new_n12184);
nor_4  g09839(new_n12188, new_n11130, new_n2895);
nand_4 g09840(new_n12189, new_n11136, new_n2862);
not_3  g09841(new_n12190, new_n12189);
nor_4  g09842(new_n12191, new_n11136, new_n2862);
nor_4  g09843(new_n12192_1, new_n12191, new_n12190);
nand_4 g09844(new_n12193, new_n11142, new_n2873);
not_3  g09845(new_n12194, new_n12193);
xnor_3 g09846(new_n12195, new_n11142, new_n2873);
nor_4  g09847(new_n12196, new_n11153, new_n2879);
xor_3  g09848(new_n12197, n25023, new_n3013);
not_3  g09849(new_n12198, new_n11150);
nor_4  g09850(new_n12199, new_n12198, new_n12197);
nor_4  g09851(new_n12200, new_n11147, new_n2886_1);
nor_4  g09852(new_n12201, new_n12200, new_n12196);
nand_4 g09853(new_n12202, new_n12201, new_n12199);
not_3  g09854(new_n12203, new_n12202);
nor_4  g09855(new_n12204, new_n12203, new_n12196);
nor_4  g09856(new_n12205, new_n12204, new_n12195);
nor_4  g09857(new_n12206, new_n12205, new_n12194);
not_3  g09858(new_n12207, new_n12206);
nand_4 g09859(new_n12208, new_n12207, new_n12192_1);
nand_4 g09860(new_n12209_1, new_n12208, new_n12189);
nor_4  g09861(new_n12210, new_n11131, new_n2857);
nor_4  g09862(new_n12211, new_n12210, new_n12188);
not_3  g09863(new_n12212, new_n12211);
nor_4  g09864(new_n12213, new_n12212, new_n12209_1);
nor_4  g09865(new_n12214, new_n12213, new_n12188);
nand_4 g09866(new_n12215, new_n12214, new_n12187);
nand_4 g09867(new_n12216, new_n12215, new_n12185);
not_3  g09868(new_n12217, new_n11086);
xnor_3 g09869(new_n12218, new_n11111, new_n12217);
nor_4  g09870(new_n12219, new_n12218, new_n2842);
nor_4  g09871(new_n12220, new_n12219, new_n12182);
nand_4 g09872(new_n12221, new_n12220, new_n12216);
nand_4 g09873(new_n12222, new_n12221, new_n12183);
nand_4 g09874(new_n12223_1, new_n12222, new_n12181);
nand_4 g09875(new_n12224, new_n12223_1, new_n12178);
nand_4 g09876(new_n12225_1, new_n12224, new_n12175);
nand_4 g09877(new_n12226, new_n12225_1, new_n12171);
not_3  g09878(new_n12227, new_n12226);
xor_3  g09879(new_n12228_1, new_n12159, new_n12144);
nor_4  g09880(new_n12229, new_n12228_1, new_n2821);
nor_4  g09881(new_n12230, new_n12229, new_n12167);
nand_4 g09882(new_n12231, new_n12230, new_n12227);
nand_4 g09883(new_n12232, new_n12231, new_n12168);
xnor_3 g09884(new_n12233, new_n12232, new_n12165);
xnor_3 g09885(new_n12234, new_n12233, new_n12142);
xor_3  g09886(new_n12235_1, new_n12140, new_n12097);
xnor_3 g09887(new_n12236, new_n12230, new_n12226);
nor_4  g09888(new_n12237, new_n12236, new_n12235_1);
xnor_3 g09889(new_n12238, new_n12236, new_n12235_1);
xor_3  g09890(new_n12239, new_n12137, new_n12099);
xnor_3 g09891(new_n12240, new_n12224, new_n12175);
nor_4  g09892(new_n12241, new_n12240, new_n12239);
not_3  g09893(new_n12242, new_n12239);
xnor_3 g09894(new_n12243, new_n12240, new_n12242);
xnor_3 g09895(new_n12244, new_n12135, new_n12101);
xnor_3 g09896(new_n12245, new_n12222, new_n12181);
not_3  g09897(new_n12246, new_n12245);
nand_4 g09898(new_n12247, new_n12246, new_n12244);
xnor_3 g09899(new_n12248, new_n12245, new_n12244);
not_3  g09900(new_n12249, new_n12105);
xor_3  g09901(new_n12250, new_n12133, new_n12249);
xnor_3 g09902(new_n12251, new_n12220, new_n12216);
not_3  g09903(new_n12252, new_n12251);
nand_4 g09904(new_n12253, new_n12252, new_n12250);
xnor_3 g09905(new_n12254, new_n12251, new_n12250);
xor_3  g09906(new_n12255, new_n12131_1, new_n12109);
not_3  g09907(new_n12256, new_n12255);
not_3  g09908(new_n12257, new_n12214);
xnor_3 g09909(new_n12258, new_n12257, new_n12187);
nand_4 g09910(new_n12259, new_n12258, new_n12256);
xor_3  g09911(new_n12260, new_n12128, new_n12112);
not_3  g09912(new_n12261, new_n12260);
xnor_3 g09913(new_n12262, new_n12212, new_n12209_1);
nand_4 g09914(new_n12263, new_n12262, new_n12261);
xnor_3 g09915(new_n12264, new_n12262, new_n12260);
xnor_3 g09916(new_n12265, new_n12206, new_n12192_1);
xor_3  g09917(new_n12266, new_n12126, new_n12114);
not_3  g09918(new_n12267, new_n12266);
nand_4 g09919(new_n12268, new_n12267, new_n12265);
xnor_3 g09920(new_n12269, new_n12204, new_n12195);
not_3  g09921(new_n12270, new_n12123);
nor_4  g09922(new_n12271, new_n12116, new_n12115);
xor_3  g09923(new_n12272, new_n12271, new_n12270);
not_3  g09924(new_n12273, new_n12272);
nor_4  g09925(new_n12274, new_n12273, new_n12269);
not_3  g09926(new_n12275, new_n12274);
not_3  g09927(new_n12276, new_n12269);
nor_4  g09928(new_n12277, new_n12272, new_n12276);
nor_4  g09929(new_n12278, new_n12277, new_n12274);
nor_4  g09930(new_n12279, new_n11150, new_n2883);
nor_4  g09931(new_n12280, new_n12279, new_n12199);
not_3  g09932(new_n12281, n13714);
xor_3  g09933(new_n12282, n18151, new_n12281);
nor_4  g09934(new_n12283, new_n12282, new_n12280);
not_3  g09935(new_n12284, new_n12283);
nor_4  g09936(new_n12285, new_n12119, new_n12118);
xor_3  g09937(new_n12286, new_n12285, new_n12120);
nor_4  g09938(new_n12287, new_n12286, new_n12284);
nor_4  g09939(new_n12288, new_n12201, new_n12199);
nor_4  g09940(new_n12289, new_n12288, new_n12203);
not_3  g09941(new_n12290, new_n12286);
xor_3  g09942(new_n12291, new_n12290, new_n12284);
nor_4  g09943(new_n12292, new_n12291, new_n12289);
nor_4  g09944(new_n12293, new_n12292, new_n12287);
nand_4 g09945(new_n12294, new_n12293, new_n12278);
nand_4 g09946(new_n12295, new_n12294, new_n12275);
not_3  g09947(new_n12296, new_n12268);
nor_4  g09948(new_n12297, new_n12267, new_n12265);
nor_4  g09949(new_n12298, new_n12297, new_n12296);
nand_4 g09950(new_n12299, new_n12298, new_n12295);
nand_4 g09951(new_n12300, new_n12299, new_n12268);
nand_4 g09952(new_n12301, new_n12300, new_n12264);
nand_4 g09953(new_n12302_1, new_n12301, new_n12263);
xnor_3 g09954(new_n12303, new_n12258, new_n12255);
nand_4 g09955(new_n12304_1, new_n12303, new_n12302_1);
nand_4 g09956(new_n12305, new_n12304_1, new_n12259);
nand_4 g09957(new_n12306, new_n12305, new_n12254);
nand_4 g09958(new_n12307, new_n12306, new_n12253);
nand_4 g09959(new_n12308, new_n12307, new_n12248);
nand_4 g09960(new_n12309, new_n12308, new_n12247);
nand_4 g09961(new_n12310, new_n12309, new_n12243);
not_3  g09962(new_n12311, new_n12310);
nor_4  g09963(new_n12312, new_n12311, new_n12241);
nor_4  g09964(new_n12313, new_n12312, new_n12238);
nor_4  g09965(new_n12314, new_n12313, new_n12237);
xnor_3 g09966(n1332, new_n12314, new_n12234);
nor_4  g09967(new_n12316, new_n6432, n14692);
not_3  g09968(new_n12317, new_n12316);
xnor_3 g09969(new_n12318, new_n6432, n14692);
not_3  g09970(new_n12319, new_n12318);
not_3  g09971(new_n12320, n4100);
nand_4 g09972(new_n12321, new_n6519, new_n12320);
not_3  g09973(new_n12322, new_n12321);
nor_4  g09974(new_n12323, new_n6519, new_n12320);
nor_4  g09975(new_n12324_1, new_n12323, new_n12322);
nor_4  g09976(new_n12325_1, new_n6529, n21957);
not_3  g09977(new_n12326, new_n12325_1);
xnor_3 g09978(new_n12327, new_n6524, n21957);
not_3  g09979(new_n12328, n15761);
nand_4 g09980(new_n12329_1, new_n6531, new_n12328);
xnor_3 g09981(new_n12330_1, new_n6531, n15761);
nor_4  g09982(new_n12331, new_n6544, n11201);
not_3  g09983(new_n12332, new_n12331);
not_3  g09984(new_n12333, n11201);
nor_4  g09985(new_n12334, new_n6537, new_n12333);
nor_4  g09986(new_n12335, new_n12334, new_n12331);
nor_4  g09987(new_n12336, new_n6547, n18690);
not_3  g09988(new_n12337, new_n12336);
not_3  g09989(new_n12338, n18690);
nor_4  g09990(new_n12339, new_n6546, new_n12338);
nor_4  g09991(new_n12340, new_n12339, new_n12336);
not_3  g09992(new_n12341_1, new_n6555);
nor_4  g09993(new_n12342, new_n12341_1, n12153);
not_3  g09994(new_n12343, new_n12342);
not_3  g09995(new_n12344, n12153);
nor_4  g09996(new_n12345, new_n6555, new_n12344);
nor_4  g09997(new_n12346_1, new_n12345, new_n12342);
not_3  g09998(new_n12347, n13044);
nor_4  g09999(new_n12348, new_n6566, new_n12347);
nor_4  g10000(new_n12349_1, new_n6565, n13044);
nor_4  g10001(new_n12350, new_n6790_1, new_n6785_1);
not_3  g10002(new_n12351, new_n12350);
nor_4  g10003(new_n12352, new_n12351, new_n12349_1);
nor_4  g10004(new_n12353, new_n12352, new_n12348);
nand_4 g10005(new_n12354, new_n12353, new_n12346_1);
nand_4 g10006(new_n12355, new_n12354, new_n12343);
nand_4 g10007(new_n12356, new_n12355, new_n12340);
nand_4 g10008(new_n12357, new_n12356, new_n12337);
nand_4 g10009(new_n12358, new_n12357, new_n12335);
nand_4 g10010(new_n12359, new_n12358, new_n12332);
nand_4 g10011(new_n12360, new_n12359, new_n12330_1);
nand_4 g10012(new_n12361, new_n12360, new_n12329_1);
nand_4 g10013(new_n12362, new_n12361, new_n12327);
nand_4 g10014(new_n12363, new_n12362, new_n12326);
nand_4 g10015(new_n12364_1, new_n12363, new_n12324_1);
nand_4 g10016(new_n12365, new_n12364_1, new_n12321);
nand_4 g10017(new_n12366, new_n12365, new_n12319);
nand_4 g10018(new_n12367, new_n12366, new_n12317);
nor_4  g10019(new_n12368, new_n12367, new_n6431_1);
not_3  g10020(new_n12369, new_n12368);
nor_4  g10021(new_n12370, new_n6807, n11302);
not_3  g10022(new_n12371, new_n12370);
nor_4  g10023(new_n12372, new_n12371, n10405);
not_3  g10024(new_n12373, new_n12372);
nor_4  g10025(new_n12374, new_n12373, n7693);
not_3  g10026(new_n12375, new_n12374);
nor_4  g10027(new_n12376, new_n12375, n20151);
not_3  g10028(new_n12377, new_n12376);
nor_4  g10029(new_n12378, new_n12377, n8964);
not_3  g10030(new_n12379, new_n12378);
nor_4  g10031(new_n12380_1, new_n12379, n27037);
not_3  g10032(new_n12381, new_n12380_1);
nor_4  g10033(new_n12382, new_n12381, n15182);
not_3  g10034(new_n12383_1, new_n12382);
nor_4  g10035(new_n12384_1, new_n12383_1, n8614);
not_3  g10036(new_n12385, n23039);
not_3  g10037(new_n12386, n18926);
nor_4  g10038(new_n12387, n25926, n7657);
nand_4 g10039(new_n12388, new_n12387, new_n4401_1);
nor_4  g10040(new_n12389, new_n12388, n5451);
nand_4 g10041(new_n12390, new_n12389, new_n12386);
nor_4  g10042(new_n12391, new_n12390, n13677);
nand_4 g10043(new_n12392, new_n12391, new_n12385);
nor_4  g10044(new_n12393, new_n12392, n7692);
not_3  g10045(new_n12394, new_n12393);
nor_4  g10046(new_n12395, new_n12394, n25629);
not_3  g10047(new_n12396, new_n12395);
nor_4  g10048(new_n12397_1, new_n12396, n15766);
not_3  g10049(new_n12398_1, new_n12397_1);
xor_3  g10050(new_n12399, new_n12395, n15766);
nand_4 g10051(new_n12400, new_n12399, new_n6319);
xor_3  g10052(new_n12401, new_n12394, n25629);
not_3  g10053(new_n12402, new_n12401);
nand_4 g10054(new_n12403, new_n12402, new_n6324);
xnor_3 g10055(new_n12404, new_n12401, new_n6324);
not_3  g10056(new_n12405, new_n12392);
xor_3  g10057(new_n12406, new_n12405, n7692);
nand_4 g10058(new_n12407, new_n12406, new_n6330_1);
xor_3  g10059(new_n12408_1, new_n12392, n7692);
xnor_3 g10060(new_n12409, new_n12408_1, new_n6330_1);
nor_4  g10061(new_n12410, new_n12391, new_n12385);
nor_4  g10062(new_n12411, new_n12410, new_n12405);
nor_4  g10063(new_n12412, new_n12411, n23200);
not_3  g10064(new_n12413, new_n12412);
xor_3  g10065(new_n12414, new_n12411, n23200);
nand_4 g10066(new_n12415, new_n12390, n13677);
not_3  g10067(new_n12416, new_n12415);
nor_4  g10068(new_n12417, new_n12416, new_n12391);
nor_4  g10069(new_n12418, new_n12417, n17959);
not_3  g10070(new_n12419, new_n12418);
not_3  g10071(new_n12420, new_n12390);
nor_4  g10072(new_n12421, new_n12389, new_n12386);
nor_4  g10073(new_n12422, new_n12421, new_n12420);
nor_4  g10074(new_n12423, new_n12422, n7566);
not_3  g10075(new_n12424, new_n12423);
not_3  g10076(new_n12425, new_n12422);
nor_4  g10077(new_n12426, new_n12425, new_n6339_1);
nor_4  g10078(new_n12427, new_n12426, new_n12423);
nand_4 g10079(new_n12428, new_n12388, n5451);
not_3  g10080(new_n12429, new_n12428);
nor_4  g10081(new_n12430, new_n12429, new_n12389);
not_3  g10082(new_n12431, new_n12430);
nor_4  g10083(new_n12432, new_n12431, new_n6343);
nor_4  g10084(new_n12433, new_n12430, n7731);
xnor_3 g10085(new_n12434, new_n12387, new_n4401_1);
nor_4  g10086(new_n12435, new_n12434, new_n6348);
xnor_3 g10087(new_n12436, new_n12434, new_n6348);
nor_4  g10088(new_n12437, new_n6797, new_n6351);
nor_4  g10089(new_n12438, new_n6801, new_n12437);
nor_4  g10090(new_n12439, new_n12438, new_n12436);
nor_4  g10091(new_n12440, new_n12439, new_n12435);
nor_4  g10092(new_n12441, new_n12440, new_n12433);
nor_4  g10093(new_n12442, new_n12441, new_n12432);
nand_4 g10094(new_n12443, new_n12442, new_n12427);
nand_4 g10095(new_n12444, new_n12443, new_n12424);
xor_3  g10096(new_n12445, new_n12417, n17959);
nand_4 g10097(new_n12446_1, new_n12445, new_n12444);
nand_4 g10098(new_n12447, new_n12446_1, new_n12419);
nand_4 g10099(new_n12448, new_n12447, new_n12414);
nand_4 g10100(new_n12449_1, new_n12448, new_n12413);
nand_4 g10101(new_n12450, new_n12449_1, new_n12409);
nand_4 g10102(new_n12451, new_n12450, new_n12407);
nand_4 g10103(new_n12452, new_n12451, new_n12404);
nand_4 g10104(new_n12453, new_n12452, new_n12403);
not_3  g10105(new_n12454, new_n12399);
nand_4 g10106(new_n12455, new_n12454, n23895);
nand_4 g10107(new_n12456, new_n12455, new_n12453);
nand_4 g10108(new_n12457, new_n12456, new_n12400);
nand_4 g10109(new_n12458, new_n12457, new_n12398_1);
not_3  g10110(new_n12459, new_n12458);
nor_4  g10111(new_n12460, new_n12459, new_n12384_1);
not_3  g10112(new_n12461_1, new_n12460);
xor_3  g10113(new_n12462_1, new_n12382, new_n6321);
nand_4 g10114(new_n12463, new_n12455, new_n12400);
not_3  g10115(new_n12464, new_n12463);
xnor_3 g10116(new_n12465, new_n12464, new_n12453);
nand_4 g10117(new_n12466, new_n12465, new_n12462_1);
xor_3  g10118(new_n12467_1, new_n12380_1, new_n6326);
not_3  g10119(new_n12468, new_n12467_1);
not_3  g10120(new_n12469_1, new_n12404);
xnor_3 g10121(new_n12470, new_n12451, new_n12469_1);
nand_4 g10122(new_n12471, new_n12470, new_n12468);
xnor_3 g10123(new_n12472, new_n12470, new_n12467_1);
xor_3  g10124(new_n12473, new_n12378, new_n6328);
not_3  g10125(new_n12474, new_n12473);
not_3  g10126(new_n12475, new_n12449_1);
xnor_3 g10127(new_n12476, new_n12475, new_n12409);
nand_4 g10128(new_n12477, new_n12476, new_n12474);
xnor_3 g10129(new_n12478, new_n12476, new_n12473);
xor_3  g10130(new_n12479, new_n12376, new_n6332);
not_3  g10131(new_n12480, new_n12414);
not_3  g10132(new_n12481, new_n12444);
xor_3  g10133(new_n12482, new_n12417, new_n6335);
nor_4  g10134(new_n12483, new_n12482, new_n12481);
nor_4  g10135(new_n12484, new_n12483, new_n12418);
nor_4  g10136(new_n12485, new_n12484, new_n12480);
nor_4  g10137(new_n12486, new_n12447, new_n12414);
nor_4  g10138(new_n12487, new_n12486, new_n12485);
not_3  g10139(new_n12488, new_n12487);
nor_4  g10140(new_n12489, new_n12488, new_n12479);
not_3  g10141(new_n12490, new_n12489);
not_3  g10142(new_n12491, new_n12479);
xnor_3 g10143(new_n12492, new_n12487, new_n12491);
not_3  g10144(new_n12493, new_n12492);
xor_3  g10145(new_n12494, new_n12374, new_n7279);
nor_4  g10146(new_n12495_1, new_n12445, new_n12444);
nor_4  g10147(new_n12496, new_n12495_1, new_n12483);
not_3  g10148(new_n12497, new_n12496);
nor_4  g10149(new_n12498, new_n12497, new_n12494);
not_3  g10150(new_n12499, new_n12498);
not_3  g10151(new_n12500, new_n12494);
xnor_3 g10152(new_n12501, new_n12496, new_n12500);
not_3  g10153(new_n12502, new_n12501);
xor_3  g10154(new_n12503, new_n12372, new_n4447);
not_3  g10155(new_n12504, new_n12443);
not_3  g10156(new_n12505, new_n12427);
not_3  g10157(new_n12506, new_n12442);
nand_4 g10158(new_n12507_1, new_n12506, new_n12505);
not_3  g10159(new_n12508, new_n12507_1);
nor_4  g10160(new_n12509, new_n12508, new_n12504);
not_3  g10161(new_n12510, new_n12509);
nor_4  g10162(new_n12511, new_n12510, new_n12503);
not_3  g10163(new_n12512, new_n12511);
not_3  g10164(new_n12513, new_n12503);
nor_4  g10165(new_n12514, new_n12509, new_n12513);
nor_4  g10166(new_n12515_1, new_n12514, new_n12511);
xor_3  g10167(new_n12516_1, new_n12370, new_n4451_1);
not_3  g10168(new_n12517, new_n12440);
nor_4  g10169(new_n12518, new_n12433, new_n12432);
xnor_3 g10170(new_n12519, new_n12518, new_n12517);
not_3  g10171(new_n12520, new_n12519);
nor_4  g10172(new_n12521, new_n12520, new_n12516_1);
not_3  g10173(new_n12522, new_n12521);
not_3  g10174(new_n12523, new_n12516_1);
nor_4  g10175(new_n12524, new_n12519, new_n12523);
nor_4  g10176(new_n12525, new_n12524, new_n12521);
xnor_3 g10177(new_n12526, new_n12438, new_n12436);
xor_3  g10178(new_n12527, new_n6806, new_n6346);
not_3  g10179(new_n12528, new_n12527);
nand_4 g10180(new_n12529, new_n12528, new_n12526);
xnor_3 g10181(new_n12530, new_n12527, new_n12526);
nor_4  g10182(new_n12531, new_n6813, new_n6802_1);
nor_4  g10183(new_n12532, new_n12531, new_n6811);
not_3  g10184(new_n12533, new_n12532);
nand_4 g10185(new_n12534, new_n12533, new_n12530);
nand_4 g10186(new_n12535, new_n12534, new_n12529);
nand_4 g10187(new_n12536, new_n12535, new_n12525);
nand_4 g10188(new_n12537, new_n12536, new_n12522);
nand_4 g10189(new_n12538, new_n12537, new_n12515_1);
nand_4 g10190(new_n12539, new_n12538, new_n12512);
nand_4 g10191(new_n12540_1, new_n12539, new_n12502);
nand_4 g10192(new_n12541, new_n12540_1, new_n12499);
nand_4 g10193(new_n12542, new_n12541, new_n12493);
nand_4 g10194(new_n12543, new_n12542, new_n12490);
nand_4 g10195(new_n12544, new_n12543, new_n12478);
nand_4 g10196(new_n12545_1, new_n12544, new_n12477);
nand_4 g10197(new_n12546_1, new_n12545_1, new_n12472);
nand_4 g10198(new_n12547, new_n12546_1, new_n12471);
not_3  g10199(new_n12548, new_n12547);
not_3  g10200(new_n12549, new_n12466);
nor_4  g10201(new_n12550, new_n12465, new_n12462_1);
nor_4  g10202(new_n12551, new_n12550, new_n12549);
nand_4 g10203(new_n12552_1, new_n12551, new_n12548);
nand_4 g10204(new_n12553, new_n12552_1, new_n12466);
nor_4  g10205(new_n12554, new_n12553, new_n12461_1);
nor_4  g10206(new_n12555, new_n12554, new_n12369);
not_3  g10207(new_n12556, new_n12554);
nor_4  g10208(new_n12557, new_n12556, new_n12368);
nor_4  g10209(new_n12558, new_n12557, new_n12555);
xnor_3 g10210(new_n12559, new_n12367, new_n6430);
xor_3  g10211(new_n12560, new_n12459, new_n12384_1);
xnor_3 g10212(new_n12561, new_n12560, new_n12553);
nor_4  g10213(new_n12562_1, new_n12561, new_n12559);
xnor_3 g10214(new_n12563, new_n12561, new_n12559);
xnor_3 g10215(new_n12564, new_n12365, new_n12318);
xnor_3 g10216(new_n12565, new_n12551, new_n12547);
not_3  g10217(new_n12566_1, new_n12565);
nor_4  g10218(new_n12567, new_n12566_1, new_n12564);
not_3  g10219(new_n12568, new_n12567);
xnor_3 g10220(new_n12569_1, new_n12365, new_n12319);
nor_4  g10221(new_n12570, new_n12565, new_n12569_1);
nor_4  g10222(new_n12571, new_n12570, new_n12567);
xnor_3 g10223(new_n12572, new_n12545_1, new_n12472);
not_3  g10224(new_n12573, new_n12572);
not_3  g10225(new_n12574, new_n12362);
nor_4  g10226(new_n12575, new_n12574, new_n12325_1);
xnor_3 g10227(new_n12576, new_n12575, new_n12324_1);
nor_4  g10228(new_n12577, new_n12576, new_n12573);
xnor_3 g10229(new_n12578, new_n12543, new_n12478);
xnor_3 g10230(new_n12579, new_n12361, new_n12327);
nor_4  g10231(new_n12580, new_n12579, new_n12578);
not_3  g10232(new_n12581, new_n12580);
xnor_3 g10233(new_n12582, new_n12579, new_n12578);
not_3  g10234(new_n12583, new_n12582);
xnor_3 g10235(new_n12584, new_n12541, new_n12492);
xnor_3 g10236(new_n12585, new_n6531, new_n12328);
xnor_3 g10237(new_n12586, new_n12359, new_n12585);
nor_4  g10238(new_n12587_1, new_n12586, new_n12584);
xnor_3 g10239(new_n12588, new_n12539, new_n12501);
xnor_3 g10240(new_n12589, new_n6537, new_n12333);
xnor_3 g10241(new_n12590, new_n12357, new_n12589);
nand_4 g10242(new_n12591, new_n12590, new_n12588);
xnor_3 g10243(new_n12592, new_n12590, new_n12588);
not_3  g10244(new_n12593_1, new_n12592);
xnor_3 g10245(new_n12594, new_n12537, new_n12515_1);
not_3  g10246(new_n12595, new_n12594);
xnor_3 g10247(new_n12596, new_n12355, new_n12340);
not_3  g10248(new_n12597, new_n12596);
nor_4  g10249(new_n12598, new_n12597, new_n12595);
xnor_3 g10250(new_n12599, new_n12596, new_n12594);
xnor_3 g10251(new_n12600, new_n12535, new_n12525);
xnor_3 g10252(new_n12601, new_n12353, new_n12346_1);
nor_4  g10253(new_n12602, new_n12601, new_n12600);
not_3  g10254(new_n12603, new_n12602);
not_3  g10255(new_n12604, new_n12600);
not_3  g10256(new_n12605, new_n12601);
nor_4  g10257(new_n12606, new_n12605, new_n12604);
nor_4  g10258(new_n12607_1, new_n12606, new_n12602);
xnor_3 g10259(new_n12608, new_n12533, new_n12530);
nor_4  g10260(new_n12609, new_n12349_1, new_n12348);
xnor_3 g10261(new_n12610, new_n12609, new_n12350);
not_3  g10262(new_n12611, new_n12610);
nor_4  g10263(new_n12612, new_n12611, new_n12608);
nor_4  g10264(new_n12613, new_n6814_1, new_n6794_1);
nor_4  g10265(new_n12614, new_n6815, new_n6783);
nor_4  g10266(new_n12615, new_n12614, new_n12613);
not_3  g10267(new_n12616, new_n12608);
nor_4  g10268(new_n12617, new_n12610, new_n12616);
nor_4  g10269(new_n12618, new_n12617, new_n12612);
not_3  g10270(new_n12619, new_n12618);
nor_4  g10271(new_n12620_1, new_n12619, new_n12615);
nor_4  g10272(new_n12621_1, new_n12620_1, new_n12612);
not_3  g10273(new_n12622, new_n12621_1);
nand_4 g10274(new_n12623, new_n12622, new_n12607_1);
nand_4 g10275(new_n12624, new_n12623, new_n12603);
nor_4  g10276(new_n12625, new_n12624, new_n12599);
nor_4  g10277(new_n12626_1, new_n12625, new_n12598);
nand_4 g10278(new_n12627, new_n12626_1, new_n12593_1);
nand_4 g10279(new_n12628, new_n12627, new_n12591);
xnor_3 g10280(new_n12629, new_n12586, new_n12584);
nor_4  g10281(new_n12630, new_n12629, new_n12628);
nor_4  g10282(new_n12631, new_n12630, new_n12587_1);
nand_4 g10283(new_n12632, new_n12631, new_n12583);
nand_4 g10284(new_n12633, new_n12632, new_n12581);
xnor_3 g10285(new_n12634, new_n12363, new_n12324_1);
xnor_3 g10286(new_n12635, new_n12634, new_n12572);
nor_4  g10287(new_n12636, new_n12635, new_n12633);
nor_4  g10288(new_n12637, new_n12636, new_n12577);
not_3  g10289(new_n12638, new_n12637);
nand_4 g10290(new_n12639, new_n12638, new_n12571);
nand_4 g10291(new_n12640, new_n12639, new_n12568);
nor_4  g10292(new_n12641, new_n12640, new_n12563);
nor_4  g10293(new_n12642, new_n12641, new_n12562_1);
xnor_3 g10294(n1357, new_n12642, new_n12558);
xor_3  g10295(new_n12644, new_n9455, new_n8503);
nor_4  g10296(new_n12645, new_n9461, n10125);
not_3  g10297(new_n12646, new_n12645);
xor_3  g10298(new_n12647, new_n9463, new_n8506);
nor_4  g10299(new_n12648, new_n9468, n8067);
not_3  g10300(new_n12649, new_n12648);
xor_3  g10301(new_n12650_1, new_n9470, new_n8509);
nor_4  g10302(new_n12651, new_n9475, n20923);
not_3  g10303(new_n12652, new_n12651);
not_3  g10304(new_n12653, n20923);
xor_3  g10305(new_n12654_1, new_n9477, new_n12653);
nor_4  g10306(new_n12655, new_n9481, n18157);
not_3  g10307(new_n12656, new_n12655);
nand_4 g10308(new_n12657_1, new_n10060, new_n10051);
nand_4 g10309(new_n12658, new_n12657_1, new_n10049);
nand_4 g10310(new_n12659, new_n12658, new_n12656);
nand_4 g10311(new_n12660, new_n12659, new_n12654_1);
nand_4 g10312(new_n12661, new_n12660, new_n12652);
nand_4 g10313(new_n12662, new_n12661, new_n12650_1);
nand_4 g10314(new_n12663, new_n12662, new_n12649);
nand_4 g10315(new_n12664, new_n12663, new_n12647);
nand_4 g10316(new_n12665_1, new_n12664, new_n12646);
xnor_3 g10317(new_n12666, new_n12665_1, new_n12644);
not_3  g10318(new_n12667, new_n12666);
not_3  g10319(new_n12668, n5077);
xor_3  g10320(new_n12669, n6381, n1099);
nor_4  g10321(new_n12670_1, n14345, n2113);
not_3  g10322(new_n12671, new_n12670_1);
xor_3  g10323(new_n12672, n14345, n2113);
nor_4  g10324(new_n12673, n21134, n11356);
not_3  g10325(new_n12674, new_n12673);
xor_3  g10326(new_n12675, n21134, n11356);
nand_4 g10327(new_n12676, n6369, n3164);
not_3  g10328(new_n12677, new_n12676);
nor_4  g10329(new_n12678, n6369, n3164);
nor_4  g10330(new_n12679, n25797, n10611);
not_3  g10331(new_n12680, new_n12679);
nand_4 g10332(new_n12681, new_n7747, new_n12680);
nor_4  g10333(new_n12682, new_n12681, new_n12678);
nor_4  g10334(new_n12683, new_n12682, new_n12677);
nand_4 g10335(new_n12684, new_n12683, new_n12675);
nand_4 g10336(new_n12685, new_n12684, new_n12674);
nand_4 g10337(new_n12686, new_n12685, new_n12672);
nand_4 g10338(new_n12687, new_n12686, new_n12671);
xnor_3 g10339(new_n12688, new_n12687, new_n12669);
xnor_3 g10340(new_n12689, new_n12688, new_n12668);
xnor_3 g10341(new_n12690, new_n12685, new_n12672);
nand_4 g10342(new_n12691, new_n12690, n15546);
not_3  g10343(new_n12692, n15546);
xnor_3 g10344(new_n12693, new_n12690, new_n12692);
xnor_3 g10345(new_n12694, new_n12683, new_n12675);
nor_4  g10346(new_n12695, new_n12694, n26452);
nor_4  g10347(new_n12696, new_n12678, new_n12677);
xnor_3 g10348(new_n12697, new_n12696, new_n12681);
nand_4 g10349(new_n12698, new_n12697, n19905);
xnor_3 g10350(new_n12699, new_n12697, new_n4668);
not_3  g10351(new_n12700, new_n10094);
nand_4 g10352(new_n12701, new_n10101_1, new_n12700);
nand_4 g10353(new_n12702_1, new_n12701, new_n12699);
nand_4 g10354(new_n12703, new_n12702_1, new_n12698);
xnor_3 g10355(new_n12704, new_n12694, n26452);
nor_4  g10356(new_n12705, new_n12704, new_n12703);
nor_4  g10357(new_n12706, new_n12705, new_n12695);
nand_4 g10358(new_n12707_1, new_n12706, new_n12693);
nand_4 g10359(new_n12708, new_n12707_1, new_n12691);
xnor_3 g10360(new_n12709, new_n12708, new_n12689);
not_3  g10361(new_n12710, new_n12709);
nor_4  g10362(new_n12711, new_n12710, new_n12667);
nor_4  g10363(new_n12712, new_n12709, new_n12666);
nor_4  g10364(new_n12713, new_n12712, new_n12711);
not_3  g10365(new_n12714, new_n12647);
xnor_3 g10366(new_n12715, new_n12663, new_n12714);
xnor_3 g10367(new_n12716, new_n12706, new_n12693);
not_3  g10368(new_n12717, new_n12716);
nand_4 g10369(new_n12718, new_n12717, new_n12715);
xnor_3 g10370(new_n12719, new_n12716, new_n12715);
xnor_3 g10371(new_n12720, new_n12661, new_n12650_1);
not_3  g10372(new_n12721, new_n12720);
xnor_3 g10373(new_n12722, new_n12704, new_n12703);
nand_4 g10374(new_n12723, new_n12722, new_n12721);
xnor_3 g10375(new_n12724, new_n12722, new_n12720);
xor_3  g10376(new_n12725_1, new_n9477, n20923);
xnor_3 g10377(new_n12726, new_n12659, new_n12725_1);
xnor_3 g10378(new_n12727_1, new_n12701, new_n12699);
not_3  g10379(new_n12728, new_n12727_1);
nand_4 g10380(new_n12729, new_n12728, new_n12726);
not_3  g10381(new_n12730, new_n12729);
nor_4  g10382(new_n12731, new_n12728, new_n12726);
nor_4  g10383(new_n12732, new_n12731, new_n12730);
nor_4  g10384(new_n12733, new_n10092, new_n10062);
nor_4  g10385(new_n12734, new_n10104, new_n10093);
nor_4  g10386(new_n12735, new_n12734, new_n12733);
nand_4 g10387(new_n12736, new_n12735, new_n12732);
nand_4 g10388(new_n12737, new_n12736, new_n12729);
nand_4 g10389(new_n12738, new_n12737, new_n12724);
nand_4 g10390(new_n12739, new_n12738, new_n12723);
nand_4 g10391(new_n12740_1, new_n12739, new_n12719);
nand_4 g10392(new_n12741, new_n12740_1, new_n12718);
xnor_3 g10393(n1371, new_n12741, new_n12713);
xor_3  g10394(new_n12743, n17250, new_n4922);
nor_4  g10395(new_n12744, new_n9090_1, n7678);
not_3  g10396(new_n12745, new_n12744);
not_3  g10397(new_n12746_1, n16524);
nor_4  g10398(new_n12747, new_n12746_1, n3785);
not_3  g10399(new_n12748, new_n12747);
xor_3  g10400(new_n12749, n16524, new_n4935);
nor_4  g10401(new_n12750, new_n4943, n11056);
nor_4  g10402(new_n12751, n15271, new_n4947_1);
xor_3  g10403(new_n12752, n15271, n5822);
not_3  g10404(new_n12753, new_n6739);
nand_4 g10405(new_n12754, new_n6740, new_n6724);
nand_4 g10406(new_n12755, new_n12754, new_n12753);
not_3  g10407(new_n12756_1, new_n12755);
nor_4  g10408(new_n12757, new_n12756_1, new_n12752);
nor_4  g10409(new_n12758, new_n12757, new_n12751);
xor_3  g10410(new_n12759, n20250, new_n9098);
not_3  g10411(new_n12760, new_n12759);
nor_4  g10412(new_n12761, new_n12760, new_n12758);
nor_4  g10413(new_n12762, new_n12761, new_n12750);
nand_4 g10414(new_n12763, new_n12762, new_n12749);
nand_4 g10415(new_n12764, new_n12763, new_n12748);
not_3  g10416(new_n12765, n7678);
xor_3  g10417(new_n12766, n23160, new_n12765);
nand_4 g10418(new_n12767, new_n12766, new_n12764);
nand_4 g10419(new_n12768, new_n12767, new_n12745);
xnor_3 g10420(new_n12769, new_n12768, new_n12743);
xor_3  g10421(new_n12770, new_n11607_1, new_n8849_1);
not_3  g10422(new_n12771, new_n12770);
nor_4  g10423(new_n12772, new_n11613, n26660);
not_3  g10424(new_n12773, new_n12772);
xnor_3 g10425(new_n12774, new_n11613, n26660);
not_3  g10426(new_n12775, new_n12774);
nor_4  g10427(new_n12776, new_n11616, new_n9045);
nor_4  g10428(new_n12777, new_n11615_1, n3018);
nor_4  g10429(new_n12778, new_n11342, new_n11326_1);
not_3  g10430(new_n12779, new_n12778);
nor_4  g10431(new_n12780, new_n12779, new_n12777);
nor_4  g10432(new_n12781, new_n12780, new_n12776);
nand_4 g10433(new_n12782, new_n12781, new_n12775);
nand_4 g10434(new_n12783_1, new_n12782, new_n12773);
xnor_3 g10435(new_n12784, new_n12783_1, new_n12771);
xnor_3 g10436(new_n12785, new_n12784, new_n12769);
xnor_3 g10437(new_n12786, new_n12781, new_n12774);
not_3  g10438(new_n12787, new_n12749);
not_3  g10439(new_n12788, new_n12750);
not_3  g10440(new_n12789, new_n12751);
not_3  g10441(new_n12790, new_n12752);
nand_4 g10442(new_n12791, new_n12755, new_n12790);
nand_4 g10443(new_n12792, new_n12791, new_n12789);
nand_4 g10444(new_n12793, new_n12759, new_n12792);
nand_4 g10445(new_n12794, new_n12793, new_n12788);
nor_4  g10446(new_n12795, new_n12794, new_n12787);
nor_4  g10447(new_n12796, new_n12795, new_n12747);
not_3  g10448(new_n12797, new_n12766);
xnor_3 g10449(new_n12798, new_n12797, new_n12796);
nor_4  g10450(new_n12799, new_n12798, new_n12786);
xnor_3 g10451(new_n12800, new_n12798, new_n12786);
xnor_3 g10452(new_n12801_1, new_n12794, new_n12787);
not_3  g10453(new_n12802, new_n12801_1);
xor_3  g10454(new_n12803, new_n11616, new_n9045);
nand_4 g10455(new_n12804, new_n12803, new_n12778);
xor_3  g10456(new_n12805, new_n11616, n3018);
nand_4 g10457(new_n12806, new_n12805, new_n12779);
nand_4 g10458(new_n12807, new_n12806, new_n12804);
not_3  g10459(new_n12808, new_n12807);
nor_4  g10460(new_n12809, new_n12808, new_n12802);
not_3  g10461(new_n12810, new_n12809);
xnor_3 g10462(new_n12811_1, new_n12807, new_n12802);
xnor_3 g10463(new_n12812_1, new_n12759, new_n12792);
nor_4  g10464(new_n12813, new_n12812_1, new_n11349);
not_3  g10465(new_n12814, new_n12813);
xnor_3 g10466(new_n12815, new_n12812_1, new_n11349);
not_3  g10467(new_n12816_1, new_n12815);
xnor_3 g10468(new_n12817, new_n12756_1, new_n12752);
not_3  g10469(new_n12818, new_n12817);
nor_4  g10470(new_n12819, new_n12818, new_n11352_1);
xnor_3 g10471(new_n12820, new_n12817, new_n11356_1);
not_3  g10472(new_n12821_1, new_n6743);
nand_4 g10473(new_n12822, new_n6760, new_n12821_1);
not_3  g10474(new_n12823, new_n12822);
nor_4  g10475(new_n12824, new_n12823, new_n12820);
nor_4  g10476(new_n12825, new_n12824, new_n12819);
nand_4 g10477(new_n12826, new_n12825, new_n12816_1);
nand_4 g10478(new_n12827, new_n12826, new_n12814);
nand_4 g10479(new_n12828, new_n12827, new_n12811_1);
nand_4 g10480(new_n12829, new_n12828, new_n12810);
nor_4  g10481(new_n12830, new_n12829, new_n12800);
nor_4  g10482(new_n12831, new_n12830, new_n12799);
nor_4  g10483(new_n12832, new_n12831, new_n12785);
nand_4 g10484(new_n12833, new_n12831, new_n12785);
not_3  g10485(new_n12834, new_n12833);
nor_4  g10486(new_n12835, new_n12834, new_n12832);
xnor_3 g10487(new_n12836, new_n12835, new_n6535);
xnor_3 g10488(new_n12837, new_n12829, new_n12800);
not_3  g10489(new_n12838, new_n12837);
nor_4  g10490(new_n12839, new_n12838, new_n6544);
not_3  g10491(new_n12840, new_n12839);
nor_4  g10492(new_n12841, new_n12837, new_n6537);
nor_4  g10493(new_n12842, new_n12841, new_n12839);
xnor_3 g10494(new_n12843_1, new_n12827, new_n12811_1);
not_3  g10495(new_n12844, new_n12843_1);
nor_4  g10496(new_n12845, new_n12844, new_n6546);
not_3  g10497(new_n12846, new_n12819);
not_3  g10498(new_n12847, new_n12824);
nand_4 g10499(new_n12848, new_n12847, new_n12846);
xnor_3 g10500(new_n12849, new_n12848, new_n12815);
nor_4  g10501(new_n12850, new_n12849, new_n12341_1);
not_3  g10502(new_n12851, new_n12850);
xnor_3 g10503(new_n12852, new_n12849, new_n12341_1);
not_3  g10504(new_n12853, new_n12852);
xnor_3 g10505(new_n12854, new_n12823, new_n12820);
nor_4  g10506(new_n12855, new_n12854, new_n6566);
nor_4  g10507(new_n12856, new_n6732, new_n6573);
nor_4  g10508(new_n12857, new_n6764, new_n6734);
nor_4  g10509(new_n12858, new_n12857, new_n12856);
xnor_3 g10510(new_n12859, new_n12854, new_n6566);
nor_4  g10511(new_n12860, new_n12859, new_n12858);
nor_4  g10512(new_n12861_1, new_n12860, new_n12855);
nand_4 g10513(new_n12862, new_n12861_1, new_n12853);
nand_4 g10514(new_n12863, new_n12862, new_n12851);
xnor_3 g10515(new_n12864_1, new_n12843_1, new_n6547);
nor_4  g10516(new_n12865_1, new_n12864_1, new_n12863);
nor_4  g10517(new_n12866, new_n12865_1, new_n12845);
nand_4 g10518(new_n12867, new_n12866, new_n12842);
nand_4 g10519(new_n12868, new_n12867, new_n12840);
xor_3  g10520(n1385, new_n12868, new_n12836);
not_3  g10521(new_n12870_1, new_n10931);
not_3  g10522(new_n12871_1, new_n9446);
nand_4 g10523(new_n12872, n26808, n24732);
not_3  g10524(new_n12873_1, new_n12872);
nor_4  g10525(new_n12874, n26808, n24732);
nor_4  g10526(new_n12875_1, new_n12874, new_n12873_1);
xnor_3 g10527(new_n12876, n7339, n6631);
xnor_3 g10528(new_n12877, new_n12876, new_n12872);
not_3  g10529(new_n12878, new_n12877);
nor_4  g10530(new_n12879, new_n12878, new_n12875_1);
not_3  g10531(new_n12880, new_n12879);
xnor_3 g10532(new_n12881, n14684, n1667);
not_3  g10533(new_n12882, new_n12881);
nor_4  g10534(new_n12883, n7339, n6631);
not_3  g10535(new_n12884, new_n12883);
not_3  g10536(new_n12885, new_n12876);
nand_4 g10537(new_n12886, new_n12885, new_n12872);
nand_4 g10538(new_n12887, new_n12886, new_n12884);
xnor_3 g10539(new_n12888, new_n12887, new_n12882);
nor_4  g10540(new_n12889, new_n12888, new_n12880);
xor_3  g10541(new_n12890, n17035, n2680);
nor_4  g10542(new_n12891, n14684, n1667);
not_3  g10543(new_n12892_1, new_n12891);
nand_4 g10544(new_n12893, new_n12887, new_n12882);
nand_4 g10545(new_n12894, new_n12893, new_n12892_1);
nor_4  g10546(new_n12895, new_n12894, new_n12890);
nand_4 g10547(new_n12896, new_n12894, new_n12890);
not_3  g10548(new_n12897, new_n12896);
nor_4  g10549(new_n12898, new_n12897, new_n12895);
nand_4 g10550(new_n12899, new_n12898, new_n12889);
not_3  g10551(new_n12900_1, new_n12899);
xor_3  g10552(new_n12901, n19905, n2547);
nor_4  g10553(new_n12902, n17035, n2680);
not_3  g10554(new_n12903, new_n12902);
nand_4 g10555(new_n12904_1, new_n12896, new_n12903);
nor_4  g10556(new_n12905, new_n12904_1, new_n12901);
nand_4 g10557(new_n12906, new_n12904_1, new_n12901);
not_3  g10558(new_n12907, new_n12906);
nor_4  g10559(new_n12908, new_n12907, new_n12905);
nand_4 g10560(new_n12909, new_n12908, new_n12900_1);
xor_3  g10561(new_n12910, n26452, n2999);
nor_4  g10562(new_n12911, n19905, n2547);
not_3  g10563(new_n12912, new_n12911);
nand_4 g10564(new_n12913, new_n12906, new_n12912);
nor_4  g10565(new_n12914, new_n12913, new_n12910);
nand_4 g10566(new_n12915, new_n12913, new_n12910);
not_3  g10567(new_n12916, new_n12915);
nor_4  g10568(new_n12917_1, new_n12916, new_n12914);
not_3  g10569(new_n12918, new_n12917_1);
nor_4  g10570(new_n12919, new_n12918, new_n12909);
xor_3  g10571(new_n12920, n15546, n14702);
nor_4  g10572(new_n12921, n26452, n2999);
not_3  g10573(new_n12922, new_n12921);
nand_4 g10574(new_n12923, new_n12915, new_n12922);
xnor_3 g10575(new_n12924, new_n12923, new_n12920);
not_3  g10576(new_n12925, new_n12924);
nand_4 g10577(new_n12926, new_n12925, new_n12919);
xor_3  g10578(new_n12927, n13914, n5077);
nand_4 g10579(new_n12928, new_n12692, new_n10949);
nand_4 g10580(new_n12929, new_n12923, new_n12920);
nand_4 g10581(new_n12930, new_n12929, new_n12928);
nor_4  g10582(new_n12931, new_n12930, new_n12927);
not_3  g10583(new_n12932, new_n12927);
not_3  g10584(new_n12933, new_n12930);
nor_4  g10585(new_n12934, new_n12933, new_n12932);
nor_4  g10586(new_n12935, new_n12934, new_n12931);
not_3  g10587(new_n12936, new_n12935);
nor_4  g10588(new_n12937, new_n12936, new_n12926);
not_3  g10589(new_n12938, new_n12937);
xor_3  g10590(new_n12939, n18035, n3279);
nor_4  g10591(new_n12940, n13914, n5077);
nor_4  g10592(new_n12941_1, new_n12934, new_n12940);
xnor_3 g10593(new_n12942_1, new_n12941_1, new_n12939);
not_3  g10594(new_n12943, new_n12942_1);
nor_4  g10595(new_n12944, new_n12943, new_n12938);
xor_3  g10596(new_n12945, n8827, n4306);
not_3  g10597(new_n12946, new_n12945);
nor_4  g10598(new_n12947, n18035, n3279);
not_3  g10599(new_n12948, new_n12939);
nor_4  g10600(new_n12949, new_n12941_1, new_n12948);
nor_4  g10601(new_n12950, new_n12949, new_n12947);
xnor_3 g10602(new_n12951, new_n12950, new_n12946);
not_3  g10603(new_n12952, new_n12951);
xnor_3 g10604(new_n12953, new_n12952, new_n12944);
xnor_3 g10605(new_n12954, new_n12953, new_n12871_1);
xnor_3 g10606(new_n12955, new_n12942_1, new_n12937);
nand_4 g10607(new_n12956_1, new_n12955, new_n9451_1);
not_3  g10608(new_n12957, new_n9451_1);
xnor_3 g10609(new_n12958, new_n12955, new_n12957);
xnor_3 g10610(new_n12959, new_n12936, new_n12926);
nand_4 g10611(new_n12960, new_n12959, new_n9455);
xnor_3 g10612(new_n12961, new_n12959, new_n9454);
xnor_3 g10613(new_n12962, new_n12925, new_n12919);
nand_4 g10614(new_n12963, new_n12962, new_n9463);
xnor_3 g10615(new_n12964, new_n12962, new_n9461);
xnor_3 g10616(new_n12965, new_n12918, new_n12909);
nand_4 g10617(new_n12966, new_n12965, new_n9470);
xnor_3 g10618(new_n12967, new_n12965, new_n9468);
xnor_3 g10619(new_n12968, new_n12908, new_n12900_1);
nand_4 g10620(new_n12969, new_n12968, new_n9477);
xnor_3 g10621(new_n12970, new_n12968, new_n9475);
xnor_3 g10622(new_n12971, new_n12898, new_n12889);
nand_4 g10623(new_n12972, new_n12971, new_n9482);
xnor_3 g10624(new_n12973, new_n12971, new_n9481);
xnor_3 g10625(new_n12974, new_n12888, new_n12880);
not_3  g10626(new_n12975, new_n12974);
nor_4  g10627(new_n12976, new_n12975, new_n9489);
nor_4  g10628(new_n12977, new_n12974, new_n10050);
nor_4  g10629(new_n12978_1, new_n12977, new_n12976);
not_3  g10630(new_n12979, new_n12875_1);
nor_4  g10631(new_n12980_1, new_n12979, new_n2593);
not_3  g10632(new_n12981, new_n12980_1);
nand_4 g10633(new_n12982, new_n12981, new_n9496);
not_3  g10634(new_n12983, new_n12982);
nor_4  g10635(new_n12984, new_n12876, new_n12979);
nor_4  g10636(new_n12985_1, new_n12984, new_n12879);
nand_4 g10637(new_n12986, new_n12980_1, new_n9424);
nand_4 g10638(new_n12987_1, new_n12986, new_n12982);
nor_4  g10639(new_n12988, new_n12987_1, new_n12985_1);
nor_4  g10640(new_n12989, new_n12988, new_n12983);
not_3  g10641(new_n12990, new_n12989);
nand_4 g10642(new_n12991, new_n12990, new_n12978_1);
not_3  g10643(new_n12992_1, new_n12991);
nor_4  g10644(new_n12993, new_n12992_1, new_n12976);
not_3  g10645(new_n12994, new_n12993);
nand_4 g10646(new_n12995, new_n12994, new_n12973);
nand_4 g10647(new_n12996, new_n12995, new_n12972);
nand_4 g10648(new_n12997, new_n12996, new_n12970);
nand_4 g10649(new_n12998, new_n12997, new_n12969);
nand_4 g10650(new_n12999, new_n12998, new_n12967);
nand_4 g10651(new_n13000, new_n12999, new_n12966);
nand_4 g10652(new_n13001, new_n13000, new_n12964);
nand_4 g10653(new_n13002, new_n13001, new_n12963);
nand_4 g10654(new_n13003, new_n13002, new_n12961);
nand_4 g10655(new_n13004, new_n13003, new_n12960);
nand_4 g10656(new_n13005_1, new_n13004, new_n12958);
nand_4 g10657(new_n13006, new_n13005_1, new_n12956_1);
xnor_3 g10658(new_n13007, new_n13006, new_n12954);
nor_4  g10659(new_n13008, new_n13007, new_n12870_1);
not_3  g10660(new_n13009, new_n13007);
nor_4  g10661(new_n13010, new_n13009, new_n10931);
nor_4  g10662(new_n13011, new_n13010, new_n13008);
xnor_3 g10663(new_n13012, new_n13004, new_n12958);
nor_4  g10664(new_n13013, new_n13012, new_n10936);
not_3  g10665(new_n13014, new_n13013);
not_3  g10666(new_n13015, new_n13012);
nor_4  g10667(new_n13016, new_n13015, new_n10939);
nor_4  g10668(new_n13017, new_n13016, new_n13013);
xnor_3 g10669(new_n13018, new_n13002, new_n12961);
nor_4  g10670(new_n13019, new_n13018, new_n10944);
not_3  g10671(new_n13020, new_n13019);
not_3  g10672(new_n13021, new_n13018);
nor_4  g10673(new_n13022, new_n13021, new_n10945);
nor_4  g10674(new_n13023, new_n13022, new_n13019);
not_3  g10675(new_n13024, new_n12964);
xnor_3 g10676(new_n13025, new_n13000, new_n13024);
nand_4 g10677(new_n13026_1, new_n13025, new_n10952);
xnor_3 g10678(new_n13027, new_n13025, new_n10951);
not_3  g10679(new_n13028, new_n12967);
xnor_3 g10680(new_n13029, new_n12998, new_n13028);
nand_4 g10681(new_n13030, new_n13029, new_n10961_1);
xnor_3 g10682(new_n13031, new_n13029, new_n10960);
not_3  g10683(new_n13032, new_n12970);
xnor_3 g10684(new_n13033, new_n12996, new_n13032);
nand_4 g10685(new_n13034, new_n13033, new_n10973);
xnor_3 g10686(new_n13035, new_n13033, new_n10977);
xnor_3 g10687(new_n13036, new_n12994, new_n12973);
nor_4  g10688(new_n13037, new_n13036, new_n10984);
not_3  g10689(new_n13038, new_n13037);
xnor_3 g10690(new_n13039, new_n12990, new_n12978_1);
nor_4  g10691(new_n13040, new_n13039, new_n10990);
not_3  g10692(new_n13041, new_n13040);
not_3  g10693(new_n13042, new_n13039);
nor_4  g10694(new_n13043_1, new_n13042, new_n10989);
nor_4  g10695(new_n13044_1, new_n13043_1, new_n13040);
xor_3  g10696(new_n13045, n22843, new_n10912);
xor_3  g10697(new_n13046, new_n12979, new_n2593);
nor_4  g10698(new_n13047, new_n13046, new_n13045);
not_3  g10699(new_n13048_1, new_n13047);
nor_4  g10700(new_n13049, new_n13048_1, new_n10996);
not_3  g10701(new_n13050, new_n13049);
xor_3  g10702(new_n13051, new_n13048_1, new_n10996);
xor_3  g10703(new_n13052, new_n12987_1, new_n12985_1);
nand_4 g10704(new_n13053, new_n13052, new_n13051);
nand_4 g10705(new_n13054_1, new_n13053, new_n13050);
nand_4 g10706(new_n13055, new_n13054_1, new_n13044_1);
nand_4 g10707(new_n13056, new_n13055, new_n13041);
not_3  g10708(new_n13057, new_n13036);
nor_4  g10709(new_n13058, new_n13057, new_n10983);
nor_4  g10710(new_n13059, new_n13058, new_n13037);
nand_4 g10711(new_n13060, new_n13059, new_n13056);
nand_4 g10712(new_n13061, new_n13060, new_n13038);
nand_4 g10713(new_n13062, new_n13061, new_n13035);
nand_4 g10714(new_n13063, new_n13062, new_n13034);
nand_4 g10715(new_n13064, new_n13063, new_n13031);
nand_4 g10716(new_n13065, new_n13064, new_n13030);
nand_4 g10717(new_n13066, new_n13065, new_n13027);
nand_4 g10718(new_n13067, new_n13066, new_n13026_1);
nand_4 g10719(new_n13068, new_n13067, new_n13023);
nand_4 g10720(new_n13069, new_n13068, new_n13020);
nand_4 g10721(new_n13070, new_n13069, new_n13017);
nand_4 g10722(new_n13071, new_n13070, new_n13014);
xnor_3 g10723(n1498, new_n13071, new_n13011);
xnor_3 g10724(new_n13073, n20658, n9090);
xor_3  g10725(new_n13074_1, new_n13073, new_n6985_1);
xor_3  g10726(n1501, new_n13074_1, new_n5719);
not_3  g10727(new_n13076, n752);
not_3  g10728(new_n13077, n25094);
not_3  g10729(new_n13078, n5131);
nor_4  g10730(new_n13079, n15506, n11473);
nand_4 g10731(new_n13080, new_n13079, new_n13078);
nor_4  g10732(new_n13081, new_n13080, n21538);
nand_4 g10733(new_n13082_1, new_n13081, new_n13077);
nor_4  g10734(new_n13083, new_n13082_1, n1611);
xor_3  g10735(new_n13084, new_n13083, new_n13076);
xnor_3 g10736(new_n13085, new_n13084, new_n11653);
not_3  g10737(new_n13086, new_n13085);
xor_3  g10738(new_n13087, new_n13082_1, n1611);
not_3  g10739(new_n13088, new_n13087);
nand_4 g10740(new_n13089, new_n13088, new_n11658);
not_3  g10741(new_n13090, new_n13089);
xnor_3 g10742(new_n13091, new_n13088, new_n11658);
not_3  g10743(new_n13092, new_n13082_1);
nor_4  g10744(new_n13093, new_n13081, new_n13077);
nor_4  g10745(new_n13094, new_n13093, new_n13092);
nor_4  g10746(new_n13095, new_n13094, new_n11663);
xnor_3 g10747(new_n13096_1, new_n13094, new_n11663);
nand_4 g10748(new_n13097, new_n13080, n21538);
not_3  g10749(new_n13098, new_n13097);
nor_4  g10750(new_n13099, new_n13098, new_n13081);
nor_4  g10751(new_n13100, new_n13099, new_n11670);
not_3  g10752(new_n13101, new_n13080);
nor_4  g10753(new_n13102, new_n13079, new_n13078);
nor_4  g10754(new_n13103, new_n13102, new_n13101);
nor_4  g10755(new_n13104, new_n13103, new_n11681);
xnor_3 g10756(new_n13105, new_n13103, new_n11681);
not_3  g10757(new_n13106, n15506);
nor_4  g10758(new_n13107, new_n11691, new_n13106);
xnor_3 g10759(new_n13108, n15506, n11473);
not_3  g10760(new_n13109, new_n13108);
nor_4  g10761(new_n13110_1, new_n13109, new_n13107);
not_3  g10762(new_n13111, n11473);
nand_4 g10763(new_n13112, new_n13107, new_n13111);
not_3  g10764(new_n13113, new_n13112);
nor_4  g10765(new_n13114, new_n13113, new_n13110_1);
not_3  g10766(new_n13115, new_n13114);
nor_4  g10767(new_n13116_1, new_n13115, new_n11688);
nor_4  g10768(new_n13117, new_n13116_1, new_n13110_1);
nor_4  g10769(new_n13118, new_n13117, new_n13105);
nor_4  g10770(new_n13119, new_n13118, new_n13104);
xnor_3 g10771(new_n13120, new_n13099, new_n11670);
nor_4  g10772(new_n13121, new_n13120, new_n13119);
nor_4  g10773(new_n13122_1, new_n13121, new_n13100);
nor_4  g10774(new_n13123, new_n13122_1, new_n13096_1);
nor_4  g10775(new_n13124, new_n13123, new_n13095);
nor_4  g10776(new_n13125, new_n13124, new_n13091);
nor_4  g10777(new_n13126, new_n13125, new_n13090);
xnor_3 g10778(new_n13127, new_n13126, new_n13086);
xor_3  g10779(new_n13128, n20470, n3366);
nand_4 g10780(new_n13129, n26565, n21222);
not_3  g10781(new_n13130, new_n13129);
nor_4  g10782(new_n13131, n26565, n21222);
nor_4  g10783(new_n13132, n9832, n3959);
not_3  g10784(new_n13133, new_n13132);
nand_4 g10785(new_n13134, new_n11437, new_n13133);
nor_4  g10786(new_n13135, new_n13134, new_n13131);
nor_4  g10787(new_n13136, new_n13135, new_n13130);
xnor_3 g10788(new_n13137_1, new_n13136, new_n13128);
not_3  g10789(new_n13138, new_n13137_1);
xnor_3 g10790(new_n13139, new_n13138, new_n13127);
not_3  g10791(new_n13140, new_n13091);
not_3  g10792(new_n13141_1, new_n13095);
not_3  g10793(new_n13142, new_n13096_1);
not_3  g10794(new_n13143, new_n13100);
not_3  g10795(new_n13144_1, new_n13104);
not_3  g10796(new_n13145, new_n13118);
nand_4 g10797(new_n13146, new_n13145, new_n13144_1);
not_3  g10798(new_n13147, new_n13120);
nand_4 g10799(new_n13148, new_n13147, new_n13146);
nand_4 g10800(new_n13149, new_n13148, new_n13143);
nand_4 g10801(new_n13150, new_n13149, new_n13142);
nand_4 g10802(new_n13151, new_n13150, new_n13141_1);
xnor_3 g10803(new_n13152, new_n13151, new_n13140);
not_3  g10804(new_n13153, new_n13134);
nor_4  g10805(new_n13154, new_n13131, new_n13130);
xor_3  g10806(new_n13155, new_n13154, new_n13153);
not_3  g10807(new_n13156, new_n13155);
nor_4  g10808(new_n13157, new_n13156, new_n13152);
not_3  g10809(new_n13158, new_n13157);
xnor_3 g10810(new_n13159, new_n13155, new_n13152);
xnor_3 g10811(new_n13160, new_n13149, new_n13142);
nor_4  g10812(new_n13161, new_n13160, new_n11439_1);
not_3  g10813(new_n13162, new_n13161);
not_3  g10814(new_n13163, new_n13160);
nor_4  g10815(new_n13164, new_n13163, new_n11440);
nor_4  g10816(new_n13165, new_n13164, new_n13161);
xnor_3 g10817(new_n13166, new_n13120, new_n13119);
nor_4  g10818(new_n13167, new_n13166, new_n11520);
not_3  g10819(new_n13168_1, new_n13167);
not_3  g10820(new_n13169, new_n13166);
nor_4  g10821(new_n13170, new_n13169, new_n11521);
nor_4  g10822(new_n13171, new_n13170, new_n13167);
xnor_3 g10823(new_n13172, new_n13117, new_n13105);
not_3  g10824(new_n13173, new_n13172);
nor_4  g10825(new_n13174, new_n13173, new_n11529);
xnor_3 g10826(new_n13175, new_n13114, new_n11687);
nor_4  g10827(new_n13176, new_n13175, new_n11535);
xor_3  g10828(new_n13177, new_n11691, new_n13106);
nor_4  g10829(new_n13178, new_n13177, new_n11538_1);
not_3  g10830(new_n13179, new_n13178);
not_3  g10831(new_n13180, new_n13175);
nor_4  g10832(new_n13181, new_n13180, new_n11540);
nor_4  g10833(new_n13182, new_n13181, new_n13176);
not_3  g10834(new_n13183, new_n13182);
nor_4  g10835(new_n13184, new_n13183, new_n13179);
nor_4  g10836(new_n13185, new_n13184, new_n13176);
not_3  g10837(new_n13186, new_n13185);
not_3  g10838(new_n13187, new_n11529);
xnor_3 g10839(new_n13188, new_n13172, new_n13187);
nor_4  g10840(new_n13189, new_n13188, new_n13186);
nor_4  g10841(new_n13190_1, new_n13189, new_n13174);
nand_4 g10842(new_n13191, new_n13190_1, new_n13171);
nand_4 g10843(new_n13192, new_n13191, new_n13168_1);
nand_4 g10844(new_n13193, new_n13192, new_n13165);
nand_4 g10845(new_n13194, new_n13193, new_n13162);
nand_4 g10846(new_n13195, new_n13194, new_n13159);
nand_4 g10847(new_n13196, new_n13195, new_n13158);
not_3  g10848(new_n13197, new_n13196);
xor_3  g10849(n1518, new_n13197, new_n13139);
not_3  g10850(new_n13199_1, n17458);
nor_4  g10851(new_n13200, new_n13199_1, n14826);
xor_3  g10852(new_n13201, n17458, new_n11929);
not_3  g10853(new_n13202, new_n13201);
nor_4  g10854(new_n13203, n23493, new_n8501);
xor_3  g10855(new_n13204_1, n23493, new_n8501);
nand_4 g10856(new_n13205, n25240, new_n11919);
xor_3  g10857(new_n13206, n25240, new_n11919);
nand_4 g10858(new_n13207, new_n9403_1, n10125);
xor_3  g10859(new_n13208, n15146, new_n8506);
nand_4 g10860(new_n13209_1, new_n11885, n8067);
xor_3  g10861(new_n13210, n11579, new_n8509);
nor_4  g10862(new_n13211, new_n12653, n21);
not_3  g10863(new_n13212, new_n13211);
xor_3  g10864(new_n13213, n20923, new_n11887);
nor_4  g10865(new_n13214, new_n8519_1, n1682);
not_3  g10866(new_n13215, new_n13214);
xor_3  g10867(new_n13216, n18157, new_n11891);
nor_4  g10868(new_n13217, n12161, new_n11896);
nor_4  g10869(new_n13218, new_n7792, n7963);
nor_4  g10870(new_n13219, new_n11898_1, n5026);
nor_4  g10871(new_n13220, n10017, new_n8524);
nand_4 g10872(new_n13221, new_n8626, n3618);
nor_4  g10873(new_n13222, new_n13221, new_n13220);
nor_4  g10874(new_n13223, new_n13222, new_n13219);
nor_4  g10875(new_n13224, new_n13223, new_n13218);
nor_4  g10876(new_n13225, new_n13224, new_n13217);
nand_4 g10877(new_n13226, new_n13225, new_n13216);
nand_4 g10878(new_n13227, new_n13226, new_n13215);
nand_4 g10879(new_n13228, new_n13227, new_n13213);
nand_4 g10880(new_n13229, new_n13228, new_n13212);
nand_4 g10881(new_n13230, new_n13229, new_n13210);
nand_4 g10882(new_n13231, new_n13230, new_n13209_1);
nand_4 g10883(new_n13232, new_n13231, new_n13208);
nand_4 g10884(new_n13233, new_n13232, new_n13207);
nand_4 g10885(new_n13234, new_n13233, new_n13206);
nand_4 g10886(new_n13235, new_n13234, new_n13205);
nand_4 g10887(new_n13236, new_n13235, new_n13204_1);
not_3  g10888(new_n13237, new_n13236);
nor_4  g10889(new_n13238, new_n13237, new_n13203);
nor_4  g10890(new_n13239, new_n13238, new_n13202);
nor_4  g10891(new_n13240, new_n13239, new_n13200);
not_3  g10892(new_n13241, new_n13240);
nor_4  g10893(new_n13242, new_n4704, n12821);
not_3  g10894(new_n13243, new_n13242);
nor_4  g10895(new_n13244, new_n13243, n22492);
nand_4 g10896(new_n13245, new_n13244, new_n2985_1);
nor_4  g10897(new_n13246, new_n13245, n767);
not_3  g10898(new_n13247, new_n13246);
nor_4  g10899(new_n13248, new_n13247, n2944);
not_3  g10900(new_n13249, new_n13248);
not_3  g10901(new_n13250, n2944);
xor_3  g10902(new_n13251, new_n13246, new_n13250);
nor_4  g10903(new_n13252, new_n13251, n19282);
not_3  g10904(new_n13253, new_n13252);
not_3  g10905(new_n13254, new_n13245);
xor_3  g10906(new_n13255, new_n13254, new_n2983);
not_3  g10907(new_n13256, new_n13255);
nand_4 g10908(new_n13257, new_n13256, new_n8553);
xor_3  g10909(new_n13258, new_n13256, new_n8553);
xor_3  g10910(new_n13259, new_n13244, new_n2985_1);
not_3  g10911(new_n13260, new_n13259);
nor_4  g10912(new_n13261, new_n13260, new_n8555);
xor_3  g10913(new_n13262, new_n13260, n17077);
xor_3  g10914(new_n13263_1, new_n13242, new_n2781);
not_3  g10915(new_n13264, new_n13263_1);
nor_4  g10916(new_n13265, new_n13264, new_n3081);
xor_3  g10917(new_n13266, new_n13264, new_n3081);
not_3  g10918(new_n13267, new_n13266);
xor_3  g10919(new_n13268, new_n4704, n12821);
not_3  g10920(new_n13269, new_n13268);
nor_4  g10921(new_n13270_1, new_n13269, new_n4187);
nor_4  g10922(new_n13271, new_n13268, n23068);
nand_4 g10923(new_n13272, new_n4742, new_n4711);
not_3  g10924(new_n13273_1, new_n13272);
nor_4  g10925(new_n13274, new_n13273_1, new_n4709);
nor_4  g10926(new_n13275, new_n13274, new_n13271);
nor_4  g10927(new_n13276, new_n13275, new_n13270_1);
nor_4  g10928(new_n13277, new_n13276, new_n13267);
nor_4  g10929(new_n13278, new_n13277, new_n13265);
nor_4  g10930(new_n13279, new_n13278, new_n13262);
nor_4  g10931(new_n13280, new_n13279, new_n13261);
nand_4 g10932(new_n13281, new_n13280, new_n13258);
nand_4 g10933(new_n13282, new_n13281, new_n13257);
not_3  g10934(new_n13283, new_n13251);
nor_4  g10935(new_n13284, new_n13283, new_n8549);
not_3  g10936(new_n13285_1, new_n13284);
nand_4 g10937(new_n13286, new_n13285_1, new_n13282);
nand_4 g10938(new_n13287, new_n13286, new_n13253);
nand_4 g10939(new_n13288, new_n13287, new_n13249);
nand_4 g10940(new_n13289, new_n13288, new_n13241);
xor_3  g10941(new_n13290, new_n13238, new_n13202);
nor_4  g10942(new_n13291, new_n13284, new_n13252);
xnor_3 g10943(new_n13292, new_n13291, new_n13282);
nor_4  g10944(new_n13293, new_n13292, new_n13290);
not_3  g10945(new_n13294, new_n13290);
not_3  g10946(new_n13295, new_n13292);
nor_4  g10947(new_n13296, new_n13295, new_n13294);
nor_4  g10948(new_n13297, new_n13296, new_n13293);
xnor_3 g10949(new_n13298, new_n13235, new_n13204_1);
xnor_3 g10950(new_n13299, new_n13280, new_n13258);
not_3  g10951(new_n13300, new_n13299);
nand_4 g10952(new_n13301, new_n13300, new_n13298);
not_3  g10953(new_n13302, new_n13298);
nor_4  g10954(new_n13303, new_n13299, new_n13302);
nor_4  g10955(new_n13304, new_n13300, new_n13298);
nor_4  g10956(new_n13305, new_n13304, new_n13303);
xnor_3 g10957(new_n13306, new_n13233, new_n13206);
xnor_3 g10958(new_n13307, new_n13278, new_n13262);
nand_4 g10959(new_n13308, new_n13307, new_n13306);
not_3  g10960(new_n13309, new_n13306);
xnor_3 g10961(new_n13310, new_n13307, new_n13309);
xnor_3 g10962(new_n13311, new_n13231, new_n13208);
xnor_3 g10963(new_n13312, new_n13276, new_n13266);
not_3  g10964(new_n13313, new_n13312);
nand_4 g10965(new_n13314, new_n13313, new_n13311);
xnor_3 g10966(new_n13315, new_n13312, new_n13311);
xnor_3 g10967(new_n13316, new_n13229, new_n13210);
not_3  g10968(new_n13317, new_n13316);
nor_4  g10969(new_n13318, new_n13271, new_n13270_1);
xnor_3 g10970(new_n13319_1, new_n13318, new_n13274);
nor_4  g10971(new_n13320, new_n13319_1, new_n13317);
not_3  g10972(new_n13321, new_n13320);
not_3  g10973(new_n13322, new_n13319_1);
nor_4  g10974(new_n13323, new_n13322, new_n13316);
nor_4  g10975(new_n13324, new_n13323, new_n13320);
not_3  g10976(new_n13325, new_n13213);
xnor_3 g10977(new_n13326, new_n13227, new_n13325);
nor_4  g10978(new_n13327, new_n13326, new_n4781);
not_3  g10979(new_n13328, new_n13327);
not_3  g10980(new_n13329, new_n13225);
xnor_3 g10981(new_n13330, new_n13329, new_n13216);
nor_4  g10982(new_n13331, new_n13330, new_n4792);
not_3  g10983(new_n13332, new_n13331);
not_3  g10984(new_n13333_1, new_n13330);
nor_4  g10985(new_n13334, new_n13333_1, new_n4786);
nor_4  g10986(new_n13335, new_n13334, new_n13331);
nor_4  g10987(new_n13336, new_n13218, new_n13217);
xor_3  g10988(new_n13337, new_n13336, new_n13223);
not_3  g10989(new_n13338_1, new_n13337);
nand_4 g10990(new_n13339, new_n13338_1, new_n4811);
xnor_3 g10991(new_n13340, new_n13337, new_n4811);
xor_3  g10992(new_n13341, n8581, n3618);
nand_4 g10993(new_n13342, new_n13341, new_n4841);
nor_4  g10994(new_n13343, new_n13220, new_n13219);
xnor_3 g10995(new_n13344, new_n13343, new_n13221);
nand_4 g10996(new_n13345, new_n13344, new_n13342);
not_3  g10997(new_n13346, new_n13345);
nor_4  g10998(new_n13347, new_n13344, new_n13342);
nor_4  g10999(new_n13348, new_n13347, new_n13346);
nand_4 g11000(new_n13349, new_n13348, new_n4797);
nand_4 g11001(new_n13350, new_n13349, new_n13345);
nand_4 g11002(new_n13351, new_n13350, new_n13340);
nand_4 g11003(new_n13352, new_n13351, new_n13339);
nand_4 g11004(new_n13353, new_n13352, new_n13335);
nand_4 g11005(new_n13354, new_n13353, new_n13332);
not_3  g11006(new_n13355, new_n13326);
nor_4  g11007(new_n13356, new_n13355, new_n4743);
nor_4  g11008(new_n13357, new_n13356, new_n13327);
nand_4 g11009(new_n13358, new_n13357, new_n13354);
nand_4 g11010(new_n13359, new_n13358, new_n13328);
nand_4 g11011(new_n13360, new_n13359, new_n13324);
nand_4 g11012(new_n13361, new_n13360, new_n13321);
nand_4 g11013(new_n13362, new_n13361, new_n13315);
nand_4 g11014(new_n13363, new_n13362, new_n13314);
nand_4 g11015(new_n13364, new_n13363, new_n13310);
nand_4 g11016(new_n13365, new_n13364, new_n13308);
nand_4 g11017(new_n13366, new_n13365, new_n13305);
nand_4 g11018(new_n13367_1, new_n13366, new_n13301);
nand_4 g11019(new_n13368, new_n13367_1, new_n13297);
not_3  g11020(new_n13369, new_n13368);
nor_4  g11021(new_n13370, new_n13369, new_n13293);
not_3  g11022(new_n13371, new_n13289);
nor_4  g11023(new_n13372, new_n13288, new_n13241);
nor_4  g11024(new_n13373, new_n13372, new_n13371);
nand_4 g11025(new_n13374, new_n13373, new_n13370);
nand_4 g11026(new_n13375, new_n13374, new_n13289);
nor_4  g11027(new_n13376, n20040, new_n8789);
nor_4  g11028(new_n13377, new_n10420_1, new_n10377);
nor_4  g11029(new_n13378, new_n13377, new_n13376);
not_3  g11030(new_n13379, new_n13378);
xnor_3 g11031(new_n13380, new_n13379, new_n13375);
xnor_3 g11032(new_n13381, new_n13373, new_n13370);
nand_4 g11033(new_n13382, new_n13381, new_n13379);
xnor_3 g11034(new_n13383, new_n13367_1, new_n13297);
nor_4  g11035(new_n13384, new_n13383, new_n10421);
not_3  g11036(new_n13385, new_n13384);
nor_4  g11037(new_n13386, new_n13367_1, new_n13297);
nor_4  g11038(new_n13387, new_n13386, new_n13369);
nor_4  g11039(new_n13388, new_n13387, new_n10422);
nor_4  g11040(new_n13389, new_n13388, new_n13384);
not_3  g11041(new_n13390, new_n10510);
xnor_3 g11042(new_n13391, new_n13365, new_n13305);
nor_4  g11043(new_n13392, new_n13391, new_n13390);
not_3  g11044(new_n13393, new_n13392);
not_3  g11045(new_n13394, new_n13305);
xnor_3 g11046(new_n13395, new_n13365, new_n13394);
nor_4  g11047(new_n13396, new_n13395, new_n10510);
nor_4  g11048(new_n13397, new_n13396, new_n13392);
xnor_3 g11049(new_n13398, new_n13363, new_n13310);
nor_4  g11050(new_n13399, new_n13398, new_n10522);
not_3  g11051(new_n13400, new_n13399);
xnor_3 g11052(new_n13401, new_n13398, new_n10517);
not_3  g11053(new_n13402, new_n13361);
xnor_3 g11054(new_n13403, new_n13402, new_n13315);
nand_4 g11055(new_n13404, new_n13403, new_n10524);
xnor_3 g11056(new_n13405, new_n13403, new_n10527);
xnor_3 g11057(new_n13406, new_n13359, new_n13324);
nor_4  g11058(new_n13407_1, new_n13406, new_n10533);
not_3  g11059(new_n13408, new_n13407_1);
not_3  g11060(new_n13409_1, new_n13324);
xnor_3 g11061(new_n13410, new_n13359, new_n13409_1);
nor_4  g11062(new_n13411, new_n13410, new_n10529);
nor_4  g11063(new_n13412, new_n13411, new_n13407_1);
xnor_3 g11064(new_n13413, new_n13357, new_n13354);
nor_4  g11065(new_n13414, new_n13413, new_n10539);
not_3  g11066(new_n13415, new_n13414);
xnor_3 g11067(new_n13416, new_n13352, new_n13335);
nor_4  g11068(new_n13417, new_n13416, new_n10542);
not_3  g11069(new_n13418, new_n13417);
not_3  g11070(new_n13419_1, new_n13335);
xnor_3 g11071(new_n13420, new_n13352, new_n13419_1);
nor_4  g11072(new_n13421, new_n13420, new_n10541);
nor_4  g11073(new_n13422, new_n13421, new_n13417);
not_3  g11074(new_n13423, new_n13350);
xnor_3 g11075(new_n13424_1, new_n13423, new_n13340);
nand_4 g11076(new_n13425, new_n13424_1, new_n10552);
xnor_3 g11077(new_n13426, new_n13341, new_n4841);
nor_4  g11078(new_n13427, new_n13426, new_n10560);
not_3  g11079(new_n13428, new_n13427);
nor_4  g11080(new_n13429, new_n13428, new_n10558);
xnor_3 g11081(new_n13430, new_n13348, new_n4797);
not_3  g11082(new_n13431, new_n13430);
xor_3  g11083(new_n13432, new_n13428, new_n10565);
nor_4  g11084(new_n13433, new_n13432, new_n13431);
nor_4  g11085(new_n13434, new_n13433, new_n13429);
xnor_3 g11086(new_n13435, new_n13350, new_n13340);
xnor_3 g11087(new_n13436, new_n13435, new_n10552);
nand_4 g11088(new_n13437, new_n13436, new_n13434);
nand_4 g11089(new_n13438, new_n13437, new_n13425);
nand_4 g11090(new_n13439, new_n13438, new_n13422);
nand_4 g11091(new_n13440, new_n13439, new_n13418);
not_3  g11092(new_n13441, new_n13357);
xnor_3 g11093(new_n13442, new_n13441, new_n13354);
nor_4  g11094(new_n13443, new_n13442, new_n10535);
nor_4  g11095(new_n13444, new_n13443, new_n13414);
nand_4 g11096(new_n13445, new_n13444, new_n13440);
nand_4 g11097(new_n13446, new_n13445, new_n13415);
nand_4 g11098(new_n13447, new_n13446, new_n13412);
nand_4 g11099(new_n13448, new_n13447, new_n13408);
nand_4 g11100(new_n13449, new_n13448, new_n13405);
nand_4 g11101(new_n13450, new_n13449, new_n13404);
nand_4 g11102(new_n13451, new_n13450, new_n13401);
nand_4 g11103(new_n13452, new_n13451, new_n13400);
nand_4 g11104(new_n13453_1, new_n13452, new_n13397);
nand_4 g11105(new_n13454, new_n13453_1, new_n13393);
nand_4 g11106(new_n13455, new_n13454, new_n13389);
nand_4 g11107(new_n13456_1, new_n13455, new_n13385);
xnor_3 g11108(new_n13457_1, new_n13381, new_n13378);
nand_4 g11109(new_n13458, new_n13457_1, new_n13456_1);
nand_4 g11110(new_n13459, new_n13458, new_n13382);
not_3  g11111(new_n13460_1, new_n13459);
xnor_3 g11112(n1527, new_n13460_1, new_n13380);
not_3  g11113(new_n13462, n23463);
xor_3  g11114(new_n13463, n25345, new_n13462);
nand_4 g11115(new_n13464, n13074, new_n6385_1);
xor_3  g11116(new_n13465, n13074, new_n6385_1);
nand_4 g11117(new_n13466, new_n7988, n10739);
not_3  g11118(new_n13467, n10739);
xor_3  g11119(new_n13468, n13490, new_n13467);
not_3  g11120(new_n13469, n22660);
nand_4 g11121(new_n13470, new_n13469, n21753);
xor_3  g11122(new_n13471, n22660, new_n2354);
nor_4  g11123(new_n13472, new_n2356, n1777);
not_3  g11124(new_n13473, new_n13472);
xor_3  g11125(new_n13474, n21832, new_n6391);
nor_4  g11126(new_n13475, new_n2361_1, n8745);
not_3  g11127(new_n13476, new_n13475);
nor_4  g11128(new_n13477_1, n16223, new_n6401);
nor_4  g11129(new_n13478, new_n11726, new_n11720);
nor_4  g11130(new_n13479, new_n13478, new_n13477_1);
xor_3  g11131(new_n13480, n26913, new_n6395);
nand_4 g11132(new_n13481, new_n13480, new_n13479);
nand_4 g11133(new_n13482, new_n13481, new_n13476);
nand_4 g11134(new_n13483, new_n13482, new_n13474);
nand_4 g11135(new_n13484_1, new_n13483, new_n13473);
nand_4 g11136(new_n13485, new_n13484_1, new_n13471);
nand_4 g11137(new_n13486_1, new_n13485, new_n13470);
nand_4 g11138(new_n13487_1, new_n13486_1, new_n13468);
nand_4 g11139(new_n13488, new_n13487_1, new_n13466);
nand_4 g11140(new_n13489, new_n13488, new_n13465);
nand_4 g11141(new_n13490_1, new_n13489, new_n13464);
xnor_3 g11142(new_n13491, new_n13490_1, new_n13463);
nor_4  g11143(new_n13492, new_n13491, new_n9323_1);
not_3  g11144(new_n13493, new_n13491);
nor_4  g11145(new_n13494_1, new_n13493, new_n9322);
nor_4  g11146(new_n13495, new_n13494_1, new_n13492);
xnor_3 g11147(new_n13496, new_n13488, new_n13465);
not_3  g11148(new_n13497, new_n13496);
nor_4  g11149(new_n13498, new_n13497, new_n9328);
nor_4  g11150(new_n13499, new_n13496, new_n9329);
nor_4  g11151(new_n13500_1, new_n13499, new_n13498);
xnor_3 g11152(new_n13501_1, new_n13486_1, new_n13468);
nand_4 g11153(new_n13502, new_n13501_1, new_n9335);
xnor_3 g11154(new_n13503, new_n13501_1, new_n9334);
xnor_3 g11155(new_n13504, new_n13484_1, new_n13471);
nand_4 g11156(new_n13505, new_n13504, new_n9343);
not_3  g11157(new_n13506_1, new_n13504);
xnor_3 g11158(new_n13507, new_n13506_1, new_n9343);
not_3  g11159(new_n13508, new_n13474);
xor_3  g11160(new_n13509, new_n13482, new_n13508);
nand_4 g11161(new_n13510, new_n13509, new_n9351);
xor_3  g11162(new_n13511, new_n13482, new_n13474);
xnor_3 g11163(new_n13512, new_n13511, new_n9351);
xnor_3 g11164(new_n13513, new_n13480, new_n13479);
nand_4 g11165(new_n13514, new_n13513, new_n9355);
nand_4 g11166(new_n13515, new_n11727, new_n9360);
nand_4 g11167(new_n13516, new_n11740, new_n11728);
nand_4 g11168(new_n13517, new_n13516, new_n13515);
not_3  g11169(new_n13518, new_n13514);
nor_4  g11170(new_n13519, new_n13513, new_n9355);
nor_4  g11171(new_n13520, new_n13519, new_n13518);
nand_4 g11172(new_n13521, new_n13520, new_n13517);
nand_4 g11173(new_n13522, new_n13521, new_n13514);
nand_4 g11174(new_n13523, new_n13522, new_n13512);
nand_4 g11175(new_n13524, new_n13523, new_n13510);
nand_4 g11176(new_n13525, new_n13524, new_n13507);
nand_4 g11177(new_n13526, new_n13525, new_n13505);
nand_4 g11178(new_n13527, new_n13526, new_n13503);
nand_4 g11179(new_n13528, new_n13527, new_n13502);
nand_4 g11180(new_n13529, new_n13528, new_n13500_1);
not_3  g11181(new_n13530, new_n13529);
nor_4  g11182(new_n13531, new_n13530, new_n13498);
xor_3  g11183(n1580, new_n13531, new_n13495);
xor_3  g11184(new_n13533, n18962, new_n3506_1);
nor_4  g11185(new_n13534, new_n13533, new_n8758);
nor_4  g11186(new_n13535, new_n8997, n12315);
not_3  g11187(new_n13536, n3952);
xor_3  g11188(new_n13537, n10158, new_n13536);
not_3  g11189(new_n13538, new_n13537);
xor_3  g11190(new_n13539, new_n13538, new_n13535);
xnor_3 g11191(new_n13540, new_n13539, new_n13534);
xor_3  g11192(n1586, new_n13540, new_n8765);
not_3  g11193(new_n13542, n1483);
xor_3  g11194(new_n13543, n19539, new_n13542);
not_3  g11195(new_n13544, new_n13543);
not_3  g11196(new_n13545, n8194);
nor_4  g11197(new_n13546, n24093, new_n13545);
xor_3  g11198(new_n13547, n24093, new_n13545);
not_3  g11199(new_n13548_1, n23035);
nand_4 g11200(new_n13549_1, n23657, new_n13548_1);
xor_3  g11201(new_n13550, n23657, new_n13548_1);
nand_4 g11202(new_n13551_1, n16911, new_n7525);
nand_4 g11203(new_n13552, new_n7559, new_n7526);
nand_4 g11204(new_n13553, new_n13552, new_n13551_1);
nand_4 g11205(new_n13554, new_n13553, new_n13550);
nand_4 g11206(new_n13555, new_n13554, new_n13549_1);
nand_4 g11207(new_n13556, new_n13555, new_n13547);
not_3  g11208(new_n13557, new_n13556);
nor_4  g11209(new_n13558, new_n13557, new_n13546);
and_4  g11210(new_n13559, new_n13558, new_n13544);
nor_4  g11211(new_n13560, new_n13558, new_n13544);
nor_4  g11212(new_n13561, new_n13560, new_n13559);
not_3  g11213(new_n13562, new_n13561);
xor_3  g11214(new_n13563, n25494, new_n9766);
nor_4  g11215(new_n13564, n10117, new_n9770);
xor_3  g11216(new_n13565, n10117, new_n9770);
not_3  g11217(new_n13566, n13460);
nand_4 g11218(new_n13567, n22335, new_n13566);
xor_3  g11219(new_n13568, n22335, new_n13566);
not_3  g11220(new_n13569, n6104);
nand_4 g11221(new_n13570, n24048, new_n13569);
nand_4 g11222(new_n13571, new_n3693, n1525);
nand_4 g11223(new_n13572, new_n5285, new_n5261);
nand_4 g11224(new_n13573, new_n13572, new_n13571);
xor_3  g11225(new_n13574, n24048, new_n13569);
nand_4 g11226(new_n13575, new_n13574, new_n13573);
nand_4 g11227(new_n13576, new_n13575, new_n13570);
nand_4 g11228(new_n13577, new_n13576, new_n13568);
nand_4 g11229(new_n13578, new_n13577, new_n13567);
nand_4 g11230(new_n13579, new_n13578, new_n13565);
not_3  g11231(new_n13580, new_n13579);
nor_4  g11232(new_n13581, new_n13580, new_n13564);
xor_3  g11233(new_n13582, new_n13581, new_n13563);
not_3  g11234(new_n13583, new_n13582);
not_3  g11235(new_n13584, n25296);
xor_3  g11236(new_n13585, new_n13584, n23717);
not_3  g11237(new_n13586, new_n13585);
not_3  g11238(new_n13587, n7788);
nor_4  g11239(new_n13588, n20013, new_n13587);
xor_3  g11240(new_n13589, n20013, new_n13587);
not_3  g11241(new_n13590, n1320);
nand_4 g11242(new_n13591, n5443, new_n13590);
xor_3  g11243(new_n13592, n5443, new_n13590);
nand_4 g11244(new_n13593, new_n7519, n18584);
nand_4 g11245(new_n13594, new_n7523, new_n7520);
nand_4 g11246(new_n13595, new_n13594, new_n13593);
nand_4 g11247(new_n13596, new_n13595, new_n13592);
nand_4 g11248(new_n13597, new_n13596, new_n13591);
nand_4 g11249(new_n13598, new_n13597, new_n13589);
not_3  g11250(new_n13599, new_n13598);
nor_4  g11251(new_n13600, new_n13599, new_n13588);
xor_3  g11252(new_n13601, new_n13600, new_n13586);
nor_4  g11253(new_n13602_1, new_n13601, new_n13583);
not_3  g11254(new_n13603, new_n13601);
nor_4  g11255(new_n13604, new_n13603, new_n13582);
nor_4  g11256(new_n13605, new_n13604, new_n13602_1);
xnor_3 g11257(new_n13606, new_n13578, new_n13565);
nor_4  g11258(new_n13607, new_n13597, new_n13589);
nor_4  g11259(new_n13608, new_n13607, new_n13599);
not_3  g11260(new_n13609, new_n13608);
nor_4  g11261(new_n13610, new_n13609, new_n13606);
not_3  g11262(new_n13611, new_n13610);
not_3  g11263(new_n13612, new_n13606);
xnor_3 g11264(new_n13613, new_n13608, new_n13612);
not_3  g11265(new_n13614, new_n13613);
xnor_3 g11266(new_n13615, new_n13576, new_n13568);
not_3  g11267(new_n13616, new_n13615);
xnor_3 g11268(new_n13617, new_n13595, new_n13592);
not_3  g11269(new_n13618, new_n13617);
nor_4  g11270(new_n13619, new_n13618, new_n13616);
xnor_3 g11271(new_n13620, new_n13617, new_n13615);
not_3  g11272(new_n13621, new_n13574);
xnor_3 g11273(new_n13622, new_n13621, new_n13573);
not_3  g11274(new_n13623, new_n13622);
nor_4  g11275(new_n13624, new_n13623, new_n7524_1);
not_3  g11276(new_n13625, new_n13624);
not_3  g11277(new_n13626_1, new_n7524_1);
nor_4  g11278(new_n13627, new_n13622, new_n13626_1);
nor_4  g11279(new_n13628, new_n13627, new_n13624);
not_3  g11280(new_n13629, new_n5319);
nand_4 g11281(new_n13630, new_n5371, new_n5322);
nand_4 g11282(new_n13631, new_n13630, new_n13629);
nand_4 g11283(new_n13632, new_n13631, new_n13628);
nand_4 g11284(new_n13633, new_n13632, new_n13625);
nor_4  g11285(new_n13634, new_n13633, new_n13620);
nor_4  g11286(new_n13635, new_n13634, new_n13619);
nand_4 g11287(new_n13636, new_n13635, new_n13614);
nand_4 g11288(new_n13637, new_n13636, new_n13611);
xnor_3 g11289(new_n13638, new_n13637, new_n13605);
xnor_3 g11290(new_n13639, new_n13638, new_n13562);
nor_4  g11291(new_n13640, new_n13555, new_n13547);
nor_4  g11292(new_n13641, new_n13640, new_n13557);
xnor_3 g11293(new_n13642, new_n13635, new_n13613);
nor_4  g11294(new_n13643, new_n13642, new_n13641);
not_3  g11295(new_n13644, new_n13643);
not_3  g11296(new_n13645, new_n13641);
xnor_3 g11297(new_n13646, new_n13635, new_n13614);
nor_4  g11298(new_n13647, new_n13646, new_n13645);
nor_4  g11299(new_n13648, new_n13647, new_n13643);
not_3  g11300(new_n13649, new_n13550);
xnor_3 g11301(new_n13650, new_n13553, new_n13649);
xnor_3 g11302(new_n13651, new_n13633, new_n13620);
nor_4  g11303(new_n13652, new_n13651, new_n13650);
not_3  g11304(new_n13653, new_n13652);
not_3  g11305(new_n13654, new_n13650);
not_3  g11306(new_n13655, new_n13620);
xnor_3 g11307(new_n13656, new_n13633, new_n13655);
nor_4  g11308(new_n13657, new_n13656, new_n13654);
nor_4  g11309(new_n13658, new_n13657, new_n13652);
not_3  g11310(new_n13659, new_n7560);
xnor_3 g11311(new_n13660, new_n13631, new_n13628);
not_3  g11312(new_n13661, new_n13660);
nor_4  g11313(new_n13662, new_n13661, new_n13659);
not_3  g11314(new_n13663, new_n13662);
nor_4  g11315(new_n13664, new_n13660, new_n7560);
nor_4  g11316(new_n13665, new_n13664, new_n13662);
nor_4  g11317(new_n13666, new_n7627, new_n5373);
not_3  g11318(new_n13667, new_n13666);
nor_4  g11319(new_n13668_1, new_n7637, new_n5377);
not_3  g11320(new_n13669, new_n13668_1);
nor_4  g11321(new_n13670, new_n7636, new_n5381);
nor_4  g11322(new_n13671, new_n13670, new_n13668_1);
nor_4  g11323(new_n13672, new_n7647_1, new_n5384);
not_3  g11324(new_n13673, new_n13672);
nor_4  g11325(new_n13674, new_n7653, new_n5389);
not_3  g11326(new_n13675, new_n13674);
not_3  g11327(new_n13676, new_n7653);
nor_4  g11328(new_n13677_1, new_n13676, new_n5388);
nor_4  g11329(new_n13678, new_n13677_1, new_n13674);
nor_4  g11330(new_n13679, new_n7662, new_n5397);
nor_4  g11331(new_n13680, new_n13679, new_n7665);
not_3  g11332(new_n13681, new_n13680);
not_3  g11333(new_n13682, new_n5403_1);
not_3  g11334(new_n13683_1, new_n7665);
not_3  g11335(new_n13684, new_n13679);
xor_3  g11336(new_n13685, new_n13684, new_n13683_1);
nand_4 g11337(new_n13686, new_n13685, new_n13682);
nand_4 g11338(new_n13687, new_n13686, new_n13681);
nand_4 g11339(new_n13688, new_n13687, new_n13678);
nand_4 g11340(new_n13689, new_n13688, new_n13675);
not_3  g11341(new_n13690, new_n7647_1);
nor_4  g11342(new_n13691, new_n13690, new_n5410);
nor_4  g11343(new_n13692, new_n13691, new_n13672);
nand_4 g11344(new_n13693, new_n13692, new_n13689);
nand_4 g11345(new_n13694, new_n13693, new_n13673);
nand_4 g11346(new_n13695, new_n13694, new_n13671);
nand_4 g11347(new_n13696, new_n13695, new_n13669);
nor_4  g11348(new_n13697, new_n7626, new_n5372);
nor_4  g11349(new_n13698, new_n13697, new_n13666);
nand_4 g11350(new_n13699, new_n13698, new_n13696);
nand_4 g11351(new_n13700, new_n13699, new_n13667);
nand_4 g11352(new_n13701, new_n13700, new_n13665);
nand_4 g11353(new_n13702, new_n13701, new_n13663);
nand_4 g11354(new_n13703, new_n13702, new_n13658);
nand_4 g11355(new_n13704, new_n13703, new_n13653);
nand_4 g11356(new_n13705, new_n13704, new_n13648);
nand_4 g11357(new_n13706, new_n13705, new_n13644);
nor_4  g11358(new_n13707, new_n13706, new_n13639);
and_4  g11359(new_n13708_1, new_n13706, new_n13639);
nor_4  g11360(n1590, new_n13708_1, new_n13707);
not_3  g11361(new_n13710_1, new_n9012_1);
xor_3  g11362(n1602, new_n13710_1, new_n8988);
xor_3  g11363(n1634, new_n2979_1, new_n2916);
not_3  g11364(new_n13713, new_n13704);
xor_3  g11365(n1636, new_n13713, new_n13648);
nor_4  g11366(new_n13715, n10514, n4514);
xor_3  g11367(new_n13716, n10514, n4514);
not_3  g11368(new_n13717, new_n13716);
nor_4  g11369(new_n13718, n18649, n3984);
xor_3  g11370(new_n13719_1, n18649, n3984);
nand_4 g11371(new_n13720, n19652, n6218);
not_3  g11372(new_n13721, new_n13720);
nor_4  g11373(new_n13722_1, n19652, n6218);
not_3  g11374(new_n13723, n3366);
not_3  g11375(new_n13724, n20470);
nand_4 g11376(new_n13725, new_n13724, new_n13723);
nand_4 g11377(new_n13726, new_n13136, new_n13128);
nand_4 g11378(new_n13727, new_n13726, new_n13725);
nor_4  g11379(new_n13728, new_n13727, new_n13722_1);
nor_4  g11380(new_n13729, new_n13728, new_n13721);
nand_4 g11381(new_n13730, new_n13729, new_n13719_1);
not_3  g11382(new_n13731, new_n13730);
nor_4  g11383(new_n13732, new_n13731, new_n13718);
nor_4  g11384(new_n13733, new_n13732, new_n13717);
nor_4  g11385(new_n13734, new_n13733, new_n13715);
not_3  g11386(new_n13735, new_n13734);
xor_3  g11387(new_n13736, n18880, n2978);
not_3  g11388(new_n13737, new_n13736);
nor_4  g11389(new_n13738, n25475, n23697);
nor_4  g11390(new_n13739, new_n7976, new_n7933);
nor_4  g11391(new_n13740, new_n13739, new_n13738);
xnor_3 g11392(new_n13741, new_n13740, new_n13737);
nand_4 g11393(new_n13742, new_n13741, n20040);
not_3  g11394(new_n13743, new_n13742);
nor_4  g11395(new_n13744, new_n13741, n20040);
nor_4  g11396(new_n13745, new_n13744, new_n13743);
nand_4 g11397(new_n13746, new_n7977, n19531);
not_3  g11398(new_n13747, new_n13746);
nor_4  g11399(new_n13748, new_n7977, n19531);
nor_4  g11400(new_n13749, new_n13748, new_n13747);
nor_4  g11401(new_n13750, new_n7982, n18345);
xnor_3 g11402(new_n13751, new_n7982, n18345);
nor_4  g11403(new_n13752, new_n7989, n13190);
xnor_3 g11404(new_n13753, new_n7989, n13190);
nand_4 g11405(new_n13754_1, new_n7995, n3460);
nand_4 g11406(new_n13755, new_n7997, n5226);
nand_4 g11407(new_n13756, new_n11467, new_n11447);
nand_4 g11408(new_n13757, new_n13756, new_n13755);
xnor_3 g11409(new_n13758, new_n7995, new_n10386);
nand_4 g11410(new_n13759, new_n13758, new_n13757);
nand_4 g11411(new_n13760, new_n13759, new_n13754_1);
nor_4  g11412(new_n13761, new_n13760, new_n13753);
nor_4  g11413(new_n13762, new_n13761, new_n13752);
nor_4  g11414(new_n13763, new_n13762, new_n13751);
nor_4  g11415(new_n13764_1, new_n13763, new_n13750);
nand_4 g11416(new_n13765, new_n13764_1, new_n13749);
nand_4 g11417(new_n13766, new_n13765, new_n13746);
nand_4 g11418(new_n13767, new_n13766, new_n13745);
nand_4 g11419(new_n13768, new_n13767, new_n13742);
nor_4  g11420(new_n13769, n18880, n2978);
nor_4  g11421(new_n13770, new_n13740, new_n13737);
nor_4  g11422(new_n13771, new_n13770, new_n13769);
nor_4  g11423(new_n13772, new_n13771, new_n13768);
nand_4 g11424(new_n13773, new_n13771, new_n13768);
not_3  g11425(new_n13774, new_n13773);
nor_4  g11426(new_n13775_1, new_n13774, new_n13772);
not_3  g11427(new_n13776, new_n11445);
nor_4  g11428(new_n13777, new_n13776, n19575);
not_3  g11429(new_n13778, new_n13777);
nor_4  g11430(new_n13779, new_n13778, n26512);
not_3  g11431(new_n13780, new_n13779);
nor_4  g11432(new_n13781_1, new_n13780, n26191);
not_3  g11433(new_n13782, new_n13781_1);
nor_4  g11434(new_n13783_1, new_n13782, n5386);
not_3  g11435(new_n13784, new_n13783_1);
nor_4  g11436(new_n13785, new_n13784, n17037);
not_3  g11437(new_n13786, new_n13785);
nor_4  g11438(new_n13787, new_n13786, n7569);
not_3  g11439(new_n13788, new_n13787);
nor_4  g11440(new_n13789, new_n13788, new_n13775_1);
not_3  g11441(new_n13790, new_n13775_1);
nor_4  g11442(new_n13791, new_n13787, new_n13790);
nor_4  g11443(new_n13792, new_n13791, new_n13789);
xnor_3 g11444(new_n13793, new_n13766, new_n13745);
not_3  g11445(new_n13794, new_n13793);
not_3  g11446(new_n13795, n7569);
xor_3  g11447(new_n13796, new_n13785, new_n13795);
nor_4  g11448(new_n13797, new_n13796, new_n13794);
not_3  g11449(new_n13798_1, new_n13797);
not_3  g11450(new_n13799, new_n13796);
nor_4  g11451(new_n13800, new_n13799, new_n13793);
nor_4  g11452(new_n13801, new_n13800, new_n13797);
xnor_3 g11453(new_n13802, new_n13764_1, new_n13749);
not_3  g11454(new_n13803, new_n13802);
not_3  g11455(new_n13804, n17037);
xor_3  g11456(new_n13805, new_n13783_1, new_n13804);
nor_4  g11457(new_n13806, new_n13805, new_n13803);
not_3  g11458(new_n13807, new_n13806);
not_3  g11459(new_n13808, new_n13805);
nor_4  g11460(new_n13809, new_n13808, new_n13802);
nor_4  g11461(new_n13810, new_n13809, new_n13806);
xnor_3 g11462(new_n13811, new_n13762, new_n13751);
not_3  g11463(new_n13812, n5386);
xor_3  g11464(new_n13813, new_n13781_1, new_n13812);
nor_4  g11465(new_n13814, new_n13813, new_n13811);
not_3  g11466(new_n13815, new_n13814);
not_3  g11467(new_n13816, new_n13811);
not_3  g11468(new_n13817, new_n13813);
nor_4  g11469(new_n13818, new_n13817, new_n13816);
nor_4  g11470(new_n13819, new_n13818, new_n13814);
xnor_3 g11471(new_n13820, new_n13760, new_n13753);
not_3  g11472(new_n13821, n26191);
xor_3  g11473(new_n13822, new_n13779, new_n13821);
nor_4  g11474(new_n13823, new_n13822, new_n13820);
not_3  g11475(new_n13824, new_n13823);
not_3  g11476(new_n13825, n26512);
xor_3  g11477(new_n13826, new_n13777, new_n13825);
not_3  g11478(new_n13827, new_n13826);
xnor_3 g11479(new_n13828, new_n13758, new_n13757);
nor_4  g11480(new_n13829, new_n13828, new_n13827);
xnor_3 g11481(new_n13830, new_n13828, new_n13827);
nor_4  g11482(new_n13831, new_n11471, new_n11446);
nor_4  g11483(new_n13832, new_n11513, new_n13831);
not_3  g11484(new_n13833, new_n13832);
nor_4  g11485(new_n13834, new_n13833, new_n13830);
nor_4  g11486(new_n13835_1, new_n13834, new_n13829);
not_3  g11487(new_n13836, new_n13820);
not_3  g11488(new_n13837, new_n13822);
nor_4  g11489(new_n13838, new_n13837, new_n13836);
nor_4  g11490(new_n13839, new_n13838, new_n13823);
nand_4 g11491(new_n13840, new_n13839, new_n13835_1);
nand_4 g11492(new_n13841, new_n13840, new_n13824);
nand_4 g11493(new_n13842, new_n13841, new_n13819);
nand_4 g11494(new_n13843, new_n13842, new_n13815);
nand_4 g11495(new_n13844, new_n13843, new_n13810);
nand_4 g11496(new_n13845, new_n13844, new_n13807);
nand_4 g11497(new_n13846, new_n13845, new_n13801);
nand_4 g11498(new_n13847, new_n13846, new_n13798_1);
not_3  g11499(new_n13848, new_n13847);
xnor_3 g11500(new_n13849, new_n13848, new_n13792);
xnor_3 g11501(new_n13850_1, new_n13849, new_n13735);
not_3  g11502(new_n13851_1, new_n13846);
nor_4  g11503(new_n13852, new_n13845, new_n13801);
nor_4  g11504(new_n13853, new_n13852, new_n13851_1);
xor_3  g11505(new_n13854, new_n13732, new_n13717);
not_3  g11506(new_n13855, new_n13854);
nand_4 g11507(new_n13856, new_n13855, new_n13853);
xnor_3 g11508(new_n13857, new_n13854, new_n13853);
not_3  g11509(new_n13858, new_n13844);
nor_4  g11510(new_n13859, new_n13843, new_n13810);
nor_4  g11511(new_n13860, new_n13859, new_n13858);
xnor_3 g11512(new_n13861, new_n13729, new_n13719_1);
nand_4 g11513(new_n13862, new_n13861, new_n13860);
not_3  g11514(new_n13863, new_n13861);
xnor_3 g11515(new_n13864, new_n13863, new_n13860);
not_3  g11516(new_n13865, new_n13842);
nor_4  g11517(new_n13866, new_n13841, new_n13819);
nor_4  g11518(new_n13867, new_n13866, new_n13865);
nor_4  g11519(new_n13868, new_n13722_1, new_n13721);
xnor_3 g11520(new_n13869, new_n13868, new_n13727);
nand_4 g11521(new_n13870, new_n13869, new_n13867);
not_3  g11522(new_n13871, new_n13869);
xnor_3 g11523(new_n13872, new_n13871, new_n13867);
xnor_3 g11524(new_n13873, new_n13839, new_n13835_1);
nor_4  g11525(new_n13874, new_n13873, new_n13138);
not_3  g11526(new_n13875, new_n13874);
not_3  g11527(new_n13876, new_n13873);
nor_4  g11528(new_n13877, new_n13876, new_n13137_1);
nor_4  g11529(new_n13878, new_n13877, new_n13874);
xnor_3 g11530(new_n13879, new_n13832, new_n13830);
not_3  g11531(new_n13880, new_n13879);
nor_4  g11532(new_n13881, new_n13880, new_n13155);
nor_4  g11533(new_n13882, new_n13879, new_n13156);
nor_4  g11534(new_n13883, new_n11514, new_n11440);
nor_4  g11535(new_n13884, new_n11548_1, new_n11515_1);
nor_4  g11536(new_n13885, new_n13884, new_n13883);
nor_4  g11537(new_n13886, new_n13885, new_n13882);
nor_4  g11538(new_n13887, new_n13886, new_n13881);
nand_4 g11539(new_n13888, new_n13887, new_n13878);
nand_4 g11540(new_n13889, new_n13888, new_n13875);
nand_4 g11541(new_n13890, new_n13889, new_n13872);
nand_4 g11542(new_n13891, new_n13890, new_n13870);
nand_4 g11543(new_n13892, new_n13891, new_n13864);
nand_4 g11544(new_n13893, new_n13892, new_n13862);
nand_4 g11545(new_n13894, new_n13893, new_n13857);
nand_4 g11546(new_n13895, new_n13894, new_n13856);
xnor_3 g11547(n1684, new_n13895, new_n13850_1);
not_3  g11548(new_n13897, n4514);
nor_4  g11549(new_n13898, new_n7255, new_n13897);
not_3  g11550(new_n13899, new_n13898);
nor_4  g11551(new_n13900, new_n7260, n4514);
nor_4  g11552(new_n13901, new_n7263, n3984);
not_3  g11553(new_n13902, new_n13901);
not_3  g11554(new_n13903, n3984);
nor_4  g11555(new_n13904, new_n7266, new_n13903);
nor_4  g11556(new_n13905, new_n13904, new_n13901);
not_3  g11557(new_n13906, new_n13905);
not_3  g11558(new_n13907, n19652);
not_3  g11559(new_n13908, new_n7270);
nand_4 g11560(new_n13909, new_n13908, new_n13907);
not_3  g11561(new_n13910, new_n13909);
xor_3  g11562(new_n13911, new_n13908, n19652);
nor_4  g11563(new_n13912_1, new_n7276, n3366);
xnor_3 g11564(new_n13913, new_n7276, n3366);
nor_4  g11565(new_n13914_1, new_n4445, n26565);
not_3  g11566(new_n13915, n26565);
nor_4  g11567(new_n13916, new_n7280_1, new_n13915);
nor_4  g11568(new_n13917, new_n13916, new_n13914_1);
xnor_3 g11569(new_n13918, new_n4440, n15424);
nor_4  g11570(new_n13919, new_n13918, n3959);
not_3  g11571(new_n13920, new_n13919);
not_3  g11572(new_n13921, n3959);
nor_4  g11573(new_n13922_1, new_n4448, new_n13921);
nor_4  g11574(new_n13923_1, new_n13922_1, new_n13919);
nor_4  g11575(new_n13924, new_n4454, n11566);
not_3  g11576(new_n13925, new_n13924);
not_3  g11577(new_n13926, n11566);
nor_4  g11578(new_n13927, new_n4455, new_n13926);
nor_4  g11579(new_n13928, new_n13927, new_n13924);
nor_4  g11580(new_n13929, new_n4465, n26744);
not_3  g11581(new_n13930, new_n13929);
not_3  g11582(new_n13931, n26744);
not_3  g11583(new_n13932, new_n4465);
nor_4  g11584(new_n13933, new_n13932, new_n13931);
nor_4  g11585(new_n13934, new_n13933, new_n13929);
not_3  g11586(new_n13935, n26625);
nand_4 g11587(new_n13936, new_n4471, new_n13935);
nand_4 g11588(new_n13937, n19922, n14230);
not_3  g11589(new_n13938, new_n13936);
nor_4  g11590(new_n13939, new_n4471, new_n13935);
nor_4  g11591(new_n13940, new_n13939, new_n13938);
nand_4 g11592(new_n13941, new_n13940, new_n13937);
nand_4 g11593(new_n13942, new_n13941, new_n13936);
nand_4 g11594(new_n13943, new_n13942, new_n13934);
nand_4 g11595(new_n13944, new_n13943, new_n13930);
nand_4 g11596(new_n13945, new_n13944, new_n13928);
nand_4 g11597(new_n13946, new_n13945, new_n13925);
nand_4 g11598(new_n13947, new_n13946, new_n13923_1);
nand_4 g11599(new_n13948, new_n13947, new_n13920);
nand_4 g11600(new_n13949, new_n13948, new_n13917);
not_3  g11601(new_n13950, new_n13949);
nor_4  g11602(new_n13951_1, new_n13950, new_n13914_1);
nor_4  g11603(new_n13952, new_n13951_1, new_n13913);
nor_4  g11604(new_n13953, new_n13952, new_n13912_1);
nor_4  g11605(new_n13954, new_n13953, new_n13911);
nor_4  g11606(new_n13955, new_n13954, new_n13910);
nor_4  g11607(new_n13956, new_n13955, new_n13906);
not_3  g11608(new_n13957, new_n13956);
nand_4 g11609(new_n13958, new_n13957, new_n13902);
nor_4  g11610(new_n13959, new_n13958, new_n13900);
nor_4  g11611(new_n13960, new_n13959, new_n7258);
nand_4 g11612(new_n13961, new_n13960, new_n13899);
not_3  g11613(new_n13962, new_n13961);
not_3  g11614(new_n13963, new_n13911);
not_3  g11615(new_n13964, new_n13912_1);
nor_4  g11616(new_n13965, new_n7273, new_n13723);
nor_4  g11617(new_n13966, new_n13965, new_n13912_1);
not_3  g11618(new_n13967, new_n13951_1);
nand_4 g11619(new_n13968, new_n13967, new_n13966);
nand_4 g11620(new_n13969, new_n13968, new_n13964);
nand_4 g11621(new_n13970, new_n13969, new_n13963);
nand_4 g11622(new_n13971, new_n13970, new_n13909);
nor_4  g11623(new_n13972, new_n13971, new_n13905);
nor_4  g11624(new_n13973, new_n13972, new_n13956);
nand_4 g11625(new_n13974, new_n13973, n13026);
not_3  g11626(new_n13975, n13026);
xnor_3 g11627(new_n13976, new_n13955, new_n13906);
nand_4 g11628(new_n13977, new_n13976, new_n13975);
nor_4  g11629(new_n13978, new_n13969, new_n13963);
nor_4  g11630(new_n13979, new_n13978, new_n13954);
nand_4 g11631(new_n13980, new_n13979, n2175);
not_3  g11632(new_n13981, n2175);
xnor_3 g11633(new_n13982, new_n13953, new_n13911);
nand_4 g11634(new_n13983, new_n13982, new_n13981);
xnor_3 g11635(new_n13984, new_n13951_1, new_n13913);
not_3  g11636(new_n13985, new_n13984);
nand_4 g11637(new_n13986, new_n13985, n752);
nand_4 g11638(new_n13987, new_n13984, new_n13076);
not_3  g11639(new_n13988, n1611);
xnor_3 g11640(new_n13989, new_n13948, new_n13917);
nor_4  g11641(new_n13990, new_n13989, new_n13988);
not_3  g11642(new_n13991, new_n13990);
not_3  g11643(new_n13992, new_n13989);
nor_4  g11644(new_n13993, new_n13992, n1611);
not_3  g11645(new_n13994, new_n13993);
not_3  g11646(new_n13995, new_n13947);
nor_4  g11647(new_n13996, new_n13946, new_n13923_1);
nor_4  g11648(new_n13997, new_n13996, new_n13995);
nand_4 g11649(new_n13998, new_n13997, n25094);
not_3  g11650(new_n13999, new_n13997);
nand_4 g11651(new_n14000, new_n13999, new_n13077);
xnor_3 g11652(new_n14001, new_n13944, new_n13928);
not_3  g11653(new_n14002, new_n14001);
nand_4 g11654(new_n14003, new_n14002, n21538);
not_3  g11655(new_n14004_1, n21538);
nand_4 g11656(new_n14005, new_n14001, new_n14004_1);
xnor_3 g11657(new_n14006, new_n13942, new_n13934);
not_3  g11658(new_n14007, new_n14006);
nand_4 g11659(new_n14008, new_n14007, n5131);
nand_4 g11660(new_n14009, new_n14006, new_n13078);
xnor_3 g11661(new_n14010, new_n13940, new_n13937);
nor_4  g11662(new_n14011, new_n14010, new_n13111);
not_3  g11663(new_n14012, new_n14011);
nand_4 g11664(new_n14013, new_n14010, new_n13111);
xor_3  g11665(new_n14014, n19922, n14230);
nor_4  g11666(new_n14015, new_n14014, new_n13106);
nand_4 g11667(new_n14016, new_n14015, new_n14013);
nand_4 g11668(new_n14017, new_n14016, new_n14012);
nand_4 g11669(new_n14018, new_n14017, new_n14009);
nand_4 g11670(new_n14019, new_n14018, new_n14008);
nand_4 g11671(new_n14020, new_n14019, new_n14005);
nand_4 g11672(new_n14021, new_n14020, new_n14003);
nand_4 g11673(new_n14022, new_n14021, new_n14000);
nand_4 g11674(new_n14023, new_n14022, new_n13998);
nand_4 g11675(new_n14024, new_n14023, new_n13994);
nand_4 g11676(new_n14025, new_n14024, new_n13991);
nand_4 g11677(new_n14026, new_n14025, new_n13987);
nand_4 g11678(new_n14027, new_n14026, new_n13986);
nand_4 g11679(new_n14028, new_n14027, new_n13983);
nand_4 g11680(new_n14029, new_n14028, new_n13980);
nand_4 g11681(new_n14030, new_n14029, new_n13977);
nand_4 g11682(new_n14031, new_n14030, new_n13974);
nor_4  g11683(new_n14032, new_n14031, n23912);
nand_4 g11684(new_n14033, new_n14031, n23912);
not_3  g11685(new_n14034, new_n14033);
nor_4  g11686(new_n14035, new_n13900, new_n13898);
not_3  g11687(new_n14036_1, new_n14035);
xnor_3 g11688(new_n14037, new_n14036_1, new_n13958);
nor_4  g11689(new_n14038, new_n14037, new_n14034);
nor_4  g11690(new_n14039, new_n14038, new_n14032);
nor_4  g11691(new_n14040, new_n14039, new_n13962);
nor_4  g11692(new_n14041, new_n5043, n15766);
not_3  g11693(new_n14042, new_n14041);
not_3  g11694(new_n14043, n15766);
nor_4  g11695(new_n14044, new_n5038, new_n14043);
nor_4  g11696(new_n14045, new_n14044, new_n14041);
nor_4  g11697(new_n14046, new_n5048, n25629);
not_3  g11698(new_n14047, new_n14046);
nor_4  g11699(new_n14048, new_n5051, new_n7394);
nor_4  g11700(new_n14049, new_n14048, new_n14046);
nor_4  g11701(new_n14050, new_n5057, n7692);
not_3  g11702(new_n14051, new_n14050);
not_3  g11703(new_n14052, n7692);
xnor_3 g11704(new_n14053, new_n5026_1, new_n5015);
nor_4  g11705(new_n14054, new_n14053, new_n14052);
nor_4  g11706(new_n14055, new_n14054, new_n14050);
nor_4  g11707(new_n14056, new_n5062_1, n23039);
not_3  g11708(new_n14057, new_n14056);
nor_4  g11709(new_n14058, new_n5067, new_n12385);
nor_4  g11710(new_n14059_1, new_n14058, new_n14056);
not_3  g11711(new_n14060, new_n4391);
nand_4 g11712(new_n14061, new_n4424_1, new_n4392);
nand_4 g11713(new_n14062, new_n14061, new_n14060);
nand_4 g11714(new_n14063, new_n14062, new_n14059_1);
nand_4 g11715(new_n14064, new_n14063, new_n14057);
nand_4 g11716(new_n14065, new_n14064, new_n14055);
nand_4 g11717(new_n14066, new_n14065, new_n14051);
nand_4 g11718(new_n14067, new_n14066, new_n14049);
nand_4 g11719(new_n14068, new_n14067, new_n14047);
nand_4 g11720(new_n14069, new_n14068, new_n14045);
nand_4 g11721(new_n14070, new_n14069, new_n14042);
nor_4  g11722(new_n14071_1, new_n14070, new_n5133);
xnor_3 g11723(new_n14072, new_n14070, new_n5125);
not_3  g11724(new_n14073, new_n14072);
xnor_3 g11725(new_n14074, new_n14039, new_n13962);
nand_4 g11726(new_n14075, new_n14074, new_n14073);
xnor_3 g11727(new_n14076, new_n14074, new_n14072);
xnor_3 g11728(new_n14077, new_n14068, new_n14045);
not_3  g11729(new_n14078, new_n14077);
not_3  g11730(new_n14079, n23912);
xnor_3 g11731(new_n14080, new_n14031, new_n14079);
xnor_3 g11732(new_n14081_1, new_n14080, new_n14037);
not_3  g11733(new_n14082, new_n14081_1);
nor_4  g11734(new_n14083, new_n14082, new_n14078);
nor_4  g11735(new_n14084, new_n14081_1, new_n14077);
xnor_3 g11736(new_n14085, new_n14066, new_n14049);
not_3  g11737(new_n14086, new_n14085);
nand_4 g11738(new_n14087, new_n13977, new_n13974);
xnor_3 g11739(new_n14088, new_n14087, new_n14029);
nand_4 g11740(new_n14089, new_n14088, new_n14086);
xnor_3 g11741(new_n14090_1, new_n14088, new_n14085);
xnor_3 g11742(new_n14091, new_n14064, new_n14055);
not_3  g11743(new_n14092, new_n14091);
nand_4 g11744(new_n14093, new_n13983, new_n13980);
xnor_3 g11745(new_n14094, new_n14093, new_n14027);
nand_4 g11746(new_n14095_1, new_n14094, new_n14092);
xnor_3 g11747(new_n14096, new_n14094, new_n14091);
xnor_3 g11748(new_n14097, new_n14062, new_n14059_1);
not_3  g11749(new_n14098, new_n14097);
nand_4 g11750(new_n14099, new_n13987, new_n13986);
xnor_3 g11751(new_n14100, new_n14099, new_n14025);
nand_4 g11752(new_n14101, new_n14100, new_n14098);
xnor_3 g11753(new_n14102, new_n14100, new_n14097);
nor_4  g11754(new_n14103, new_n13993, new_n13990);
xnor_3 g11755(new_n14104, new_n14103, new_n14023);
nor_4  g11756(new_n14105, new_n14104, new_n4425);
not_3  g11757(new_n14106, new_n14105);
not_3  g11758(new_n14107_1, new_n4392);
nor_4  g11759(new_n14108, new_n4423, new_n14107_1);
nor_4  g11760(new_n14109, new_n4424_1, new_n4392);
nor_4  g11761(new_n14110, new_n14109, new_n14108);
not_3  g11762(new_n14111, new_n14104);
nor_4  g11763(new_n14112, new_n14111, new_n14110);
nor_4  g11764(new_n14113, new_n14112, new_n14105);
nand_4 g11765(new_n14114, new_n14000, new_n13998);
xnor_3 g11766(new_n14115, new_n14114, new_n14021);
nand_4 g11767(new_n14116, new_n14115, new_n4547);
nand_4 g11768(new_n14117, new_n14005, new_n14003);
xnor_3 g11769(new_n14118, new_n14117, new_n14019);
nand_4 g11770(new_n14119, new_n14118, new_n4559);
xnor_3 g11771(new_n14120, new_n14118, new_n4558);
nand_4 g11772(new_n14121_1, new_n14009, new_n14008);
xnor_3 g11773(new_n14122, new_n14121_1, new_n14017);
nand_4 g11774(new_n14123, new_n14122, new_n4563);
xnor_3 g11775(new_n14124, new_n14010, n11473);
xnor_3 g11776(new_n14125, new_n14124, new_n14015);
nor_4  g11777(new_n14126_1, new_n14125, new_n4572);
not_3  g11778(new_n14127, new_n14126_1);
xnor_3 g11779(new_n14128, new_n14014, new_n13106);
nand_4 g11780(new_n14129, new_n14128, new_n2609);
not_3  g11781(new_n14130_1, new_n14125);
nor_4  g11782(new_n14131, new_n14130_1, new_n4571);
nor_4  g11783(new_n14132, new_n14131, new_n14126_1);
nand_4 g11784(new_n14133, new_n14132, new_n14129);
nand_4 g11785(new_n14134, new_n14133, new_n14127);
not_3  g11786(new_n14135, new_n14123);
nor_4  g11787(new_n14136_1, new_n14122, new_n4563);
nor_4  g11788(new_n14137, new_n14136_1, new_n14135);
nand_4 g11789(new_n14138, new_n14137, new_n14134);
nand_4 g11790(new_n14139, new_n14138, new_n14123);
nand_4 g11791(new_n14140, new_n14139, new_n14120);
nand_4 g11792(new_n14141, new_n14140, new_n14119);
xnor_3 g11793(new_n14142, new_n14115, new_n4546);
nand_4 g11794(new_n14143, new_n14142, new_n14141);
nand_4 g11795(new_n14144, new_n14143, new_n14116);
nand_4 g11796(new_n14145, new_n14144, new_n14113);
nand_4 g11797(new_n14146, new_n14145, new_n14106);
nand_4 g11798(new_n14147_1, new_n14146, new_n14102);
nand_4 g11799(new_n14148_1, new_n14147_1, new_n14101);
nand_4 g11800(new_n14149, new_n14148_1, new_n14096);
nand_4 g11801(new_n14150, new_n14149, new_n14095_1);
nand_4 g11802(new_n14151, new_n14150, new_n14090_1);
nand_4 g11803(new_n14152, new_n14151, new_n14089);
nor_4  g11804(new_n14153, new_n14152, new_n14084);
nor_4  g11805(new_n14154, new_n14153, new_n14083);
nand_4 g11806(new_n14155, new_n14154, new_n14076);
nand_4 g11807(new_n14156, new_n14155, new_n14075);
xnor_3 g11808(new_n14157, new_n14156, new_n14071_1);
xnor_3 g11809(n1701, new_n14157, new_n14040);
not_3  g11810(new_n14159, new_n4292);
xor_3  g11811(n1703, new_n4330, new_n14159);
xor_3  g11812(n1721, new_n5221, new_n5149);
nor_4  g11813(new_n14162, new_n9127, new_n4905);
nor_4  g11814(new_n14163, new_n10726, new_n10724);
nor_4  g11815(new_n14164, new_n14163, new_n14162);
nor_4  g11816(new_n14165, new_n14164, new_n10784);
not_3  g11817(new_n14166, new_n10727);
nor_4  g11818(new_n14167, new_n10783, new_n14166);
nor_4  g11819(new_n14168, new_n10866, new_n10785);
nor_4  g11820(new_n14169, new_n14168, new_n14167);
nor_4  g11821(new_n14170, new_n14169, new_n14165);
not_3  g11822(new_n14171, new_n14164);
nor_4  g11823(new_n14172, new_n14171, new_n10783);
nor_4  g11824(new_n14173, new_n14172, new_n14168);
nor_4  g11825(n1760, new_n14173, new_n14170);
not_3  g11826(new_n14175, new_n4583);
xor_3  g11827(n1791, new_n14175, new_n4566);
xor_3  g11828(n1808, new_n3614, new_n3613);
nand_4 g11829(new_n14178, new_n9127, new_n9075);
nand_4 g11830(new_n14179, new_n9244, new_n9128);
nand_4 g11831(new_n14180, new_n14179, new_n14178);
not_3  g11832(new_n14181, n4319);
nor_4  g11833(new_n14182, n13494, new_n14181);
xor_3  g11834(new_n14183, n13494, n4319);
nor_4  g11835(new_n14184, n25345, new_n13462);
nand_4 g11836(new_n14185, new_n13490_1, new_n13463);
not_3  g11837(new_n14186, new_n14185);
nor_4  g11838(new_n14187, new_n14186, new_n14184);
nor_4  g11839(new_n14188, new_n14187, new_n14183);
nor_4  g11840(new_n14189, new_n14188, new_n14182);
not_3  g11841(new_n14190_1, new_n14189);
nor_4  g11842(new_n14191, new_n14190_1, new_n14180);
nor_4  g11843(new_n14192, new_n14189, new_n9245);
xnor_3 g11844(new_n14193, new_n14189, new_n9245);
xor_3  g11845(new_n14194, new_n14187, new_n14183);
nand_4 g11846(new_n14195, new_n14194, new_n9320);
xnor_3 g11847(new_n14196, new_n14194, new_n9316);
not_3  g11848(new_n14197, new_n13492);
nand_4 g11849(new_n14198, new_n13531, new_n13495);
nand_4 g11850(new_n14199, new_n14198, new_n14197);
nand_4 g11851(new_n14200, new_n14199, new_n14196);
nand_4 g11852(new_n14201, new_n14200, new_n14195);
nor_4  g11853(new_n14202, new_n14201, new_n14193);
nor_4  g11854(new_n14203, new_n14202, new_n14192);
nor_4  g11855(new_n14204, new_n14203, new_n14191);
not_3  g11856(new_n14205, new_n14180);
nor_4  g11857(new_n14206, new_n14189, new_n14205);
nor_4  g11858(new_n14207, new_n14206, new_n14202);
nor_4  g11859(n1821, new_n14207, new_n14204);
xor_3  g11860(n1832, new_n8180, new_n8177);
not_3  g11861(new_n14210, n2160);
xor_3  g11862(new_n14211_1, n9934, n2272);
not_3  g11863(new_n14212, new_n14211_1);
nor_4  g11864(new_n14213, n25331, n18496);
xor_3  g11865(new_n14214, n25331, n18496);
not_3  g11866(new_n14215, new_n14214);
nor_4  g11867(new_n14216, n26224, n18483);
xor_3  g11868(new_n14217, n26224, n18483);
not_3  g11869(new_n14218, new_n14217);
nand_4 g11870(new_n14219, new_n8210, new_n5426);
xor_3  g11871(new_n14220, n21934, n19327);
nor_4  g11872(new_n14221, n22597, n18901);
not_3  g11873(new_n14222_1, new_n14221);
xor_3  g11874(new_n14223, n22597, n18901);
nor_4  g11875(new_n14224, n26107, n4376);
not_3  g11876(new_n14225, new_n14224);
xor_3  g11877(new_n14226, n26107, n4376);
nor_4  g11878(new_n14227, n14570, n342);
not_3  g11879(new_n14228, new_n14227);
xor_3  g11880(new_n14229, n14570, n342);
nor_4  g11881(new_n14230_1, n26553, n23775);
not_3  g11882(new_n14231, new_n14230_1);
xor_3  g11883(new_n14232, n26553, n23775);
nand_4 g11884(new_n14233, new_n8229, new_n4116);
nand_4 g11885(new_n14234, n11479, n7876);
xor_3  g11886(new_n14235, n8259, n4964);
nand_4 g11887(new_n14236, new_n14235, new_n14234);
nand_4 g11888(new_n14237, new_n14236, new_n14233);
nand_4 g11889(new_n14238, new_n14237, new_n14232);
nand_4 g11890(new_n14239, new_n14238, new_n14231);
nand_4 g11891(new_n14240, new_n14239, new_n14229);
nand_4 g11892(new_n14241, new_n14240, new_n14228);
nand_4 g11893(new_n14242, new_n14241, new_n14226);
nand_4 g11894(new_n14243, new_n14242, new_n14225);
nand_4 g11895(new_n14244, new_n14243, new_n14223);
nand_4 g11896(new_n14245, new_n14244, new_n14222_1);
nand_4 g11897(new_n14246, new_n14245, new_n14220);
nand_4 g11898(new_n14247, new_n14246, new_n14219);
not_3  g11899(new_n14248, new_n14247);
nor_4  g11900(new_n14249, new_n14248, new_n14218);
nor_4  g11901(new_n14250, new_n14249, new_n14216);
nor_4  g11902(new_n14251, new_n14250, new_n14215);
nor_4  g11903(new_n14252, new_n14251, new_n14213);
xor_3  g11904(new_n14253, new_n14252, new_n14212);
xnor_3 g11905(new_n14254, new_n14253, new_n14210);
not_3  g11906(new_n14255, new_n14254);
xor_3  g11907(new_n14256, new_n14250, new_n14215);
nor_4  g11908(new_n14257, new_n14256, n10763);
not_3  g11909(new_n14258, new_n14257);
xnor_3 g11910(new_n14259, new_n14256, n10763);
not_3  g11911(new_n14260, new_n14259);
not_3  g11912(new_n14261, n7437);
xnor_3 g11913(new_n14262, new_n14247, new_n14217);
nor_4  g11914(new_n14263, new_n14262, new_n14261);
xnor_3 g11915(new_n14264, new_n14262, n7437);
xnor_3 g11916(new_n14265, new_n14245, new_n14220);
not_3  g11917(new_n14266, new_n14265);
nand_4 g11918(new_n14267_1, new_n14266, n20700);
xnor_3 g11919(new_n14268, new_n14265, n20700);
xnor_3 g11920(new_n14269, new_n14243, new_n14223);
not_3  g11921(new_n14270, new_n14269);
nand_4 g11922(new_n14271_1, new_n14270, n7099);
xnor_3 g11923(new_n14272, new_n14269, n7099);
xnor_3 g11924(new_n14273, new_n14241, new_n14226);
not_3  g11925(new_n14274, new_n14273);
nand_4 g11926(new_n14275_1, new_n14274, n12811);
xnor_3 g11927(new_n14276, new_n14273, n12811);
not_3  g11928(new_n14277_1, new_n14229);
xnor_3 g11929(new_n14278, new_n14239, new_n14277_1);
nand_4 g11930(new_n14279, new_n14278, n1118);
not_3  g11931(new_n14280, n1118);
xnor_3 g11932(new_n14281, new_n14278, new_n14280);
not_3  g11933(new_n14282, new_n14232);
xnor_3 g11934(new_n14283, new_n14237, new_n14282);
nand_4 g11935(new_n14284, new_n14283, n25974);
not_3  g11936(new_n14285, n25974);
xnor_3 g11937(new_n14286, new_n14283, new_n14285);
not_3  g11938(new_n14287, n1630);
xor_3  g11939(new_n14288, n11479, new_n4168);
nand_4 g11940(new_n14289, new_n14288, n1451);
nand_4 g11941(new_n14290, new_n14289, new_n14287);
not_3  g11942(new_n14291, new_n14290);
not_3  g11943(new_n14292, new_n14234);
xnor_3 g11944(new_n14293, new_n14235, new_n14292);
xnor_3 g11945(new_n14294_1, new_n14289, new_n14287);
nor_4  g11946(new_n14295, new_n14294_1, new_n14293);
nor_4  g11947(new_n14296, new_n14295, new_n14291);
nand_4 g11948(new_n14297, new_n14296, new_n14286);
nand_4 g11949(new_n14298, new_n14297, new_n14284);
nand_4 g11950(new_n14299, new_n14298, new_n14281);
nand_4 g11951(new_n14300, new_n14299, new_n14279);
nand_4 g11952(new_n14301, new_n14300, new_n14276);
nand_4 g11953(new_n14302, new_n14301, new_n14275_1);
nand_4 g11954(new_n14303, new_n14302, new_n14272);
nand_4 g11955(new_n14304, new_n14303, new_n14271_1);
nand_4 g11956(new_n14305, new_n14304, new_n14268);
nand_4 g11957(new_n14306, new_n14305, new_n14267_1);
nand_4 g11958(new_n14307, new_n14306, new_n14264);
not_3  g11959(new_n14308, new_n14307);
nor_4  g11960(new_n14309, new_n14308, new_n14263);
nand_4 g11961(new_n14310_1, new_n14309, new_n14260);
nand_4 g11962(new_n14311, new_n14310_1, new_n14258);
xnor_3 g11963(new_n14312, new_n14311, new_n14255);
not_3  g11964(new_n14313, n21784);
not_3  g11965(new_n14314, new_n4227);
nor_4  g11966(new_n14315, new_n14314, n4325);
not_3  g11967(new_n14316, new_n14315);
nor_4  g11968(new_n14317, new_n14316, n11926);
not_3  g11969(new_n14318, new_n14317);
nor_4  g11970(new_n14319, new_n14318, n5521);
xor_3  g11971(new_n14320, new_n14319, new_n14313);
xnor_3 g11972(new_n14321, new_n14320, new_n8573);
not_3  g11973(new_n14322, new_n14321);
not_3  g11974(new_n14323_1, n5521);
xor_3  g11975(new_n14324, new_n14317, new_n14323_1);
nor_4  g11976(new_n14325, new_n14324, new_n8580);
not_3  g11977(new_n14326_1, new_n14325);
not_3  g11978(new_n14327, new_n14324);
nor_4  g11979(new_n14328, new_n14327, new_n8584);
nor_4  g11980(new_n14329, new_n14328, new_n14325);
not_3  g11981(new_n14330, n11926);
xor_3  g11982(new_n14331, new_n14315, new_n14330);
nor_4  g11983(new_n14332, new_n14331, new_n8590);
not_3  g11984(new_n14333, new_n14332);
not_3  g11985(new_n14334, new_n14331);
xor_3  g11986(new_n14335, new_n14334, new_n8590);
not_3  g11987(new_n14336, new_n14335);
not_3  g11988(new_n14337, new_n4228);
nand_4 g11989(new_n14338, new_n14337, new_n4218);
nand_4 g11990(new_n14339, new_n4281, new_n4229);
nand_4 g11991(new_n14340, new_n14339, new_n14338);
nand_4 g11992(new_n14341, new_n14340, new_n14336);
nand_4 g11993(new_n14342_1, new_n14341, new_n14333);
nand_4 g11994(new_n14343, new_n14342_1, new_n14329);
nand_4 g11995(new_n14344, new_n14343, new_n14326_1);
xnor_3 g11996(new_n14345_1, new_n14344, new_n14322);
xnor_3 g11997(new_n14346, new_n14345_1, new_n14312);
xnor_3 g11998(new_n14347, new_n14309, new_n14259);
xnor_3 g11999(new_n14348, new_n14342_1, new_n14329);
nor_4  g12000(new_n14349, new_n14348, new_n14347);
xnor_3 g12001(new_n14350, new_n14348, new_n14347);
xnor_3 g12002(new_n14351, new_n14306, new_n14264);
not_3  g12003(new_n14352, new_n14351);
not_3  g12004(new_n14353_1, new_n14340);
xnor_3 g12005(new_n14354, new_n14353_1, new_n14335);
not_3  g12006(new_n14355, new_n14354);
nand_4 g12007(new_n14356, new_n14355, new_n14352);
xnor_3 g12008(new_n14357, new_n14355, new_n14351);
xnor_3 g12009(new_n14358, new_n14304, new_n14268);
not_3  g12010(new_n14359, new_n14358);
nand_4 g12011(new_n14360, new_n14359, new_n4283);
xnor_3 g12012(new_n14361, new_n14358, new_n4283);
xnor_3 g12013(new_n14362, new_n14302, new_n14272);
not_3  g12014(new_n14363, new_n14362);
nand_4 g12015(new_n14364_1, new_n14363, new_n4291);
xnor_3 g12016(new_n14365, new_n14362, new_n4291);
not_3  g12017(new_n14366, new_n14276);
xnor_3 g12018(new_n14367, new_n14300, new_n14366);
nand_4 g12019(new_n14368, new_n14367, new_n4294);
xnor_3 g12020(new_n14369, new_n14367, new_n4293);
not_3  g12021(new_n14370, new_n14281);
xnor_3 g12022(new_n14371, new_n14298, new_n14370);
nand_4 g12023(new_n14372, new_n14371, new_n4299);
xnor_3 g12024(new_n14373, new_n14371, new_n4298);
xnor_3 g12025(new_n14374, new_n14296, new_n14286);
not_3  g12026(new_n14375_1, new_n14374);
nand_4 g12027(new_n14376, new_n14375_1, new_n4306_1);
xnor_3 g12028(new_n14377, new_n14374, new_n4306_1);
xnor_3 g12029(new_n14378, new_n14288, n1451);
nand_4 g12030(new_n14379, new_n14378, new_n4318);
xnor_3 g12031(new_n14380, new_n14294_1, new_n14293);
nor_4  g12032(new_n14381, new_n14380, new_n14379);
xnor_3 g12033(new_n14382, new_n14380, new_n14379);
nor_4  g12034(new_n14383, new_n14382, new_n4311);
nor_4  g12035(new_n14384, new_n14383, new_n14381);
nand_4 g12036(new_n14385, new_n14384, new_n14377);
nand_4 g12037(new_n14386, new_n14385, new_n14376);
nand_4 g12038(new_n14387, new_n14386, new_n14373);
nand_4 g12039(new_n14388, new_n14387, new_n14372);
nand_4 g12040(new_n14389, new_n14388, new_n14369);
nand_4 g12041(new_n14390, new_n14389, new_n14368);
nand_4 g12042(new_n14391, new_n14390, new_n14365);
nand_4 g12043(new_n14392, new_n14391, new_n14364_1);
nand_4 g12044(new_n14393, new_n14392, new_n14361);
nand_4 g12045(new_n14394, new_n14393, new_n14360);
nand_4 g12046(new_n14395, new_n14394, new_n14357);
nand_4 g12047(new_n14396, new_n14395, new_n14356);
not_3  g12048(new_n14397, new_n14396);
nor_4  g12049(new_n14398, new_n14397, new_n14350);
nor_4  g12050(new_n14399, new_n14398, new_n14349);
xnor_3 g12051(n1859, new_n14399, new_n14346);
nor_4  g12052(new_n14401, new_n6000, new_n5974);
xor_3  g12053(n1860, new_n14401, new_n5971);
nand_4 g12054(new_n14403, new_n10327_1, new_n6326);
nand_4 g12055(new_n14404, new_n8072, new_n8044);
nand_4 g12056(new_n14405, new_n14404, new_n14403);
not_3  g12057(new_n14406, new_n14405);
nor_4  g12058(new_n14407, n25972, n8614);
nand_4 g12059(new_n14408, n25972, n8614);
not_3  g12060(new_n14409, new_n14408);
nor_4  g12061(new_n14410, new_n14409, new_n14407);
not_3  g12062(new_n14411, new_n14410);
xor_3  g12063(new_n14412_1, new_n14411, new_n14406);
nor_4  g12064(new_n14413, new_n14412_1, new_n10324);
not_3  g12065(new_n14414_1, new_n14413);
not_3  g12066(new_n14415, new_n14412_1);
nor_4  g12067(new_n14416, new_n14415, n10250);
nor_4  g12068(new_n14417, new_n14416, new_n14413);
nor_4  g12069(new_n14418, new_n8074, new_n10329);
not_3  g12070(new_n14419, new_n14418);
xor_3  g12071(new_n14420, new_n8074, new_n10329);
nand_4 g12072(new_n14421, new_n8078, n6397);
xor_3  g12073(new_n14422, new_n8077, new_n10331);
nor_4  g12074(new_n14423, new_n8084, new_n7209);
not_3  g12075(new_n14424, new_n14423);
nor_4  g12076(new_n14425, new_n8087, n19196);
nor_4  g12077(new_n14426, new_n14425, new_n14423);
not_3  g12078(new_n14427, n23586);
nor_4  g12079(new_n14428, new_n8092, new_n14427);
not_3  g12080(new_n14429, new_n14428);
nor_4  g12081(new_n14430, new_n8102, n21226);
not_3  g12082(new_n14431, n21226);
nor_4  g12083(new_n14432, new_n8099, new_n14431);
nor_4  g12084(new_n14433, new_n14432, new_n14430);
not_3  g12085(new_n14434, new_n14433);
not_3  g12086(new_n14435, n4426);
nor_4  g12087(new_n14436, new_n8107, new_n14435);
not_3  g12088(new_n14437, new_n14436);
xor_3  g12089(new_n14438, new_n8107, new_n14435);
nor_4  g12090(new_n14439, new_n8119, n20036);
nor_4  g12091(new_n14440_1, new_n4618, new_n4607);
not_3  g12092(new_n14441, new_n14440_1);
nor_4  g12093(new_n14442, new_n8179_1, new_n4609);
nor_4  g12094(new_n14443, new_n4629, n11192);
nor_4  g12095(new_n14444, new_n14443, new_n14440_1);
nand_4 g12096(new_n14445, new_n14444, new_n14442);
nand_4 g12097(new_n14446, new_n14445, new_n14441);
xnor_3 g12098(new_n14447, new_n4603, new_n10346);
nor_4  g12099(new_n14448, new_n14447, new_n14446);
nor_4  g12100(new_n14449, new_n14448, new_n14439);
nand_4 g12101(new_n14450, new_n14449, new_n14438);
nand_4 g12102(new_n14451, new_n14450, new_n14437);
nor_4  g12103(new_n14452, new_n14451, new_n14434);
nor_4  g12104(new_n14453, new_n14452, new_n14430);
nor_4  g12105(new_n14454, new_n8095_1, n23586);
nor_4  g12106(new_n14455, new_n14454, new_n14428);
nand_4 g12107(new_n14456, new_n14455, new_n14453);
nand_4 g12108(new_n14457_1, new_n14456, new_n14429);
nand_4 g12109(new_n14458, new_n14457_1, new_n14426);
nand_4 g12110(new_n14459, new_n14458, new_n14424);
nand_4 g12111(new_n14460, new_n14459, new_n14422);
nand_4 g12112(new_n14461, new_n14460, new_n14421);
nand_4 g12113(new_n14462, new_n14461, new_n14420);
nand_4 g12114(new_n14463, new_n14462, new_n14419);
nand_4 g12115(new_n14464_1, new_n14463, new_n14417);
nand_4 g12116(new_n14465, new_n14464_1, new_n14414_1);
not_3  g12117(new_n14466, new_n14407);
nand_4 g12118(new_n14467, new_n14466, new_n14406);
nand_4 g12119(new_n14468, new_n14467, new_n14408);
nand_4 g12120(new_n14469, new_n14468, new_n14465);
nand_4 g12121(new_n14470, new_n14469, new_n13774);
xnor_3 g12122(new_n14471_1, new_n14469, new_n13773);
xnor_3 g12123(new_n14472, new_n14468, new_n14465);
nand_4 g12124(new_n14473, new_n14472, new_n13775_1);
xnor_3 g12125(new_n14474, new_n14472, new_n13790);
xnor_3 g12126(new_n14475_1, new_n14463, new_n14417);
nand_4 g12127(new_n14476, new_n14475_1, new_n13794);
xnor_3 g12128(new_n14477, new_n14475_1, new_n13793);
xnor_3 g12129(new_n14478, new_n14461, new_n14420);
nand_4 g12130(new_n14479, new_n14478, new_n13803);
xnor_3 g12131(new_n14480, new_n14478, new_n13802);
xnor_3 g12132(new_n14481, new_n14459, new_n14422);
nand_4 g12133(new_n14482, new_n14481, new_n13811);
xnor_3 g12134(new_n14483, new_n14481, new_n13816);
xnor_3 g12135(new_n14484, new_n14457_1, new_n14426);
nand_4 g12136(new_n14485, new_n14484, new_n13820);
xnor_3 g12137(new_n14486, new_n14484, new_n13836);
not_3  g12138(new_n14487, new_n13828);
xnor_3 g12139(new_n14488, new_n14455, new_n14453);
nand_4 g12140(new_n14489, new_n14488, new_n14487);
xnor_3 g12141(new_n14490, new_n14488, new_n13828);
not_3  g12142(new_n14491, new_n11471);
xnor_3 g12143(new_n14492, new_n14451, new_n14434);
nor_4  g12144(new_n14493, new_n14492, new_n14491);
not_3  g12145(new_n14494, new_n14493);
xnor_3 g12146(new_n14495, new_n14451, new_n14433);
nor_4  g12147(new_n14496, new_n14495, new_n11471);
nor_4  g12148(new_n14497, new_n14496, new_n14493);
not_3  g12149(new_n14498, new_n11486_1);
xor_3  g12150(new_n14499, new_n8107, n4426);
xnor_3 g12151(new_n14500, new_n14449, new_n14499);
nor_4  g12152(new_n14501, new_n14500, new_n14498);
not_3  g12153(new_n14502, new_n14501);
xnor_3 g12154(new_n14503, new_n14449, new_n14438);
nor_4  g12155(new_n14504, new_n14503, new_n11486_1);
nor_4  g12156(new_n14505, new_n14504, new_n14501);
not_3  g12157(new_n14506, new_n14442);
xnor_3 g12158(new_n14507, new_n4618, new_n4607);
nor_4  g12159(new_n14508, new_n14507, new_n14506);
nor_4  g12160(new_n14509, new_n14508, new_n14440_1);
xnor_3 g12161(new_n14510_1, new_n14447, new_n14509);
nand_4 g12162(new_n14511, new_n14510_1, new_n11491);
not_3  g12163(new_n14512, new_n14511);
nor_4  g12164(new_n14513, new_n14510_1, new_n11491);
nor_4  g12165(new_n14514, new_n14513, new_n14512);
not_3  g12166(new_n14515, new_n11496_1);
xnor_3 g12167(new_n14516, new_n14507, new_n14506);
nand_4 g12168(new_n14517, new_n14516, new_n14515);
xor_3  g12169(new_n14518, new_n8179_1, new_n4609);
nor_4  g12170(new_n14519, new_n14518, new_n8492);
not_3  g12171(new_n14520, new_n14517);
nor_4  g12172(new_n14521, new_n14516, new_n14515);
nor_4  g12173(new_n14522, new_n14521, new_n14520);
nand_4 g12174(new_n14523, new_n14522, new_n14519);
nand_4 g12175(new_n14524, new_n14523, new_n14517);
nand_4 g12176(new_n14525, new_n14524, new_n14514);
nand_4 g12177(new_n14526, new_n14525, new_n14511);
nand_4 g12178(new_n14527, new_n14526, new_n14505);
nand_4 g12179(new_n14528, new_n14527, new_n14502);
nand_4 g12180(new_n14529, new_n14528, new_n14497);
nand_4 g12181(new_n14530, new_n14529, new_n14494);
nand_4 g12182(new_n14531, new_n14530, new_n14490);
nand_4 g12183(new_n14532, new_n14531, new_n14489);
nand_4 g12184(new_n14533, new_n14532, new_n14486);
nand_4 g12185(new_n14534, new_n14533, new_n14485);
nand_4 g12186(new_n14535, new_n14534, new_n14483);
nand_4 g12187(new_n14536, new_n14535, new_n14482);
nand_4 g12188(new_n14537, new_n14536, new_n14480);
nand_4 g12189(new_n14538, new_n14537, new_n14479);
nand_4 g12190(new_n14539, new_n14538, new_n14477);
nand_4 g12191(new_n14540, new_n14539, new_n14476);
nand_4 g12192(new_n14541_1, new_n14540, new_n14474);
nand_4 g12193(new_n14542, new_n14541_1, new_n14473);
nand_4 g12194(new_n14543, new_n14542, new_n14471_1);
nand_4 g12195(n1861, new_n14543, new_n14470);
nor_4  g12196(new_n14545, n13714, n12593);
nand_4 g12197(new_n14546_1, new_n14545, new_n10474);
nor_4  g12198(new_n14547_1, new_n14546_1, n8309);
not_3  g12199(new_n14548, new_n14547_1);
nor_4  g12200(new_n14549, new_n14548, n19081);
nand_4 g12201(new_n14550, new_n14549, new_n12106);
xor_3  g12202(new_n14551, new_n14550, n26318);
xnor_3 g12203(new_n14552, new_n14551, new_n6167);
xor_3  g12204(new_n14553, new_n14549, new_n12106);
not_3  g12205(new_n14554, new_n14553);
nand_4 g12206(new_n14555, new_n14554, new_n6172);
xor_3  g12207(new_n14556, new_n14547_1, n19081);
nand_4 g12208(new_n14557, new_n14556, new_n6228);
xnor_3 g12209(new_n14558, new_n14556, new_n6227);
xor_3  g12210(new_n14559, new_n14546_1, n8309);
nor_4  g12211(new_n14560, new_n14559, new_n6180);
not_3  g12212(new_n14561, new_n14560);
xor_3  g12213(new_n14562, new_n14545, new_n10474);
nor_4  g12214(new_n14563, new_n14562, new_n6211);
not_3  g12215(new_n14564, new_n14563);
xnor_3 g12216(new_n14565, new_n14562, new_n6191);
nand_4 g12217(new_n14566, new_n6203, n13714);
xnor_3 g12218(new_n14567, new_n14566, n12593);
not_3  g12219(new_n14568, new_n14567);
nor_4  g12220(new_n14569, new_n14568, new_n6196);
nor_4  g12221(new_n14570_1, new_n6203, new_n12281);
not_3  g12222(new_n14571, new_n14570_1);
nor_4  g12223(new_n14572, new_n14571, n12593);
nor_4  g12224(new_n14573, new_n14572, new_n14569);
nand_4 g12225(new_n14574, new_n14573, new_n14565);
nand_4 g12226(new_n14575_1, new_n14574, new_n14564);
not_3  g12227(new_n14576_1, new_n14559);
nor_4  g12228(new_n14577, new_n14576_1, new_n6179);
nor_4  g12229(new_n14578, new_n14577, new_n14560);
nand_4 g12230(new_n14579, new_n14578, new_n14575_1);
nand_4 g12231(new_n14580, new_n14579, new_n14561);
nand_4 g12232(new_n14581, new_n14580, new_n14558);
nand_4 g12233(new_n14582, new_n14581, new_n14557);
xnor_3 g12234(new_n14583, new_n14553, new_n6172);
nand_4 g12235(new_n14584, new_n14583, new_n14582);
nand_4 g12236(new_n14585, new_n14584, new_n14555);
xnor_3 g12237(new_n14586, new_n14585, new_n14552);
nor_4  g12238(new_n14587, new_n10229, n20179);
xor_3  g12239(new_n14588, new_n14587, new_n7937_1);
nand_4 g12240(new_n14589, new_n14588, new_n8596);
not_3  g12241(new_n14590, new_n14589);
nor_4  g12242(new_n14591, new_n14588, new_n8596);
nor_4  g12243(new_n14592, new_n14591, new_n14590);
nand_4 g12244(new_n14593_1, new_n10229, n20179);
not_3  g12245(new_n14594, new_n14593_1);
nor_4  g12246(new_n14595, new_n14594, new_n14587);
nand_4 g12247(new_n14596, new_n14595, new_n8602);
not_3  g12248(new_n14597, new_n14596);
nor_4  g12249(new_n14598, new_n14595, new_n8602);
nor_4  g12250(new_n14599, new_n14598, new_n14597);
nor_4  g12251(new_n14600, new_n10232, new_n8604);
xnor_3 g12252(new_n14601, new_n10232, new_n8604);
nor_4  g12253(new_n14602, new_n10237, new_n8611);
xnor_3 g12254(new_n14603_1, new_n10238, new_n8610);
nand_4 g12255(new_n14604, new_n10245, new_n8618);
not_3  g12256(new_n14605, new_n10245);
nand_4 g12257(new_n14606, new_n14605, new_n8617);
nor_4  g12258(new_n14607, new_n10251, new_n8629);
not_3  g12259(new_n14608, new_n8627);
nor_4  g12260(new_n14609, new_n14608, new_n8997);
xnor_3 g12261(new_n14610, new_n10255, new_n8624);
nor_4  g12262(new_n14611, new_n14610, new_n14609);
nor_4  g12263(new_n14612, new_n14611, new_n14607);
nand_4 g12264(new_n14613, new_n14612, new_n14606);
nand_4 g12265(new_n14614, new_n14613, new_n14604);
nor_4  g12266(new_n14615, new_n14614, new_n14603_1);
nor_4  g12267(new_n14616, new_n14615, new_n14602);
nor_4  g12268(new_n14617, new_n14616, new_n14601);
nor_4  g12269(new_n14618, new_n14617, new_n14600);
nand_4 g12270(new_n14619, new_n14618, new_n14599);
nand_4 g12271(new_n14620, new_n14619, new_n14596);
nand_4 g12272(new_n14621, new_n14620, new_n14592);
not_3  g12273(new_n14622, new_n14621);
nor_4  g12274(new_n14623, new_n14620, new_n14592);
nor_4  g12275(new_n14624, new_n14623, new_n14622);
nor_4  g12276(new_n14625, new_n14624, new_n14586);
not_3  g12277(new_n14626, new_n14552);
xnor_3 g12278(new_n14627, new_n14585, new_n14626);
not_3  g12279(new_n14628, new_n14624);
nor_4  g12280(new_n14629, new_n14628, new_n14627);
nor_4  g12281(new_n14630, new_n14629, new_n14625);
xnor_3 g12282(new_n14631, new_n14618, new_n14599);
xnor_3 g12283(new_n14632, new_n14583, new_n14582);
not_3  g12284(new_n14633_1, new_n14632);
nand_4 g12285(new_n14634, new_n14633_1, new_n14631);
xnor_3 g12286(new_n14635, new_n14632, new_n14631);
not_3  g12287(new_n14636_1, new_n14558);
xnor_3 g12288(new_n14637, new_n14580, new_n14636_1);
xnor_3 g12289(new_n14638, new_n14616, new_n14601);
not_3  g12290(new_n14639, new_n14638);
nand_4 g12291(new_n14640, new_n14639, new_n14637);
xnor_3 g12292(new_n14641, new_n14638, new_n14637);
xnor_3 g12293(new_n14642, new_n14578, new_n14575_1);
not_3  g12294(new_n14643, new_n14642);
not_3  g12295(new_n14644, new_n14603_1);
not_3  g12296(new_n14645, new_n14614);
nor_4  g12297(new_n14646, new_n14645, new_n14644);
nor_4  g12298(new_n14647, new_n14646, new_n14615);
nand_4 g12299(new_n14648, new_n14647, new_n14643);
xnor_3 g12300(new_n14649, new_n14647, new_n14642);
xnor_3 g12301(new_n14650, new_n14573, new_n14565);
nand_4 g12302(new_n14651, new_n14606, new_n14604);
xnor_3 g12303(new_n14652, new_n14651, new_n14612);
nor_4  g12304(new_n14653, new_n14652, new_n14650);
not_3  g12305(new_n14654, new_n14653);
not_3  g12306(new_n14655, new_n14650);
not_3  g12307(new_n14656, new_n14652);
nor_4  g12308(new_n14657, new_n14656, new_n14655);
nor_4  g12309(new_n14658, new_n14657, new_n14653);
not_3  g12310(new_n14659, new_n14609);
not_3  g12311(new_n14660, new_n14610);
nor_4  g12312(new_n14661, new_n14660, new_n14659);
nor_4  g12313(new_n14662, new_n14661, new_n14611);
not_3  g12314(new_n14663, new_n14662);
nor_4  g12315(new_n14664, new_n14567, new_n6206);
nor_4  g12316(new_n14665, new_n14664, new_n14569);
nor_4  g12317(new_n14666, new_n14665, new_n14663);
not_3  g12318(new_n14667, new_n14666);
xor_3  g12319(new_n14668, new_n8627, n18962);
xor_3  g12320(new_n14669, new_n6203, new_n12281);
nand_4 g12321(new_n14670, new_n14669, new_n14668);
not_3  g12322(new_n14671, new_n14665);
nor_4  g12323(new_n14672, new_n14671, new_n14662);
nor_4  g12324(new_n14673, new_n14672, new_n14666);
nand_4 g12325(new_n14674, new_n14673, new_n14670);
nand_4 g12326(new_n14675, new_n14674, new_n14667);
nand_4 g12327(new_n14676, new_n14675, new_n14658);
nand_4 g12328(new_n14677, new_n14676, new_n14654);
nand_4 g12329(new_n14678, new_n14677, new_n14649);
nand_4 g12330(new_n14679, new_n14678, new_n14648);
nand_4 g12331(new_n14680_1, new_n14679, new_n14641);
nand_4 g12332(new_n14681, new_n14680_1, new_n14640);
nand_4 g12333(new_n14682, new_n14681, new_n14635);
nand_4 g12334(new_n14683, new_n14682, new_n14634);
xnor_3 g12335(n1891, new_n14683, new_n14630);
xor_3  g12336(new_n14685, n20169, n1949);
nor_4  g12337(new_n14686, new_n4437, n8285);
not_3  g12338(new_n14687, new_n14686);
not_3  g12339(new_n14688, n8285);
nor_4  g12340(new_n14689, n9323, new_n14688);
not_3  g12341(new_n14690, new_n14689);
nor_4  g12342(new_n14691, new_n4460, n6729);
not_3  g12343(new_n14692_1, new_n14691);
not_3  g12344(new_n14693, n6729);
nor_4  g12345(new_n14694, n10792, new_n14693);
not_3  g12346(new_n14695, new_n14694);
nor_4  g12347(new_n14696, n21687, new_n4461);
nand_4 g12348(new_n14697, new_n14696, new_n14695);
nand_4 g12349(new_n14698, new_n14697, new_n14692_1);
nand_4 g12350(new_n14699, new_n14698, new_n14690);
nand_4 g12351(new_n14700, new_n14699, new_n14687);
not_3  g12352(new_n14701_1, new_n14700);
xor_3  g12353(new_n14702_1, new_n14701_1, new_n14685);
xnor_3 g12354(new_n14703, new_n14702_1, new_n7699);
nor_4  g12355(new_n14704_1, new_n14689, new_n14686);
xor_3  g12356(new_n14705, new_n14704_1, new_n14698);
not_3  g12357(new_n14706, new_n14705);
nor_4  g12358(new_n14707, new_n14706, new_n7705);
not_3  g12359(new_n14708, new_n14707);
nor_4  g12360(new_n14709, new_n14705, new_n7708_1);
nor_4  g12361(new_n14710, new_n14709, new_n14707);
xor_3  g12362(new_n14711, n21687, new_n4461);
nor_4  g12363(new_n14712, new_n14711, new_n7711);
nor_4  g12364(new_n14713, new_n14694, new_n14691);
xor_3  g12365(new_n14714, new_n14713, new_n14696);
not_3  g12366(new_n14715, new_n14714);
nor_4  g12367(new_n14716, new_n14715, new_n14712);
not_3  g12368(new_n14717, new_n14716);
not_3  g12369(new_n14718, new_n14712);
nor_4  g12370(new_n14719, new_n14714, new_n14718);
nor_4  g12371(new_n14720, new_n14719, new_n14716);
nand_4 g12372(new_n14721, new_n14720, new_n7715);
nand_4 g12373(new_n14722, new_n14721, new_n14717);
nand_4 g12374(new_n14723, new_n14722, new_n14710);
nand_4 g12375(new_n14724, new_n14723, new_n14708);
not_3  g12376(new_n14725, new_n14724);
xor_3  g12377(n1925, new_n14725, new_n14703);
not_3  g12378(new_n14727, new_n8977);
xor_3  g12379(n1942, new_n9016, new_n14727);
xnor_3 g12380(n1972, new_n7513, new_n7436);
nor_4  g12381(new_n14730, new_n10507, new_n10422);
nor_4  g12382(new_n14731, new_n10580, new_n10515);
nor_4  g12383(new_n14732, new_n14731, new_n10513);
nor_4  g12384(new_n14733, new_n14732, new_n10508);
nor_4  g12385(new_n14734_1, new_n14733, new_n14730);
not_3  g12386(new_n14735, new_n10432_1);
nor_4  g12387(new_n14736, new_n14735, n22764);
not_3  g12388(new_n14737, new_n10435);
not_3  g12389(new_n14738, new_n10436);
nand_4 g12390(new_n14739, new_n10506, new_n14738);
nand_4 g12391(new_n14740, new_n14739, new_n14737);
nor_4  g12392(new_n14741, new_n14740, new_n14736);
nand_4 g12393(new_n14742, new_n14741, new_n13379);
not_3  g12394(new_n14743, new_n14742);
nand_4 g12395(new_n14744, new_n14743, new_n14734_1);
not_3  g12396(new_n14745, new_n14730);
nand_4 g12397(new_n14746_1, new_n10583, new_n10509);
nand_4 g12398(new_n14747, new_n14746_1, new_n14745);
nor_4  g12399(new_n14748, new_n14741, new_n13379);
nand_4 g12400(new_n14749, new_n14748, new_n14747);
nand_4 g12401(new_n14750, new_n14749, new_n14744);
nor_4  g12402(new_n14751, new_n14750, new_n13240);
not_3  g12403(new_n14752, new_n14750);
nor_4  g12404(new_n14753, new_n14752, new_n13241);
nor_4  g12405(new_n14754, new_n14753, new_n14751);
not_3  g12406(new_n14755, new_n14754);
nor_4  g12407(new_n14756, new_n14748, new_n14743);
xnor_3 g12408(new_n14757, new_n14756, new_n14747);
nor_4  g12409(new_n14758, new_n14757, new_n13240);
not_3  g12410(new_n14759, new_n14758);
xnor_3 g12411(new_n14760, new_n14756, new_n14734_1);
nor_4  g12412(new_n14761, new_n14760, new_n13241);
nor_4  g12413(new_n14762, new_n14761, new_n14758);
not_3  g12414(new_n14763_1, new_n10584);
nor_4  g12415(new_n14764, new_n13290, new_n14763_1);
not_3  g12416(new_n14765, new_n14764);
nand_4 g12417(new_n14766, new_n13298, new_n10588_1);
xnor_3 g12418(new_n14767, new_n13302, new_n10588_1);
nand_4 g12419(new_n14768, new_n13306, new_n10597);
nor_4  g12420(new_n14769, new_n13309, new_n10593_1);
nor_4  g12421(new_n14770, new_n13306, new_n10597);
nor_4  g12422(new_n14771, new_n14770, new_n14769);
nand_4 g12423(new_n14772_1, new_n13311, new_n10602);
xnor_3 g12424(new_n14773, new_n13311, new_n10601);
nand_4 g12425(new_n14774, new_n13316, new_n10608);
xnor_3 g12426(new_n14775, new_n13317, new_n10608);
nand_4 g12427(new_n14776, new_n13355, new_n10614_1);
xnor_3 g12428(new_n14777, new_n13326, new_n10614_1);
nand_4 g12429(new_n14778, new_n13333_1, new_n10619);
xnor_3 g12430(new_n14779, new_n13330, new_n10619);
nor_4  g12431(new_n14780, new_n13337, new_n10627);
not_3  g12432(new_n14781, new_n14780);
nor_4  g12433(new_n14782, new_n13338_1, new_n10628_1);
nor_4  g12434(new_n14783, new_n14782, new_n14780);
not_3  g12435(new_n14784, new_n13344);
xor_3  g12436(new_n14785, n8581, new_n11981);
nor_4  g12437(new_n14786, new_n14785, new_n10635);
nor_4  g12438(new_n14787, new_n14786, new_n14784);
not_3  g12439(new_n14788, new_n14787);
not_3  g12440(new_n14789, new_n14786);
xor_3  g12441(new_n14790_1, new_n14789, new_n13344);
nand_4 g12442(new_n14791, new_n14790_1, new_n10643);
nand_4 g12443(new_n14792, new_n14791, new_n14788);
nand_4 g12444(new_n14793, new_n14792, new_n14783);
nand_4 g12445(new_n14794, new_n14793, new_n14781);
nand_4 g12446(new_n14795, new_n14794, new_n14779);
nand_4 g12447(new_n14796, new_n14795, new_n14778);
nand_4 g12448(new_n14797, new_n14796, new_n14777);
nand_4 g12449(new_n14798, new_n14797, new_n14776);
nand_4 g12450(new_n14799, new_n14798, new_n14775);
nand_4 g12451(new_n14800, new_n14799, new_n14774);
nand_4 g12452(new_n14801_1, new_n14800, new_n14773);
nand_4 g12453(new_n14802, new_n14801_1, new_n14772_1);
nand_4 g12454(new_n14803, new_n14802, new_n14771);
nand_4 g12455(new_n14804, new_n14803, new_n14768);
nand_4 g12456(new_n14805, new_n14804, new_n14767);
nand_4 g12457(new_n14806, new_n14805, new_n14766);
nor_4  g12458(new_n14807, new_n13294, new_n10584);
nor_4  g12459(new_n14808, new_n14807, new_n14764);
nand_4 g12460(new_n14809, new_n14808, new_n14806);
nand_4 g12461(new_n14810, new_n14809, new_n14765);
nand_4 g12462(new_n14811, new_n14810, new_n14762);
nand_4 g12463(new_n14812, new_n14811, new_n14759);
nor_4  g12464(new_n14813, new_n14812, new_n14755);
nor_4  g12465(n1981, new_n14813, new_n14751);
xnor_3 g12466(n2004, new_n14808, new_n14806);
not_3  g12467(new_n14816, n5140);
nor_4  g12468(new_n14817, n6105, new_n14816);
xor_3  g12469(new_n14818, n6105, new_n14816);
not_3  g12470(new_n14819_1, new_n14818);
not_3  g12471(new_n14820, n6204);
nor_4  g12472(new_n14821, new_n14820, n3795);
xor_3  g12473(new_n14822, n6204, new_n7393);
not_3  g12474(new_n14823, n25464);
nand_4 g12475(new_n14824, new_n14823, n3349);
not_3  g12476(new_n14825, n3349);
xor_3  g12477(new_n14826_1, n25464, new_n14825);
not_3  g12478(new_n14827_1, n4590);
nand_4 g12479(new_n14828, new_n14827_1, n1742);
not_3  g12480(new_n14829, n1742);
xor_3  g12481(new_n14830, n4590, new_n14829);
not_3  g12482(new_n14831, n26752);
nand_4 g12483(new_n14832, new_n14831, n4858);
xor_3  g12484(new_n14833, n26752, new_n7579);
nor_4  g12485(new_n14834, new_n7583, n6513);
not_3  g12486(new_n14835, new_n14834);
not_3  g12487(new_n14836, n6513);
xor_3  g12488(new_n14837, n8244, new_n14836);
nor_4  g12489(new_n14838, new_n7614, n3918);
not_3  g12490(new_n14839_1, new_n14838);
not_3  g12491(new_n14840, n3918);
xor_3  g12492(new_n14841, n9493, new_n14840);
not_3  g12493(new_n14842, n919);
nor_4  g12494(new_n14843, n15167, new_n14842);
nor_4  g12495(new_n14844, new_n7599, n919);
not_3  g12496(new_n14845, n25316);
nor_4  g12497(new_n14846, new_n14845, n21095);
nor_4  g12498(new_n14847, n25316, new_n7602);
not_3  g12499(new_n14848, n8656);
nand_4 g12500(new_n14849_1, n20385, new_n14848);
nor_4  g12501(new_n14850, new_n14849_1, new_n14847);
nor_4  g12502(new_n14851, new_n14850, new_n14846);
nor_4  g12503(new_n14852, new_n14851, new_n14844);
nor_4  g12504(new_n14853, new_n14852, new_n14843);
nand_4 g12505(new_n14854, new_n14853, new_n14841);
nand_4 g12506(new_n14855, new_n14854, new_n14839_1);
nand_4 g12507(new_n14856, new_n14855, new_n14837);
nand_4 g12508(new_n14857, new_n14856, new_n14835);
nand_4 g12509(new_n14858, new_n14857, new_n14833);
nand_4 g12510(new_n14859, new_n14858, new_n14832);
nand_4 g12511(new_n14860, new_n14859, new_n14830);
nand_4 g12512(new_n14861, new_n14860, new_n14828);
nand_4 g12513(new_n14862, new_n14861, new_n14826_1);
nand_4 g12514(new_n14863, new_n14862, new_n14824);
nand_4 g12515(new_n14864, new_n14863, new_n14822);
not_3  g12516(new_n14865, new_n14864);
nor_4  g12517(new_n14866, new_n14865, new_n14821);
nor_4  g12518(new_n14867, new_n14866, new_n14819_1);
nor_4  g12519(new_n14868, new_n14867, new_n14817);
nor_4  g12520(new_n14869, new_n7255, n10018);
not_3  g12521(new_n14870, n10018);
nor_4  g12522(new_n14871, new_n7260, new_n14870);
nor_4  g12523(new_n14872, new_n7266, n2184);
not_3  g12524(new_n14873, n2184);
nor_4  g12525(new_n14874, new_n7263, new_n14873);
nor_4  g12526(new_n14875, new_n14874, new_n14872);
not_3  g12527(new_n14876, n3541);
nand_4 g12528(new_n14877, new_n7270, new_n14876);
xnor_3 g12529(new_n14878, new_n7270, n3541);
nand_4 g12530(new_n14879, new_n7276, new_n7561);
xnor_3 g12531(new_n14880, new_n7276, n16818);
not_3  g12532(new_n14881, n1269);
nand_4 g12533(new_n14882, new_n4445, new_n14881);
xor_3  g12534(new_n14883, new_n4445, new_n14881);
nor_4  g12535(new_n14884, new_n4448, n14576);
not_3  g12536(new_n14885, new_n14884);
xor_3  g12537(new_n14886, new_n13918, new_n7562);
not_3  g12538(new_n14887, n2985);
nor_4  g12539(new_n14888, new_n4454, new_n14887);
xnor_3 g12540(new_n14889, new_n4454, new_n14887);
nand_4 g12541(new_n14890, new_n4465, new_n7563);
not_3  g12542(new_n14891_1, n15652);
nor_4  g12543(new_n14892, new_n4472, new_n14891_1);
nand_4 g12544(new_n14893, new_n4461, n4939);
xnor_3 g12545(new_n14894, new_n4471, n15652);
nor_4  g12546(new_n14895, new_n14894, new_n14893);
nor_4  g12547(new_n14896, new_n14895, new_n14892);
not_3  g12548(new_n14897, new_n14890);
nor_4  g12549(new_n14898, new_n4465, new_n7563);
nor_4  g12550(new_n14899_1, new_n14898, new_n14897);
nand_4 g12551(new_n14900, new_n14899_1, new_n14896);
nand_4 g12552(new_n14901, new_n14900, new_n14890);
nor_4  g12553(new_n14902, new_n14901, new_n14889);
nor_4  g12554(new_n14903, new_n14902, new_n14888);
nand_4 g12555(new_n14904, new_n14903, new_n14886);
nand_4 g12556(new_n14905, new_n14904, new_n14885);
nand_4 g12557(new_n14906, new_n14905, new_n14883);
nand_4 g12558(new_n14907, new_n14906, new_n14882);
nand_4 g12559(new_n14908, new_n14907, new_n14880);
nand_4 g12560(new_n14909, new_n14908, new_n14879);
nand_4 g12561(new_n14910, new_n14909, new_n14878);
nand_4 g12562(new_n14911, new_n14910, new_n14877);
nand_4 g12563(new_n14912, new_n14911, new_n14875);
not_3  g12564(new_n14913, new_n14912);
nor_4  g12565(new_n14914, new_n14913, new_n14872);
nor_4  g12566(new_n14915, new_n14914, new_n14871);
xnor_3 g12567(new_n14916, new_n14915, new_n7259);
nor_4  g12568(new_n14917, new_n14916, new_n14869);
nand_4 g12569(new_n14918, new_n14917, new_n7247);
nor_4  g12570(new_n14919, new_n14917, new_n7247);
not_3  g12571(new_n14920, new_n14919);
nand_4 g12572(new_n14921, new_n14920, new_n14918);
nor_4  g12573(new_n14922, new_n14871, new_n14869);
xnor_3 g12574(new_n14923, new_n14922, new_n14914);
not_3  g12575(new_n14924, new_n14923);
nand_4 g12576(new_n14925, new_n14924, new_n7307);
xnor_3 g12577(new_n14926, new_n14923, new_n7307);
xor_3  g12578(new_n14927, new_n7304, new_n7300);
xnor_3 g12579(new_n14928, new_n14911, new_n14875);
nand_4 g12580(new_n14929, new_n14928, new_n14927);
xnor_3 g12581(new_n14930, new_n14928, new_n14927);
not_3  g12582(new_n14931_1, new_n14930);
xor_3  g12583(new_n14932, new_n7302, new_n7301);
xnor_3 g12584(new_n14933, new_n14909, new_n14878);
nand_4 g12585(new_n14934, new_n14933, new_n14932);
xnor_3 g12586(new_n14935, new_n14933, new_n7318);
xnor_3 g12587(new_n14936, new_n14907, new_n14880);
nand_4 g12588(new_n14937, new_n14936, new_n7326);
xnor_3 g12589(new_n14938, new_n14905, new_n14883);
nand_4 g12590(new_n14939, new_n14938, new_n7330_1);
xnor_3 g12591(new_n14940, new_n14938, new_n7332);
xnor_3 g12592(new_n14941, new_n7235, new_n7218);
xnor_3 g12593(new_n14942, new_n14903, new_n14886);
not_3  g12594(new_n14943, new_n14942);
nor_4  g12595(new_n14944_1, new_n14943, new_n14941);
not_3  g12596(new_n14945, new_n14944_1);
nor_4  g12597(new_n14946, new_n14942, new_n7335_1);
nor_4  g12598(new_n14947, new_n14946, new_n14944_1);
xnor_3 g12599(new_n14948, new_n14901, new_n14889);
nor_4  g12600(new_n14949, new_n14948, new_n7343);
not_3  g12601(new_n14950, new_n14900);
nor_4  g12602(new_n14951, new_n14899_1, new_n14896);
nor_4  g12603(new_n14952, new_n14951, new_n14950);
not_3  g12604(new_n14953, new_n14952);
nor_4  g12605(new_n14954_1, new_n14953, new_n7346_1);
not_3  g12606(new_n14955, new_n14954_1);
xnor_3 g12607(new_n14956, new_n14952, new_n7345);
not_3  g12608(new_n14957, new_n14956);
xnor_3 g12609(new_n14958, new_n14894, new_n14893);
not_3  g12610(new_n14959, new_n14958);
nor_4  g12611(new_n14960, new_n14959, new_n7351);
not_3  g12612(new_n14961, new_n14960);
xor_3  g12613(new_n14962, n19922, n4939);
nand_4 g12614(new_n14963, new_n14962, new_n7354);
not_3  g12615(new_n14964, new_n14963);
nor_4  g12616(new_n14965, new_n14958, new_n7357);
nor_4  g12617(new_n14966, new_n14965, new_n14960);
nand_4 g12618(new_n14967, new_n14966, new_n14964);
nand_4 g12619(new_n14968, new_n14967, new_n14961);
nand_4 g12620(new_n14969, new_n14968, new_n14957);
nand_4 g12621(new_n14970, new_n14969, new_n14955);
xnor_3 g12622(new_n14971, new_n14948, new_n7343);
nor_4  g12623(new_n14972, new_n14971, new_n14970);
nor_4  g12624(new_n14973, new_n14972, new_n14949);
not_3  g12625(new_n14974, new_n14973);
nand_4 g12626(new_n14975, new_n14974, new_n14947);
nand_4 g12627(new_n14976, new_n14975, new_n14945);
nand_4 g12628(new_n14977_1, new_n14976, new_n14940);
nand_4 g12629(new_n14978, new_n14977_1, new_n14939);
xnor_3 g12630(new_n14979, new_n14936, new_n7374);
nand_4 g12631(new_n14980, new_n14979, new_n14978);
nand_4 g12632(new_n14981, new_n14980, new_n14937);
nand_4 g12633(new_n14982, new_n14981, new_n14935);
nand_4 g12634(new_n14983, new_n14982, new_n14934);
nand_4 g12635(new_n14984, new_n14983, new_n14931_1);
nand_4 g12636(new_n14985, new_n14984, new_n14929);
nand_4 g12637(new_n14986, new_n14985, new_n14926);
nand_4 g12638(new_n14987, new_n14986, new_n14925);
xnor_3 g12639(new_n14988, new_n14987, new_n14921);
not_3  g12640(new_n14989_1, new_n14988);
nor_4  g12641(new_n14990, new_n14989_1, new_n14868);
not_3  g12642(new_n14991, new_n14990);
not_3  g12643(new_n14992, new_n14868);
nor_4  g12644(new_n14993, new_n14988, new_n14992);
nor_4  g12645(new_n14994, new_n14993, new_n14990);
xor_3  g12646(new_n14995, new_n14866, new_n14819_1);
not_3  g12647(new_n14996, new_n14926);
not_3  g12648(new_n14997, new_n14929);
not_3  g12649(new_n14998, new_n14983);
nor_4  g12650(new_n14999, new_n14998, new_n14930);
nor_4  g12651(new_n15000, new_n14999, new_n14997);
xnor_3 g12652(new_n15001, new_n15000, new_n14996);
nor_4  g12653(new_n15002_1, new_n15001, new_n14995);
not_3  g12654(new_n15003, new_n15002_1);
not_3  g12655(new_n15004_1, new_n14995);
xnor_3 g12656(new_n15005, new_n15001, new_n15004_1);
xnor_3 g12657(new_n15006, new_n14863, new_n14822);
not_3  g12658(new_n15007, new_n15006);
xnor_3 g12659(new_n15008, new_n14983, new_n14931_1);
nor_4  g12660(new_n15009, new_n15008, new_n15007);
not_3  g12661(new_n15010, new_n15009);
xnor_3 g12662(new_n15011_1, new_n15008, new_n15006);
xnor_3 g12663(new_n15012, new_n14861, new_n14826_1);
xnor_3 g12664(new_n15013, new_n14981, new_n14935);
not_3  g12665(new_n15014, new_n15013);
nand_4 g12666(new_n15015, new_n15014, new_n15012);
xnor_3 g12667(new_n15016, new_n15013, new_n15012);
xnor_3 g12668(new_n15017, new_n14859, new_n14830);
not_3  g12669(new_n15018, new_n14979);
xnor_3 g12670(new_n15019_1, new_n15018, new_n14978);
nand_4 g12671(new_n15020, new_n15019_1, new_n15017);
not_3  g12672(new_n15021, new_n15017);
xnor_3 g12673(new_n15022, new_n15019_1, new_n15021);
xnor_3 g12674(new_n15023, new_n14857, new_n14833);
not_3  g12675(new_n15024, new_n14940);
xnor_3 g12676(new_n15025, new_n14976, new_n15024);
nand_4 g12677(new_n15026, new_n15025, new_n15023);
not_3  g12678(new_n15027, new_n15023);
xnor_3 g12679(new_n15028, new_n15025, new_n15027);
not_3  g12680(new_n15029, new_n14855);
xnor_3 g12681(new_n15030, new_n15029, new_n14837);
xnor_3 g12682(new_n15031_1, new_n14974, new_n14947);
nor_4  g12683(new_n15032, new_n15031_1, new_n15030);
not_3  g12684(new_n15033_1, new_n15032);
not_3  g12685(new_n15034, new_n15030);
xnor_3 g12686(new_n15035, new_n14973, new_n14947);
nor_4  g12687(new_n15036, new_n15035, new_n15034);
nor_4  g12688(new_n15037, new_n15036, new_n15032);
not_3  g12689(new_n15038, new_n14854);
nor_4  g12690(new_n15039, new_n14853, new_n14841);
nor_4  g12691(new_n15040, new_n15039, new_n15038);
not_3  g12692(new_n15041, new_n15040);
not_3  g12693(new_n15042, new_n14971);
xnor_3 g12694(new_n15043, new_n15042, new_n14970);
nand_4 g12695(new_n15044, new_n15043, new_n15041);
xnor_3 g12696(new_n15045, new_n15043, new_n15040);
xnor_3 g12697(new_n15046, new_n14968, new_n14956);
nor_4  g12698(new_n15047, new_n14844, new_n14843);
not_3  g12699(new_n15048, new_n15047);
xnor_3 g12700(new_n15049, new_n15048, new_n14851);
nor_4  g12701(new_n15050, new_n15049, new_n15046);
not_3  g12702(new_n15051, new_n15050);
not_3  g12703(new_n15052_1, new_n15046);
not_3  g12704(new_n15053_1, new_n15049);
nor_4  g12705(new_n15054, new_n15053_1, new_n15052_1);
nor_4  g12706(new_n15055, new_n15054, new_n15050);
xnor_3 g12707(new_n15056, new_n14962, new_n7354);
xor_3  g12708(new_n15057, n20385, new_n14848);
nor_4  g12709(new_n15058, new_n15057, new_n15056);
not_3  g12710(new_n15059, new_n14849_1);
nor_4  g12711(new_n15060, new_n14847, new_n14846);
xnor_3 g12712(new_n15061, new_n15060, new_n15059);
nor_4  g12713(new_n15062, new_n15061, new_n15058);
not_3  g12714(new_n15063, new_n15062);
xnor_3 g12715(new_n15064, new_n14966, new_n14964);
not_3  g12716(new_n15065, new_n15058);
not_3  g12717(new_n15066, new_n15061);
xor_3  g12718(new_n15067, new_n15066, new_n15065);
nand_4 g12719(new_n15068, new_n15067, new_n15064);
nand_4 g12720(new_n15069, new_n15068, new_n15063);
nand_4 g12721(new_n15070, new_n15069, new_n15055);
nand_4 g12722(new_n15071, new_n15070, new_n15051);
nand_4 g12723(new_n15072, new_n15071, new_n15045);
nand_4 g12724(new_n15073, new_n15072, new_n15044);
nand_4 g12725(new_n15074, new_n15073, new_n15037);
nand_4 g12726(new_n15075, new_n15074, new_n15033_1);
nand_4 g12727(new_n15076, new_n15075, new_n15028);
nand_4 g12728(new_n15077_1, new_n15076, new_n15026);
nand_4 g12729(new_n15078, new_n15077_1, new_n15022);
nand_4 g12730(new_n15079, new_n15078, new_n15020);
nand_4 g12731(new_n15080, new_n15079, new_n15016);
nand_4 g12732(new_n15081, new_n15080, new_n15015);
nand_4 g12733(new_n15082_1, new_n15081, new_n15011_1);
nand_4 g12734(new_n15083, new_n15082_1, new_n15010);
nand_4 g12735(new_n15084, new_n15083, new_n15005);
nand_4 g12736(new_n15085, new_n15084, new_n15003);
nand_4 g12737(new_n15086, new_n15085, new_n14994);
nand_4 g12738(new_n15087, new_n15086, new_n14991);
not_3  g12739(new_n15088, new_n15087);
and_4  g12740(new_n15089, new_n14915, new_n7258);
not_3  g12741(new_n15090, new_n15089);
not_3  g12742(new_n15091, new_n14987);
nand_4 g12743(new_n15092, new_n15091, new_n14918);
nand_4 g12744(new_n15093, new_n15092, new_n15090);
nor_4  g12745(new_n15094_1, new_n15093, new_n14919);
not_3  g12746(new_n15095, new_n15094_1);
nor_4  g12747(n2007, new_n15095, new_n15088);
not_3  g12748(new_n15097, new_n10648);
xor_3  g12749(n2061, new_n15097, new_n10632);
xnor_3 g12750(new_n15099, new_n13606, new_n8395);
nand_4 g12751(new_n15100, new_n13615, new_n8402);
xnor_3 g12752(new_n15101, new_n13615, new_n8401);
nand_4 g12753(new_n15102, new_n13623, new_n8408_1);
nand_4 g12754(new_n15103, new_n8414, new_n5286);
xnor_3 g12755(new_n15104, new_n8414, new_n5320);
nand_4 g12756(new_n15105, new_n8420, new_n5323);
xnor_3 g12757(new_n15106, new_n8420, new_n5327);
not_3  g12758(new_n15107, new_n5332);
nand_4 g12759(new_n15108, new_n8424, new_n15107);
nand_4 g12760(new_n15109, new_n8429, new_n5346);
xnor_3 g12761(new_n15110, new_n8428, new_n5346);
nor_4  g12762(new_n15111, new_n8435, new_n5357);
not_3  g12763(new_n15112, new_n15111);
nor_4  g12764(new_n15113, new_n15112, new_n5351_1);
xor_3  g12765(new_n15114, new_n15112, new_n5360);
nor_4  g12766(new_n15115, new_n15114, new_n8443);
nor_4  g12767(new_n15116, new_n15115, new_n15113);
nand_4 g12768(new_n15117, new_n15116, new_n15110);
nand_4 g12769(new_n15118_1, new_n15117, new_n15109);
xnor_3 g12770(new_n15119, new_n8424, new_n5332);
nand_4 g12771(new_n15120, new_n15119, new_n15118_1);
nand_4 g12772(new_n15121, new_n15120, new_n15108);
nand_4 g12773(new_n15122, new_n15121, new_n15106);
nand_4 g12774(new_n15123, new_n15122, new_n15105);
nand_4 g12775(new_n15124, new_n15123, new_n15104);
nand_4 g12776(new_n15125, new_n15124, new_n15103);
xnor_3 g12777(new_n15126, new_n13623, new_n8407);
nand_4 g12778(new_n15127, new_n15126, new_n15125);
nand_4 g12779(new_n15128_1, new_n15127, new_n15102);
nand_4 g12780(new_n15129, new_n15128_1, new_n15101);
nand_4 g12781(new_n15130, new_n15129, new_n15100);
not_3  g12782(new_n15131, new_n15130);
xor_3  g12783(n2092, new_n15131, new_n15099);
xor_3  g12784(new_n15133, n22253, n10650);
nor_4  g12785(new_n15134, n12900, n1255);
xor_3  g12786(new_n15135, n12900, n1255);
not_3  g12787(new_n15136, new_n15135);
nor_4  g12788(new_n15137, n20411, n9512);
xor_3  g12789(new_n15138, n20411, n9512);
not_3  g12790(new_n15139_1, new_n15138);
not_3  g12791(new_n15140, n17069);
nand_4 g12792(new_n15141, new_n15140, new_n8257);
xor_3  g12793(new_n15142, n17069, n16608);
nor_4  g12794(new_n15143, n21735, n15918);
not_3  g12795(new_n15144, new_n15143);
xor_3  g12796(new_n15145_1, n21735, n15918);
nor_4  g12797(new_n15146_1, n24085, n17784);
not_3  g12798(new_n15147, new_n15146_1);
xor_3  g12799(new_n15148, n24085, n17784);
nor_4  g12800(new_n15149, n14323, n14071);
not_3  g12801(new_n15150, new_n15149);
xor_3  g12802(new_n15151, n14323, n14071);
nor_4  g12803(new_n15152, n2886, n1738);
not_3  g12804(new_n15153, new_n15152);
xor_3  g12805(new_n15154, n2886, n1738);
nor_4  g12806(new_n15155, n12152, n1040);
not_3  g12807(new_n15156, new_n15155);
nand_4 g12808(new_n15157, n19107, n9090);
nand_4 g12809(new_n15158, n12152, n1040);
not_3  g12810(new_n15159, new_n15158);
nor_4  g12811(new_n15160, new_n15159, new_n15155);
nand_4 g12812(new_n15161, new_n15160, new_n15157);
nand_4 g12813(new_n15162, new_n15161, new_n15156);
nand_4 g12814(new_n15163, new_n15162, new_n15154);
nand_4 g12815(new_n15164, new_n15163, new_n15153);
nand_4 g12816(new_n15165_1, new_n15164, new_n15151);
nand_4 g12817(new_n15166, new_n15165_1, new_n15150);
nand_4 g12818(new_n15167_1, new_n15166, new_n15148);
nand_4 g12819(new_n15168, new_n15167_1, new_n15147);
nand_4 g12820(new_n15169, new_n15168, new_n15145_1);
nand_4 g12821(new_n15170, new_n15169, new_n15144);
nand_4 g12822(new_n15171, new_n15170, new_n15142);
nand_4 g12823(new_n15172, new_n15171, new_n15141);
not_3  g12824(new_n15173, new_n15172);
nor_4  g12825(new_n15174, new_n15173, new_n15139_1);
nor_4  g12826(new_n15175, new_n15174, new_n15137);
nor_4  g12827(new_n15176_1, new_n15175, new_n15136);
nor_4  g12828(new_n15177, new_n15176_1, new_n15134);
xor_3  g12829(new_n15178, new_n15177, new_n15133);
nor_4  g12830(new_n15179, new_n15178, new_n8200);
not_3  g12831(new_n15180_1, new_n15133);
nor_4  g12832(new_n15181, new_n15177, new_n15180_1);
and_4  g12833(new_n15182_1, new_n15177, new_n15180_1);
nor_4  g12834(new_n15183, new_n15182_1, new_n15181);
xnor_3 g12835(new_n15184, new_n15183, n2272);
and_4  g12836(new_n15185, new_n15175, new_n15136);
nor_4  g12837(new_n15186, new_n15185, new_n15176_1);
not_3  g12838(new_n15187, new_n15186);
nor_4  g12839(new_n15188, new_n15187, new_n8203);
xnor_3 g12840(new_n15189, new_n15186, n25331);
not_3  g12841(new_n15190, n18483);
xnor_3 g12842(new_n15191, new_n15172, new_n15138);
nor_4  g12843(new_n15192, new_n15191, new_n15190);
not_3  g12844(new_n15193, new_n15191);
nor_4  g12845(new_n15194, new_n15193, n18483);
nor_4  g12846(new_n15195, new_n15194, new_n15192);
not_3  g12847(new_n15196, new_n15170);
xnor_3 g12848(new_n15197, new_n15196, new_n15142);
nand_4 g12849(new_n15198, new_n15197, n21934);
xnor_3 g12850(new_n15199, new_n15197, new_n8210);
xnor_3 g12851(new_n15200, new_n15168, new_n15145_1);
nor_4  g12852(new_n15201, new_n15200, new_n8214);
not_3  g12853(new_n15202, new_n15201);
not_3  g12854(new_n15203, new_n15200);
nor_4  g12855(new_n15204, new_n15203, n18901);
nor_4  g12856(new_n15205_1, new_n15204, new_n15201);
xnor_3 g12857(new_n15206, new_n15166, new_n15148);
nor_4  g12858(new_n15207, new_n15206, new_n8218);
not_3  g12859(new_n15208, new_n15207);
not_3  g12860(new_n15209, new_n15206);
nor_4  g12861(new_n15210, new_n15209, n4376);
nor_4  g12862(new_n15211, new_n15210, new_n15207);
not_3  g12863(new_n15212, new_n15151);
xnor_3 g12864(new_n15213, new_n15164, new_n15212);
nand_4 g12865(new_n15214, new_n15213, n14570);
xnor_3 g12866(new_n15215, new_n15213, new_n8222);
not_3  g12867(new_n15216, new_n15162);
xnor_3 g12868(new_n15217, new_n15216, new_n15154);
nand_4 g12869(new_n15218, new_n15217, n23775);
not_3  g12870(new_n15219, new_n15218);
nor_4  g12871(new_n15220, new_n15217, n23775);
nor_4  g12872(new_n15221, new_n15220, new_n15219);
xnor_3 g12873(new_n15222, n19107, n9090);
nand_4 g12874(new_n15223, new_n15222, n11479);
nand_4 g12875(new_n15224, new_n15223, new_n8229);
not_3  g12876(new_n15225, new_n15224);
xor_3  g12877(new_n15226, new_n15160, new_n15157);
xor_3  g12878(new_n15227, new_n15223, n8259);
nor_4  g12879(new_n15228, new_n15227, new_n15226);
nor_4  g12880(new_n15229, new_n15228, new_n15225);
nand_4 g12881(new_n15230_1, new_n15229, new_n15221);
nand_4 g12882(new_n15231, new_n15230_1, new_n15218);
nand_4 g12883(new_n15232, new_n15231, new_n15215);
nand_4 g12884(new_n15233, new_n15232, new_n15214);
nand_4 g12885(new_n15234, new_n15233, new_n15211);
nand_4 g12886(new_n15235, new_n15234, new_n15208);
nand_4 g12887(new_n15236, new_n15235, new_n15205_1);
nand_4 g12888(new_n15237, new_n15236, new_n15202);
nand_4 g12889(new_n15238, new_n15237, new_n15199);
nand_4 g12890(new_n15239, new_n15238, new_n15198);
nand_4 g12891(new_n15240, new_n15239, new_n15195);
not_3  g12892(new_n15241_1, new_n15240);
nor_4  g12893(new_n15242, new_n15241_1, new_n15192);
nor_4  g12894(new_n15243, new_n15242, new_n15189);
nor_4  g12895(new_n15244, new_n15243, new_n15188);
nor_4  g12896(new_n15245, new_n15244, new_n15184);
nor_4  g12897(new_n15246, new_n15245, new_n15179);
nor_4  g12898(new_n15247, n22253, n10650);
nor_4  g12899(new_n15248, new_n15181, new_n15247);
nor_4  g12900(new_n15249, new_n15248, new_n15246);
not_3  g12901(new_n15250, n9934);
nor_4  g12902(new_n15251, n7876, n4964);
nand_4 g12903(new_n15252, new_n15251, new_n4107);
nor_4  g12904(new_n15253, new_n15252, n342);
not_3  g12905(new_n15254, new_n15253);
nor_4  g12906(new_n15255_1, new_n15254, n26107);
not_3  g12907(new_n15256, new_n15255_1);
nor_4  g12908(new_n15257, new_n15256, n22597);
not_3  g12909(new_n15258_1, new_n15257);
nor_4  g12910(new_n15259, new_n15258_1, n19327);
not_3  g12911(new_n15260, new_n15259);
nor_4  g12912(new_n15261, new_n15260, n26224);
not_3  g12913(new_n15262, new_n15261);
nor_4  g12914(new_n15263, new_n15262, n18496);
xor_3  g12915(new_n15264, new_n15263, new_n15250);
not_3  g12916(new_n15265, new_n15264);
nor_4  g12917(new_n15266, n18409, n5704);
nand_4 g12918(new_n15267, new_n15266, new_n4201);
nor_4  g12919(new_n15268, new_n15267, n19911);
nand_4 g12920(new_n15269, new_n15268, new_n4190);
nor_4  g12921(new_n15270, new_n15269, n18907);
nand_4 g12922(new_n15271_1, new_n15270, new_n4185);
nor_4  g12923(new_n15272, new_n15271_1, n4256);
not_3  g12924(new_n15273, new_n15272);
xor_3  g12925(new_n15274, new_n15273, n21287);
nor_4  g12926(new_n15275_1, new_n15274, n12861);
not_3  g12927(new_n15276, new_n15274);
xor_3  g12928(new_n15277, new_n15276, n12861);
xor_3  g12929(new_n15278, new_n15271_1, n4256);
nor_4  g12930(new_n15279, new_n15278, n13333);
not_3  g12931(new_n15280, new_n15278);
xor_3  g12932(new_n15281, new_n15280, n13333);
xor_3  g12933(new_n15282, new_n15270, new_n4185);
nor_4  g12934(new_n15283, new_n15282, n2210);
not_3  g12935(new_n15284, new_n15282);
xor_3  g12936(new_n15285, new_n15284, n2210);
xor_3  g12937(new_n15286, new_n15269, n18907);
nor_4  g12938(new_n15287, new_n15286, n20604);
not_3  g12939(new_n15288, new_n15286);
xor_3  g12940(new_n15289_1, new_n15288, n20604);
xnor_3 g12941(new_n15290, new_n15268, n2731);
nor_4  g12942(new_n15291, new_n15290, n16158);
not_3  g12943(new_n15292, new_n15290);
nor_4  g12944(new_n15293, new_n15292, new_n5234);
nor_4  g12945(new_n15294, new_n15293, new_n15291);
nand_4 g12946(new_n15295, new_n15267, n19911);
not_3  g12947(new_n15296, new_n15295);
nor_4  g12948(new_n15297, new_n15296, new_n15268);
nor_4  g12949(new_n15298, new_n15297, n5752);
not_3  g12950(new_n15299, new_n15298);
xnor_3 g12951(new_n15300_1, new_n15266, n13708);
nor_4  g12952(new_n15301, new_n15300_1, n18171);
not_3  g12953(new_n15302, new_n15301);
not_3  g12954(new_n15303, new_n15300_1);
nor_4  g12955(new_n15304, new_n15303, new_n5240);
nor_4  g12956(new_n15305, new_n15304, new_n15301);
xnor_3 g12957(new_n15306, n18409, n5704);
nand_4 g12958(new_n15307_1, new_n15306, new_n5244);
nand_4 g12959(new_n15308, n22309, n5704);
xnor_3 g12960(new_n15309, new_n15306, n25073);
nand_4 g12961(new_n15310, new_n15309, new_n15308);
nand_4 g12962(new_n15311, new_n15310, new_n15307_1);
nand_4 g12963(new_n15312, new_n15311, new_n15305);
nand_4 g12964(new_n15313, new_n15312, new_n15302);
not_3  g12965(new_n15314, n5752);
not_3  g12966(new_n15315, new_n15297);
nor_4  g12967(new_n15316, new_n15315, new_n15314);
nor_4  g12968(new_n15317, new_n15316, new_n15298);
nand_4 g12969(new_n15318, new_n15317, new_n15313);
nand_4 g12970(new_n15319, new_n15318, new_n15299);
nand_4 g12971(new_n15320, new_n15319, new_n15294);
not_3  g12972(new_n15321, new_n15320);
nor_4  g12973(new_n15322, new_n15321, new_n15291);
nor_4  g12974(new_n15323, new_n15322, new_n15289_1);
nor_4  g12975(new_n15324, new_n15323, new_n15287);
nor_4  g12976(new_n15325, new_n15324, new_n15285);
nor_4  g12977(new_n15326, new_n15325, new_n15283);
nor_4  g12978(new_n15327_1, new_n15326, new_n15281);
nor_4  g12979(new_n15328, new_n15327_1, new_n15279);
nor_4  g12980(new_n15329, new_n15328, new_n15277);
nor_4  g12981(new_n15330, new_n15329, new_n15275_1);
not_3  g12982(new_n15331, n8305);
nor_4  g12983(new_n15332_1, new_n15273, n21287);
xor_3  g12984(new_n15333, new_n15332_1, new_n8547);
not_3  g12985(new_n15334, new_n15333);
nor_4  g12986(new_n15335, new_n15334, new_n15331);
nor_4  g12987(new_n15336, new_n15333, n8305);
nor_4  g12988(new_n15337, new_n15336, new_n15335);
xnor_3 g12989(new_n15338, new_n15337, new_n15330);
nor_4  g12990(new_n15339, new_n15338, new_n15265);
not_3  g12991(new_n15340, new_n15339);
xnor_3 g12992(new_n15341, new_n15338, new_n15265);
not_3  g12993(new_n15342, new_n15341);
not_3  g12994(new_n15343, n18496);
xor_3  g12995(new_n15344, new_n15261, new_n15343);
not_3  g12996(new_n15345_1, new_n15344);
not_3  g12997(new_n15346, new_n15328);
xnor_3 g12998(new_n15347, new_n15346, new_n15277);
nor_4  g12999(new_n15348, new_n15347, new_n15345_1);
not_3  g13000(new_n15349, new_n15348);
xnor_3 g13001(new_n15350, new_n15347, new_n15345_1);
not_3  g13002(new_n15351, new_n15350);
not_3  g13003(new_n15352, n26224);
xor_3  g13004(new_n15353_1, new_n15259, new_n15352);
not_3  g13005(new_n15354, new_n15353_1);
not_3  g13006(new_n15355, new_n15326);
xnor_3 g13007(new_n15356, new_n15355, new_n15281);
nor_4  g13008(new_n15357, new_n15356, new_n15354);
not_3  g13009(new_n15358, new_n15357);
xnor_3 g13010(new_n15359, new_n15356, new_n15354);
not_3  g13011(new_n15360, new_n15359);
xor_3  g13012(new_n15361, new_n15257, new_n5426);
xnor_3 g13013(new_n15362, new_n15324, new_n15285);
nand_4 g13014(new_n15363, new_n15362, new_n15361);
xnor_3 g13015(new_n15364, new_n15362, new_n15361);
not_3  g13016(new_n15365, new_n15364);
xor_3  g13017(new_n15366_1, new_n15255_1, n22597);
not_3  g13018(new_n15367, new_n15322);
xnor_3 g13019(new_n15368, new_n15367, new_n15289_1);
nor_4  g13020(new_n15369, new_n15368, new_n15366_1);
not_3  g13021(new_n15370, new_n15369);
xnor_3 g13022(new_n15371, new_n15368, new_n15366_1);
not_3  g13023(new_n15372, new_n15371);
xor_3  g13024(new_n15373, new_n15253, new_n4093);
xnor_3 g13025(new_n15374, new_n15319, new_n15294);
nand_4 g13026(new_n15375, new_n15374, new_n15373);
not_3  g13027(new_n15376, new_n15374);
xnor_3 g13028(new_n15377, new_n15376, new_n15373);
xor_3  g13029(new_n15378_1, new_n15252, new_n4123_1);
xnor_3 g13030(new_n15379, new_n15317, new_n15313);
not_3  g13031(new_n15380, new_n15379);
nor_4  g13032(new_n15381, new_n15380, new_n15378_1);
not_3  g13033(new_n15382_1, new_n15381);
not_3  g13034(new_n15383, new_n15378_1);
nor_4  g13035(new_n15384, new_n15379, new_n15383);
nor_4  g13036(new_n15385, new_n15384, new_n15381);
xnor_3 g13037(new_n15386, new_n15311, new_n15305);
xor_3  g13038(new_n15387, new_n15251, new_n4107);
nand_4 g13039(new_n15388, new_n15387, new_n15386);
not_3  g13040(new_n15389, new_n15386);
xnor_3 g13041(new_n15390, new_n15387, new_n15389);
xor_3  g13042(new_n15391, n7876, n4964);
xnor_3 g13043(new_n15392, new_n15309, new_n15308);
nand_4 g13044(new_n15393, new_n15392, new_n15391);
xor_3  g13045(new_n15394, n22309, n5704);
not_3  g13046(new_n15395, new_n15394);
nor_4  g13047(new_n15396, new_n15395, new_n4168);
not_3  g13048(new_n15397, new_n15392);
xnor_3 g13049(new_n15398, new_n15397, new_n15391);
nand_4 g13050(new_n15399, new_n15398, new_n15396);
nand_4 g13051(new_n15400, new_n15399, new_n15393);
nand_4 g13052(new_n15401, new_n15400, new_n15390);
nand_4 g13053(new_n15402, new_n15401, new_n15388);
nand_4 g13054(new_n15403, new_n15402, new_n15385);
nand_4 g13055(new_n15404, new_n15403, new_n15382_1);
nand_4 g13056(new_n15405, new_n15404, new_n15377);
nand_4 g13057(new_n15406, new_n15405, new_n15375);
nand_4 g13058(new_n15407_1, new_n15406, new_n15372);
nand_4 g13059(new_n15408, new_n15407_1, new_n15370);
nand_4 g13060(new_n15409, new_n15408, new_n15365);
nand_4 g13061(new_n15410, new_n15409, new_n15363);
nand_4 g13062(new_n15411, new_n15410, new_n15360);
nand_4 g13063(new_n15412, new_n15411, new_n15358);
nand_4 g13064(new_n15413, new_n15412, new_n15351);
nand_4 g13065(new_n15414, new_n15413, new_n15349);
nand_4 g13066(new_n15415, new_n15414, new_n15342);
nand_4 g13067(new_n15416, new_n15415, new_n15340);
not_3  g13068(new_n15417, new_n15263);
nor_4  g13069(new_n15418, new_n15417, n9934);
not_3  g13070(new_n15419, new_n15336);
nand_4 g13071(new_n15420, new_n15419, new_n15330);
not_3  g13072(new_n15421, new_n15332_1);
nor_4  g13073(new_n15422, new_n15421, n26986);
nor_4  g13074(new_n15423, new_n15335, new_n15422);
nand_4 g13075(new_n15424_1, new_n15423, new_n15420);
not_3  g13076(new_n15425, new_n15424_1);
nor_4  g13077(new_n15426, new_n15425, new_n15418);
not_3  g13078(new_n15427, new_n15426);
nor_4  g13079(new_n15428_1, new_n15427, new_n15416);
not_3  g13080(new_n15429, new_n15428_1);
xnor_3 g13081(new_n15430, new_n15429, new_n15249);
xnor_3 g13082(new_n15431, new_n15248, new_n15246);
not_3  g13083(new_n15432, new_n15418);
nor_4  g13084(new_n15433, new_n15424_1, new_n15432);
nor_4  g13085(new_n15434, new_n15433, new_n15426);
xnor_3 g13086(new_n15435_1, new_n15434, new_n15416);
nor_4  g13087(new_n15436, new_n15435_1, new_n15431);
not_3  g13088(new_n15437, new_n15436);
not_3  g13089(new_n15438_1, new_n15431);
not_3  g13090(new_n15439, new_n15435_1);
nor_4  g13091(new_n15440, new_n15439, new_n15438_1);
nor_4  g13092(new_n15441, new_n15440, new_n15436);
xnor_3 g13093(new_n15442, new_n15244, new_n15184);
xnor_3 g13094(new_n15443, new_n15414, new_n15341);
nor_4  g13095(new_n15444, new_n15443, new_n15442);
not_3  g13096(new_n15445, new_n15444);
xnor_3 g13097(new_n15446, new_n15443, new_n15442);
not_3  g13098(new_n15447, new_n15446);
not_3  g13099(new_n15448, new_n15192);
nand_4 g13100(new_n15449, new_n15240, new_n15448);
xnor_3 g13101(new_n15450, new_n15449, new_n15189);
not_3  g13102(new_n15451, new_n15450);
xnor_3 g13103(new_n15452, new_n15412, new_n15350);
nor_4  g13104(new_n15453, new_n15452, new_n15451);
not_3  g13105(new_n15454, new_n15453);
not_3  g13106(new_n15455, new_n15452);
xnor_3 g13107(new_n15456, new_n15455, new_n15450);
xnor_3 g13108(new_n15457, new_n15239, new_n15195);
xnor_3 g13109(new_n15458, new_n15410, new_n15360);
not_3  g13110(new_n15459, new_n15458);
nor_4  g13111(new_n15460, new_n15459, new_n15457);
not_3  g13112(new_n15461, new_n15457);
xnor_3 g13113(new_n15462, new_n15458, new_n15461);
xnor_3 g13114(new_n15463, new_n15237, new_n15199);
xnor_3 g13115(new_n15464, new_n15408, new_n15364);
nor_4  g13116(new_n15465_1, new_n15464, new_n15463);
xnor_3 g13117(new_n15466, new_n15464, new_n15463);
xnor_3 g13118(new_n15467_1, new_n15235, new_n15205_1);
not_3  g13119(new_n15468, new_n15467_1);
xnor_3 g13120(new_n15469, new_n15406, new_n15372);
nand_4 g13121(new_n15470_1, new_n15469, new_n15468);
xnor_3 g13122(new_n15471, new_n15469, new_n15467_1);
not_3  g13123(new_n15472, new_n15211);
xnor_3 g13124(new_n15473, new_n15233, new_n15472);
xnor_3 g13125(new_n15474, new_n15404, new_n15377);
nand_4 g13126(new_n15475, new_n15474, new_n15473);
not_3  g13127(new_n15476, new_n15474);
xnor_3 g13128(new_n15477_1, new_n15476, new_n15473);
xnor_3 g13129(new_n15478, new_n15231, new_n15215);
not_3  g13130(new_n15479, new_n15478);
xnor_3 g13131(new_n15480, new_n15402, new_n15385);
nand_4 g13132(new_n15481_1, new_n15480, new_n15479);
xnor_3 g13133(new_n15482, new_n15480, new_n15478);
not_3  g13134(new_n15483, new_n15221);
xnor_3 g13135(new_n15484, new_n15229, new_n15483);
not_3  g13136(new_n15485, new_n15390);
xnor_3 g13137(new_n15486, new_n15400, new_n15485);
not_3  g13138(new_n15487, new_n15486);
nand_4 g13139(new_n15488, new_n15487, new_n15484);
xnor_3 g13140(new_n15489, new_n15486, new_n15484);
xnor_3 g13141(new_n15490_1, new_n15398, new_n15396);
xnor_3 g13142(new_n15491, new_n15227, new_n15226);
nor_4  g13143(new_n15492, new_n15491, new_n15490_1);
xor_3  g13144(new_n15493, new_n15222, n11479);
not_3  g13145(new_n15494, new_n15493);
nor_4  g13146(new_n15495, new_n15394, n7876);
nor_4  g13147(new_n15496_1, new_n15495, new_n15396);
nand_4 g13148(new_n15497, new_n15496_1, new_n15494);
xnor_3 g13149(new_n15498, new_n15491, new_n15490_1);
nor_4  g13150(new_n15499, new_n15498, new_n15497);
nor_4  g13151(new_n15500, new_n15499, new_n15492);
nand_4 g13152(new_n15501_1, new_n15500, new_n15489);
nand_4 g13153(new_n15502, new_n15501_1, new_n15488);
nand_4 g13154(new_n15503, new_n15502, new_n15482);
nand_4 g13155(new_n15504, new_n15503, new_n15481_1);
nand_4 g13156(new_n15505, new_n15504, new_n15477_1);
nand_4 g13157(new_n15506_1, new_n15505, new_n15475);
nand_4 g13158(new_n15507, new_n15506_1, new_n15471);
nand_4 g13159(new_n15508_1, new_n15507, new_n15470_1);
not_3  g13160(new_n15509, new_n15508_1);
nor_4  g13161(new_n15510, new_n15509, new_n15466);
nor_4  g13162(new_n15511, new_n15510, new_n15465_1);
nor_4  g13163(new_n15512, new_n15511, new_n15462);
nor_4  g13164(new_n15513, new_n15512, new_n15460);
nor_4  g13165(new_n15514, new_n15513, new_n15456);
not_3  g13166(new_n15515, new_n15514);
nand_4 g13167(new_n15516, new_n15515, new_n15454);
nand_4 g13168(new_n15517, new_n15516, new_n15447);
nand_4 g13169(new_n15518, new_n15517, new_n15445);
nand_4 g13170(new_n15519, new_n15518, new_n15441);
nand_4 g13171(new_n15520, new_n15519, new_n15437);
xnor_3 g13172(n2095, new_n15520, new_n15430);
not_3  g13173(new_n15522, new_n13698);
xor_3  g13174(n2105, new_n15522, new_n13696);
not_3  g13175(new_n15524, new_n7126);
xor_3  g13176(new_n15525, n23166, n11898);
nand_4 g13177(new_n15526, n19941, n10577);
not_3  g13178(new_n15527, new_n15526);
nor_4  g13179(new_n15528, n19941, n10577);
nor_4  g13180(new_n15529, n6381, n1099);
not_3  g13181(new_n15530, new_n15529);
nand_4 g13182(new_n15531, new_n12687, new_n12669);
nand_4 g13183(new_n15532, new_n15531, new_n15530);
nor_4  g13184(new_n15533, new_n15532, new_n15528);
nor_4  g13185(new_n15534, new_n15533, new_n15527);
xnor_3 g13186(new_n15535, new_n15534, new_n15525);
not_3  g13187(new_n15536, new_n15535);
xor_3  g13188(new_n15537, new_n15536, n8827);
not_3  g13189(new_n15538, n18035);
not_3  g13190(new_n15539_1, new_n15532);
nor_4  g13191(new_n15540, new_n15528, new_n15527);
nor_4  g13192(new_n15541, new_n15540, new_n15539_1);
not_3  g13193(new_n15542, new_n15540);
nor_4  g13194(new_n15543, new_n15542, new_n15532);
nor_4  g13195(new_n15544, new_n15543, new_n15541);
not_3  g13196(new_n15545, new_n15544);
nor_4  g13197(new_n15546_1, new_n15545, new_n15538);
not_3  g13198(new_n15547, new_n15546_1);
nor_4  g13199(new_n15548, new_n15544, n18035);
nor_4  g13200(new_n15549, new_n15548, new_n15546_1);
nand_4 g13201(new_n15550, new_n12688, n5077);
nand_4 g13202(new_n15551, new_n12708, new_n12689);
nand_4 g13203(new_n15552, new_n15551, new_n15550);
nand_4 g13204(new_n15553, new_n15552, new_n15549);
nand_4 g13205(new_n15554, new_n15553, new_n15547);
xnor_3 g13206(new_n15555_1, new_n15554, new_n15537);
nor_4  g13207(new_n15556, new_n15555_1, new_n15524);
not_3  g13208(new_n15557, n8827);
xor_3  g13209(new_n15558_1, new_n15536, new_n15557);
xnor_3 g13210(new_n15559_1, new_n15554, new_n15558_1);
nor_4  g13211(new_n15560, new_n15559_1, new_n7126);
nor_4  g13212(new_n15561, new_n15560, new_n15556);
xnor_3 g13213(new_n15562, new_n15552, new_n15549);
nor_4  g13214(new_n15563, new_n15562, new_n7128);
not_3  g13215(new_n15564, new_n15563);
not_3  g13216(new_n15565, new_n7128);
not_3  g13217(new_n15566, new_n15562);
nor_4  g13218(new_n15567, new_n15566, new_n15565);
nor_4  g13219(new_n15568, new_n15567, new_n15563);
not_3  g13220(new_n15569, new_n7136);
nor_4  g13221(new_n15570_1, new_n12709, new_n15569);
not_3  g13222(new_n15571, new_n15570_1);
nor_4  g13223(new_n15572, new_n12710, new_n7136);
nor_4  g13224(new_n15573_1, new_n15572, new_n15570_1);
not_3  g13225(new_n15574, new_n7141);
nor_4  g13226(new_n15575, new_n12716, new_n15574);
not_3  g13227(new_n15576, new_n15575);
nor_4  g13228(new_n15577, new_n12717, new_n7141);
nor_4  g13229(new_n15578, new_n15577, new_n15575);
nand_4 g13230(new_n15579, new_n12722, new_n7150);
xnor_3 g13231(new_n15580, new_n12722, new_n7146);
nor_4  g13232(new_n15581, new_n12727_1, new_n7157);
not_3  g13233(new_n15582, new_n15581);
nor_4  g13234(new_n15583, new_n12728, new_n7155);
nor_4  g13235(new_n15584, new_n15583, new_n15581);
nand_4 g13236(new_n15585, new_n10104, new_n7161);
not_3  g13237(new_n15586, new_n7161);
xnor_3 g13238(new_n15587, new_n10104, new_n15586);
nand_4 g13239(new_n15588_1, new_n10074, new_n7169);
not_3  g13240(new_n15589, new_n15588_1);
nor_4  g13241(new_n15590_1, new_n10074, new_n7169);
nor_4  g13242(new_n15591, new_n15590_1, new_n15589);
not_3  g13243(new_n15592, new_n7175);
not_3  g13244(new_n15593, new_n10079);
nor_4  g13245(new_n15594, new_n15593, new_n15592);
not_3  g13246(new_n15595, new_n15594);
nor_4  g13247(new_n15596, new_n10083, new_n6771);
nor_4  g13248(new_n15597, new_n10079, new_n7175);
nor_4  g13249(new_n15598_1, new_n15597, new_n15594);
nand_4 g13250(new_n15599, new_n15598_1, new_n15596);
nand_4 g13251(new_n15600, new_n15599, new_n15595);
nand_4 g13252(new_n15601, new_n15600, new_n15591);
nand_4 g13253(new_n15602_1, new_n15601, new_n15588_1);
nand_4 g13254(new_n15603, new_n15602_1, new_n15587);
nand_4 g13255(new_n15604, new_n15603, new_n15585);
nand_4 g13256(new_n15605, new_n15604, new_n15584);
nand_4 g13257(new_n15606, new_n15605, new_n15582);
nand_4 g13258(new_n15607, new_n15606, new_n15580);
nand_4 g13259(new_n15608, new_n15607, new_n15579);
nand_4 g13260(new_n15609, new_n15608, new_n15578);
nand_4 g13261(new_n15610, new_n15609, new_n15576);
nand_4 g13262(new_n15611, new_n15610, new_n15573_1);
nand_4 g13263(new_n15612, new_n15611, new_n15571);
nand_4 g13264(new_n15613, new_n15612, new_n15568);
nand_4 g13265(new_n15614_1, new_n15613, new_n15564);
xnor_3 g13266(n2122, new_n15614_1, new_n15561);
not_3  g13267(new_n15616, new_n2971_1);
xor_3  g13268(n2147, new_n15616, new_n2941);
xor_3  g13269(n2209, new_n12631, new_n12582);
not_3  g13270(new_n15619, new_n6731);
xor_3  g13271(n2214, new_n15619, new_n6577);
nor_4  g13272(new_n15621, new_n13442, new_n4699);
not_3  g13273(new_n15622, new_n4699);
nor_4  g13274(new_n15623, new_n13413, new_n15622);
nor_4  g13275(new_n15624, new_n15623, new_n15621);
not_3  g13276(new_n15625, new_n4823);
nor_4  g13277(new_n15626, new_n13416, new_n15625);
xnor_3 g13278(new_n15627, new_n13416, new_n15625);
nor_4  g13279(new_n15628, new_n13424_1, new_n4829);
not_3  g13280(new_n15629, new_n15628);
nor_4  g13281(new_n15630, new_n13435, new_n4828);
nor_4  g13282(new_n15631, new_n15630, new_n15628);
nor_4  g13283(new_n15632, new_n13430, new_n4837);
nor_4  g13284(new_n15633, new_n13426, new_n4840);
xnor_3 g13285(new_n15634, new_n13430, new_n4837);
nor_4  g13286(new_n15635, new_n15634, new_n15633);
nor_4  g13287(new_n15636_1, new_n15635, new_n15632);
nand_4 g13288(new_n15637, new_n15636_1, new_n15631);
nand_4 g13289(new_n15638, new_n15637, new_n15629);
nor_4  g13290(new_n15639, new_n15638, new_n15627);
nor_4  g13291(new_n15640, new_n15639, new_n15626);
xor_3  g13292(n2238, new_n15640, new_n15624);
not_3  g13293(new_n15642, new_n13444);
xor_3  g13294(n2327, new_n15642, new_n13440);
not_3  g13295(new_n15644, new_n6663);
xor_3  g13296(n2343, new_n6707_1, new_n15644);
xnor_3 g13297(new_n15646, new_n12697, new_n9246_1);
nor_4  g13298(new_n15647, new_n7749, new_n7733);
not_3  g13299(new_n15648, new_n15647);
not_3  g13300(new_n15649, new_n7750);
not_3  g13301(new_n15650, new_n7775);
nand_4 g13302(new_n15651, new_n15650, new_n15649);
nand_4 g13303(new_n15652_1, new_n15651, new_n15648);
xnor_3 g13304(new_n15653, new_n15652_1, new_n15646);
not_3  g13305(new_n15654, new_n15653);
xor_3  g13306(new_n15655, n20923, n16524);
not_3  g13307(new_n15656, new_n15655);
nor_4  g13308(new_n15657, n18157, n11056);
nor_4  g13309(new_n15658, new_n7800, new_n15657);
xnor_3 g13310(new_n15659, new_n15658, new_n15656);
nor_4  g13311(new_n15660, new_n15659, n3785);
not_3  g13312(new_n15661, new_n15659);
nor_4  g13313(new_n15662_1, new_n15661, new_n4935);
nor_4  g13314(new_n15663, new_n15662_1, new_n15660);
nand_4 g13315(new_n15664, new_n7824, new_n7805);
nand_4 g13316(new_n15665, new_n15664, new_n7802);
xnor_3 g13317(new_n15666, new_n15665, new_n15663);
xnor_3 g13318(new_n15667, new_n15666, new_n15654);
xnor_3 g13319(new_n15668, new_n7801, new_n4943);
not_3  g13320(new_n15669, new_n7808);
nor_4  g13321(new_n15670, new_n7836, new_n7814);
nor_4  g13322(new_n15671, new_n15670, new_n7810);
xor_3  g13323(new_n15672, new_n7821, new_n4947_1);
nor_4  g13324(new_n15673, new_n15672, new_n15671);
nor_4  g13325(new_n15674, new_n15673, new_n15669);
nor_4  g13326(new_n15675, new_n15674, new_n15668);
nor_4  g13327(new_n15676, new_n7824, new_n7805);
nor_4  g13328(new_n15677, new_n15676, new_n15675);
nand_4 g13329(new_n15678, new_n15677, new_n7777);
nand_4 g13330(new_n15679, new_n7849, new_n7826);
nand_4 g13331(new_n15680, new_n15679, new_n15678);
not_3  g13332(new_n15681, new_n15680);
xor_3  g13333(n2361, new_n15681, new_n15667);
xor_3  g13334(n2363, new_n4051, new_n4047);
not_3  g13335(new_n15684, new_n5172);
xor_3  g13336(n2374, new_n5214, new_n15684);
not_3  g13337(new_n15686, new_n5547);
xor_3  g13338(new_n15687, n7305, n1204);
not_3  g13339(new_n15688, new_n6819);
nand_4 g13340(new_n15689, new_n6830, new_n6822);
nand_4 g13341(new_n15690, new_n15689, new_n15688);
nor_4  g13342(new_n15691, new_n15690, new_n15687);
nand_4 g13343(new_n15692, new_n15690, new_n15687);
not_3  g13344(new_n15693, new_n15692);
nor_4  g13345(new_n15694, new_n15693, new_n15691);
nand_4 g13346(new_n15695, new_n15694, new_n15686);
xnor_3 g13347(new_n15696, new_n15694, new_n5547);
nor_4  g13348(new_n15697, new_n6836, new_n6818);
nor_4  g13349(new_n15698, new_n6845, new_n6837);
nor_4  g13350(new_n15699, new_n15698, new_n15697);
nand_4 g13351(new_n15700, new_n15699, new_n15696);
nand_4 g13352(new_n15701, new_n15700, new_n15695);
xor_3  g13353(new_n15702, n20826, n626);
nor_4  g13354(new_n15703, n7305, n1204);
not_3  g13355(new_n15704, new_n15703);
nand_4 g13356(new_n15705, new_n15692, new_n15704);
xnor_3 g13357(new_n15706, new_n15705, new_n15702);
not_3  g13358(new_n15707, new_n15706);
xnor_3 g13359(new_n15708, new_n15707, new_n15701);
xnor_3 g13360(new_n15709, new_n15708, new_n5541);
xnor_3 g13361(new_n15710, new_n15709, new_n4143);
not_3  g13362(new_n15711, new_n15700);
nor_4  g13363(new_n15712, new_n15699, new_n15696);
nor_4  g13364(new_n15713, new_n15712, new_n15711);
nand_4 g13365(new_n15714, new_n15713, new_n4150_1);
nor_4  g13366(new_n15715, new_n6846, new_n4157);
nor_4  g13367(new_n15716_1, new_n6859, new_n6847);
nor_4  g13368(new_n15717, new_n15716_1, new_n15715);
not_3  g13369(new_n15718, new_n15714);
nor_4  g13370(new_n15719, new_n15713, new_n4150_1);
nor_4  g13371(new_n15720, new_n15719, new_n15718);
nand_4 g13372(new_n15721, new_n15720, new_n15717);
nand_4 g13373(new_n15722, new_n15721, new_n15714);
xor_3  g13374(n2388, new_n15722, new_n15710);
xor_3  g13375(new_n15724, n7335, n2160);
nor_4  g13376(new_n15725, n10763, n5696);
not_3  g13377(new_n15726, new_n6113);
nor_4  g13378(new_n15727, new_n6154, new_n15726);
nor_4  g13379(new_n15728, new_n15727, new_n15725);
xnor_3 g13380(new_n15729, new_n15728, new_n15724);
xor_3  g13381(new_n15730, n11220, n3425);
not_3  g13382(new_n15731, new_n15730);
nor_4  g13383(new_n15732, n22379, n9967);
nor_4  g13384(new_n15733, new_n6110, new_n15732);
xnor_3 g13385(new_n15734, new_n15733, new_n15731);
xnor_3 g13386(new_n15735, new_n15734, new_n15729);
nand_4 g13387(new_n15736, new_n6155, new_n6111);
nand_4 g13388(new_n15737, new_n6237, new_n6156);
nand_4 g13389(new_n15738, new_n15737, new_n15736);
xnor_3 g13390(new_n15739, new_n15738, new_n15735);
not_3  g13391(new_n15740, n5025);
not_3  g13392(new_n15741, n7593);
nor_4  g13393(new_n15742, new_n6015, n337);
xor_3  g13394(new_n15743_1, new_n15742, new_n15741);
not_3  g13395(new_n15744, new_n15743_1);
nor_4  g13396(new_n15745, new_n15744, new_n15740);
nor_4  g13397(new_n15746, new_n15743_1, n5025);
nor_4  g13398(new_n15747, new_n15746, new_n15745);
not_3  g13399(new_n15748, new_n15747);
nor_4  g13400(new_n15749_1, new_n6016, n6485);
not_3  g13401(new_n15750, new_n15749_1);
not_3  g13402(new_n15751, new_n6020);
not_3  g13403(new_n15752, new_n6061);
nand_4 g13404(new_n15753, new_n15752, new_n15751);
nand_4 g13405(new_n15754, new_n15753, new_n6017);
nand_4 g13406(new_n15755, new_n15754, new_n15750);
xnor_3 g13407(new_n15756, new_n15755, new_n15748);
xnor_3 g13408(new_n15757, new_n15756, new_n15739);
not_3  g13409(new_n15758, new_n6063);
nor_4  g13410(new_n15759, new_n6238, new_n15758);
not_3  g13411(new_n15760, new_n15759);
nand_4 g13412(new_n15761_1, new_n6315, new_n15760);
nand_4 g13413(new_n15762_1, new_n15761_1, new_n15757);
not_3  g13414(new_n15763, new_n15762_1);
nor_4  g13415(new_n15764, new_n15761_1, new_n15757);
nor_4  g13416(n2440, new_n15764, new_n15763);
not_3  g13417(new_n15766_1, new_n13889);
xor_3  g13418(n2444, new_n15766_1, new_n13872);
not_3  g13419(new_n15768, new_n5851);
xor_3  g13420(n2513, new_n15768, new_n3510);
not_3  g13421(new_n15770, n14323);
nor_4  g13422(new_n15771, new_n6970, new_n15770);
nor_4  g13423(new_n15772, new_n6969, n14323);
nor_4  g13424(new_n15773, new_n15772, new_n15771);
not_3  g13425(new_n15774, n2886);
nor_4  g13426(new_n15775, new_n6981, new_n15774);
xnor_3 g13427(new_n15776, new_n6980, n2886);
not_3  g13428(new_n15777, new_n15776);
not_3  g13429(new_n15778, n1040);
nor_4  g13430(new_n15779, new_n6996, new_n15778);
not_3  g13431(new_n15780_1, new_n15779);
nand_4 g13432(new_n15781, n20658, n9090);
not_3  g13433(new_n15782, new_n15781);
xnor_3 g13434(new_n15783, new_n6996, n1040);
nand_4 g13435(new_n15784, new_n15783, new_n15782);
nand_4 g13436(new_n15785, new_n15784, new_n15780_1);
nand_4 g13437(new_n15786, new_n15785, new_n15777);
not_3  g13438(new_n15787, new_n15786);
nor_4  g13439(new_n15788, new_n15787, new_n15775);
not_3  g13440(new_n15789, new_n15788);
xnor_3 g13441(new_n15790, new_n15789, new_n15773);
not_3  g13442(new_n15791, new_n15790);
nor_4  g13443(new_n15792, new_n15791, n12562);
not_3  g13444(new_n15793_1, n12562);
nor_4  g13445(new_n15794, new_n15790, new_n15793_1);
nor_4  g13446(new_n15795, new_n15794, new_n15792);
not_3  g13447(new_n15796, new_n15795);
nor_4  g13448(new_n15797, new_n15785, new_n15777);
nor_4  g13449(new_n15798, new_n15797, new_n15787);
nor_4  g13450(new_n15799, new_n15798, n7949);
not_3  g13451(new_n15800, new_n15799);
not_3  g13452(new_n15801, n7949);
not_3  g13453(new_n15802, new_n15798);
nor_4  g13454(new_n15803, new_n15802, new_n15801);
nor_4  g13455(new_n15804, new_n15803, new_n15799);
not_3  g13456(new_n15805, n14575);
nor_4  g13457(new_n15806, new_n13073, new_n15805);
nor_4  g13458(new_n15807, new_n15806, n24374);
not_3  g13459(new_n15808, new_n15807);
xnor_3 g13460(new_n15809, new_n6996, new_n15778);
xnor_3 g13461(new_n15810, new_n15809, new_n15781);
xor_3  g13462(new_n15811, new_n15806, n24374);
nand_4 g13463(new_n15812_1, new_n15811, new_n15810);
nand_4 g13464(new_n15813, new_n15812_1, new_n15808);
nand_4 g13465(new_n15814, new_n15813, new_n15804);
nand_4 g13466(new_n15815_1, new_n15814, new_n15800);
nor_4  g13467(new_n15816_1, new_n15815_1, new_n15796);
not_3  g13468(new_n15817, new_n15804);
not_3  g13469(new_n15818, new_n15810);
not_3  g13470(new_n15819, n24374);
xor_3  g13471(new_n15820, new_n15806, new_n15819);
nor_4  g13472(new_n15821, new_n15820, new_n15818);
nor_4  g13473(new_n15822, new_n15821, new_n15807);
nor_4  g13474(new_n15823, new_n15822, new_n15817);
nor_4  g13475(new_n15824, new_n15823, new_n15799);
nor_4  g13476(new_n15825, new_n15824, new_n15795);
nor_4  g13477(new_n15826, new_n15825, new_n15816_1);
xnor_3 g13478(new_n15827, new_n15826, new_n15480);
not_3  g13479(new_n15828, new_n15827);
nor_4  g13480(new_n15829, new_n15813, new_n15804);
nor_4  g13481(new_n15830, new_n15829, new_n15823);
nand_4 g13482(new_n15831_1, new_n15830, new_n15487);
xnor_3 g13483(new_n15832, new_n15830, new_n15486);
nor_4  g13484(new_n15833, new_n15811, new_n15810);
nor_4  g13485(new_n15834, new_n15833, new_n15821);
nand_4 g13486(new_n15835, new_n15834, new_n15490_1);
not_3  g13487(new_n15836, new_n15496_1);
xor_3  g13488(new_n15837, new_n13073, new_n15805);
not_3  g13489(new_n15838, new_n15837);
nor_4  g13490(new_n15839, new_n15838, new_n15836);
not_3  g13491(new_n15840, new_n15839);
not_3  g13492(new_n15841, new_n15835);
nor_4  g13493(new_n15842, new_n15834, new_n15490_1);
nor_4  g13494(new_n15843, new_n15842, new_n15841);
nand_4 g13495(new_n15844, new_n15843, new_n15840);
nand_4 g13496(new_n15845, new_n15844, new_n15835);
nand_4 g13497(new_n15846_1, new_n15845, new_n15832);
nand_4 g13498(new_n15847, new_n15846_1, new_n15831_1);
xor_3  g13499(n2515, new_n15847, new_n15828);
xnor_3 g13500(n2533, new_n13065, new_n13027);
nor_4  g13501(new_n15850, n26986, new_n3330);
xor_3  g13502(new_n15851, n26986, new_n3330);
not_3  g13503(new_n15852, new_n15851);
nor_4  g13504(new_n15853, n21287, new_n3464);
xor_3  g13505(new_n15854, n21287, new_n3464);
nor_4  g13506(new_n15855, new_n8884_1, n4256);
not_3  g13507(new_n15856, new_n15855);
xor_3  g13508(new_n15857, n20946, new_n8207);
nor_4  g13509(new_n15858, n22332, new_n3475);
not_3  g13510(new_n15859_1, new_n15858);
xor_3  g13511(new_n15860, n22332, new_n3475);
nor_4  g13512(new_n15861, new_n3482, n18907);
not_3  g13513(new_n15862, new_n15861);
xor_3  g13514(new_n15863, n26823, new_n2443);
not_3  g13515(new_n15864, n4812);
nor_4  g13516(new_n15865, new_n15864, n2731);
not_3  g13517(new_n15866, new_n15865);
not_3  g13518(new_n15867, new_n10001);
nor_4  g13519(new_n15868, new_n10017_1, new_n15867);
not_3  g13520(new_n15869_1, new_n15868);
nand_4 g13521(new_n15870, new_n15869_1, new_n15866);
nand_4 g13522(new_n15871, new_n15870, new_n15863);
nand_4 g13523(new_n15872, new_n15871, new_n15862);
nand_4 g13524(new_n15873, new_n15872, new_n15860);
nand_4 g13525(new_n15874, new_n15873, new_n15859_1);
nand_4 g13526(new_n15875, new_n15874, new_n15857);
nand_4 g13527(new_n15876, new_n15875, new_n15856);
nand_4 g13528(new_n15877, new_n15876, new_n15854);
not_3  g13529(new_n15878, new_n15877);
nor_4  g13530(new_n15879, new_n15878, new_n15853);
nor_4  g13531(new_n15880, new_n15879, new_n15852);
nor_4  g13532(new_n15881, new_n15880, new_n15850);
not_3  g13533(new_n15882, new_n15881);
not_3  g13534(new_n15883, new_n8472);
nand_4 g13535(new_n15884_1, new_n5905, new_n5896);
nor_4  g13536(new_n15885_1, new_n8324_1, new_n15884_1);
nand_4 g13537(new_n15886, new_n15885_1, new_n8319);
nor_4  g13538(new_n15887, new_n15886, new_n8309_1);
nand_4 g13539(new_n15888, new_n15887, new_n8385);
nor_4  g13540(new_n15889_1, new_n15888, new_n15883);
nand_4 g13541(new_n15890, new_n15888, new_n8475);
not_3  g13542(new_n15891, new_n15890);
nor_4  g13543(new_n15892, new_n15891, new_n15889_1);
not_3  g13544(new_n15893, new_n15892);
nor_4  g13545(new_n15894, new_n15893, new_n3547);
nor_4  g13546(new_n15895, new_n15892, new_n3546);
not_3  g13547(new_n15896, new_n3381);
xnor_3 g13548(new_n15897, new_n15887, new_n8385);
not_3  g13549(new_n15898, new_n15897);
nor_4  g13550(new_n15899, new_n15898, new_n15896);
not_3  g13551(new_n15900, new_n15899);
xnor_3 g13552(new_n15901, new_n15897, new_n3381);
not_3  g13553(new_n15902, new_n15901);
xnor_3 g13554(new_n15903, new_n15886, new_n8309_1);
not_3  g13555(new_n15904, new_n15903);
nor_4  g13556(new_n15905, new_n15904, new_n3383);
not_3  g13557(new_n15906, new_n15905);
nor_4  g13558(new_n15907, new_n15903, new_n3384);
nor_4  g13559(new_n15908, new_n15907, new_n15905);
xnor_3 g13560(new_n15909, new_n15885_1, new_n8319);
nand_4 g13561(new_n15910, new_n15909, new_n3391);
not_3  g13562(new_n15911, new_n15910);
nor_4  g13563(new_n15912, new_n15909, new_n3391);
nor_4  g13564(new_n15913, new_n15912, new_n15911);
xnor_3 g13565(new_n15914, new_n8324_1, new_n15884_1);
nand_4 g13566(new_n15915, new_n15914, new_n3398);
xnor_3 g13567(new_n15916, new_n15914, new_n3397);
nand_4 g13568(new_n15917_1, new_n5906, new_n3406);
nand_4 g13569(new_n15918_1, new_n5938, new_n5907);
nand_4 g13570(new_n15919, new_n15918_1, new_n15917_1);
nand_4 g13571(new_n15920, new_n15919, new_n15916);
nand_4 g13572(new_n15921, new_n15920, new_n15915);
nand_4 g13573(new_n15922_1, new_n15921, new_n15913);
nand_4 g13574(new_n15923, new_n15922_1, new_n15910);
nand_4 g13575(new_n15924, new_n15923, new_n15908);
nand_4 g13576(new_n15925, new_n15924, new_n15906);
nand_4 g13577(new_n15926, new_n15925, new_n15902);
nand_4 g13578(new_n15927, new_n15926, new_n15900);
nor_4  g13579(new_n15928, new_n15927, new_n15895);
nor_4  g13580(new_n15929, new_n15928, new_n15889_1);
not_3  g13581(new_n15930, new_n15929);
nor_4  g13582(new_n15931, new_n15930, new_n15894);
xnor_3 g13583(new_n15932, new_n15931, new_n15882);
nor_4  g13584(new_n15933, new_n15895, new_n15894);
xnor_3 g13585(new_n15934, new_n15933, new_n15927);
nor_4  g13586(new_n15935, new_n15934, new_n15881);
not_3  g13587(new_n15936_1, new_n15935);
not_3  g13588(new_n15937, new_n15934);
nor_4  g13589(new_n15938, new_n15937, new_n15882);
nor_4  g13590(new_n15939, new_n15938, new_n15935);
xor_3  g13591(new_n15940, new_n15879, new_n15852);
xnor_3 g13592(new_n15941, new_n15925, new_n15901);
not_3  g13593(new_n15942, new_n15941);
nor_4  g13594(new_n15943, new_n15942, new_n15940);
not_3  g13595(new_n15944, new_n15943);
not_3  g13596(new_n15945, new_n15940);
nor_4  g13597(new_n15946, new_n15941, new_n15945);
nor_4  g13598(new_n15947_1, new_n15946, new_n15943);
xnor_3 g13599(new_n15948, new_n15876, new_n15854);
xnor_3 g13600(new_n15949, new_n15923, new_n15908);
not_3  g13601(new_n15950, new_n15949);
nand_4 g13602(new_n15951, new_n15950, new_n15948);
xnor_3 g13603(new_n15952, new_n15949, new_n15948);
not_3  g13604(new_n15953, new_n15857);
xor_3  g13605(new_n15954, new_n15874, new_n15953);
xnor_3 g13606(new_n15955, new_n15921, new_n15913);
not_3  g13607(new_n15956_1, new_n15955);
nand_4 g13608(new_n15957, new_n15956_1, new_n15954);
xnor_3 g13609(new_n15958_1, new_n15955, new_n15954);
not_3  g13610(new_n15959, new_n15860);
xor_3  g13611(new_n15960, new_n15872, new_n15959);
xnor_3 g13612(new_n15961, new_n15919, new_n15916);
not_3  g13613(new_n15962, new_n15961);
nand_4 g13614(new_n15963, new_n15962, new_n15960);
not_3  g13615(new_n15964, new_n15963);
nor_4  g13616(new_n15965, new_n15962, new_n15960);
nor_4  g13617(new_n15966, new_n15965, new_n15964);
not_3  g13618(new_n15967_1, new_n5939);
not_3  g13619(new_n15968, new_n15863);
xor_3  g13620(new_n15969, new_n15870, new_n15968);
nor_4  g13621(new_n15970, new_n15969, new_n15967_1);
xnor_3 g13622(new_n15971, new_n15969, new_n15967_1);
nor_4  g13623(new_n15972, new_n10018_1, new_n10000);
nor_4  g13624(new_n15973, new_n10047, new_n10019_1);
nor_4  g13625(new_n15974, new_n15973, new_n15972);
nor_4  g13626(new_n15975, new_n15974, new_n15971);
nor_4  g13627(new_n15976, new_n15975, new_n15970);
nand_4 g13628(new_n15977, new_n15976, new_n15966);
nand_4 g13629(new_n15978, new_n15977, new_n15963);
nand_4 g13630(new_n15979_1, new_n15978, new_n15958_1);
nand_4 g13631(new_n15980, new_n15979_1, new_n15957);
nand_4 g13632(new_n15981, new_n15980, new_n15952);
nand_4 g13633(new_n15982, new_n15981, new_n15951);
nand_4 g13634(new_n15983, new_n15982, new_n15947_1);
nand_4 g13635(new_n15984, new_n15983, new_n15944);
nand_4 g13636(new_n15985, new_n15984, new_n15939);
nand_4 g13637(new_n15986_1, new_n15985, new_n15936_1);
xnor_3 g13638(n2535, new_n15986_1, new_n15932);
nor_4  g13639(new_n15988, n20259, n3925);
nand_4 g13640(new_n15989, new_n15988, new_n5625);
nor_4  g13641(new_n15990, new_n15989, n7305);
nand_4 g13642(new_n15991, new_n15990, new_n5641);
nor_4  g13643(new_n15992, new_n15991, n22198);
nand_4 g13644(new_n15993, new_n15991, n22198);
not_3  g13645(new_n15994, new_n15993);
nor_4  g13646(new_n15995, new_n15994, new_n15992);
not_3  g13647(new_n15996, new_n15995);
nor_4  g13648(new_n15997, new_n15996, new_n3838);
nor_4  g13649(new_n15998, new_n15995, n21674);
nor_4  g13650(new_n15999, new_n15998, new_n15997);
not_3  g13651(new_n16000, new_n15999);
not_3  g13652(new_n16001, new_n15991);
nor_4  g13653(new_n16002, new_n15990, new_n5641);
nor_4  g13654(new_n16003, new_n16002, new_n16001);
nor_4  g13655(new_n16004, new_n16003, n17251);
not_3  g13656(new_n16005, new_n16003);
nor_4  g13657(new_n16006, new_n16005, new_n9754);
nor_4  g13658(new_n16007, new_n16006, new_n16004);
nand_4 g13659(new_n16008, new_n15989, n7305);
not_3  g13660(new_n16009, new_n16008);
nor_4  g13661(new_n16010, new_n16009, new_n15990);
nor_4  g13662(new_n16011, new_n16010, n14790);
not_3  g13663(new_n16012, new_n16011);
xnor_3 g13664(new_n16013_1, new_n15988, new_n5625);
nand_4 g13665(new_n16014, new_n16013_1, new_n3850_1);
xnor_3 g13666(new_n16015, new_n16013_1, n10096);
xnor_3 g13667(new_n16016, n20259, n3925);
nand_4 g13668(new_n16017, new_n16016, new_n3854);
nand_4 g13669(new_n16018, n9246, n3925);
xnor_3 g13670(new_n16019, new_n16016, n16994);
nand_4 g13671(new_n16020, new_n16019, new_n16018);
nand_4 g13672(new_n16021, new_n16020, new_n16017);
nand_4 g13673(new_n16022, new_n16021, new_n16015);
nand_4 g13674(new_n16023, new_n16022, new_n16014);
not_3  g13675(new_n16024, n14790);
not_3  g13676(new_n16025, new_n16010);
nor_4  g13677(new_n16026, new_n16025, new_n16024);
nor_4  g13678(new_n16027, new_n16026, new_n16011);
nand_4 g13679(new_n16028, new_n16027, new_n16023);
nand_4 g13680(new_n16029_1, new_n16028, new_n16012);
nand_4 g13681(new_n16030, new_n16029_1, new_n16007);
not_3  g13682(new_n16031, new_n16030);
nor_4  g13683(new_n16032, new_n16031, new_n16004);
xnor_3 g13684(new_n16033, new_n16032, new_n16000);
xnor_3 g13685(new_n16034, new_n16033, new_n9182_1);
not_3  g13686(new_n16035, new_n16034);
xnor_3 g13687(new_n16036, new_n16029_1, new_n16007);
nor_4  g13688(new_n16037, new_n16036, new_n9188);
xnor_3 g13689(new_n16038, new_n16036, new_n9188);
xnor_3 g13690(new_n16039, new_n16027, new_n16023);
nor_4  g13691(new_n16040, new_n16039, new_n9197);
xnor_3 g13692(new_n16041, new_n16039, new_n9197);
not_3  g13693(new_n16042, new_n9206);
xnor_3 g13694(new_n16043, new_n16021, new_n16015);
nand_4 g13695(new_n16044, new_n16043, new_n16042);
not_3  g13696(new_n16045, new_n16044);
nor_4  g13697(new_n16046, new_n16043, new_n16042);
nor_4  g13698(new_n16047, new_n16046, new_n16045);
xnor_3 g13699(new_n16048, new_n16019, new_n16018);
nand_4 g13700(new_n16049, new_n16048, new_n9224);
nor_4  g13701(new_n16050, new_n11714, new_n9221);
not_3  g13702(new_n16051, new_n16049);
nor_4  g13703(new_n16052, new_n16048, new_n9224);
nor_4  g13704(new_n16053, new_n16052, new_n16051);
nand_4 g13705(new_n16054, new_n16053, new_n16050);
nand_4 g13706(new_n16055, new_n16054, new_n16049);
nand_4 g13707(new_n16056, new_n16055, new_n16047);
nand_4 g13708(new_n16057, new_n16056, new_n16044);
nor_4  g13709(new_n16058, new_n16057, new_n16041);
nor_4  g13710(new_n16059, new_n16058, new_n16040);
nor_4  g13711(new_n16060_1, new_n16059, new_n16038);
nor_4  g13712(new_n16061, new_n16060_1, new_n16037);
nor_4  g13713(new_n16062_1, new_n16061, new_n16035);
not_3  g13714(new_n16063, new_n16061);
nor_4  g13715(new_n16064, new_n16063, new_n16034);
nor_4  g13716(new_n16065, new_n16064, new_n16062_1);
not_3  g13717(new_n16066, new_n16065);
xor_3  g13718(new_n16067, n1163, new_n9849);
nor_4  g13719(new_n16068_1, new_n9857, n18537);
not_3  g13720(new_n16069, new_n16068_1);
xor_3  g13721(new_n16070, n24170, new_n10143);
nor_4  g13722(new_n16071, n7057, new_n9858);
not_3  g13723(new_n16072, new_n16071);
xor_3  g13724(new_n16073, n7057, new_n9858);
nor_4  g13725(new_n16074, n8869, new_n5757);
nor_4  g13726(new_n16075, new_n9864, n8381);
nor_4  g13727(new_n16076, new_n5778, n10372);
nand_4 g13728(new_n16077, n12495, new_n9869);
nor_4  g13729(new_n16078, n20235, new_n8273);
nor_4  g13730(new_n16079, new_n16078, new_n16077);
nor_4  g13731(new_n16080_1, new_n16079, new_n16076);
nor_4  g13732(new_n16081, new_n16080_1, new_n16075);
nor_4  g13733(new_n16082, new_n16081, new_n16074);
nand_4 g13734(new_n16083, new_n16082, new_n16073);
nand_4 g13735(new_n16084, new_n16083, new_n16072);
nand_4 g13736(new_n16085, new_n16084, new_n16070);
nand_4 g13737(new_n16086, new_n16085, new_n16069);
xor_3  g13738(new_n16087, new_n16086, new_n16067);
xnor_3 g13739(new_n16088, new_n16087, new_n16066);
xor_3  g13740(new_n16089, new_n16084, new_n16070);
not_3  g13741(new_n16090, new_n16038);
not_3  g13742(new_n16091, new_n16059);
nor_4  g13743(new_n16092, new_n16091, new_n16090);
nor_4  g13744(new_n16093, new_n16092, new_n16060_1);
not_3  g13745(new_n16094, new_n16093);
nor_4  g13746(new_n16095, new_n16094, new_n16089);
not_3  g13747(new_n16096, new_n16095);
not_3  g13748(new_n16097, new_n16089);
nor_4  g13749(new_n16098_1, new_n16093, new_n16097);
nor_4  g13750(new_n16099, new_n16098_1, new_n16095);
not_3  g13751(new_n16100, new_n16041);
not_3  g13752(new_n16101, new_n16057);
nor_4  g13753(new_n16102, new_n16101, new_n16100);
nor_4  g13754(new_n16103, new_n16102, new_n16058);
not_3  g13755(new_n16104, new_n16103);
xor_3  g13756(new_n16105, new_n16082, new_n16073);
nor_4  g13757(new_n16106, new_n16105, new_n16104);
not_3  g13758(new_n16107, new_n16106);
not_3  g13759(new_n16108, new_n16105);
nor_4  g13760(new_n16109, new_n16108, new_n16103);
nor_4  g13761(new_n16110_1, new_n16109, new_n16106);
not_3  g13762(new_n16111, new_n16056);
nor_4  g13763(new_n16112, new_n16055, new_n16047);
nor_4  g13764(new_n16113, new_n16112, new_n16111);
nor_4  g13765(new_n16114, new_n16075, new_n16074);
xor_3  g13766(new_n16115, new_n16114, new_n16080_1);
nor_4  g13767(new_n16116, new_n16115, new_n16113);
not_3  g13768(new_n16117, new_n16116);
xnor_3 g13769(new_n16118, new_n16115, new_n16113);
not_3  g13770(new_n16119, new_n16118);
nor_4  g13771(new_n16120, new_n11717, new_n11716);
nor_4  g13772(new_n16121, new_n16078, new_n16076);
xor_3  g13773(new_n16122, new_n16121, new_n16077);
nor_4  g13774(new_n16123, new_n16122, new_n16120);
not_3  g13775(new_n16124, new_n16123);
xnor_3 g13776(new_n16125, new_n16053, new_n16050);
not_3  g13777(new_n16126, new_n16125);
xnor_3 g13778(new_n16127, new_n16122, new_n16120);
nor_4  g13779(new_n16128, new_n16127, new_n16126);
not_3  g13780(new_n16129, new_n16128);
nand_4 g13781(new_n16130, new_n16129, new_n16124);
nand_4 g13782(new_n16131, new_n16130, new_n16119);
nand_4 g13783(new_n16132, new_n16131, new_n16117);
nand_4 g13784(new_n16133, new_n16132, new_n16110_1);
nand_4 g13785(new_n16134, new_n16133, new_n16107);
nand_4 g13786(new_n16135, new_n16134, new_n16099);
nand_4 g13787(new_n16136, new_n16135, new_n16096);
xor_3  g13788(n2537, new_n16136, new_n16088);
nor_4  g13789(new_n16138, new_n13269, new_n3134);
not_3  g13790(new_n16139, new_n3086);
xnor_3 g13791(new_n16140, new_n3111, new_n16139);
nor_4  g13792(new_n16141, new_n13268, new_n16140);
nor_4  g13793(new_n16142_1, new_n16141, new_n16138);
not_3  g13794(new_n16143, new_n16142_1);
nor_4  g13795(new_n16144, new_n4708, new_n3139);
not_3  g13796(new_n16145, new_n3089_1);
xnor_3 g13797(new_n16146, new_n3109, new_n16145);
nor_4  g13798(new_n16147, new_n4707, new_n16146);
nor_4  g13799(new_n16148, new_n16147, new_n16144);
not_3  g13800(new_n16149, new_n16148);
nor_4  g13801(new_n16150, new_n4714, new_n3145);
not_3  g13802(new_n16151, new_n16150);
nor_4  g13803(new_n16152, new_n4715, new_n3146);
nor_4  g13804(new_n16153, new_n16152, new_n16150);
nor_4  g13805(new_n16154, new_n4723, new_n3156);
nor_4  g13806(new_n16155, new_n4722_1, new_n3155);
nor_4  g13807(new_n16156, new_n16155, new_n16154);
not_3  g13808(new_n16157, new_n16156);
nor_4  g13809(new_n16158_1, new_n4730, new_n3162);
not_3  g13810(new_n16159, new_n16158_1);
nor_4  g13811(new_n16160, new_n3167, n1152);
xnor_3 g13812(new_n16161, new_n4730, new_n3162);
not_3  g13813(new_n16162, new_n16161);
nand_4 g13814(new_n16163, new_n16162, new_n16160);
nand_4 g13815(new_n16164, new_n16163, new_n16159);
nor_4  g13816(new_n16165, new_n16164, new_n16157);
nor_4  g13817(new_n16166, new_n16165, new_n16154);
nand_4 g13818(new_n16167_1, new_n16166, new_n16153);
nand_4 g13819(new_n16168, new_n16167_1, new_n16151);
nor_4  g13820(new_n16169, new_n16168, new_n16149);
nor_4  g13821(new_n16170, new_n16169, new_n16144);
xnor_3 g13822(new_n16171, new_n16170, new_n16143);
xnor_3 g13823(new_n16172, new_n16171, new_n14487);
not_3  g13824(new_n16173, new_n16172);
xnor_3 g13825(new_n16174, new_n16168, new_n16149);
nand_4 g13826(new_n16175, new_n16174, new_n14491);
xnor_3 g13827(new_n16176, new_n16174, new_n11471);
not_3  g13828(new_n16177, new_n16167_1);
nor_4  g13829(new_n16178, new_n16166, new_n16153);
nor_4  g13830(new_n16179, new_n16178, new_n16177);
nand_4 g13831(new_n16180, new_n16179, new_n14498);
not_3  g13832(new_n16181, new_n16180);
nor_4  g13833(new_n16182, new_n16179, new_n14498);
nor_4  g13834(new_n16183, new_n16182, new_n16181);
not_3  g13835(new_n16184, new_n16164);
nor_4  g13836(new_n16185_1, new_n16184, new_n16156);
nor_4  g13837(new_n16186, new_n16185_1, new_n16165);
not_3  g13838(new_n16187, new_n16186);
nor_4  g13839(new_n16188, new_n16187, new_n11490);
xnor_3 g13840(new_n16189, new_n16186, new_n11491);
not_3  g13841(new_n16190, new_n16163);
nor_4  g13842(new_n16191, new_n16162, new_n16160);
nor_4  g13843(new_n16192, new_n16191, new_n16190);
nand_4 g13844(new_n16193, new_n16192, new_n11496_1);
xor_3  g13845(new_n16194, new_n3167, new_n3013);
not_3  g13846(new_n16195, new_n16194);
nor_4  g13847(new_n16196_1, new_n16195, new_n8492);
not_3  g13848(new_n16197, new_n16196_1);
not_3  g13849(new_n16198, new_n16193);
nor_4  g13850(new_n16199, new_n16192, new_n11496_1);
nor_4  g13851(new_n16200, new_n16199, new_n16198);
nand_4 g13852(new_n16201, new_n16200, new_n16197);
nand_4 g13853(new_n16202, new_n16201, new_n16193);
nor_4  g13854(new_n16203, new_n16202, new_n16189);
nor_4  g13855(new_n16204, new_n16203, new_n16188);
nand_4 g13856(new_n16205, new_n16204, new_n16183);
nand_4 g13857(new_n16206_1, new_n16205, new_n16180);
nand_4 g13858(new_n16207, new_n16206_1, new_n16176);
nand_4 g13859(new_n16208, new_n16207, new_n16175);
xor_3  g13860(n2553, new_n16208, new_n16173);
not_3  g13861(new_n16210, new_n14369);
xor_3  g13862(n2555, new_n14388, new_n16210);
not_3  g13863(new_n16212, n12892);
xor_3  g13864(new_n16213, new_n12875_1, new_n16212);
not_3  g13865(new_n16214, new_n16213);
nand_4 g13866(new_n16215_1, new_n16214, new_n12071);
not_3  g13867(new_n16216, new_n12067);
nor_4  g13868(new_n16217_1, new_n12979, new_n16212);
not_3  g13869(new_n16218_1, new_n16217_1);
not_3  g13870(new_n16219_1, n12209);
xnor_3 g13871(new_n16220, new_n12877, new_n16219_1);
not_3  g13872(new_n16221, new_n16220);
nor_4  g13873(new_n16222, new_n16221, new_n16218_1);
nor_4  g13874(new_n16223_1, new_n16220, new_n16217_1);
nor_4  g13875(new_n16224, new_n16223_1, new_n16222);
not_3  g13876(new_n16225, new_n16224);
nor_4  g13877(new_n16226, new_n16225, new_n16216);
nor_4  g13878(new_n16227, new_n16224, new_n12067);
nor_4  g13879(new_n16228, new_n16227, new_n16226);
xor_3  g13880(n2560, new_n16228, new_n16215_1);
nor_4  g13881(new_n16230_1, n26180, n10650);
xor_3  g13882(new_n16231, n26180, n10650);
not_3  g13883(new_n16232, new_n16231);
nor_4  g13884(new_n16233, n24004, n12900);
xor_3  g13885(new_n16234, n24004, n12900);
not_3  g13886(new_n16235, new_n16234);
nor_4  g13887(new_n16236, n20411, n12871);
xor_3  g13888(new_n16237, n20411, n12871);
not_3  g13889(new_n16238, new_n16237);
nand_4 g13890(new_n16239, new_n3764, new_n15140);
xor_3  g13891(new_n16240, n23304, n17069);
nor_4  g13892(new_n16241, n19361, n15918);
not_3  g13893(new_n16242, new_n16241);
xor_3  g13894(new_n16243_1, n19361, n15918);
nor_4  g13895(new_n16244, n17784, n1437);
not_3  g13896(new_n16245, new_n16244);
xor_3  g13897(new_n16246, n17784, n1437);
nor_4  g13898(new_n16247_1, n14323, n4722);
not_3  g13899(new_n16248, new_n16247_1);
xor_3  g13900(new_n16249, n14323, n4722);
nor_4  g13901(new_n16250, n14633, n2886);
not_3  g13902(new_n16251, new_n16250);
xor_3  g13903(new_n16252, n14633, n2886);
nand_4 g13904(new_n16253, new_n3797, new_n15778);
nand_4 g13905(new_n16254, n18578, n9090);
xor_3  g13906(new_n16255, n8721, n1040);
nand_4 g13907(new_n16256, new_n16255, new_n16254);
nand_4 g13908(new_n16257, new_n16256, new_n16253);
nand_4 g13909(new_n16258, new_n16257, new_n16252);
nand_4 g13910(new_n16259, new_n16258, new_n16251);
nand_4 g13911(new_n16260, new_n16259, new_n16249);
nand_4 g13912(new_n16261, new_n16260, new_n16248);
nand_4 g13913(new_n16262, new_n16261, new_n16246);
nand_4 g13914(new_n16263, new_n16262, new_n16245);
nand_4 g13915(new_n16264, new_n16263, new_n16243_1);
nand_4 g13916(new_n16265, new_n16264, new_n16242);
nand_4 g13917(new_n16266, new_n16265, new_n16240);
nand_4 g13918(new_n16267, new_n16266, new_n16239);
not_3  g13919(new_n16268, new_n16267);
nor_4  g13920(new_n16269, new_n16268, new_n16238);
nor_4  g13921(new_n16270, new_n16269, new_n16236);
nor_4  g13922(new_n16271, new_n16270, new_n16235);
nor_4  g13923(new_n16272, new_n16271, new_n16233);
nor_4  g13924(new_n16273, new_n16272, new_n16232);
nor_4  g13925(new_n16274, new_n16273, new_n16230_1);
nor_4  g13926(new_n16275_1, n9259, n6456);
nor_4  g13927(new_n16276, new_n6924, new_n6878);
nor_4  g13928(new_n16277, new_n16276, new_n16275_1);
not_3  g13929(new_n16278, new_n16277);
nor_4  g13930(new_n16279_1, new_n16278, new_n16274);
xor_3  g13931(new_n16280, new_n16277, new_n16274);
not_3  g13932(new_n16281, new_n6925);
xor_3  g13933(new_n16282, new_n16272, new_n16232);
not_3  g13934(new_n16283, new_n16282);
nor_4  g13935(new_n16284, new_n16283, new_n16281);
xnor_3 g13936(new_n16285, new_n16282, new_n6925);
xor_3  g13937(new_n16286, new_n16270, new_n16234);
nor_4  g13938(new_n16287, new_n16286, new_n6933);
xor_3  g13939(new_n16288, new_n16270, new_n16235);
xnor_3 g13940(new_n16289, new_n16288, new_n6930);
xor_3  g13941(new_n16290, new_n16268, new_n16237);
nor_4  g13942(new_n16291, new_n16290, new_n6938);
not_3  g13943(new_n16292, new_n16291);
xnor_3 g13944(new_n16293, new_n16290, new_n6937);
xnor_3 g13945(new_n16294, new_n16265, new_n16240);
not_3  g13946(new_n16295, new_n16294);
nand_4 g13947(new_n16296, new_n16295, new_n6945);
xnor_3 g13948(new_n16297, new_n16294, new_n6945);
xnor_3 g13949(new_n16298, new_n16263, new_n16243_1);
nor_4  g13950(new_n16299, new_n16298, new_n6955);
not_3  g13951(new_n16300, new_n16299);
xnor_3 g13952(new_n16301, new_n16298, new_n6952);
not_3  g13953(new_n16302, new_n16246);
xnor_3 g13954(new_n16303, new_n16261, new_n16302);
nand_4 g13955(new_n16304, new_n16303, new_n6960);
xnor_3 g13956(new_n16305, new_n16303, new_n6963);
not_3  g13957(new_n16306, new_n16249);
xnor_3 g13958(new_n16307, new_n16259, new_n16306);
nor_4  g13959(new_n16308, new_n16307, new_n6971_1);
xnor_3 g13960(new_n16309, new_n16307, new_n6971_1);
xor_3  g13961(new_n16310, n14633, new_n15774);
xnor_3 g13962(new_n16311, new_n16257, new_n16310);
nor_4  g13963(new_n16312, new_n16311, new_n6982);
xnor_3 g13964(new_n16313, new_n16311, new_n6982);
not_3  g13965(new_n16314, new_n6993);
xor_3  g13966(new_n16315, n18578, n9090);
nor_4  g13967(new_n16316, new_n16315, new_n6985_1);
nor_4  g13968(new_n16317, new_n16316, new_n16314);
not_3  g13969(new_n16318, new_n16254);
xnor_3 g13970(new_n16319, n8721, n1040);
xor_3  g13971(new_n16320, new_n16319, new_n16318);
not_3  g13972(new_n16321, new_n16317);
nand_4 g13973(new_n16322_1, new_n16316, new_n6907);
nand_4 g13974(new_n16323, new_n16322_1, new_n16321);
nor_4  g13975(new_n16324, new_n16323, new_n16320);
nor_4  g13976(new_n16325, new_n16324, new_n16317);
nor_4  g13977(new_n16326, new_n16325, new_n16313);
nor_4  g13978(new_n16327_1, new_n16326, new_n16312);
nor_4  g13979(new_n16328, new_n16327_1, new_n16309);
nor_4  g13980(new_n16329, new_n16328, new_n16308);
nand_4 g13981(new_n16330, new_n16329, new_n16305);
nand_4 g13982(new_n16331, new_n16330, new_n16304);
nand_4 g13983(new_n16332, new_n16331, new_n16301);
nand_4 g13984(new_n16333, new_n16332, new_n16300);
nand_4 g13985(new_n16334, new_n16333, new_n16297);
nand_4 g13986(new_n16335, new_n16334, new_n16296);
nand_4 g13987(new_n16336, new_n16335, new_n16293);
nand_4 g13988(new_n16337, new_n16336, new_n16292);
not_3  g13989(new_n16338, new_n16337);
nor_4  g13990(new_n16339, new_n16338, new_n16289);
nor_4  g13991(new_n16340, new_n16339, new_n16287);
nor_4  g13992(new_n16341, new_n16340, new_n16285);
nor_4  g13993(new_n16342, new_n16341, new_n16284);
nor_4  g13994(new_n16343, new_n16342, new_n16280);
nor_4  g13995(new_n16344, new_n16343, new_n16279_1);
xnor_3 g13996(new_n16345, new_n16342, new_n16280);
nor_4  g13997(new_n16346, n3506, new_n3825);
nor_4  g13998(new_n16347, new_n3876, new_n3827);
nor_4  g13999(new_n16348, new_n16347, new_n16346);
not_3  g14000(new_n16349, new_n16348);
nor_4  g14001(new_n16350_1, new_n16349, new_n16345);
not_3  g14002(new_n16351, new_n16350_1);
xnor_3 g14003(new_n16352, new_n16348, new_n16345);
not_3  g14004(new_n16353, new_n3877);
xnor_3 g14005(new_n16354, new_n16340, new_n16285);
nor_4  g14006(new_n16355, new_n16354, new_n16353);
not_3  g14007(new_n16356, new_n16355);
not_3  g14008(new_n16357, new_n16285);
xnor_3 g14009(new_n16358, new_n16340, new_n16357);
nor_4  g14010(new_n16359, new_n16358, new_n3877);
nor_4  g14011(new_n16360, new_n16359, new_n16355);
not_3  g14012(new_n16361, new_n16289);
xnor_3 g14013(new_n16362, new_n16338, new_n16361);
not_3  g14014(new_n16363, new_n16362);
nor_4  g14015(new_n16364, new_n16363, new_n3896);
not_3  g14016(new_n16365, new_n16364);
xnor_3 g14017(new_n16366, new_n16362, new_n3896);
xnor_3 g14018(new_n16367_1, new_n16335, new_n16293);
not_3  g14019(new_n16368, new_n16367_1);
nand_4 g14020(new_n16369, new_n16368, new_n3904);
xnor_3 g14021(new_n16370, new_n16367_1, new_n3904);
xnor_3 g14022(new_n16371, new_n16333, new_n16297);
not_3  g14023(new_n16372, new_n16371);
nand_4 g14024(new_n16373, new_n16372, new_n3912);
xnor_3 g14025(new_n16374, new_n16371, new_n3912);
xnor_3 g14026(new_n16375, new_n16331, new_n16301);
not_3  g14027(new_n16376_1, new_n16375);
nand_4 g14028(new_n16377, new_n16376_1, new_n3924);
xnor_3 g14029(new_n16378, new_n16375, new_n3924);
not_3  g14030(new_n16379_1, new_n16308);
not_3  g14031(new_n16380, new_n16309);
not_3  g14032(new_n16381, new_n16312);
not_3  g14033(new_n16382, new_n16313);
not_3  g14034(new_n16383, new_n16325);
nand_4 g14035(new_n16384, new_n16383, new_n16382);
nand_4 g14036(new_n16385, new_n16384, new_n16381);
nand_4 g14037(new_n16386, new_n16385, new_n16380);
nand_4 g14038(new_n16387, new_n16386, new_n16379_1);
xnor_3 g14039(new_n16388, new_n16387, new_n16305);
nand_4 g14040(new_n16389, new_n16388, new_n3932_1);
xnor_3 g14041(new_n16390, new_n16388, new_n3935);
xnor_3 g14042(new_n16391, new_n16327_1, new_n16309);
nand_4 g14043(new_n16392, new_n16391, new_n3940);
xnor_3 g14044(new_n16393, new_n16391, new_n3939);
xnor_3 g14045(new_n16394, new_n16325, new_n16313);
nand_4 g14046(new_n16395, new_n16394, new_n3947);
not_3  g14047(new_n16396_1, new_n16395);
nor_4  g14048(new_n16397, new_n16394, new_n3947);
nor_4  g14049(new_n16398_1, new_n16397, new_n16396_1);
xnor_3 g14050(new_n16399, new_n16323, new_n16320);
nand_4 g14051(new_n16400, new_n16399, new_n3961);
not_3  g14052(new_n16401, new_n16315);
xor_3  g14053(new_n16402, new_n16401, new_n6985_1);
nor_4  g14054(new_n16403, new_n16402, new_n3958);
not_3  g14055(new_n16404, new_n16400);
nor_4  g14056(new_n16405, new_n16399, new_n3961);
nor_4  g14057(new_n16406_1, new_n16405, new_n16404);
nand_4 g14058(new_n16407_1, new_n16406_1, new_n16403);
nand_4 g14059(new_n16408, new_n16407_1, new_n16400);
nand_4 g14060(new_n16409, new_n16408, new_n16398_1);
nand_4 g14061(new_n16410, new_n16409, new_n16395);
nand_4 g14062(new_n16411, new_n16410, new_n16393);
nand_4 g14063(new_n16412, new_n16411, new_n16392);
nand_4 g14064(new_n16413, new_n16412, new_n16390);
nand_4 g14065(new_n16414, new_n16413, new_n16389);
nand_4 g14066(new_n16415, new_n16414, new_n16378);
nand_4 g14067(new_n16416, new_n16415, new_n16377);
nand_4 g14068(new_n16417, new_n16416, new_n16374);
nand_4 g14069(new_n16418, new_n16417, new_n16373);
nand_4 g14070(new_n16419_1, new_n16418, new_n16370);
nand_4 g14071(new_n16420, new_n16419_1, new_n16369);
nand_4 g14072(new_n16421, new_n16420, new_n16366);
nand_4 g14073(new_n16422, new_n16421, new_n16365);
nand_4 g14074(new_n16423, new_n16422, new_n16360);
nand_4 g14075(new_n16424_1, new_n16423, new_n16356);
nand_4 g14076(new_n16425, new_n16424_1, new_n16352);
nand_4 g14077(new_n16426, new_n16425, new_n16351);
xnor_3 g14078(n2561, new_n16426, new_n16344);
xor_3  g14079(n2573, new_n10038, new_n10035);
xor_3  g14080(new_n16429, n18558, n10411);
nor_4  g14081(new_n16430, new_n2760, n7149);
nor_4  g14082(new_n16431, n16971, new_n3005);
nor_4  g14083(new_n16432, n14148, new_n12117);
nor_4  g14084(new_n16433_1, new_n3009, n11503);
nand_4 g14085(new_n16434, n18151, new_n3013);
nor_4  g14086(new_n16435, new_n16434, new_n16433_1);
nor_4  g14087(new_n16436, new_n16435, new_n16432);
nor_4  g14088(new_n16437, new_n16436, new_n16431);
nor_4  g14089(new_n16438, new_n16437, new_n16430);
xnor_3 g14090(new_n16439_1, new_n16438, new_n16429);
not_3  g14091(new_n16440_1, new_n16439_1);
not_3  g14092(new_n16441, new_n11961);
not_3  g14093(new_n16442, new_n11967);
not_3  g14094(new_n16443, new_n11966);
not_3  g14095(new_n16444, new_n11974);
nand_4 g14096(new_n16445_1, new_n11899, n10017);
nand_4 g14097(new_n16446, new_n11980_1, new_n16445_1);
nand_4 g14098(new_n16447, new_n16446, new_n16444);
nand_4 g14099(new_n16448, new_n16447, new_n16443);
nand_4 g14100(new_n16449, new_n16448, new_n16442);
xnor_3 g14101(new_n16450, new_n16449, new_n16441);
nor_4  g14102(new_n16451, new_n16450, new_n16440_1);
not_3  g14103(new_n16452, new_n16450);
nor_4  g14104(new_n16453, new_n16452, new_n16439_1);
nor_4  g14105(new_n16454, new_n16453, new_n16451);
nor_4  g14106(new_n16455, new_n16431, new_n16430);
xnor_3 g14107(new_n16456, new_n16455, new_n16436);
nor_4  g14108(new_n16457, new_n16447, new_n11969);
not_3  g14109(new_n16458, new_n16446);
nor_4  g14110(new_n16459, new_n16458, new_n11974);
nor_4  g14111(new_n16460_1, new_n16459, new_n11968);
nor_4  g14112(new_n16461, new_n16460_1, new_n16457);
not_3  g14113(new_n16462, new_n16461);
nor_4  g14114(new_n16463, new_n16462, new_n16456);
not_3  g14115(new_n16464, new_n16463);
not_3  g14116(new_n16465, new_n16456);
nor_4  g14117(new_n16466, new_n16461, new_n16465);
nor_4  g14118(new_n16467, new_n16466, new_n16463);
not_3  g14119(new_n16468, new_n16434);
nor_4  g14120(new_n16469, n18151, new_n3013);
nor_4  g14121(new_n16470, new_n16469, new_n16468);
nor_4  g14122(new_n16471, new_n16470, new_n11983);
nor_4  g14123(new_n16472, new_n16433_1, new_n16432);
xnor_3 g14124(new_n16473, new_n16472, new_n16434);
not_3  g14125(new_n16474, new_n16473);
nor_4  g14126(new_n16475, new_n16474, new_n16471);
not_3  g14127(new_n16476_1, new_n16471);
nor_4  g14128(new_n16477, new_n16473, new_n16476_1);
nor_4  g14129(new_n16478, new_n16477, new_n16475);
not_3  g14130(new_n16479, new_n16478);
not_3  g14131(new_n16480, new_n11980_1);
xor_3  g14132(new_n16481_1, new_n16480, new_n11975);
nor_4  g14133(new_n16482_1, new_n16481_1, new_n16479);
nor_4  g14134(new_n16483, new_n16482_1, new_n16475);
nand_4 g14135(new_n16484, new_n16483, new_n16467);
nand_4 g14136(new_n16485, new_n16484, new_n16464);
xnor_3 g14137(new_n16486, new_n16485, new_n16454);
xor_3  g14138(new_n16487, n19515, n17035);
not_3  g14139(new_n16488, n22588);
nor_4  g14140(new_n16489, new_n16488, n14684);
nor_4  g14141(new_n16490, n22588, new_n4669);
nor_4  g14142(new_n16491, new_n16219_1, n6631);
nor_4  g14143(new_n16492, n12209, new_n4688);
not_3  g14144(new_n16493_1, n24732);
nand_4 g14145(new_n16494, new_n16493_1, n12892);
nor_4  g14146(new_n16495, new_n16494, new_n16492);
nor_4  g14147(new_n16496, new_n16495, new_n16491);
nor_4  g14148(new_n16497, new_n16496, new_n16490);
nor_4  g14149(new_n16498, new_n16497, new_n16489);
xor_3  g14150(new_n16499, new_n16498, new_n16487);
not_3  g14151(new_n16500, new_n16499);
xnor_3 g14152(new_n16501, new_n16500, new_n16486);
not_3  g14153(new_n16502_1, new_n16501);
not_3  g14154(new_n16503, new_n16467);
not_3  g14155(new_n16504, new_n16475);
xor_3  g14156(new_n16505, new_n11980_1, new_n11975);
nand_4 g14157(new_n16506_1, new_n16505, new_n16478);
nand_4 g14158(new_n16507_1, new_n16506_1, new_n16504);
xnor_3 g14159(new_n16508, new_n16507_1, new_n16503);
not_3  g14160(new_n16509, new_n16496);
nor_4  g14161(new_n16510, new_n16490, new_n16489);
xor_3  g14162(new_n16511, new_n16510, new_n16509);
nand_4 g14163(new_n16512, new_n16511, new_n16508);
xor_3  g14164(new_n16513, n24732, new_n16212);
not_3  g14165(new_n16514, new_n11983);
xor_3  g14166(new_n16515, new_n16470, new_n16514);
nor_4  g14167(new_n16516_1, new_n16515, new_n16513);
not_3  g14168(new_n16517_1, new_n16516_1);
not_3  g14169(new_n16518, new_n16494);
nor_4  g14170(new_n16519, new_n16492, new_n16491);
xor_3  g14171(new_n16520, new_n16519, new_n16518);
nand_4 g14172(new_n16521_1, new_n16520, new_n16517_1);
xnor_3 g14173(new_n16522, new_n16520, new_n16516_1);
nor_4  g14174(new_n16523, new_n16505, new_n16478);
nor_4  g14175(new_n16524_1, new_n16523, new_n16482_1);
nand_4 g14176(new_n16525, new_n16524_1, new_n16522);
nand_4 g14177(new_n16526, new_n16525, new_n16521_1);
not_3  g14178(new_n16527_1, new_n16512);
nor_4  g14179(new_n16528, new_n16511, new_n16508);
nor_4  g14180(new_n16529, new_n16528, new_n16527_1);
nand_4 g14181(new_n16530, new_n16529, new_n16526);
nand_4 g14182(new_n16531, new_n16530, new_n16512);
xor_3  g14183(n2578, new_n16531, new_n16502_1);
nor_4  g14184(new_n16533, new_n14180, new_n9313);
xnor_3 g14185(new_n16534, new_n14180, new_n9313);
not_3  g14186(new_n16535, new_n9245);
not_3  g14187(new_n16536, new_n9313);
nor_4  g14188(new_n16537, new_n16536, new_n16535);
nor_4  g14189(new_n16538, new_n9394, new_n9314);
nor_4  g14190(new_n16539, new_n16538, new_n16537);
nor_4  g14191(new_n16540, new_n16539, new_n16534);
nor_4  g14192(n2582, new_n16540, new_n16533);
xor_3  g14193(n2602, new_n4846, new_n4831);
nor_4  g14194(new_n16543, n22201, n2420);
nand_4 g14195(new_n16544_1, new_n16543, new_n9612);
nor_4  g14196(new_n16545, new_n16544_1, n21078);
not_3  g14197(new_n16546, new_n16545);
nor_4  g14198(new_n16547, new_n16546, n12546);
xor_3  g14199(new_n16548, new_n16547, new_n9592);
not_3  g14200(new_n16549, new_n16548);
nor_4  g14201(new_n16550, new_n16549, new_n4389);
nor_4  g14202(new_n16551, new_n16548, new_n4388);
nor_4  g14203(new_n16552, new_n16551, new_n16550);
xor_3  g14204(new_n16553, new_n16545, new_n9600);
nor_4  g14205(new_n16554_1, new_n16553, new_n4393);
not_3  g14206(new_n16555, new_n16554_1);
xor_3  g14207(new_n16556, new_n16544_1, new_n9608);
nand_4 g14208(new_n16557, new_n16556, new_n5081);
xnor_3 g14209(new_n16558, new_n16556, new_n4396);
xor_3  g14210(new_n16559, new_n16543, n24485);
nor_4  g14211(new_n16560, new_n16559, new_n4403);
not_3  g14212(new_n16561, new_n16559);
nor_4  g14213(new_n16562, new_n16561, new_n4402);
nor_4  g14214(new_n16563, new_n16562, new_n16560);
not_3  g14215(new_n16564, new_n16563);
xor_3  g14216(new_n16565, n22201, n2420);
nor_4  g14217(new_n16566, new_n16565, new_n4409_1);
not_3  g14218(new_n16567, new_n16566);
not_3  g14219(new_n16568, new_n2605);
nor_4  g14220(new_n16569, new_n16568, new_n2596);
not_3  g14221(new_n16570, new_n16569);
not_3  g14222(new_n16571, new_n16565);
nor_4  g14223(new_n16572, new_n16571, new_n4410);
nor_4  g14224(new_n16573, new_n16572, new_n16566);
nand_4 g14225(new_n16574, new_n16573, new_n16570);
nand_4 g14226(new_n16575, new_n16574, new_n16567);
nor_4  g14227(new_n16576, new_n16575, new_n16564);
nor_4  g14228(new_n16577, new_n16576, new_n16560);
nand_4 g14229(new_n16578, new_n16577, new_n16558);
nand_4 g14230(new_n16579, new_n16578, new_n16557);
not_3  g14231(new_n16580, new_n16553);
nor_4  g14232(new_n16581, new_n16580, new_n5102);
nor_4  g14233(new_n16582, new_n16581, new_n16554_1);
nand_4 g14234(new_n16583_1, new_n16582, new_n16579);
nand_4 g14235(new_n16584_1, new_n16583_1, new_n16555);
xnor_3 g14236(new_n16585, new_n16584_1, new_n16552);
xnor_3 g14237(new_n16586, new_n9593, new_n12765);
nor_4  g14238(new_n16587, new_n9597, n3785);
not_3  g14239(new_n16588, new_n16587);
nor_4  g14240(new_n16589_1, new_n9601, new_n4935);
nor_4  g14241(new_n16590, new_n16589_1, new_n16587);
nand_4 g14242(new_n16591, new_n9609, new_n4943);
xor_3  g14243(new_n16592, new_n9609, new_n4943);
nor_4  g14244(new_n16593, new_n9616_1, new_n4947_1);
nor_4  g14245(new_n16594, new_n9615, n5822);
nor_4  g14246(new_n16595, new_n9623, n26443);
not_3  g14247(new_n16596_1, new_n16595);
nand_4 g14248(new_n16597, new_n2597, n1681);
nor_4  g14249(new_n16598, new_n9622_1, new_n4961);
nor_4  g14250(new_n16599, new_n16598, new_n16595);
nand_4 g14251(new_n16600, new_n16599, new_n16597);
nand_4 g14252(new_n16601, new_n16600, new_n16596_1);
nor_4  g14253(new_n16602, new_n16601, new_n16594);
nor_4  g14254(new_n16603, new_n16602, new_n16593);
nand_4 g14255(new_n16604, new_n16603, new_n16592);
nand_4 g14256(new_n16605, new_n16604, new_n16591);
nand_4 g14257(new_n16606, new_n16605, new_n16590);
nand_4 g14258(new_n16607, new_n16606, new_n16588);
xnor_3 g14259(new_n16608_1, new_n16607, new_n16586);
xnor_3 g14260(new_n16609, new_n16608_1, new_n16585);
not_3  g14261(new_n16610, new_n16609);
xnor_3 g14262(new_n16611, new_n16605, new_n16590);
not_3  g14263(new_n16612, new_n16611);
not_3  g14264(new_n16613, new_n16582);
xnor_3 g14265(new_n16614, new_n16613, new_n16579);
nand_4 g14266(new_n16615, new_n16614, new_n16612);
xnor_3 g14267(new_n16616, new_n16614, new_n16611);
xnor_3 g14268(new_n16617_1, new_n16577, new_n16558);
not_3  g14269(new_n16618, new_n16617_1);
not_3  g14270(new_n16619, new_n16603);
xnor_3 g14271(new_n16620, new_n16619, new_n16592);
nand_4 g14272(new_n16621, new_n16620, new_n16618);
xnor_3 g14273(new_n16622, new_n16620, new_n16617_1);
xnor_3 g14274(new_n16623, new_n16575, new_n16564);
nor_4  g14275(new_n16624, new_n16594, new_n16593);
not_3  g14276(new_n16625, new_n16624);
xnor_3 g14277(new_n16626, new_n16625, new_n16601);
nor_4  g14278(new_n16627, new_n16626, new_n16623);
xnor_3 g14279(new_n16628, new_n16573, new_n16570);
not_3  g14280(new_n16629, new_n16600);
nor_4  g14281(new_n16630_1, new_n16599, new_n16597);
nor_4  g14282(new_n16631, new_n16630_1, new_n16629);
not_3  g14283(new_n16632, new_n16631);
nor_4  g14284(new_n16633, new_n16632, new_n16628);
not_3  g14285(new_n16634, new_n16633);
not_3  g14286(new_n16635, new_n16597);
nor_4  g14287(new_n16636, new_n2597, n1681);
nor_4  g14288(new_n16637, new_n16636, new_n16635);
not_3  g14289(new_n16638, new_n16637);
nor_4  g14290(new_n16639, new_n2605, n22201);
nor_4  g14291(new_n16640_1, new_n16639, new_n16569);
not_3  g14292(new_n16641, new_n16640_1);
nor_4  g14293(new_n16642, new_n16641, new_n16638);
not_3  g14294(new_n16643, new_n16642);
not_3  g14295(new_n16644, new_n16628);
nor_4  g14296(new_n16645, new_n16631, new_n16644);
nor_4  g14297(new_n16646, new_n16645, new_n16633);
nand_4 g14298(new_n16647, new_n16646, new_n16643);
nand_4 g14299(new_n16648, new_n16647, new_n16634);
xnor_3 g14300(new_n16649, new_n16626, new_n16623);
nor_4  g14301(new_n16650, new_n16649, new_n16648);
nor_4  g14302(new_n16651, new_n16650, new_n16627);
nand_4 g14303(new_n16652, new_n16651, new_n16622);
nand_4 g14304(new_n16653, new_n16652, new_n16621);
nand_4 g14305(new_n16654, new_n16653, new_n16616);
nand_4 g14306(new_n16655, new_n16654, new_n16615);
xor_3  g14307(n2619, new_n16655, new_n16610);
nor_4  g14308(new_n16657, new_n6928, n12900);
not_3  g14309(new_n16658, new_n16657);
not_3  g14310(new_n16659, n12900);
xor_3  g14311(new_n16660, new_n6929, new_n16659);
nor_4  g14312(new_n16661, new_n6936, n20411);
not_3  g14313(new_n16662, new_n16661);
not_3  g14314(new_n16663, n20411);
xor_3  g14315(new_n16664, new_n6940, new_n16663);
nor_4  g14316(new_n16665, new_n6943, n17069);
not_3  g14317(new_n16666, new_n16665);
xor_3  g14318(new_n16667, new_n6944, new_n15140);
not_3  g14319(new_n16668, n15918);
nand_4 g14320(new_n16669, new_n6951, new_n16668);
nor_4  g14321(new_n16670, new_n6962, n17784);
not_3  g14322(new_n16671, new_n16670);
xor_3  g14323(new_n16672, new_n6962, n17784);
nor_4  g14324(new_n16673, new_n15788, new_n15772);
nor_4  g14325(new_n16674_1, new_n16673, new_n15771);
nand_4 g14326(new_n16675, new_n16674_1, new_n16672);
nand_4 g14327(new_n16676, new_n16675, new_n16671);
not_3  g14328(new_n16677, new_n16669);
nor_4  g14329(new_n16678, new_n6951, new_n16668);
nor_4  g14330(new_n16679, new_n16678, new_n16677);
nand_4 g14331(new_n16680, new_n16679, new_n16676);
nand_4 g14332(new_n16681, new_n16680, new_n16669);
nand_4 g14333(new_n16682_1, new_n16681, new_n16667);
nand_4 g14334(new_n16683, new_n16682_1, new_n16666);
nand_4 g14335(new_n16684_1, new_n16683, new_n16664);
nand_4 g14336(new_n16685, new_n16684_1, new_n16662);
nand_4 g14337(new_n16686, new_n16685, new_n16660);
nand_4 g14338(new_n16687, new_n16686, new_n16658);
nor_4  g14339(new_n16688_1, new_n6875, n10650);
not_3  g14340(new_n16689, n10650);
nor_4  g14341(new_n16690, new_n6876, new_n16689);
nor_4  g14342(new_n16691, new_n16690, new_n16688_1);
xnor_3 g14343(new_n16692, new_n16691, new_n16687);
nor_4  g14344(new_n16693, new_n16692, n6456);
not_3  g14345(new_n16694, new_n16693);
not_3  g14346(new_n16695, n6456);
not_3  g14347(new_n16696, new_n16692);
nor_4  g14348(new_n16697, new_n16696, new_n16695);
nor_4  g14349(new_n16698, new_n16697, new_n16693);
xnor_3 g14350(new_n16699, new_n16685, new_n16660);
nor_4  g14351(new_n16700, new_n16699, n4085);
not_3  g14352(new_n16701, new_n16700);
not_3  g14353(new_n16702, n4085);
not_3  g14354(new_n16703, new_n16699);
nor_4  g14355(new_n16704, new_n16703, new_n16702);
nor_4  g14356(new_n16705, new_n16704, new_n16700);
xnor_3 g14357(new_n16706, new_n16683, new_n16664);
nor_4  g14358(new_n16707, new_n16706, n26725);
not_3  g14359(new_n16708, new_n16707);
not_3  g14360(new_n16709, n26725);
not_3  g14361(new_n16710, new_n16706);
nor_4  g14362(new_n16711, new_n16710, new_n16709);
nor_4  g14363(new_n16712, new_n16711, new_n16707);
xnor_3 g14364(new_n16713, new_n16681, new_n16667);
nor_4  g14365(new_n16714, new_n16713, n11980);
not_3  g14366(new_n16715, new_n16714);
xnor_3 g14367(new_n16716, new_n16713, n11980);
not_3  g14368(new_n16717, new_n16716);
xnor_3 g14369(new_n16718, new_n16679, new_n16676);
nor_4  g14370(new_n16719, new_n16718, n3253);
not_3  g14371(new_n16720, new_n16719);
xnor_3 g14372(new_n16721, new_n16718, n3253);
not_3  g14373(new_n16722_1, new_n16721);
not_3  g14374(new_n16723, n7759);
not_3  g14375(new_n16724, n17784);
xor_3  g14376(new_n16725, new_n6962, new_n16724);
not_3  g14377(new_n16726, new_n16674_1);
nor_4  g14378(new_n16727, new_n16726, new_n16725);
nand_4 g14379(new_n16728, new_n16726, new_n16725);
not_3  g14380(new_n16729, new_n16728);
nor_4  g14381(new_n16730, new_n16729, new_n16727);
nor_4  g14382(new_n16731, new_n16730, new_n16723);
nand_4 g14383(new_n16732, new_n16728, new_n16675);
xnor_3 g14384(new_n16733_1, new_n16732, n7759);
nor_4  g14385(new_n16734, new_n15816_1, new_n15794);
nor_4  g14386(new_n16735, new_n16734, new_n16733_1);
nor_4  g14387(new_n16736, new_n16735, new_n16731);
nand_4 g14388(new_n16737, new_n16736, new_n16722_1);
nand_4 g14389(new_n16738, new_n16737, new_n16720);
nand_4 g14390(new_n16739, new_n16738, new_n16717);
nand_4 g14391(new_n16740, new_n16739, new_n16715);
nand_4 g14392(new_n16741, new_n16740, new_n16712);
nand_4 g14393(new_n16742, new_n16741, new_n16708);
nand_4 g14394(new_n16743_1, new_n16742, new_n16705);
nand_4 g14395(new_n16744, new_n16743_1, new_n16701);
nand_4 g14396(new_n16745, new_n16744, new_n16698);
nand_4 g14397(new_n16746, new_n16745, new_n16694);
nor_4  g14398(new_n16747, new_n16688_1, new_n16687);
not_3  g14399(new_n16748, new_n16747);
not_3  g14400(new_n16749, new_n6874);
nor_4  g14401(new_n16750, new_n16749, n2979);
nor_4  g14402(new_n16751, new_n16690, new_n16750);
nand_4 g14403(new_n16752, new_n16751, new_n16748);
nor_4  g14404(new_n16753, new_n16752, new_n16746);
nor_4  g14405(new_n16754, new_n16753, new_n15428_1);
xnor_3 g14406(new_n16755, new_n16753, new_n15429);
not_3  g14407(new_n16756, new_n16755);
xnor_3 g14408(new_n16757, new_n16752, new_n16746);
nand_4 g14409(new_n16758, new_n16757, new_n15439);
xnor_3 g14410(new_n16759, new_n16757, new_n15435_1);
not_3  g14411(new_n16760, new_n15443);
not_3  g14412(new_n16761, new_n16698);
xnor_3 g14413(new_n16762, new_n16744, new_n16761);
nand_4 g14414(new_n16763, new_n16762, new_n16760);
xnor_3 g14415(new_n16764, new_n16762, new_n15443);
not_3  g14416(new_n16765, new_n16705);
xnor_3 g14417(new_n16766, new_n16742, new_n16765);
nand_4 g14418(new_n16767, new_n16766, new_n15455);
xnor_3 g14419(new_n16768, new_n16766, new_n15452);
xnor_3 g14420(new_n16769, new_n16740, new_n16712);
nor_4  g14421(new_n16770, new_n16769, new_n15459);
not_3  g14422(new_n16771, new_n16770);
not_3  g14423(new_n16772, new_n16731);
nor_4  g14424(new_n16773, new_n16732, n7759);
nor_4  g14425(new_n16774, new_n16773, new_n16731);
not_3  g14426(new_n16775, new_n15794);
nand_4 g14427(new_n16776, new_n15824, new_n15795);
nand_4 g14428(new_n16777, new_n16776, new_n16775);
nand_4 g14429(new_n16778, new_n16777, new_n16774);
nand_4 g14430(new_n16779, new_n16778, new_n16772);
nor_4  g14431(new_n16780, new_n16779, new_n16721);
nor_4  g14432(new_n16781, new_n16780, new_n16719);
nor_4  g14433(new_n16782, new_n16781, new_n16716);
nor_4  g14434(new_n16783, new_n16782, new_n16714);
xnor_3 g14435(new_n16784, new_n16783, new_n16712);
nor_4  g14436(new_n16785, new_n16784, new_n15458);
nor_4  g14437(new_n16786, new_n16785, new_n16770);
not_3  g14438(new_n16787, new_n15464);
xnor_3 g14439(new_n16788, new_n16738, new_n16717);
not_3  g14440(new_n16789, new_n16788);
nand_4 g14441(new_n16790, new_n16789, new_n16787);
xnor_3 g14442(new_n16791, new_n16788, new_n16787);
xnor_3 g14443(new_n16792, new_n16779, new_n16721);
not_3  g14444(new_n16793, new_n16792);
nand_4 g14445(new_n16794, new_n16793, new_n15469);
xnor_3 g14446(new_n16795, new_n16792, new_n15469);
xnor_3 g14447(new_n16796, new_n16734, new_n16733_1);
nand_4 g14448(new_n16797, new_n16796, new_n15474);
xnor_3 g14449(new_n16798_1, new_n16796, new_n15476);
not_3  g14450(new_n16799, new_n15826);
nand_4 g14451(new_n16800, new_n16799, new_n15480);
nand_4 g14452(new_n16801, new_n15847, new_n15827);
nand_4 g14453(new_n16802, new_n16801, new_n16800);
nand_4 g14454(new_n16803, new_n16802, new_n16798_1);
nand_4 g14455(new_n16804, new_n16803, new_n16797);
nand_4 g14456(new_n16805, new_n16804, new_n16795);
nand_4 g14457(new_n16806, new_n16805, new_n16794);
nand_4 g14458(new_n16807, new_n16806, new_n16791);
nand_4 g14459(new_n16808, new_n16807, new_n16790);
nand_4 g14460(new_n16809, new_n16808, new_n16786);
nand_4 g14461(new_n16810, new_n16809, new_n16771);
nand_4 g14462(new_n16811, new_n16810, new_n16768);
nand_4 g14463(new_n16812_1, new_n16811, new_n16767);
nand_4 g14464(new_n16813, new_n16812_1, new_n16764);
nand_4 g14465(new_n16814, new_n16813, new_n16763);
nand_4 g14466(new_n16815, new_n16814, new_n16759);
nand_4 g14467(new_n16816, new_n16815, new_n16758);
not_3  g14468(new_n16817, new_n16816);
nor_4  g14469(new_n16818_1, new_n16817, new_n16756);
nor_4  g14470(n2661, new_n16818_1, new_n16754);
not_3  g14471(new_n16820, new_n13436);
xor_3  g14472(n2693, new_n16820, new_n13434);
nor_4  g14473(new_n16822, new_n16440_1, new_n8610);
nor_4  g14474(new_n16823, new_n16439_1, new_n8611);
nor_4  g14475(new_n16824_1, new_n16823, new_n16822);
nor_4  g14476(new_n16825, new_n16456, new_n8617);
not_3  g14477(new_n16826, new_n16825);
nor_4  g14478(new_n16827, new_n16465, new_n8618);
nor_4  g14479(new_n16828, new_n16827, new_n16825);
nor_4  g14480(new_n16829, new_n16473, new_n8624);
not_3  g14481(new_n16830, new_n16829);
nor_4  g14482(new_n16831, new_n16470, new_n14608);
xnor_3 g14483(new_n16832, new_n16473, new_n8624);
not_3  g14484(new_n16833, new_n16832);
nand_4 g14485(new_n16834_1, new_n16833, new_n16831);
nand_4 g14486(new_n16835, new_n16834_1, new_n16830);
nand_4 g14487(new_n16836, new_n16835, new_n16828);
nand_4 g14488(new_n16837_1, new_n16836, new_n16826);
xnor_3 g14489(new_n16838, new_n16837_1, new_n16824_1);
xor_3  g14490(new_n16839, n8309, n4665);
nor_4  g14491(new_n16840, new_n10474, n19005);
not_3  g14492(new_n16841_1, new_n16840);
nor_4  g14493(new_n16842, n19144, new_n3007);
not_3  g14494(new_n16843, new_n16842);
nor_4  g14495(new_n16844, new_n10483, n4326);
not_3  g14496(new_n16845, new_n16844);
nor_4  g14497(new_n16846, n12593, new_n3011);
not_3  g14498(new_n16847, new_n16846);
nor_4  g14499(new_n16848, new_n12281, n5438);
nand_4 g14500(new_n16849, new_n16848, new_n16847);
nand_4 g14501(new_n16850, new_n16849, new_n16845);
nand_4 g14502(new_n16851, new_n16850, new_n16843);
nand_4 g14503(new_n16852, new_n16851, new_n16841_1);
xor_3  g14504(new_n16853, new_n16852, new_n16839);
xnor_3 g14505(new_n16854, new_n16853, new_n16838);
not_3  g14506(new_n16855, new_n16854);
xnor_3 g14507(new_n16856, new_n16835, new_n16828);
nand_4 g14508(new_n16857, new_n16843, new_n16841_1);
xor_3  g14509(new_n16858, new_n16857, new_n16850);
not_3  g14510(new_n16859, new_n16858);
nand_4 g14511(new_n16860, new_n16859, new_n16856);
xnor_3 g14512(new_n16861, new_n16858, new_n16856);
xor_3  g14513(new_n16862, n13714, new_n6772);
xor_3  g14514(new_n16863, new_n16470, new_n8627);
nor_4  g14515(new_n16864, new_n16863, new_n16862);
nor_4  g14516(new_n16865, new_n16846, new_n16844);
xor_3  g14517(new_n16866, new_n16865, new_n16848);
not_3  g14518(new_n16867, new_n16866);
nor_4  g14519(new_n16868, new_n16867, new_n16864);
not_3  g14520(new_n16869, new_n16868);
xor_3  g14521(new_n16870, new_n16832, new_n16831);
not_3  g14522(new_n16871, new_n16864);
nor_4  g14523(new_n16872, new_n16866, new_n16871);
nor_4  g14524(new_n16873, new_n16872, new_n16868);
nand_4 g14525(new_n16874, new_n16873, new_n16870);
nand_4 g14526(new_n16875, new_n16874, new_n16869);
nand_4 g14527(new_n16876, new_n16875, new_n16861);
nand_4 g14528(new_n16877, new_n16876, new_n16860);
xor_3  g14529(n2703, new_n16877, new_n16855);
not_3  g14530(new_n16879, new_n15587);
xor_3  g14531(n2706, new_n15602_1, new_n16879);
not_3  g14532(new_n16881, n1831);
nor_4  g14533(new_n16882, n3320, new_n16881);
xor_3  g14534(new_n16883, n3320, new_n16881);
not_3  g14535(new_n16884, new_n16883);
not_3  g14536(new_n16885_1, n13137);
nor_4  g14537(new_n16886, new_n16885_1, n1288);
not_3  g14538(new_n16887, new_n16886);
xor_3  g14539(new_n16888, n13137, new_n7265);
not_3  g14540(new_n16889, n18452);
nor_4  g14541(new_n16890, new_n16889, n1752);
not_3  g14542(new_n16891, new_n16890);
xor_3  g14543(new_n16892, n18452, new_n7249);
nor_4  g14544(new_n16893, new_n7210, n13110);
not_3  g14545(new_n16894, new_n16893);
xor_3  g14546(new_n16895, n21317, new_n7250);
nor_4  g14547(new_n16896, n25694, new_n4426_1);
not_3  g14548(new_n16897, new_n16896);
xor_3  g14549(new_n16898, n25694, new_n4426_1);
not_3  g14550(new_n16899, n19789);
nor_4  g14551(new_n16900, new_n16899, n15424);
not_3  g14552(new_n16901, new_n16900);
xor_3  g14553(new_n16902, n19789, n15424);
not_3  g14554(new_n16903, new_n16902);
not_3  g14555(new_n16904, n1949);
nor_4  g14556(new_n16905_1, n20169, new_n16904);
nor_4  g14557(new_n16906, new_n14701_1, new_n14685);
nor_4  g14558(new_n16907, new_n16906, new_n16905_1);
nand_4 g14559(new_n16908, new_n16907, new_n16903);
nand_4 g14560(new_n16909, new_n16908, new_n16901);
nand_4 g14561(new_n16910, new_n16909, new_n16898);
nand_4 g14562(new_n16911_1, new_n16910, new_n16897);
nand_4 g14563(new_n16912, new_n16911_1, new_n16895);
nand_4 g14564(new_n16913, new_n16912, new_n16894);
nand_4 g14565(new_n16914, new_n16913, new_n16892);
nand_4 g14566(new_n16915, new_n16914, new_n16891);
nand_4 g14567(new_n16916, new_n16915, new_n16888);
nand_4 g14568(new_n16917, new_n16916, new_n16887);
not_3  g14569(new_n16918, new_n16917);
nor_4  g14570(new_n16919, new_n16918, new_n16884);
nor_4  g14571(new_n16920, new_n16919, new_n16882);
nor_4  g14572(new_n16921, n19539, new_n13542);
nor_4  g14573(new_n16922, new_n13560, new_n16921);
not_3  g14574(new_n16923, new_n16922);
nand_4 g14575(new_n16924, new_n7568, new_n7561);
nor_4  g14576(new_n16925, new_n16924, n3541);
xor_3  g14577(new_n16926, new_n16925, new_n14873);
nor_4  g14578(new_n16927, new_n16926, n6204);
not_3  g14579(new_n16928, new_n16926);
xor_3  g14580(new_n16929, new_n16928, n6204);
xor_3  g14581(new_n16930, new_n16924, n3541);
nor_4  g14582(new_n16931, new_n16930, n3349);
xor_3  g14583(new_n16932, new_n16924, new_n14876);
nor_4  g14584(new_n16933, new_n16932, new_n14825);
not_3  g14585(new_n16934, new_n7572_1);
nand_4 g14586(new_n16935, new_n7623, new_n7570);
nand_4 g14587(new_n16936, new_n16935, new_n16934);
not_3  g14588(new_n16937, new_n16936);
nor_4  g14589(new_n16938, new_n16937, new_n16933);
nor_4  g14590(new_n16939, new_n16938, new_n16931);
nor_4  g14591(new_n16940, new_n16939, new_n16929);
nor_4  g14592(new_n16941, new_n16940, new_n16927);
nand_4 g14593(new_n16942, new_n16925, new_n14873);
not_3  g14594(new_n16943, new_n16942);
xor_3  g14595(new_n16944, new_n16943, new_n14870);
nor_4  g14596(new_n16945, new_n16944, n5140);
not_3  g14597(new_n16946, new_n16944);
nor_4  g14598(new_n16947, new_n16946, new_n14816);
nor_4  g14599(new_n16948, new_n16947, new_n16945);
not_3  g14600(new_n16949, new_n16948);
xnor_3 g14601(new_n16950, new_n16949, new_n16941);
nor_4  g14602(new_n16951_1, new_n16950, new_n13561);
not_3  g14603(new_n16952, new_n16951_1);
xnor_3 g14604(new_n16953, new_n16950, new_n13562);
xnor_3 g14605(new_n16954_1, new_n16939, new_n16929);
nor_4  g14606(new_n16955, new_n16954_1, new_n13641);
not_3  g14607(new_n16956, new_n16955);
xnor_3 g14608(new_n16957, new_n16954_1, new_n13641);
nor_4  g14609(new_n16958, new_n16933, new_n16931);
xnor_3 g14610(new_n16959, new_n16958, new_n16936);
nand_4 g14611(new_n16960, new_n16959, new_n13650);
not_3  g14612(new_n16961, new_n16960);
nor_4  g14613(new_n16962, new_n16959, new_n13650);
nor_4  g14614(new_n16963, new_n16962, new_n16961);
nand_4 g14615(new_n16964, new_n7624, new_n13659);
nand_4 g14616(new_n16965, new_n7681, new_n7625);
nand_4 g14617(new_n16966, new_n16965, new_n16964);
nand_4 g14618(new_n16967, new_n16966, new_n16963);
nand_4 g14619(new_n16968_1, new_n16967, new_n16960);
nor_4  g14620(new_n16969, new_n16968_1, new_n16957);
not_3  g14621(new_n16970, new_n16969);
nand_4 g14622(new_n16971_1, new_n16970, new_n16956);
nand_4 g14623(new_n16972, new_n16971_1, new_n16953);
nand_4 g14624(new_n16973, new_n16972, new_n16952);
nor_4  g14625(new_n16974, new_n16942, n10018);
nor_4  g14626(new_n16975, new_n16947, new_n16941);
nor_4  g14627(new_n16976, new_n16975, new_n16945);
nor_4  g14628(new_n16977, new_n16976, new_n16974);
nor_4  g14629(new_n16978, new_n16977, new_n16973);
not_3  g14630(new_n16979, new_n16978);
nor_4  g14631(new_n16980, new_n16979, new_n16923);
nand_4 g14632(new_n16981, new_n16977, new_n16973);
nor_4  g14633(new_n16982, new_n16981, new_n16922);
nor_4  g14634(new_n16983, new_n16982, new_n16980);
nor_4  g14635(new_n16984, new_n16983, new_n16920);
not_3  g14636(new_n16985, new_n16920);
not_3  g14637(new_n16986, new_n16983);
nor_4  g14638(new_n16987, new_n16986, new_n16985);
nor_4  g14639(new_n16988_1, new_n16987, new_n16984);
not_3  g14640(new_n16989_1, new_n16977);
xnor_3 g14641(new_n16990, new_n16989_1, new_n16973);
xnor_3 g14642(new_n16991, new_n16990, new_n16923);
nor_4  g14643(new_n16992, new_n16991, new_n16985);
xnor_3 g14644(new_n16993, new_n16990, new_n16922);
nor_4  g14645(new_n16994_1, new_n16993, new_n16920);
xor_3  g14646(new_n16995, new_n16918, new_n16884);
not_3  g14647(new_n16996, new_n16995);
xnor_3 g14648(new_n16997, new_n16950, new_n13561);
xnor_3 g14649(new_n16998, new_n16971_1, new_n16997);
nand_4 g14650(new_n16999, new_n16998, new_n16996);
xnor_3 g14651(new_n17000, new_n16998, new_n16996);
not_3  g14652(new_n17001, new_n17000);
xor_3  g14653(new_n17002, new_n16915, new_n16888);
xnor_3 g14654(new_n17003, new_n16968_1, new_n16957);
nor_4  g14655(new_n17004, new_n17003, new_n17002);
not_3  g14656(new_n17005, new_n17004);
not_3  g14657(new_n17006_1, new_n17002);
not_3  g14658(new_n17007, new_n17003);
nor_4  g14659(new_n17008, new_n17007, new_n17006_1);
nor_4  g14660(new_n17009, new_n17008, new_n17004);
xor_3  g14661(new_n17010, new_n16913, new_n16892);
not_3  g14662(new_n17011, new_n17010);
xnor_3 g14663(new_n17012, new_n16966, new_n16963);
nand_4 g14664(new_n17013, new_n17012, new_n17011);
xnor_3 g14665(new_n17014, new_n17012, new_n17010);
xor_3  g14666(new_n17015, new_n16911_1, new_n16895);
not_3  g14667(new_n17016, new_n17015);
nand_4 g14668(new_n17017, new_n17016, new_n7682);
not_3  g14669(new_n17018, new_n16898);
xor_3  g14670(new_n17019, new_n16909, new_n17018);
nand_4 g14671(new_n17020, new_n17019, new_n7689);
xnor_3 g14672(new_n17021, new_n17019, new_n7686_1);
xor_3  g14673(new_n17022, new_n16907, new_n16903);
not_3  g14674(new_n17023, new_n17022);
nand_4 g14675(new_n17024, new_n17023, new_n7694);
xnor_3 g14676(new_n17025, new_n17022, new_n7694);
nand_4 g14677(new_n17026, new_n14702_1, new_n7702);
nand_4 g14678(new_n17027, new_n14724, new_n14703);
nand_4 g14679(new_n17028, new_n17027, new_n17026);
nand_4 g14680(new_n17029, new_n17028, new_n17025);
nand_4 g14681(new_n17030, new_n17029, new_n17024);
nand_4 g14682(new_n17031, new_n17030, new_n17021);
nand_4 g14683(new_n17032, new_n17031, new_n17020);
xnor_3 g14684(new_n17033, new_n17015, new_n7682);
nand_4 g14685(new_n17034, new_n17033, new_n17032);
nand_4 g14686(new_n17035_1, new_n17034, new_n17017);
nand_4 g14687(new_n17036, new_n17035_1, new_n17014);
nand_4 g14688(new_n17037_1, new_n17036, new_n17013);
nand_4 g14689(new_n17038, new_n17037_1, new_n17009);
nand_4 g14690(new_n17039, new_n17038, new_n17005);
nand_4 g14691(new_n17040, new_n17039, new_n17001);
nand_4 g14692(new_n17041, new_n17040, new_n16999);
nor_4  g14693(new_n17042, new_n17041, new_n16994_1);
nor_4  g14694(new_n17043, new_n17042, new_n16992);
not_3  g14695(new_n17044, new_n17043);
xnor_3 g14696(n2711, new_n17044, new_n16988_1);
xor_3  g14697(new_n17046, n10611, n2680);
nor_4  g14698(new_n17047, n2783, new_n10869);
not_3  g14699(new_n17048, new_n17047);
nor_4  g14700(new_n17049, new_n10907, n1667);
not_3  g14701(new_n17050, new_n17049);
not_3  g14702(new_n17051, n7339);
nor_4  g14703(new_n17052, n15490, new_n17051);
not_3  g14704(new_n17053, new_n17052);
nor_4  g14705(new_n17054, new_n10910, n7339);
not_3  g14706(new_n17055, new_n17054);
not_3  g14707(new_n17056, n26808);
nor_4  g14708(new_n17057, new_n17056, n18);
nand_4 g14709(new_n17058, new_n17057, new_n17055);
nand_4 g14710(new_n17059, new_n17058, new_n17053);
nand_4 g14711(new_n17060, new_n17059, new_n17050);
nand_4 g14712(new_n17061, new_n17060, new_n17048);
not_3  g14713(new_n17062, new_n17061);
xor_3  g14714(new_n17063, new_n17062, new_n17046);
xnor_3 g14715(new_n17064, new_n17063, new_n10819);
nand_4 g14716(new_n17065, new_n17050, new_n17048);
xor_3  g14717(new_n17066, new_n17065, new_n17059);
nor_4  g14718(new_n17067, new_n17066, new_n10825);
not_3  g14719(new_n17068_1, new_n17067);
not_3  g14720(new_n17069_1, new_n17066);
nor_4  g14721(new_n17070_1, new_n17069_1, new_n10824);
nor_4  g14722(new_n17071, new_n17070_1, new_n17067);
xor_3  g14723(new_n17072, n26808, new_n10912);
nor_4  g14724(new_n17073, new_n17072, new_n10834_1);
nor_4  g14725(new_n17074, new_n17054, new_n17052);
xor_3  g14726(new_n17075_1, new_n17074, new_n17057);
not_3  g14727(new_n17076, new_n17075_1);
nor_4  g14728(new_n17077_1, new_n17076, new_n17073);
not_3  g14729(new_n17078, new_n17077_1);
not_3  g14730(new_n17079, new_n17073);
nor_4  g14731(new_n17080, new_n17075_1, new_n17079);
nor_4  g14732(new_n17081, new_n17080, new_n17077_1);
nand_4 g14733(new_n17082, new_n17081, new_n10843);
nand_4 g14734(new_n17083, new_n17082, new_n17078);
nand_4 g14735(new_n17084_1, new_n17083, new_n17071);
nand_4 g14736(new_n17085, new_n17084_1, new_n17068_1);
not_3  g14737(new_n17086, new_n17085);
xor_3  g14738(n2761, new_n17086, new_n17064);
xor_3  g14739(new_n17088, n25120, n8526);
not_3  g14740(new_n17089, new_n17088);
nor_4  g14741(new_n17090_1, n8363, n2816);
xor_3  g14742(new_n17091, n8363, n2816);
not_3  g14743(new_n17092, new_n17091);
nor_4  g14744(new_n17093, n20359, n14680);
xor_3  g14745(new_n17094, n20359, n14680);
not_3  g14746(new_n17095_1, new_n17094);
nand_4 g14747(new_n17096, new_n9087, new_n7083);
nand_4 g14748(new_n17097, new_n11196, new_n11167);
nand_4 g14749(new_n17098, new_n17097, new_n17096);
not_3  g14750(new_n17099, new_n17098);
nor_4  g14751(new_n17100, new_n17099, new_n17095_1);
nor_4  g14752(new_n17101, new_n17100, new_n17093);
nor_4  g14753(new_n17102, new_n17101, new_n17092);
nor_4  g14754(new_n17103, new_n17102, new_n17090_1);
xnor_3 g14755(new_n17104_1, new_n17103, new_n17089);
nor_4  g14756(new_n17105, new_n17104_1, n17458);
xnor_3 g14757(new_n17106_1, new_n17104_1, n17458);
xnor_3 g14758(new_n17107, new_n17101, new_n17092);
not_3  g14759(new_n17108, new_n17107);
nor_4  g14760(new_n17109, new_n17108, new_n8501);
not_3  g14761(new_n17110, new_n17109);
nor_4  g14762(new_n17111, new_n17098, new_n17094);
nor_4  g14763(new_n17112, new_n17111, new_n17100);
not_3  g14764(new_n17113, new_n17112);
nor_4  g14765(new_n17114, new_n17113, n25240);
xnor_3 g14766(new_n17115, new_n17112, new_n8503);
nor_4  g14767(new_n17116, new_n11198, new_n8506);
not_3  g14768(new_n17117, new_n17116);
nor_4  g14769(new_n17118, new_n11197, n10125);
nor_4  g14770(new_n17119_1, new_n17118, new_n17116);
nor_4  g14771(new_n17120, new_n11203, new_n8509);
not_3  g14772(new_n17121, new_n17120);
nor_4  g14773(new_n17122, new_n11202, n8067);
nor_4  g14774(new_n17123, new_n17122, new_n17120);
nor_4  g14775(new_n17124, new_n11209, new_n12653);
not_3  g14776(new_n17125, new_n17124);
nor_4  g14777(new_n17126, new_n11208, n20923);
nor_4  g14778(new_n17127, new_n17126, new_n17124);
nand_4 g14779(new_n17128, new_n11215, n18157);
not_3  g14780(new_n17129, new_n17128);
nor_4  g14781(new_n17130_1, new_n11215, n18157);
nor_4  g14782(new_n17131, new_n17130_1, new_n17129);
nor_4  g14783(new_n17132, new_n11220_1, new_n7792);
not_3  g14784(new_n17133, new_n17132);
nor_4  g14785(new_n17134, new_n11226, n5026);
nor_4  g14786(new_n17135, new_n11228, new_n8626);
xnor_3 g14787(new_n17136, new_n11225, new_n8524);
nor_4  g14788(new_n17137, new_n17136, new_n17135);
nor_4  g14789(new_n17138_1, new_n17137, new_n17134);
not_3  g14790(new_n17139, new_n11220_1);
nor_4  g14791(new_n17140, new_n17139, n12161);
nor_4  g14792(new_n17141, new_n17140, new_n17132);
nand_4 g14793(new_n17142, new_n17141, new_n17138_1);
nand_4 g14794(new_n17143, new_n17142, new_n17133);
nand_4 g14795(new_n17144, new_n17143, new_n17131);
nand_4 g14796(new_n17145, new_n17144, new_n17128);
nand_4 g14797(new_n17146, new_n17145, new_n17127);
nand_4 g14798(new_n17147, new_n17146, new_n17125);
nand_4 g14799(new_n17148, new_n17147, new_n17123);
nand_4 g14800(new_n17149, new_n17148, new_n17121);
nand_4 g14801(new_n17150, new_n17149, new_n17119_1);
nand_4 g14802(new_n17151, new_n17150, new_n17117);
nor_4  g14803(new_n17152, new_n17151, new_n17115);
nor_4  g14804(new_n17153, new_n17152, new_n17114);
nor_4  g14805(new_n17154, new_n17107, n1222);
nor_4  g14806(new_n17155, new_n17154, new_n17109);
nand_4 g14807(new_n17156, new_n17155, new_n17153);
nand_4 g14808(new_n17157, new_n17156, new_n17110);
nor_4  g14809(new_n17158, new_n17157, new_n17106_1);
nor_4  g14810(new_n17159, new_n17158, new_n17105);
nor_4  g14811(new_n17160, n25120, n8526);
nor_4  g14812(new_n17161, new_n17103, new_n17089);
nor_4  g14813(new_n17162, new_n17161, new_n17160);
nand_4 g14814(new_n17163_1, new_n17162, new_n17159);
not_3  g14815(new_n17164, n11898);
nand_4 g14816(new_n17165, new_n4081, new_n4074);
nor_4  g14817(new_n17166, new_n17165, n1099);
not_3  g14818(new_n17167, new_n17166);
nor_4  g14819(new_n17168_1, new_n17167, n19941);
xor_3  g14820(new_n17169, new_n17168_1, new_n17164);
nor_4  g14821(new_n17170, new_n17169, new_n5518);
not_3  g14822(new_n17171, new_n17169);
nor_4  g14823(new_n17172, new_n17171, new_n5519);
nor_4  g14824(new_n17173, new_n17172, new_n17170);
not_3  g14825(new_n17174, new_n17173);
not_3  g14826(new_n17175, new_n5522);
xor_3  g14827(new_n17176, new_n17167, n19941);
nor_4  g14828(new_n17177, new_n17176, new_n17175);
not_3  g14829(new_n17178, new_n17176);
nor_4  g14830(new_n17179, new_n17178, new_n5522);
nor_4  g14831(new_n17180, new_n17179, new_n17177);
not_3  g14832(new_n17181, new_n17180);
not_3  g14833(new_n17182, new_n5527);
xor_3  g14834(new_n17183, new_n17165, n1099);
nor_4  g14835(new_n17184, new_n17183, new_n17182);
not_3  g14836(new_n17185, new_n17183);
nor_4  g14837(new_n17186, new_n17185, new_n5527);
nor_4  g14838(new_n17187, new_n17186, new_n17184);
nor_4  g14839(new_n17188, new_n5532_1, new_n4082);
not_3  g14840(new_n17189, new_n17188);
nor_4  g14841(new_n17190, new_n5531, new_n4083);
nor_4  g14842(new_n17191, new_n17190, new_n17188);
nor_4  g14843(new_n17192, new_n5537, new_n4085_1);
not_3  g14844(new_n17193, new_n17192);
nor_4  g14845(new_n17194, new_n5536, new_n4087);
nor_4  g14846(new_n17195, new_n17194, new_n17192);
nor_4  g14847(new_n17196, new_n5542, new_n4091);
not_3  g14848(new_n17197, new_n17196);
nor_4  g14849(new_n17198, new_n5541, new_n4094);
nor_4  g14850(new_n17199, new_n17198, new_n17196);
nor_4  g14851(new_n17200, new_n5547, new_n4099);
not_3  g14852(new_n17201, new_n17200);
nor_4  g14853(new_n17202_1, new_n15686, new_n4124);
nor_4  g14854(new_n17203, new_n17202_1, new_n17200);
nor_4  g14855(new_n17204, new_n5554, new_n4104);
not_3  g14856(new_n17205, new_n17204);
nor_4  g14857(new_n17206, new_n6818, new_n4108);
nor_4  g14858(new_n17207, new_n17206, new_n17204);
nand_4 g14859(new_n17208, new_n6853_1, new_n8680);
nor_4  g14860(new_n17209, new_n17208, n13319);
not_3  g14861(new_n17210, new_n17209);
nor_4  g14862(new_n17211, new_n5560, n25435);
nor_4  g14863(new_n17212, new_n17211, new_n4111);
nor_4  g14864(new_n17213, new_n17212, new_n17209);
nand_4 g14865(new_n17214, new_n17213, new_n5556);
nand_4 g14866(new_n17215, new_n17214, new_n17210);
nand_4 g14867(new_n17216, new_n17215, new_n17207);
nand_4 g14868(new_n17217, new_n17216, new_n17205);
nand_4 g14869(new_n17218, new_n17217, new_n17203);
nand_4 g14870(new_n17219_1, new_n17218, new_n17201);
nand_4 g14871(new_n17220, new_n17219_1, new_n17199);
nand_4 g14872(new_n17221, new_n17220, new_n17197);
nand_4 g14873(new_n17222, new_n17221, new_n17195);
nand_4 g14874(new_n17223, new_n17222, new_n17193);
nand_4 g14875(new_n17224, new_n17223, new_n17191);
nand_4 g14876(new_n17225, new_n17224, new_n17189);
nand_4 g14877(new_n17226, new_n17225, new_n17187);
not_3  g14878(new_n17227, new_n17226);
nor_4  g14879(new_n17228, new_n17227, new_n17184);
nor_4  g14880(new_n17229, new_n17228, new_n17181);
nor_4  g14881(new_n17230, new_n17229, new_n17177);
nor_4  g14882(new_n17231, new_n17230, new_n17174);
nor_4  g14883(new_n17232_1, new_n17231, new_n17170);
not_3  g14884(new_n17233, new_n17168_1);
nor_4  g14885(new_n17234, new_n17233, n11898);
not_3  g14886(new_n17235, new_n17234);
nor_4  g14887(new_n17236_1, new_n17235, new_n5590);
nand_4 g14888(new_n17237, new_n17236_1, new_n17232_1);
not_3  g14889(new_n17238, new_n17232_1);
not_3  g14890(new_n17239, new_n5590);
nor_4  g14891(new_n17240, new_n17234, new_n17239);
nand_4 g14892(new_n17241, new_n17240, new_n17238);
nand_4 g14893(new_n17242, new_n17241, new_n17237);
nor_4  g14894(new_n17243_1, new_n17242, new_n17163_1);
nand_4 g14895(new_n17244, new_n17242, new_n17163_1);
not_3  g14896(new_n17245, new_n17162);
xnor_3 g14897(new_n17246, new_n17245, new_n17159);
nor_4  g14898(new_n17247, new_n17240, new_n17236_1);
xnor_3 g14899(new_n17248, new_n17247, new_n17232_1);
nor_4  g14900(new_n17249, new_n17248, new_n17246);
xnor_3 g14901(new_n17250_1, new_n17248, new_n17246);
xnor_3 g14902(new_n17251_1, new_n17157, new_n17106_1);
not_3  g14903(new_n17252, new_n17230);
nor_4  g14904(new_n17253, new_n17252, new_n17173);
nor_4  g14905(new_n17254, new_n17253, new_n17231);
not_3  g14906(new_n17255, new_n17254);
nor_4  g14907(new_n17256, new_n17255, new_n17251_1);
xnor_3 g14908(new_n17257, new_n17255, new_n17251_1);
xnor_3 g14909(new_n17258, new_n17228, new_n17181);
not_3  g14910(new_n17259, new_n17155);
xnor_3 g14911(new_n17260, new_n17259, new_n17153);
nor_4  g14912(new_n17261, new_n17260, new_n17258);
xnor_3 g14913(new_n17262, new_n17260, new_n17258);
nand_4 g14914(new_n17263_1, new_n17151, new_n17115);
not_3  g14915(new_n17264, new_n17263_1);
nor_4  g14916(new_n17265, new_n17264, new_n17152);
xnor_3 g14917(new_n17266, new_n17225, new_n17187);
not_3  g14918(new_n17267, new_n17266);
nand_4 g14919(new_n17268, new_n17267, new_n17265);
xnor_3 g14920(new_n17269, new_n17266, new_n17265);
xnor_3 g14921(new_n17270, new_n17223, new_n17191);
not_3  g14922(new_n17271, new_n17270);
xnor_3 g14923(new_n17272, new_n17149, new_n17119_1);
nand_4 g14924(new_n17273, new_n17272, new_n17271);
xnor_3 g14925(new_n17274, new_n17272, new_n17270);
xnor_3 g14926(new_n17275, new_n17221, new_n17195);
not_3  g14927(new_n17276, new_n17275);
xnor_3 g14928(new_n17277, new_n17147, new_n17123);
nand_4 g14929(new_n17278, new_n17277, new_n17276);
xnor_3 g14930(new_n17279, new_n17277, new_n17275);
not_3  g14931(new_n17280, new_n17199);
xnor_3 g14932(new_n17281, new_n17219_1, new_n17280);
xnor_3 g14933(new_n17282, new_n17145, new_n17127);
nand_4 g14934(new_n17283, new_n17282, new_n17281);
not_3  g14935(new_n17284, new_n17282);
xnor_3 g14936(new_n17285_1, new_n17284, new_n17281);
xnor_3 g14937(new_n17286, new_n17217, new_n17203);
xnor_3 g14938(new_n17287, new_n17143, new_n17131);
not_3  g14939(new_n17288, new_n17287);
nor_4  g14940(new_n17289, new_n17288, new_n17286);
not_3  g14941(new_n17290, new_n17289);
not_3  g14942(new_n17291, new_n17286);
nor_4  g14943(new_n17292, new_n17287, new_n17291);
nor_4  g14944(new_n17293, new_n17292, new_n17289);
not_3  g14945(new_n17294, new_n17216);
nor_4  g14946(new_n17295, new_n17215, new_n17207);
nor_4  g14947(new_n17296, new_n17295, new_n17294);
not_3  g14948(new_n17297, new_n17142);
nor_4  g14949(new_n17298, new_n17141, new_n17138_1);
nor_4  g14950(new_n17299, new_n17298, new_n17297);
not_3  g14951(new_n17300, new_n17299);
nor_4  g14952(new_n17301, new_n17300, new_n17296);
xnor_3 g14953(new_n17302_1, new_n17300, new_n17296);
xnor_3 g14954(new_n17303, new_n17136, new_n17135);
not_3  g14955(new_n17304, new_n17303);
xor_3  g14956(new_n17305, new_n17213, new_n5556);
nand_4 g14957(new_n17306, new_n17305, new_n17304);
xor_3  g14958(new_n17307, new_n11228, new_n8626);
xor_3  g14959(new_n17308, new_n5560, n25435);
not_3  g14960(new_n17309, new_n17308);
nand_4 g14961(new_n17310, new_n17309, new_n17307);
not_3  g14962(new_n17311, new_n17306);
nor_4  g14963(new_n17312, new_n17305, new_n17304);
nor_4  g14964(new_n17313, new_n17312, new_n17311);
nand_4 g14965(new_n17314, new_n17313, new_n17310);
nand_4 g14966(new_n17315, new_n17314, new_n17306);
nor_4  g14967(new_n17316, new_n17315, new_n17302_1);
nor_4  g14968(new_n17317, new_n17316, new_n17301);
nand_4 g14969(new_n17318, new_n17317, new_n17293);
nand_4 g14970(new_n17319, new_n17318, new_n17290);
nand_4 g14971(new_n17320_1, new_n17319, new_n17285_1);
nand_4 g14972(new_n17321, new_n17320_1, new_n17283);
nand_4 g14973(new_n17322, new_n17321, new_n17279);
nand_4 g14974(new_n17323, new_n17322, new_n17278);
nand_4 g14975(new_n17324, new_n17323, new_n17274);
nand_4 g14976(new_n17325, new_n17324, new_n17273);
nand_4 g14977(new_n17326, new_n17325, new_n17269);
nand_4 g14978(new_n17327, new_n17326, new_n17268);
not_3  g14979(new_n17328, new_n17327);
nor_4  g14980(new_n17329, new_n17328, new_n17262);
nor_4  g14981(new_n17330, new_n17329, new_n17261);
nor_4  g14982(new_n17331, new_n17330, new_n17257);
nor_4  g14983(new_n17332, new_n17331, new_n17256);
nor_4  g14984(new_n17333, new_n17332, new_n17250_1);
nor_4  g14985(new_n17334, new_n17333, new_n17249);
nand_4 g14986(new_n17335, new_n17334, new_n17244);
nand_4 g14987(new_n17336, new_n17335, new_n17237);
nor_4  g14988(n2774, new_n17336, new_n17243_1);
not_3  g14989(new_n17338, n2858);
nand_4 g14990(new_n17339, new_n11297, new_n7036);
nor_4  g14991(new_n17340, new_n17339, n2421);
nand_4 g14992(new_n17341, new_n17340, new_n7030);
nor_4  g14993(new_n17342, new_n17341, n5031);
xor_3  g14994(new_n17343, new_n17342, new_n9080);
not_3  g14995(new_n17344_1, new_n17343);
nor_4  g14996(new_n17345, new_n17344_1, new_n17338);
nor_4  g14997(new_n17346, new_n17343, n2858);
nor_4  g14998(new_n17347, new_n17346, new_n17345);
xor_3  g14999(new_n17348, new_n17341, n5031);
not_3  g15000(new_n17349, new_n17348);
nor_4  g15001(new_n17350, new_n17349, new_n5602);
nor_4  g15002(new_n17351_1, new_n17348, n2659);
xor_3  g15003(new_n17352, new_n17340, new_n7030);
not_3  g15004(new_n17353, new_n17352);
nor_4  g15005(new_n17354, new_n17353, new_n5606);
nor_4  g15006(new_n17355, new_n17352, n24327);
nand_4 g15007(new_n17356, new_n17339, n2421);
not_3  g15008(new_n17357, new_n17356);
nor_4  g15009(new_n17358, new_n17357, new_n17340);
nor_4  g15010(new_n17359_1, new_n17358, n22198);
not_3  g15011(new_n17360, new_n17359_1);
xnor_3 g15012(new_n17361, new_n11297, n987);
not_3  g15013(new_n17362, new_n17361);
nor_4  g15014(new_n17363, new_n17362, new_n5641);
nor_4  g15015(new_n17364, new_n17361, n20826);
nor_4  g15016(new_n17365, new_n17364, new_n17363);
nand_4 g15017(new_n17366, new_n11300, n7305);
nand_4 g15018(new_n17367, new_n11317, new_n11301);
nand_4 g15019(new_n17368, new_n17367, new_n17366);
nand_4 g15020(new_n17369, new_n17368, new_n17365);
not_3  g15021(new_n17370, new_n17369);
nor_4  g15022(new_n17371, new_n17370, new_n17363);
not_3  g15023(new_n17372, new_n17358);
nor_4  g15024(new_n17373, new_n17372, new_n5610);
nor_4  g15025(new_n17374, new_n17373, new_n17359_1);
nand_4 g15026(new_n17375, new_n17374, new_n17371);
nand_4 g15027(new_n17376, new_n17375, new_n17360);
nor_4  g15028(new_n17377, new_n17376, new_n17355);
nor_4  g15029(new_n17378, new_n17377, new_n17354);
nor_4  g15030(new_n17379, new_n17378, new_n17351_1);
nor_4  g15031(new_n17380, new_n17379, new_n17350);
xnor_3 g15032(new_n17381, new_n17380, new_n17347);
not_3  g15033(new_n17382, new_n17381);
nor_4  g15034(new_n17383, new_n17382, new_n3750);
nor_4  g15035(new_n17384, new_n17381, new_n3747);
nor_4  g15036(new_n17385, new_n17384, new_n17383);
not_3  g15037(new_n17386, new_n17385);
nor_4  g15038(new_n17387_1, new_n17351_1, new_n17350);
xnor_3 g15039(new_n17388, new_n17387_1, new_n17378);
not_3  g15040(new_n17389, new_n17388);
nor_4  g15041(new_n17390, new_n17389, new_n3756);
not_3  g15042(new_n17391_1, new_n17390);
xor_3  g15043(new_n17392_1, new_n17353, new_n5606);
xnor_3 g15044(new_n17393, new_n17392_1, new_n17376);
nor_4  g15045(new_n17394, new_n17393, new_n3761);
not_3  g15046(new_n17395, new_n17393);
nor_4  g15047(new_n17396, new_n17395, new_n3760_1);
nor_4  g15048(new_n17397, new_n17396, new_n17394);
not_3  g15049(new_n17398, new_n17397);
xnor_3 g15050(new_n17399, new_n17374, new_n17371);
nor_4  g15051(new_n17400, new_n17399, new_n3772);
not_3  g15052(new_n17401, new_n17399);
nor_4  g15053(new_n17402, new_n17401, new_n3770);
nor_4  g15054(new_n17403, new_n17402, new_n17400);
not_3  g15055(new_n17404, new_n17403);
nor_4  g15056(new_n17405, new_n17368, new_n17365);
nor_4  g15057(new_n17406, new_n17405, new_n17370);
nor_4  g15058(new_n17407, new_n17406, new_n3776);
xnor_3 g15059(new_n17408, new_n17368, new_n17365);
nor_4  g15060(new_n17409, new_n17408, new_n3780);
nor_4  g15061(new_n17410, new_n17409, new_n17407);
not_3  g15062(new_n17411, new_n17410);
nor_4  g15063(new_n17412, new_n11318, new_n3787);
not_3  g15064(new_n17413, new_n17412);
nor_4  g15065(new_n17414, new_n11348_1, new_n3783);
nor_4  g15066(new_n17415, new_n17414, new_n17412);
nor_4  g15067(new_n17416, new_n11353, new_n3792);
not_3  g15068(new_n17417, new_n17416);
nor_4  g15069(new_n17418, new_n11357, new_n3791);
nor_4  g15070(new_n17419, new_n17418, new_n17416);
nor_4  g15071(new_n17420, new_n11360, new_n3799);
not_3  g15072(new_n17421_1, new_n17420);
nand_4 g15073(new_n17422, new_n11363, new_n3801);
nor_4  g15074(new_n17423, new_n11366, new_n3798);
nor_4  g15075(new_n17424, new_n17423, new_n17420);
not_3  g15076(new_n17425, new_n17424);
nor_4  g15077(new_n17426, new_n17425, new_n17422);
not_3  g15078(new_n17427, new_n17426);
nand_4 g15079(new_n17428, new_n17427, new_n17421_1);
nand_4 g15080(new_n17429, new_n17428, new_n17419);
nand_4 g15081(new_n17430, new_n17429, new_n17417);
nand_4 g15082(new_n17431, new_n17430, new_n17415);
nand_4 g15083(new_n17432_1, new_n17431, new_n17413);
nor_4  g15084(new_n17433, new_n17432_1, new_n17411);
nor_4  g15085(new_n17434, new_n17433, new_n17407);
nor_4  g15086(new_n17435, new_n17434, new_n17404);
nor_4  g15087(new_n17436_1, new_n17435, new_n17400);
nor_4  g15088(new_n17437, new_n17436_1, new_n17398);
nor_4  g15089(new_n17438, new_n17437, new_n17394);
not_3  g15090(new_n17439, new_n3756);
nor_4  g15091(new_n17440_1, new_n17388, new_n17439);
nor_4  g15092(new_n17441, new_n17440_1, new_n17390);
nand_4 g15093(new_n17442, new_n17441, new_n17438);
nand_4 g15094(new_n17443, new_n17442, new_n17391_1);
xnor_3 g15095(new_n17444, new_n17443, new_n17386);
nand_4 g15096(new_n17445, new_n3898, n7026);
nand_4 g15097(new_n17446, new_n3899, new_n3828_1);
nand_4 g15098(new_n17447, new_n17446, new_n17445);
nand_4 g15099(new_n17448, new_n3905, n13719);
nand_4 g15100(new_n17449, new_n3909_1, new_n3831);
nor_4  g15101(new_n17450_1, new_n3914, n442);
xor_3  g15102(new_n17451, new_n3918_1, new_n3836);
not_3  g15103(new_n17452, new_n17451);
nor_4  g15104(new_n17453, new_n3921, n9172);
xor_3  g15105(new_n17454, new_n3922, new_n3840);
not_3  g15106(new_n17455, new_n17454);
nor_4  g15107(new_n17456, new_n3929, n4913);
xor_3  g15108(new_n17457, new_n3929, n4913);
nand_4 g15109(new_n17458_1, new_n3969, new_n3846);
nor_4  g15110(new_n17459, new_n3944, n16824);
not_3  g15111(new_n17460, new_n17459);
xor_3  g15112(new_n17461_1, new_n3950, new_n3852);
nor_4  g15113(new_n17462, new_n3953, n16521);
not_3  g15114(new_n17463, new_n17462);
nand_4 g15115(new_n17464, n21993, n7139);
xor_3  g15116(new_n17465, new_n3954, new_n3856);
nand_4 g15117(new_n17466_1, new_n17465, new_n17464);
nand_4 g15118(new_n17467, new_n17466_1, new_n17463);
nand_4 g15119(new_n17468, new_n17467, new_n17461_1);
nand_4 g15120(new_n17469, new_n17468, new_n17460);
xor_3  g15121(new_n17470, new_n3969, new_n3846);
nand_4 g15122(new_n17471, new_n17470, new_n17469);
nand_4 g15123(new_n17472, new_n17471, new_n17458_1);
nand_4 g15124(new_n17473, new_n17472, new_n17457);
not_3  g15125(new_n17474, new_n17473);
nor_4  g15126(new_n17475, new_n17474, new_n17456);
nor_4  g15127(new_n17476, new_n17475, new_n17455);
nor_4  g15128(new_n17477, new_n17476, new_n17453);
nor_4  g15129(new_n17478, new_n17477, new_n17452);
nor_4  g15130(new_n17479, new_n17478, new_n17450_1);
nand_4 g15131(new_n17480, new_n17479, new_n17449);
nand_4 g15132(new_n17481, new_n17480, new_n17448);
xnor_3 g15133(new_n17482, new_n17481, new_n17447);
xnor_3 g15134(new_n17483, new_n17482, new_n17444);
not_3  g15135(new_n17484, new_n17394);
not_3  g15136(new_n17485, new_n17400);
not_3  g15137(new_n17486, new_n17434);
nand_4 g15138(new_n17487, new_n17486, new_n17403);
nand_4 g15139(new_n17488, new_n17487, new_n17485);
nand_4 g15140(new_n17489, new_n17488, new_n17397);
nand_4 g15141(new_n17490, new_n17489, new_n17484);
not_3  g15142(new_n17491, new_n17441);
nor_4  g15143(new_n17492, new_n17491, new_n17490);
nor_4  g15144(new_n17493_1, new_n17441, new_n17438);
nor_4  g15145(new_n17494, new_n17493_1, new_n17492);
not_3  g15146(new_n17495, new_n17494);
nand_4 g15147(new_n17496, new_n17449, new_n17448);
not_3  g15148(new_n17497, new_n17496);
xnor_3 g15149(new_n17498, new_n17497, new_n17479);
nor_4  g15150(new_n17499, new_n17498, new_n17495);
not_3  g15151(new_n17500_1, new_n17499);
xnor_3 g15152(new_n17501, new_n17498, new_n17494);
xnor_3 g15153(new_n17502, new_n17477, new_n17451);
not_3  g15154(new_n17503, new_n17502);
xnor_3 g15155(new_n17504, new_n17488, new_n17397);
nor_4  g15156(new_n17505, new_n17504, new_n17503);
xnor_3 g15157(new_n17506, new_n17504, new_n17503);
xnor_3 g15158(new_n17507, new_n17475, new_n17455);
xnor_3 g15159(new_n17508, new_n17486, new_n17403);
nor_4  g15160(new_n17509, new_n17508, new_n17507);
xnor_3 g15161(new_n17510, new_n17508, new_n17507);
xnor_3 g15162(new_n17511, new_n17472, new_n17457);
not_3  g15163(new_n17512, new_n17432_1);
nor_4  g15164(new_n17513, new_n17512, new_n17410);
nor_4  g15165(new_n17514, new_n17513, new_n17433);
not_3  g15166(new_n17515, new_n17514);
nand_4 g15167(new_n17516, new_n17515, new_n17511);
xnor_3 g15168(new_n17517, new_n17470, new_n17469);
not_3  g15169(new_n17518, new_n17517);
xnor_3 g15170(new_n17519, new_n17430, new_n17415);
nor_4  g15171(new_n17520, new_n17519, new_n17518);
not_3  g15172(new_n17521, new_n17520);
not_3  g15173(new_n17522, new_n17519);
nor_4  g15174(new_n17523, new_n17522, new_n17517);
nor_4  g15175(new_n17524_1, new_n17523, new_n17520);
xnor_3 g15176(new_n17525, new_n17467, new_n17461_1);
not_3  g15177(new_n17526, new_n17525);
not_3  g15178(new_n17527, new_n17419);
nor_4  g15179(new_n17528, new_n17426, new_n17420);
nor_4  g15180(new_n17529_1, new_n17528, new_n17527);
nor_4  g15181(new_n17530, new_n17428, new_n17419);
nor_4  g15182(new_n17531, new_n17530, new_n17529_1);
not_3  g15183(new_n17532, new_n17531);
nor_4  g15184(new_n17533, new_n17532, new_n17526);
not_3  g15185(new_n17534, new_n17533);
nor_4  g15186(new_n17535, new_n17531, new_n17525);
nor_4  g15187(new_n17536, new_n17535, new_n17533);
xnor_3 g15188(new_n17537, new_n17425, new_n17422);
not_3  g15189(new_n17538, new_n17537);
nor_4  g15190(new_n17539, new_n17538, new_n17465);
not_3  g15191(new_n17540, new_n17466_1);
nor_4  g15192(new_n17541, new_n17465, new_n17464);
nor_4  g15193(new_n17542, new_n17541, new_n17540);
nor_4  g15194(new_n17543, new_n17542, new_n17537);
xor_3  g15195(new_n17544, n21993, n7139);
not_3  g15196(new_n17545, new_n17544);
xnor_3 g15197(new_n17546, new_n11363, new_n3801);
nor_4  g15198(new_n17547, new_n17546, new_n17545);
nor_4  g15199(new_n17548, new_n17547, new_n17543);
nor_4  g15200(new_n17549, new_n17548, new_n17539);
nand_4 g15201(new_n17550, new_n17549, new_n17536);
nand_4 g15202(new_n17551, new_n17550, new_n17534);
nand_4 g15203(new_n17552, new_n17551, new_n17524_1);
nand_4 g15204(new_n17553, new_n17552, new_n17521);
xnor_3 g15205(new_n17554, new_n17514, new_n17511);
nand_4 g15206(new_n17555, new_n17554, new_n17553);
nand_4 g15207(new_n17556, new_n17555, new_n17516);
nor_4  g15208(new_n17557_1, new_n17556, new_n17510);
nor_4  g15209(new_n17558, new_n17557_1, new_n17509);
nor_4  g15210(new_n17559, new_n17558, new_n17506);
nor_4  g15211(new_n17560, new_n17559, new_n17505);
nand_4 g15212(new_n17561, new_n17560, new_n17501);
nand_4 g15213(new_n17562, new_n17561, new_n17500_1);
not_3  g15214(new_n17563, new_n17562);
xor_3  g15215(n2779, new_n17563, new_n17483);
not_3  g15216(new_n17565, new_n12559);
nor_4  g15217(new_n17566, new_n12401, n25751);
not_3  g15218(new_n17567, new_n17566);
xor_3  g15219(new_n17568, new_n12402, n25751);
not_3  g15220(new_n17569, new_n17568);
nor_4  g15221(new_n17570, new_n12408_1, n26053);
not_3  g15222(new_n17571, new_n17570);
not_3  g15223(new_n17572, n26053);
nor_4  g15224(new_n17573, new_n12406, new_n17572);
nor_4  g15225(new_n17574, new_n17573, new_n17570);
nor_4  g15226(new_n17575, new_n12411, n7917);
not_3  g15227(new_n17576, n7917);
not_3  g15228(new_n17577, new_n12411);
nor_4  g15229(new_n17578, new_n17577, new_n17576);
nor_4  g15230(new_n17579, new_n17578, new_n17575);
not_3  g15231(new_n17580, new_n17579);
nor_4  g15232(new_n17581, new_n12417, n17302);
xnor_3 g15233(new_n17582, new_n12417, n17302);
nor_4  g15234(new_n17583_1, new_n12422, n2013);
not_3  g15235(new_n17584, n2013);
nor_4  g15236(new_n17585, new_n12425, new_n17584);
nor_4  g15237(new_n17586, new_n17585, new_n17583_1);
nor_4  g15238(new_n17587, new_n12430, n23755);
not_3  g15239(new_n17588, new_n17587);
not_3  g15240(new_n17589, new_n12434);
nor_4  g15241(new_n17590, new_n17589, n19163);
not_3  g15242(new_n17591, new_n17590);
not_3  g15243(new_n17592_1, n19163);
nor_4  g15244(new_n17593, new_n12434, new_n17592_1);
nor_4  g15245(new_n17594, new_n17593, new_n17590);
not_3  g15246(new_n17595, n22358);
nand_4 g15247(new_n17596, new_n6797, new_n17595);
nand_4 g15248(new_n17597, n25926, n9646);
xnor_3 g15249(new_n17598, new_n6797, n22358);
nand_4 g15250(new_n17599, new_n17598, new_n17597);
nand_4 g15251(new_n17600, new_n17599, new_n17596);
nand_4 g15252(new_n17601, new_n17600, new_n17594);
nand_4 g15253(new_n17602, new_n17601, new_n17591);
not_3  g15254(new_n17603, n23755);
nor_4  g15255(new_n17604, new_n12431, new_n17603);
nor_4  g15256(new_n17605, new_n17604, new_n17587);
nand_4 g15257(new_n17606, new_n17605, new_n17602);
nand_4 g15258(new_n17607, new_n17606, new_n17588);
nand_4 g15259(new_n17608, new_n17607, new_n17586);
not_3  g15260(new_n17609, new_n17608);
nor_4  g15261(new_n17610, new_n17609, new_n17583_1);
nor_4  g15262(new_n17611, new_n17610, new_n17582);
nor_4  g15263(new_n17612, new_n17611, new_n17581);
nor_4  g15264(new_n17613, new_n17612, new_n17580);
nor_4  g15265(new_n17614, new_n17613, new_n17575);
not_3  g15266(new_n17615, new_n17614);
nand_4 g15267(new_n17616, new_n17615, new_n17574);
nand_4 g15268(new_n17617, new_n17616, new_n17571);
nand_4 g15269(new_n17618, new_n17617, new_n17569);
nand_4 g15270(new_n17619, new_n17618, new_n17567);
not_3  g15271(new_n17620, n25586);
xor_3  g15272(new_n17621, new_n12454, new_n17620);
not_3  g15273(new_n17622, new_n17621);
xnor_3 g15274(new_n17623, new_n17622, new_n17619);
xnor_3 g15275(new_n17624, new_n17623, new_n13897);
not_3  g15276(new_n17625, new_n17624);
xnor_3 g15277(new_n17626, new_n17617, new_n17568);
nor_4  g15278(new_n17627, new_n17626, n3984);
xnor_3 g15279(new_n17628, new_n17626, n3984);
xnor_3 g15280(new_n17629, new_n17614, new_n17574);
nor_4  g15281(new_n17630, new_n17629, n19652);
xnor_3 g15282(new_n17631, new_n17629, n19652);
xnor_3 g15283(new_n17632, new_n17612, new_n17579);
nor_4  g15284(new_n17633, new_n17632, n3366);
not_3  g15285(new_n17634, new_n17582);
xnor_3 g15286(new_n17635, new_n17610, new_n17634);
nor_4  g15287(new_n17636, new_n17635, n26565);
xnor_3 g15288(new_n17637, new_n17635, n26565);
xnor_3 g15289(new_n17638_1, new_n17607, new_n17586);
nand_4 g15290(new_n17639, new_n17638_1, new_n13921);
xnor_3 g15291(new_n17640, new_n17638_1, n3959);
xnor_3 g15292(new_n17641, new_n17605, new_n17602);
nand_4 g15293(new_n17642, new_n17641, new_n13926);
xnor_3 g15294(new_n17643, new_n17641, n11566);
xnor_3 g15295(new_n17644, new_n17600, new_n17594);
nand_4 g15296(new_n17645, new_n17644, new_n13931);
xnor_3 g15297(new_n17646, new_n17598, new_n17597);
nand_4 g15298(new_n17647, new_n17646, new_n13935);
not_3  g15299(new_n17648, new_n7730);
nor_4  g15300(new_n17649, new_n17648, new_n7729);
not_3  g15301(new_n17650, new_n17649);
xnor_3 g15302(new_n17651, new_n17646, n26625);
nand_4 g15303(new_n17652, new_n17651, new_n17650);
nand_4 g15304(new_n17653, new_n17652, new_n17647);
xnor_3 g15305(new_n17654, new_n17644, n26744);
nand_4 g15306(new_n17655, new_n17654, new_n17653);
nand_4 g15307(new_n17656, new_n17655, new_n17645);
nand_4 g15308(new_n17657, new_n17656, new_n17643);
nand_4 g15309(new_n17658, new_n17657, new_n17642);
nand_4 g15310(new_n17659, new_n17658, new_n17640);
nand_4 g15311(new_n17660, new_n17659, new_n17639);
not_3  g15312(new_n17661, new_n17660);
nor_4  g15313(new_n17662, new_n17661, new_n17637);
nor_4  g15314(new_n17663, new_n17662, new_n17636);
xnor_3 g15315(new_n17664_1, new_n17632, n3366);
nor_4  g15316(new_n17665, new_n17664_1, new_n17663);
nor_4  g15317(new_n17666, new_n17665, new_n17633);
nor_4  g15318(new_n17667, new_n17666, new_n17631);
nor_4  g15319(new_n17668, new_n17667, new_n17630);
nor_4  g15320(new_n17669, new_n17668, new_n17628);
nor_4  g15321(new_n17670, new_n17669, new_n17627);
xnor_3 g15322(new_n17671, new_n17670, new_n17625);
nor_4  g15323(new_n17672, new_n17671, new_n12569_1);
not_3  g15324(new_n17673, new_n17672);
xnor_3 g15325(new_n17674, new_n17670, new_n17624);
nor_4  g15326(new_n17675, new_n17674, new_n12564);
nor_4  g15327(new_n17676, new_n17675, new_n17672);
xnor_3 g15328(new_n17677, new_n17626, new_n13903);
xnor_3 g15329(new_n17678, new_n17668, new_n17677);
nor_4  g15330(new_n17679, new_n17678, new_n12634);
not_3  g15331(new_n17680, new_n17679);
xnor_3 g15332(new_n17681, new_n17668, new_n17628);
nor_4  g15333(new_n17682, new_n17681, new_n12576);
nor_4  g15334(new_n17683, new_n17682, new_n17679);
xnor_3 g15335(new_n17684, new_n17629, new_n13907);
xnor_3 g15336(new_n17685, new_n17666, new_n17684);
nor_4  g15337(new_n17686, new_n17685, new_n12579);
not_3  g15338(new_n17687_1, new_n17686);
xnor_3 g15339(new_n17688, new_n6529, n21957);
xnor_3 g15340(new_n17689, new_n12361, new_n17688);
xnor_3 g15341(new_n17690, new_n17685, new_n17689);
xnor_3 g15342(new_n17691, new_n12359, new_n12330_1);
xnor_3 g15343(new_n17692, new_n17664_1, new_n17663);
not_3  g15344(new_n17693, new_n17692);
nor_4  g15345(new_n17694, new_n17693, new_n17691);
not_3  g15346(new_n17695, new_n17694);
nor_4  g15347(new_n17696, new_n17692, new_n12586);
nor_4  g15348(new_n17697, new_n17696, new_n17694);
not_3  g15349(new_n17698, new_n17637);
nor_4  g15350(new_n17699, new_n17660, new_n17698);
nor_4  g15351(new_n17700, new_n17699, new_n17662);
not_3  g15352(new_n17701, new_n17700);
nand_4 g15353(new_n17702, new_n17701, new_n12590);
xnor_3 g15354(new_n17703, new_n17700, new_n12590);
xnor_3 g15355(new_n17704, new_n17658, new_n17640);
nand_4 g15356(new_n17705, new_n17704, new_n12597);
xnor_3 g15357(new_n17706, new_n17704, new_n12596);
xnor_3 g15358(new_n17707, new_n17656, new_n17643);
nand_4 g15359(new_n17708, new_n17707, new_n12605);
xnor_3 g15360(new_n17709, new_n17707, new_n12601);
not_3  g15361(new_n17710, new_n17654);
xnor_3 g15362(new_n17711, new_n17710, new_n17653);
nor_4  g15363(new_n17712, new_n17711, new_n12611);
not_3  g15364(new_n17713, new_n17712);
not_3  g15365(new_n17714, new_n17711);
nor_4  g15366(new_n17715, new_n17714, new_n12610);
nor_4  g15367(new_n17716, new_n17715, new_n17712);
xnor_3 g15368(new_n17717, new_n17651, new_n17649);
nor_4  g15369(new_n17718, new_n17717, new_n6788);
not_3  g15370(new_n17719, new_n17718);
nand_4 g15371(new_n17720, new_n7731_1, new_n6781);
nand_4 g15372(new_n17721_1, new_n17717, new_n6794_1);
nand_4 g15373(new_n17722, new_n17721_1, new_n17720);
nand_4 g15374(new_n17723, new_n17722, new_n17719);
nand_4 g15375(new_n17724, new_n17723, new_n17716);
nand_4 g15376(new_n17725, new_n17724, new_n17713);
nand_4 g15377(new_n17726, new_n17725, new_n17709);
nand_4 g15378(new_n17727, new_n17726, new_n17708);
nand_4 g15379(new_n17728, new_n17727, new_n17706);
nand_4 g15380(new_n17729, new_n17728, new_n17705);
nand_4 g15381(new_n17730, new_n17729, new_n17703);
nand_4 g15382(new_n17731, new_n17730, new_n17702);
nand_4 g15383(new_n17732, new_n17731, new_n17697);
nand_4 g15384(new_n17733, new_n17732, new_n17695);
nand_4 g15385(new_n17734, new_n17733, new_n17690);
nand_4 g15386(new_n17735_1, new_n17734, new_n17687_1);
nand_4 g15387(new_n17736, new_n17735_1, new_n17683);
nand_4 g15388(new_n17737, new_n17736, new_n17680);
nand_4 g15389(new_n17738_1, new_n17737, new_n17676);
nand_4 g15390(new_n17739, new_n17738_1, new_n17673);
nand_4 g15391(new_n17740, new_n17739, new_n17565);
not_3  g15392(new_n17741, new_n17740);
not_3  g15393(new_n17742, new_n17739);
nand_4 g15394(new_n17743, new_n17742, new_n12559);
not_3  g15395(new_n17744, new_n17743);
nor_4  g15396(new_n17745, new_n17744, new_n17741);
not_3  g15397(new_n17746_1, new_n17623);
nand_4 g15398(new_n17747, new_n17746_1, n4514);
nand_4 g15399(new_n17748, new_n17670, new_n17625);
nand_4 g15400(new_n17749_1, new_n17748, new_n17747);
nor_4  g15401(new_n17750, new_n12399, new_n17620);
not_3  g15402(new_n17751, new_n17750);
nor_4  g15403(new_n17752, new_n12454, n25586);
nor_4  g15404(new_n17753, new_n17752, new_n17619);
nor_4  g15405(new_n17754, new_n17753, new_n12397_1);
nand_4 g15406(new_n17755, new_n17754, new_n17751);
xnor_3 g15407(new_n17756, new_n17755, new_n17749_1);
not_3  g15408(new_n17757, new_n17756);
xnor_3 g15409(n2826, new_n17757, new_n17745);
nor_4  g15410(new_n17759, new_n7307, new_n14816);
xnor_3 g15411(new_n17760, new_n7307, new_n14816);
nor_4  g15412(new_n17761, new_n14927, new_n14820);
not_3  g15413(new_n17762, new_n17761);
nor_4  g15414(new_n17763, new_n7314, n6204);
nor_4  g15415(new_n17764, new_n17763, new_n17761);
nor_4  g15416(new_n17765, new_n14932, new_n14825);
not_3  g15417(new_n17766, new_n17765);
nor_4  g15418(new_n17767, new_n7318, n3349);
nor_4  g15419(new_n17768, new_n17767, new_n17765);
nor_4  g15420(new_n17769, new_n7326, new_n14829);
not_3  g15421(new_n17770, new_n17769);
nor_4  g15422(new_n17771, new_n7374, n1742);
nor_4  g15423(new_n17772, new_n17771, new_n17769);
nor_4  g15424(new_n17773, new_n7330_1, new_n7579);
not_3  g15425(new_n17774, new_n17773);
nor_4  g15426(new_n17775, new_n14941, n8244);
xnor_3 g15427(new_n17776, new_n14941, n8244);
nand_4 g15428(new_n17777, new_n7343, n9493);
xnor_3 g15429(new_n17778, new_n7343, n9493);
not_3  g15430(new_n17779, new_n17778);
nor_4  g15431(new_n17780, new_n7345, n15167);
nor_4  g15432(new_n17781, new_n7351, new_n7602);
not_3  g15433(new_n17782, new_n17781);
nor_4  g15434(new_n17783, new_n7355, new_n14848);
xor_3  g15435(new_n17784_1, new_n7357, n21095);
nand_4 g15436(new_n17785, new_n17784_1, new_n17783);
nand_4 g15437(new_n17786, new_n17785, new_n17782);
xor_3  g15438(new_n17787, new_n7346_1, n15167);
nor_4  g15439(new_n17788, new_n17787, new_n17786);
nor_4  g15440(new_n17789, new_n17788, new_n17780);
nand_4 g15441(new_n17790, new_n17789, new_n17779);
nand_4 g15442(new_n17791, new_n17790, new_n17777);
nor_4  g15443(new_n17792, new_n17791, new_n17776);
nor_4  g15444(new_n17793, new_n17792, new_n17775);
nor_4  g15445(new_n17794, new_n7332, n4858);
nor_4  g15446(new_n17795, new_n17794, new_n17773);
nand_4 g15447(new_n17796, new_n17795, new_n17793);
nand_4 g15448(new_n17797, new_n17796, new_n17774);
nand_4 g15449(new_n17798, new_n17797, new_n17772);
nand_4 g15450(new_n17799, new_n17798, new_n17770);
nand_4 g15451(new_n17800, new_n17799, new_n17768);
nand_4 g15452(new_n17801, new_n17800, new_n17766);
nand_4 g15453(new_n17802, new_n17801, new_n17764);
nand_4 g15454(new_n17803, new_n17802, new_n17762);
not_3  g15455(new_n17804, new_n17803);
nor_4  g15456(new_n17805, new_n17804, new_n17760);
nor_4  g15457(new_n17806, new_n17805, new_n17759);
not_3  g15458(new_n17807, new_n17806);
nand_4 g15459(new_n17808, new_n17807, new_n7248);
nor_4  g15460(new_n17809, new_n2666, new_n2611);
not_3  g15461(new_n17810, new_n17809);
nand_4 g15462(new_n17811, new_n2753, new_n17810);
not_3  g15463(new_n17812, new_n17811);
nor_4  g15464(new_n17813, n20040, n9396);
nor_4  g15465(new_n17814, new_n2665, new_n17813);
not_3  g15466(new_n17815, new_n17814);
nor_4  g15467(new_n17816, new_n17815, new_n17812);
not_3  g15468(new_n17817, new_n17816);
xnor_3 g15469(new_n17818, new_n17817, new_n17808);
xnor_3 g15470(new_n17819, new_n17806, new_n7247);
xnor_3 g15471(new_n17820_1, new_n17814, new_n17811);
not_3  g15472(new_n17821, new_n17820_1);
nand_4 g15473(new_n17822, new_n17821, new_n17819);
xnor_3 g15474(new_n17823, new_n17820_1, new_n17819);
xnor_3 g15475(new_n17824, new_n17804, new_n17760);
nand_4 g15476(new_n17825, new_n17824, new_n2756);
not_3  g15477(new_n17826, new_n2756);
xnor_3 g15478(new_n17827, new_n17824, new_n17826);
xnor_3 g15479(new_n17828, new_n17801, new_n17764);
nand_4 g15480(new_n17829, new_n17828, new_n2912);
xnor_3 g15481(new_n17830, new_n17828, new_n2913);
xnor_3 g15482(new_n17831, new_n17799, new_n17768);
nand_4 g15483(new_n17832, new_n17831, new_n2922);
xnor_3 g15484(new_n17833, new_n17831, new_n2917);
xnor_3 g15485(new_n17834, new_n17797, new_n17772);
nand_4 g15486(new_n17835, new_n17834, new_n2925);
xnor_3 g15487(new_n17836, new_n17834, new_n2924);
xnor_3 g15488(new_n17837, new_n17795, new_n17793);
nand_4 g15489(new_n17838, new_n17837, new_n2930);
xnor_3 g15490(new_n17839, new_n17837, new_n2931);
xnor_3 g15491(new_n17840, new_n17791, new_n17776);
nor_4  g15492(new_n17841, new_n17840, new_n2937);
not_3  g15493(new_n17842, new_n17841);
nor_4  g15494(new_n17843, new_n7335_1, new_n7583);
nor_4  g15495(new_n17844, new_n17843, new_n17775);
xnor_3 g15496(new_n17845, new_n17791, new_n17844);
nor_4  g15497(new_n17846, new_n17845, new_n2936);
nor_4  g15498(new_n17847, new_n17846, new_n17841);
not_3  g15499(new_n17848, new_n2944_1);
xnor_3 g15500(new_n17849, new_n17789, new_n17779);
nand_4 g15501(new_n17850, new_n17849, new_n17848);
not_3  g15502(new_n17851, new_n17850);
nor_4  g15503(new_n17852, new_n17849, new_n17848);
nor_4  g15504(new_n17853, new_n17852, new_n17851);
not_3  g15505(new_n17854, new_n17786);
xnor_3 g15506(new_n17855_1, new_n17787, new_n17854);
nand_4 g15507(new_n17856, new_n17855_1, new_n2951);
not_3  g15508(new_n17857, new_n17856);
nor_4  g15509(new_n17858, new_n17855_1, new_n2951);
nor_4  g15510(new_n17859, new_n17858, new_n17857);
xnor_3 g15511(new_n17860, new_n17784_1, new_n17783);
nand_4 g15512(new_n17861, new_n17860, new_n2959);
not_3  g15513(new_n17862, new_n2962);
xor_3  g15514(new_n17863, new_n7355, new_n14848);
nor_4  g15515(new_n17864, new_n17863, new_n17862);
not_3  g15516(new_n17865, new_n17861);
nor_4  g15517(new_n17866, new_n17860, new_n2959);
nor_4  g15518(new_n17867, new_n17866, new_n17865);
nand_4 g15519(new_n17868, new_n17867, new_n17864);
nand_4 g15520(new_n17869, new_n17868, new_n17861);
nand_4 g15521(new_n17870, new_n17869, new_n17859);
nand_4 g15522(new_n17871, new_n17870, new_n17856);
nand_4 g15523(new_n17872, new_n17871, new_n17853);
nand_4 g15524(new_n17873, new_n17872, new_n17850);
nand_4 g15525(new_n17874, new_n17873, new_n17847);
nand_4 g15526(new_n17875, new_n17874, new_n17842);
nand_4 g15527(new_n17876, new_n17875, new_n17839);
nand_4 g15528(new_n17877_1, new_n17876, new_n17838);
nand_4 g15529(new_n17878, new_n17877_1, new_n17836);
nand_4 g15530(new_n17879, new_n17878, new_n17835);
nand_4 g15531(new_n17880, new_n17879, new_n17833);
nand_4 g15532(new_n17881, new_n17880, new_n17832);
nand_4 g15533(new_n17882, new_n17881, new_n17830);
nand_4 g15534(new_n17883, new_n17882, new_n17829);
nand_4 g15535(new_n17884, new_n17883, new_n17827);
nand_4 g15536(new_n17885, new_n17884, new_n17825);
nand_4 g15537(new_n17886, new_n17885, new_n17823);
nand_4 g15538(new_n17887, new_n17886, new_n17822);
xnor_3 g15539(n2853, new_n17887, new_n17818);
xor_3  g15540(new_n17889_1, n7099, new_n2993);
not_3  g15541(new_n17890, new_n17889_1);
not_3  g15542(new_n17891, n12811);
nor_4  g15543(new_n17892, new_n17891, n5213);
not_3  g15544(new_n17893, new_n17892);
xor_3  g15545(new_n17894, n12811, new_n2997);
not_3  g15546(new_n17895, new_n17894);
nor_4  g15547(new_n17896, n4665, new_n14280);
xor_3  g15548(new_n17897, n4665, n1118);
nor_4  g15549(new_n17898, n25974, new_n3007);
nor_4  g15550(new_n17899, new_n14285, n19005);
nor_4  g15551(new_n17900, new_n3011, n1630);
nor_4  g15552(new_n17901, n4326, new_n14287);
nor_4  g15553(new_n17902, new_n6772, n1451);
not_3  g15554(new_n17903, new_n17902);
nor_4  g15555(new_n17904, new_n17903, new_n17901);
nor_4  g15556(new_n17905, new_n17904, new_n17900);
nor_4  g15557(new_n17906, new_n17905, new_n17899);
nor_4  g15558(new_n17907, new_n17906, new_n17898);
not_3  g15559(new_n17908, new_n17907);
nor_4  g15560(new_n17909, new_n17908, new_n17897);
nor_4  g15561(new_n17910, new_n17909, new_n17896);
nor_4  g15562(new_n17911_1, new_n17910, new_n17895);
not_3  g15563(new_n17912_1, new_n17911_1);
nand_4 g15564(new_n17913, new_n17912_1, new_n17893);
xor_3  g15565(new_n17914, new_n17913, new_n17890);
nand_4 g15566(new_n17915, new_n4748, new_n4744);
xor_3  g15567(new_n17916, new_n17915, n3570);
nand_4 g15568(new_n17917, new_n17916, n5337);
not_3  g15569(new_n17918, new_n17917);
nor_4  g15570(new_n17919, new_n17916, n5337);
nor_4  g15571(new_n17920, new_n17919, new_n17918);
nand_4 g15572(new_n17921, new_n4749, n626);
nand_4 g15573(new_n17922, new_n4778, new_n4750);
nand_4 g15574(new_n17923, new_n17922, new_n17921);
xnor_3 g15575(new_n17924, new_n17923, new_n17920);
xnor_3 g15576(new_n17925, new_n17924, new_n13319_1);
not_3  g15577(new_n17926, new_n4780);
nand_4 g15578(new_n17927_1, new_n4779, new_n4743);
nand_4 g15579(new_n17928, new_n4817, new_n17927_1);
nand_4 g15580(new_n17929, new_n17928, new_n17926);
xnor_3 g15581(new_n17930, new_n17929, new_n17925);
xnor_3 g15582(new_n17931_1, new_n17930, new_n17914);
xor_3  g15583(new_n17932, new_n17910, new_n17895);
not_3  g15584(new_n17933, new_n17932);
nand_4 g15585(new_n17934, new_n17933, new_n4818);
xor_3  g15586(new_n17935, new_n17908, new_n17897);
not_3  g15587(new_n17936, new_n17935);
nand_4 g15588(new_n17937, new_n17936, new_n4824);
xnor_3 g15589(new_n17938, new_n17935, new_n4824);
xor_3  g15590(new_n17939, n25974, n19005);
xor_3  g15591(new_n17940, new_n17939, new_n17905);
nand_4 g15592(new_n17941, new_n17940, new_n4827);
not_3  g15593(new_n17942, new_n17940);
xnor_3 g15594(new_n17943, new_n17942, new_n4827);
not_3  g15595(new_n17944, n1451);
xor_3  g15596(new_n17945, n5438, new_n17944);
nor_4  g15597(new_n17946, new_n17945, new_n4842);
not_3  g15598(new_n17947, new_n17946);
nor_4  g15599(new_n17948_1, new_n17901, new_n17900);
xor_3  g15600(new_n17949, new_n17948_1, new_n17903);
not_3  g15601(new_n17950, new_n17949);
nor_4  g15602(new_n17951, new_n17950, new_n17947);
xnor_3 g15603(new_n17952, new_n17949, new_n17946);
nor_4  g15604(new_n17953, new_n17952, new_n4832);
nor_4  g15605(new_n17954_1, new_n17953, new_n17951);
nand_4 g15606(new_n17955, new_n17954_1, new_n17943);
nand_4 g15607(new_n17956_1, new_n17955, new_n17941);
nand_4 g15608(new_n17957, new_n17956_1, new_n17938);
nand_4 g15609(new_n17958, new_n17957, new_n17937);
xnor_3 g15610(new_n17959_1, new_n17932, new_n4818);
nand_4 g15611(new_n17960, new_n17959_1, new_n17958);
nand_4 g15612(new_n17961, new_n17960, new_n17934);
xor_3  g15613(n2860, new_n17961, new_n17931_1);
not_3  g15614(new_n17963_1, new_n16786);
xor_3  g15615(n2887, new_n16808, new_n17963_1);
nor_4  g15616(new_n17965, new_n17915, n3570);
nand_4 g15617(new_n17966, new_n17965, new_n7083);
nor_4  g15618(new_n17967, new_n17966, n20359);
not_3  g15619(new_n17968_1, new_n17967);
nor_4  g15620(new_n17969, new_n17968_1, n2816);
xor_3  g15621(new_n17970, new_n17969, new_n7022);
nor_4  g15622(new_n17971, new_n17970, n21784);
xor_3  g15623(new_n17972, new_n17968_1, n2816);
not_3  g15624(new_n17973, new_n17972);
nor_4  g15625(new_n17974, new_n17973, new_n14323_1);
nor_4  g15626(new_n17975, new_n17972, n5521);
xor_3  g15627(new_n17976_1, new_n17966, n20359);
nor_4  g15628(new_n17977, new_n17976_1, n11926);
not_3  g15629(new_n17978, new_n17977);
not_3  g15630(new_n17979, new_n17976_1);
xor_3  g15631(new_n17980, new_n17979, new_n14330);
xor_3  g15632(new_n17981, new_n17965, new_n7083);
not_3  g15633(new_n17982, new_n17981);
nor_4  g15634(new_n17983, new_n17982, new_n4219);
nor_4  g15635(new_n17984, new_n17981, n4325);
not_3  g15636(new_n17985, new_n17984);
not_3  g15637(new_n17986, new_n17919);
nand_4 g15638(new_n17987, new_n17923, new_n17986);
nand_4 g15639(new_n17988, new_n17987, new_n17917);
nand_4 g15640(new_n17989, new_n17988, new_n17985);
not_3  g15641(new_n17990, new_n17989);
nor_4  g15642(new_n17991, new_n17990, new_n17983);
nand_4 g15643(new_n17992, new_n17991, new_n17980);
nand_4 g15644(new_n17993, new_n17992, new_n17978);
nor_4  g15645(new_n17994, new_n17993, new_n17975);
nor_4  g15646(new_n17995, new_n17994, new_n17974);
nor_4  g15647(new_n17996, new_n17995, new_n17971);
not_3  g15648(new_n17997, new_n17969);
nor_4  g15649(new_n17998_1, new_n17997, n8526);
not_3  g15650(new_n17999, new_n17970);
nor_4  g15651(new_n18000, new_n17999, new_n14313);
nor_4  g15652(new_n18001, new_n18000, new_n17998_1);
not_3  g15653(new_n18002, new_n18001);
nor_4  g15654(new_n18003, new_n18002, new_n17996);
xnor_3 g15655(new_n18004, new_n18003, new_n13288);
nor_4  g15656(new_n18005, new_n18000, new_n17971);
not_3  g15657(new_n18006, new_n18005);
xnor_3 g15658(new_n18007, new_n18006, new_n17995);
nor_4  g15659(new_n18008, new_n18007, new_n13295);
xnor_3 g15660(new_n18009, new_n18005, new_n17995);
xnor_3 g15661(new_n18010, new_n18009, new_n13292);
nor_4  g15662(new_n18011, new_n17975, new_n17974);
xnor_3 g15663(new_n18012, new_n18011, new_n17993);
nor_4  g15664(new_n18013, new_n18012, new_n13299);
not_3  g15665(new_n18014, new_n18013);
not_3  g15666(new_n18015, new_n17980);
not_3  g15667(new_n18016, new_n17983);
nand_4 g15668(new_n18017, new_n17989, new_n18016);
nor_4  g15669(new_n18018, new_n18017, new_n18015);
nor_4  g15670(new_n18019, new_n18018, new_n17977);
xnor_3 g15671(new_n18020, new_n18011, new_n18019);
nor_4  g15672(new_n18021, new_n18020, new_n13300);
nor_4  g15673(new_n18022, new_n18021, new_n18013);
nor_4  g15674(new_n18023, new_n17991, new_n17980);
nor_4  g15675(new_n18024, new_n18023, new_n18018);
nand_4 g15676(new_n18025_1, new_n18024, new_n13307);
nor_4  g15677(new_n18026, new_n17984, new_n17983);
xnor_3 g15678(new_n18027, new_n18026, new_n17988);
nor_4  g15679(new_n18028, new_n18027, new_n13313);
xnor_3 g15680(new_n18029, new_n18027, new_n13313);
nor_4  g15681(new_n18030, new_n17924, new_n13322);
nand_4 g15682(new_n18031, new_n17929, new_n17925);
not_3  g15683(new_n18032, new_n18031);
nor_4  g15684(new_n18033, new_n18032, new_n18030);
nor_4  g15685(new_n18034, new_n18033, new_n18029);
nor_4  g15686(new_n18035_1, new_n18034, new_n18028);
xnor_3 g15687(new_n18036, new_n17991, new_n17980);
xnor_3 g15688(new_n18037, new_n18036, new_n13307);
nand_4 g15689(new_n18038, new_n18037, new_n18035_1);
nand_4 g15690(new_n18039, new_n18038, new_n18025_1);
nand_4 g15691(new_n18040, new_n18039, new_n18022);
nand_4 g15692(new_n18041, new_n18040, new_n18014);
nor_4  g15693(new_n18042, new_n18041, new_n18010);
nor_4  g15694(new_n18043_1, new_n18042, new_n18008);
xnor_3 g15695(new_n18044, new_n18043_1, new_n18004);
nand_4 g15696(new_n18045_1, new_n4672, new_n4668);
nor_4  g15697(new_n18046, new_n18045_1, n26452);
nand_4 g15698(new_n18047, new_n18046, new_n12692);
nor_4  g15699(new_n18048, new_n18047, n5077);
not_3  g15700(new_n18049, new_n18048);
nor_4  g15701(new_n18050, new_n18049, n18035);
not_3  g15702(new_n18051, new_n18050);
nor_4  g15703(new_n18052, new_n18051, n8827);
xor_3  g15704(new_n18053, new_n18050, new_n15557);
nor_4  g15705(new_n18054, new_n18053, n11898);
xor_3  g15706(new_n18055, new_n18048, new_n15538);
nor_4  g15707(new_n18056, new_n18055, n19941);
not_3  g15708(new_n18057, new_n18055);
xor_3  g15709(new_n18058, new_n18057, n19941);
xor_3  g15710(new_n18059_1, new_n18047, n5077);
nor_4  g15711(new_n18060, new_n18059_1, n1099);
not_3  g15712(new_n18061_1, new_n18059_1);
xor_3  g15713(new_n18062, new_n18061_1, n1099);
xor_3  g15714(new_n18063, new_n18046, new_n12692);
nor_4  g15715(new_n18064, new_n18063, n2113);
not_3  g15716(new_n18065, n21134);
not_3  g15717(new_n18066, n26452);
xor_3  g15718(new_n18067, new_n18045_1, new_n18066);
nand_4 g15719(new_n18068, new_n18067, new_n18065);
not_3  g15720(new_n18069, new_n18045_1);
xor_3  g15721(new_n18070, new_n18069, new_n18066);
xnor_3 g15722(new_n18071_1, new_n18070, new_n18065);
xor_3  g15723(new_n18072, new_n4672, n19905);
nand_4 g15724(new_n18073, new_n18072, new_n4075);
nand_4 g15725(new_n18074, new_n4698, new_n4674_1);
nand_4 g15726(new_n18075, new_n18074, new_n18073);
nand_4 g15727(new_n18076, new_n18075, new_n18071_1);
nand_4 g15728(new_n18077, new_n18076, new_n18068);
xnor_3 g15729(new_n18078, new_n18063, new_n4074);
nand_4 g15730(new_n18079, new_n18078, new_n18077);
not_3  g15731(new_n18080, new_n18079);
nor_4  g15732(new_n18081, new_n18080, new_n18064);
nor_4  g15733(new_n18082, new_n18081, new_n18062);
nor_4  g15734(new_n18083, new_n18082, new_n18060);
nor_4  g15735(new_n18084, new_n18083, new_n18058);
nor_4  g15736(new_n18085, new_n18084, new_n18056);
not_3  g15737(new_n18086, new_n18053);
nor_4  g15738(new_n18087, new_n18086, new_n17164);
nor_4  g15739(new_n18088, new_n18087, new_n18085);
nor_4  g15740(new_n18089, new_n18088, new_n18054);
nor_4  g15741(new_n18090, new_n18089, new_n18052);
xnor_3 g15742(new_n18091, new_n18090, new_n18044);
not_3  g15743(new_n18092, new_n18010);
xnor_3 g15744(new_n18093, new_n18041, new_n18092);
nor_4  g15745(new_n18094, new_n18087, new_n18054);
xor_3  g15746(new_n18095, new_n18094, new_n18085);
nor_4  g15747(new_n18096, new_n18095, new_n18093);
not_3  g15748(new_n18097, new_n18096);
xnor_3 g15749(new_n18098, new_n18041, new_n18010);
not_3  g15750(new_n18099, new_n18095);
nor_4  g15751(new_n18100, new_n18099, new_n18098);
nor_4  g15752(new_n18101, new_n18100, new_n18096);
xor_3  g15753(new_n18102, new_n18083, new_n18058);
xnor_3 g15754(new_n18103, new_n18039, new_n18022);
not_3  g15755(new_n18104, new_n18103);
nand_4 g15756(new_n18105_1, new_n18104, new_n18102);
xnor_3 g15757(new_n18106, new_n18103, new_n18102);
xor_3  g15758(new_n18107, new_n18081, new_n18062);
not_3  g15759(new_n18108, new_n18107);
xnor_3 g15760(new_n18109, new_n18037, new_n18035_1);
nor_4  g15761(new_n18110, new_n18109, new_n18108);
not_3  g15762(new_n18111, new_n18110);
not_3  g15763(new_n18112, new_n18037);
xnor_3 g15764(new_n18113, new_n18112, new_n18035_1);
nor_4  g15765(new_n18114, new_n18113, new_n18107);
nor_4  g15766(new_n18115, new_n18114, new_n18110);
nor_4  g15767(new_n18116, new_n18026, new_n17988);
nand_4 g15768(new_n18117, new_n18026, new_n17988);
not_3  g15769(new_n18118, new_n18117);
nor_4  g15770(new_n18119, new_n18118, new_n18116);
nor_4  g15771(new_n18120, new_n18119, new_n13312);
nor_4  g15772(new_n18121, new_n18120, new_n18028);
xnor_3 g15773(new_n18122, new_n18033, new_n18121);
xnor_3 g15774(new_n18123, new_n18078, new_n18077);
nor_4  g15775(new_n18124, new_n18123, new_n18122);
not_3  g15776(new_n18125, new_n18124);
xnor_3 g15777(new_n18126, new_n18033, new_n18029);
not_3  g15778(new_n18127, new_n18123);
nor_4  g15779(new_n18128, new_n18127, new_n18126);
nor_4  g15780(new_n18129, new_n18128, new_n18124);
not_3  g15781(new_n18130, new_n18071_1);
xnor_3 g15782(new_n18131, new_n18075, new_n18130);
nand_4 g15783(new_n18132, new_n18131, new_n17930);
not_3  g15784(new_n18133, new_n18132);
nor_4  g15785(new_n18134, new_n18131, new_n17930);
nor_4  g15786(new_n18135, new_n18134, new_n18133);
nand_4 g15787(new_n18136, new_n4850_1, new_n4822);
nand_4 g15788(new_n18137, new_n18136, new_n4820);
nand_4 g15789(new_n18138, new_n18137, new_n18135);
nand_4 g15790(new_n18139, new_n18138, new_n18132);
nand_4 g15791(new_n18140, new_n18139, new_n18129);
nand_4 g15792(new_n18141, new_n18140, new_n18125);
nand_4 g15793(new_n18142, new_n18141, new_n18115);
nand_4 g15794(new_n18143_1, new_n18142, new_n18111);
nand_4 g15795(new_n18144, new_n18143_1, new_n18106);
nand_4 g15796(new_n18145_1, new_n18144, new_n18105_1);
nand_4 g15797(new_n18146, new_n18145_1, new_n18101);
nand_4 g15798(new_n18147, new_n18146, new_n18097);
nor_4  g15799(new_n18148, new_n18147, new_n18091);
nand_4 g15800(new_n18149, new_n18043_1, new_n18004);
not_3  g15801(new_n18150, new_n18149);
nor_4  g15802(new_n18151_1, new_n18043_1, new_n18004);
nor_4  g15803(new_n18152_1, new_n18151_1, new_n18150);
not_3  g15804(new_n18153, new_n18090);
nor_4  g15805(new_n18154, new_n18153, new_n18152_1);
nor_4  g15806(new_n18155, new_n18090, new_n18044);
nor_4  g15807(new_n18156, new_n18155, new_n18154);
xnor_3 g15808(new_n18157_1, new_n18095, new_n18093);
not_3  g15809(new_n18158, new_n18145_1);
nor_4  g15810(new_n18159, new_n18158, new_n18157_1);
nor_4  g15811(new_n18160, new_n18159, new_n18096);
nor_4  g15812(new_n18161, new_n18160, new_n18156);
nor_4  g15813(n2929, new_n18161, new_n18148);
xor_3  g15814(new_n18163, n22793, new_n2983);
nor_4  g15815(new_n18164, n8439, new_n2985_1);
not_3  g15816(new_n18165, new_n18164);
xor_3  g15817(new_n18166, n8439, new_n2985_1);
nor_4  g15818(new_n18167, n25523, new_n2781);
not_3  g15819(new_n18168, new_n18167);
xor_3  g15820(new_n18169, n25523, new_n2781);
not_3  g15821(new_n18170, n12821);
nor_4  g15822(new_n18171_1, new_n18170, n5579);
not_3  g15823(new_n18172, new_n18171_1);
xor_3  g15824(new_n18173, n12821, new_n2759);
nor_4  g15825(new_n18174, n23430, new_n3000);
not_3  g15826(new_n18175, new_n18174);
xor_3  g15827(new_n18176, n23430, new_n3000);
nor_4  g15828(new_n18177, n18558, new_n2860_1);
nor_4  g15829(new_n18178, new_n16438, new_n16429);
nor_4  g15830(new_n18179, new_n18178, new_n18177);
nand_4 g15831(new_n18180, new_n18179, new_n18176);
nand_4 g15832(new_n18181, new_n18180, new_n18175);
nand_4 g15833(new_n18182, new_n18181, new_n18173);
nand_4 g15834(new_n18183, new_n18182, new_n18172);
nand_4 g15835(new_n18184, new_n18183, new_n18169);
nand_4 g15836(new_n18185, new_n18184, new_n18168);
nand_4 g15837(new_n18186, new_n18185, new_n18166);
nand_4 g15838(new_n18187, new_n18186, new_n18165);
xnor_3 g15839(new_n18188, new_n18187, new_n18163);
xnor_3 g15840(new_n18189, new_n18188, new_n8578);
not_3  g15841(new_n18190, new_n18189);
xnor_3 g15842(new_n18191, new_n18185, new_n18166);
not_3  g15843(new_n18192, new_n18191);
nand_4 g15844(new_n18193_1, new_n18192, new_n8588);
xnor_3 g15845(new_n18194, new_n18191, new_n8588);
not_3  g15846(new_n18195, new_n18184);
nor_4  g15847(new_n18196, new_n18183, new_n18169);
nor_4  g15848(new_n18197, new_n18196, new_n18195);
nor_4  g15849(new_n18198, new_n18197, new_n8596);
xnor_3 g15850(new_n18199, new_n18197, new_n8596);
xnor_3 g15851(new_n18200, new_n18181, new_n18173);
not_3  g15852(new_n18201, new_n18200);
nor_4  g15853(new_n18202, new_n18201, new_n8602);
xnor_3 g15854(new_n18203, new_n18200, new_n8600);
not_3  g15855(new_n18204, new_n18180);
not_3  g15856(new_n18205, new_n18176);
not_3  g15857(new_n18206, new_n18177);
not_3  g15858(new_n18207, new_n16429);
not_3  g15859(new_n18208, new_n16438);
nand_4 g15860(new_n18209, new_n18208, new_n18207);
nand_4 g15861(new_n18210, new_n18209, new_n18206);
nand_4 g15862(new_n18211, new_n18210, new_n18205);
not_3  g15863(new_n18212, new_n18211);
nor_4  g15864(new_n18213, new_n18212, new_n18204);
nand_4 g15865(new_n18214, new_n18213, new_n8604);
xnor_3 g15866(new_n18215, new_n18213, new_n8607);
not_3  g15867(new_n18216, new_n16822);
nand_4 g15868(new_n18217, new_n16837_1, new_n16824_1);
nand_4 g15869(new_n18218, new_n18217, new_n18216);
nand_4 g15870(new_n18219, new_n18218, new_n18215);
nand_4 g15871(new_n18220, new_n18219, new_n18214);
nor_4  g15872(new_n18221, new_n18220, new_n18203);
nor_4  g15873(new_n18222, new_n18221, new_n18202);
nor_4  g15874(new_n18223, new_n18222, new_n18199);
nor_4  g15875(new_n18224, new_n18223, new_n18198);
nand_4 g15876(new_n18225, new_n18224, new_n18194);
nand_4 g15877(new_n18226, new_n18225, new_n18193_1);
xnor_3 g15878(new_n18227_1, new_n18226, new_n18190);
xor_3  g15879(new_n18228, n22379, new_n10438);
nor_4  g15880(new_n18229, n3710, new_n2987);
not_3  g15881(new_n18230, new_n18229);
xor_3  g15882(new_n18231, n3710, new_n2987);
nor_4  g15883(new_n18232_1, n26318, new_n2989);
not_3  g15884(new_n18233, new_n18232_1);
xor_3  g15885(new_n18234, n26318, new_n2989);
nor_4  g15886(new_n18235, n26054, new_n2993);
not_3  g15887(new_n18236, new_n18235);
xor_3  g15888(new_n18237, n26054, new_n2993);
nor_4  g15889(new_n18238_1, n19081, new_n2997);
not_3  g15890(new_n18239, new_n18238_1);
nor_4  g15891(new_n18240, new_n10462, n5213);
not_3  g15892(new_n18241_1, new_n18240);
nor_4  g15893(new_n18242, new_n10490, n4665);
not_3  g15894(new_n18243, new_n16852);
nor_4  g15895(new_n18244, new_n18243, new_n16839);
nor_4  g15896(new_n18245, new_n18244, new_n18242);
nand_4 g15897(new_n18246, new_n18245, new_n18241_1);
nand_4 g15898(new_n18247, new_n18246, new_n18239);
nand_4 g15899(new_n18248, new_n18247, new_n18237);
nand_4 g15900(new_n18249, new_n18248, new_n18236);
nand_4 g15901(new_n18250, new_n18249, new_n18234);
nand_4 g15902(new_n18251, new_n18250, new_n18233);
nand_4 g15903(new_n18252, new_n18251, new_n18231);
nand_4 g15904(new_n18253, new_n18252, new_n18230);
not_3  g15905(new_n18254_1, new_n18253);
xor_3  g15906(new_n18255, new_n18254_1, new_n18228);
xnor_3 g15907(new_n18256, new_n18255, new_n18227_1);
xor_3  g15908(new_n18257, new_n18251, new_n18231);
not_3  g15909(new_n18258, new_n18257);
xnor_3 g15910(new_n18259, new_n18224, new_n18194);
nand_4 g15911(new_n18260, new_n18259, new_n18258);
xnor_3 g15912(new_n18261, new_n18259, new_n18257);
xor_3  g15913(new_n18262, new_n18249, new_n18234);
not_3  g15914(new_n18263, new_n18262);
not_3  g15915(new_n18264, new_n18199);
xnor_3 g15916(new_n18265, new_n18222, new_n18264);
nand_4 g15917(new_n18266, new_n18265, new_n18263);
xnor_3 g15918(new_n18267, new_n18265, new_n18262);
xor_3  g15919(new_n18268, new_n18247, new_n18237);
not_3  g15920(new_n18269, new_n18268);
not_3  g15921(new_n18270, new_n18203);
xnor_3 g15922(new_n18271, new_n18220, new_n18270);
nand_4 g15923(new_n18272, new_n18271, new_n18269);
not_3  g15924(new_n18273, new_n18215);
xnor_3 g15925(new_n18274_1, new_n18218, new_n18273);
not_3  g15926(new_n18275, new_n18274_1);
nand_4 g15927(new_n18276, new_n18241_1, new_n18239);
xor_3  g15928(new_n18277, new_n18276, new_n18245);
nand_4 g15929(new_n18278, new_n18277, new_n18275);
xnor_3 g15930(new_n18279, new_n18277, new_n18274_1);
not_3  g15931(new_n18280, new_n16853);
nand_4 g15932(new_n18281, new_n18280, new_n16838);
nand_4 g15933(new_n18282, new_n16877, new_n16854);
nand_4 g15934(new_n18283, new_n18282, new_n18281);
nand_4 g15935(new_n18284, new_n18283, new_n18279);
nand_4 g15936(new_n18285, new_n18284, new_n18278);
xnor_3 g15937(new_n18286, new_n18271, new_n18268);
nand_4 g15938(new_n18287, new_n18286, new_n18285);
nand_4 g15939(new_n18288_1, new_n18287, new_n18272);
nand_4 g15940(new_n18289, new_n18288_1, new_n18267);
nand_4 g15941(new_n18290_1, new_n18289, new_n18266);
nand_4 g15942(new_n18291, new_n18290_1, new_n18261);
nand_4 g15943(new_n18292, new_n18291, new_n18260);
xnor_3 g15944(n2948, new_n18292, new_n18256);
xor_3  g15945(n2961, new_n17551, new_n17524_1);
xnor_3 g15946(n2971, new_n13700, new_n13665);
xor_3  g15947(n3010, new_n2585, new_n2561_1);
xor_3  g15948(n3017, new_n7925, new_n7913);
nor_4  g15949(new_n18298, new_n14172, new_n14165);
xnor_3 g15950(n3020, new_n18298, new_n14169);
not_3  g15951(new_n18300, new_n7187);
xor_3  g15952(n3067, new_n18300, new_n7158);
xor_3  g15953(new_n18302, n23541, n19234);
xor_3  g15954(new_n18303, n27134, n4588);
xnor_3 g15955(new_n18304_1, new_n18303, new_n18302);
xor_3  g15956(n3076, new_n18304_1, new_n11983);
nor_4  g15957(new_n18306, n15490, n18);
nand_4 g15958(new_n18307, new_n18306, new_n10907);
xor_3  g15959(new_n18308, new_n18307, n10611);
not_3  g15960(new_n18309, new_n18308);
nor_4  g15961(new_n18310_1, new_n18309, new_n7733);
nor_4  g15962(new_n18311_1, new_n18308, n7421);
nor_4  g15963(new_n18312, new_n18311_1, new_n18310_1);
xor_3  g15964(new_n18313, new_n18306, n2783);
nor_4  g15965(new_n18314, new_n18313, new_n7751_1);
xnor_3 g15966(new_n18315, new_n18313, new_n7751_1);
xnor_3 g15967(new_n18316, n15490, n18);
not_3  g15968(new_n18317, new_n18316);
nor_4  g15969(new_n18318, new_n18317, n2809);
not_3  g15970(new_n18319, new_n18318);
nand_4 g15971(new_n18320, n15508, n18);
xor_3  g15972(new_n18321, new_n18316, new_n7769_1);
nand_4 g15973(new_n18322, new_n18321, new_n18320);
nand_4 g15974(new_n18323_1, new_n18322, new_n18319);
nor_4  g15975(new_n18324, new_n18323_1, new_n18315);
nor_4  g15976(new_n18325, new_n18324, new_n18314);
xnor_3 g15977(new_n18326, new_n18325, new_n18312);
xnor_3 g15978(new_n18327, new_n18326, new_n12849);
xnor_3 g15979(new_n18328, new_n18323_1, new_n18315);
nor_4  g15980(new_n18329, new_n18328, new_n12854);
xnor_3 g15981(new_n18330, new_n18328, new_n12854);
nor_4  g15982(new_n18331, new_n18321, new_n6763);
not_3  g15983(new_n18332_1, new_n18331);
not_3  g15984(new_n18333, new_n18320);
not_3  g15985(new_n18334, new_n18321);
xor_3  g15986(new_n18335, new_n18334, new_n18333);
not_3  g15987(new_n18336, new_n18335);
nand_4 g15988(new_n18337, new_n18336, new_n6763);
xor_3  g15989(new_n18338, n15508, n18);
nand_4 g15990(new_n18339, new_n18338, new_n6731);
nand_4 g15991(new_n18340, new_n18339, new_n18337);
nand_4 g15992(new_n18341, new_n18340, new_n18332_1);
nor_4  g15993(new_n18342, new_n18341, new_n18330);
nor_4  g15994(new_n18343_1, new_n18342, new_n18329);
xor_3  g15995(n3089, new_n18343_1, new_n18327);
xor_3  g15996(n3125, new_n5986, new_n5984);
xor_3  g15997(new_n18346, n21839, n19282);
nor_4  g15998(new_n18347, n27089, n12657);
nor_4  g15999(new_n18348, new_n3118, new_n3076_1);
nor_4  g16000(new_n18349, new_n18348, new_n18347);
xnor_3 g16001(new_n18350_1, new_n18349, new_n18346);
nor_4  g16002(new_n18351, new_n18350_1, new_n13251);
not_3  g16003(new_n18352, new_n18346);
xnor_3 g16004(new_n18353, new_n18349, new_n18352);
nor_4  g16005(new_n18354, new_n18353, new_n13283);
nor_4  g16006(new_n18355, new_n18354, new_n18351);
not_3  g16007(new_n18356, new_n18355);
xnor_3 g16008(new_n18357, new_n3118, new_n3075);
nor_4  g16009(new_n18358, new_n13255, new_n18357);
nor_4  g16010(new_n18359, new_n13259, new_n3125_1);
nor_4  g16011(new_n18360, new_n13260, new_n3123);
nor_4  g16012(new_n18361, new_n18360, new_n18359);
nor_4  g16013(new_n18362_1, new_n13264, new_n3129);
not_3  g16014(new_n18363, new_n3110);
nor_4  g16015(new_n18364, new_n18363, new_n3087);
nor_4  g16016(new_n18365, new_n18364, new_n16139);
nor_4  g16017(new_n18366, new_n18365, new_n3084);
xnor_3 g16018(new_n18367, new_n18366, new_n3083);
nor_4  g16019(new_n18368, new_n13263_1, new_n18367);
nor_4  g16020(new_n18369, new_n18368, new_n18362_1);
not_3  g16021(new_n18370, new_n18369);
nor_4  g16022(new_n18371, new_n16170, new_n16143);
nor_4  g16023(new_n18372, new_n18371, new_n16138);
nor_4  g16024(new_n18373, new_n18372, new_n18370);
nor_4  g16025(new_n18374, new_n18373, new_n18362_1);
nand_4 g16026(new_n18375, new_n18374, new_n18361);
not_3  g16027(new_n18376, new_n18375);
nor_4  g16028(new_n18377_1, new_n18376, new_n18359);
nor_4  g16029(new_n18378, new_n13256, new_n3119);
nor_4  g16030(new_n18379, new_n18378, new_n18358);
not_3  g16031(new_n18380, new_n18379);
nor_4  g16032(new_n18381, new_n18380, new_n18377_1);
nor_4  g16033(new_n18382, new_n18381, new_n18358);
nor_4  g16034(new_n18383, new_n18382, new_n18356);
nor_4  g16035(new_n18384, new_n18383, new_n18351);
not_3  g16036(new_n18385, new_n18384);
nor_4  g16037(new_n18386, n21839, n19282);
nor_4  g16038(new_n18387, new_n18349, new_n18352);
nor_4  g16039(new_n18388, new_n18387, new_n18386);
not_3  g16040(new_n18389, new_n18388);
nand_4 g16041(new_n18390, new_n18389, new_n13248);
nor_4  g16042(new_n18391, new_n18390, new_n18385);
nand_4 g16043(new_n18392, new_n18388, new_n13249);
nor_4  g16044(new_n18393, new_n18392, new_n18384);
nor_4  g16045(new_n18394, new_n18393, new_n18391);
xnor_3 g16046(new_n18395, new_n18394, new_n13774);
nand_4 g16047(new_n18396, new_n18392, new_n18390);
xnor_3 g16048(new_n18397, new_n18396, new_n18385);
nor_4  g16049(new_n18398, new_n18397, new_n13775_1);
xnor_3 g16050(new_n18399, new_n18397, new_n13775_1);
not_3  g16051(new_n18400, new_n18382);
nor_4  g16052(new_n18401, new_n18400, new_n18355);
nor_4  g16053(new_n18402, new_n18401, new_n18383);
nand_4 g16054(new_n18403, new_n18402, new_n13793);
xnor_3 g16055(new_n18404, new_n18402, new_n13794);
xnor_3 g16056(new_n18405_1, new_n18380, new_n18377_1);
not_3  g16057(new_n18406, new_n18405_1);
nand_4 g16058(new_n18407, new_n18406, new_n13802);
nor_4  g16059(new_n18408, new_n18405_1, new_n13803);
nor_4  g16060(new_n18409_1, new_n18406, new_n13802);
nor_4  g16061(new_n18410, new_n18409_1, new_n18408);
nor_4  g16062(new_n18411, new_n18374, new_n18361);
nor_4  g16063(new_n18412, new_n18411, new_n18376);
nand_4 g16064(new_n18413, new_n18412, new_n13816);
xnor_3 g16065(new_n18414_1, new_n18412, new_n13811);
xnor_3 g16066(new_n18415, new_n18372, new_n18370);
nand_4 g16067(new_n18416, new_n18415, new_n13836);
xnor_3 g16068(new_n18417, new_n18415, new_n13820);
nand_4 g16069(new_n18418_1, new_n16171, new_n13828);
nand_4 g16070(new_n18419, new_n16208, new_n16172);
nand_4 g16071(new_n18420, new_n18419, new_n18418_1);
nand_4 g16072(new_n18421, new_n18420, new_n18417);
nand_4 g16073(new_n18422, new_n18421, new_n18416);
nand_4 g16074(new_n18423, new_n18422, new_n18414_1);
nand_4 g16075(new_n18424, new_n18423, new_n18413);
nand_4 g16076(new_n18425, new_n18424, new_n18410);
nand_4 g16077(new_n18426, new_n18425, new_n18407);
nand_4 g16078(new_n18427, new_n18426, new_n18404);
nand_4 g16079(new_n18428, new_n18427, new_n18403);
not_3  g16080(new_n18429, new_n18428);
nor_4  g16081(new_n18430, new_n18429, new_n18399);
nor_4  g16082(new_n18431, new_n18430, new_n18398);
xnor_3 g16083(n3126, new_n18431, new_n18395);
xnor_3 g16084(n3208, new_n14534, new_n14483);
not_3  g16085(new_n18434, new_n17310);
xor_3  g16086(n3219, new_n17313, new_n18434);
not_3  g16087(new_n18436, new_n17869);
xor_3  g16088(n3235, new_n18436, new_n17859);
xnor_3 g16089(n3244, new_n13524, new_n13507);
nand_4 g16090(new_n18439_1, n15146, new_n11882);
nand_4 g16091(new_n18440, n11579, new_n11884);
not_3  g16092(new_n18441, new_n11912);
nor_4  g16093(new_n18442, n23513, new_n11887);
not_3  g16094(new_n18443, new_n18442);
nor_4  g16095(new_n18444_1, new_n16459, new_n11966);
nor_4  g16096(new_n18445_1, new_n18444_1, new_n11967);
nand_4 g16097(new_n18446, new_n18445_1, new_n11961);
nor_4  g16098(new_n18447, n6427, new_n11891);
not_3  g16099(new_n18448, new_n18447);
nand_4 g16100(new_n18449, new_n18448, new_n18446);
nand_4 g16101(new_n18450, new_n18449, new_n11957);
nand_4 g16102(new_n18451, new_n18450, new_n18443);
nand_4 g16103(new_n18452_1, new_n18451, new_n18441);
nand_4 g16104(new_n18453, new_n18452_1, new_n18440);
nand_4 g16105(new_n18454, new_n18453, new_n11915);
nand_4 g16106(new_n18455, new_n18454, new_n18439_1);
xnor_3 g16107(new_n18456, new_n18455, new_n11921);
not_3  g16108(new_n18457, new_n18456);
xnor_3 g16109(new_n18458, new_n18457, new_n18191);
not_3  g16110(new_n18459, new_n18197);
xnor_3 g16111(new_n18460, new_n18453, new_n11915);
nand_4 g16112(new_n18461, new_n18460, new_n18459);
xnor_3 g16113(new_n18462, new_n18460, new_n18197);
xnor_3 g16114(new_n18463, new_n18451, new_n18441);
not_3  g16115(new_n18464, new_n18463);
nor_4  g16116(new_n18465, new_n18464, new_n18201);
not_3  g16117(new_n18466, new_n18465);
nor_4  g16118(new_n18467_1, new_n18463, new_n18200);
nor_4  g16119(new_n18468, new_n18467_1, new_n18465);
not_3  g16120(new_n18469, new_n18450);
nor_4  g16121(new_n18470, new_n18449, new_n11957);
nor_4  g16122(new_n18471, new_n18470, new_n18469);
nor_4  g16123(new_n18472, new_n18471, new_n18213);
not_3  g16124(new_n18473, new_n18472);
not_3  g16125(new_n18474, new_n18213);
not_3  g16126(new_n18475, new_n18471);
nor_4  g16127(new_n18476, new_n18475, new_n18474);
nor_4  g16128(new_n18477, new_n18476, new_n18472);
not_3  g16129(new_n18478, new_n16454);
nor_4  g16130(new_n18479, new_n16507_1, new_n16503);
nor_4  g16131(new_n18480, new_n18479, new_n16463);
nor_4  g16132(new_n18481, new_n18480, new_n18478);
nor_4  g16133(new_n18482_1, new_n18481, new_n16451);
nand_4 g16134(new_n18483_1, new_n18482_1, new_n18477);
nand_4 g16135(new_n18484, new_n18483_1, new_n18473);
nand_4 g16136(new_n18485, new_n18484, new_n18468);
nand_4 g16137(new_n18486, new_n18485, new_n18466);
nand_4 g16138(new_n18487, new_n18486, new_n18462);
nand_4 g16139(new_n18488, new_n18487, new_n18461);
xnor_3 g16140(new_n18489, new_n18488, new_n18458);
not_3  g16141(new_n18490, n26483);
nor_4  g16142(new_n18491, n23541, n16247);
nand_4 g16143(new_n18492, new_n18491, new_n2709);
nor_4  g16144(new_n18493, new_n18492, n15979);
nand_4 g16145(new_n18494, new_n18493, new_n18490);
nor_4  g16146(new_n18495, new_n18494, n24768);
nand_4 g16147(new_n18496_1, new_n18495, new_n2685);
xor_3  g16148(new_n18497, new_n18496_1, n19270);
not_3  g16149(new_n18498, new_n18497);
xor_3  g16150(new_n18499, new_n18498, new_n10381);
xor_3  g16151(new_n18500, new_n18495, new_n2685);
nor_4  g16152(new_n18501, new_n18500, n13190);
not_3  g16153(new_n18502, new_n18500);
xor_3  g16154(new_n18503, new_n18502, n13190);
nand_4 g16155(new_n18504, new_n18494, n24768);
not_3  g16156(new_n18505, new_n18504);
nor_4  g16157(new_n18506, new_n18505, new_n18495);
nor_4  g16158(new_n18507, new_n18506, n3460);
not_3  g16159(new_n18508, new_n18506);
nor_4  g16160(new_n18509_1, new_n18508, new_n10386);
nor_4  g16161(new_n18510, new_n18509_1, new_n18507);
not_3  g16162(new_n18511, new_n18510);
xnor_3 g16163(new_n18512, new_n18493, n26483);
nor_4  g16164(new_n18513_1, new_n18512, n5226);
not_3  g16165(new_n18514, new_n18512);
nor_4  g16166(new_n18515_1, new_n18514, new_n10391);
nor_4  g16167(new_n18516, new_n18515_1, new_n18513_1);
nand_4 g16168(new_n18517, new_n18492, n15979);
not_3  g16169(new_n18518, new_n18517);
nor_4  g16170(new_n18519, new_n18518, new_n18493);
nor_4  g16171(new_n18520, new_n18519, n17664);
not_3  g16172(new_n18521, new_n18520);
xnor_3 g16173(new_n18522, new_n18491, n8638);
nor_4  g16174(new_n18523, new_n18522, n23369);
not_3  g16175(new_n18524, new_n18523);
not_3  g16176(new_n18525, new_n18522);
nor_4  g16177(new_n18526, new_n18525, new_n10396);
nor_4  g16178(new_n18527, new_n18526, new_n18523);
xnor_3 g16179(new_n18528, n23541, n16247);
nand_4 g16180(new_n18529, new_n18528, new_n10399);
nand_4 g16181(new_n18530, n23541, n19234);
xnor_3 g16182(new_n18531, new_n18528, n1136);
nand_4 g16183(new_n18532, new_n18531, new_n18530);
nand_4 g16184(new_n18533, new_n18532, new_n18529);
nand_4 g16185(new_n18534, new_n18533, new_n18527);
nand_4 g16186(new_n18535, new_n18534, new_n18524);
not_3  g16187(new_n18536, new_n18519);
nor_4  g16188(new_n18537_1, new_n18536, new_n11449);
nor_4  g16189(new_n18538, new_n18537_1, new_n18520);
nand_4 g16190(new_n18539, new_n18538, new_n18535);
nand_4 g16191(new_n18540, new_n18539, new_n18521);
nand_4 g16192(new_n18541, new_n18540, new_n18516);
not_3  g16193(new_n18542, new_n18541);
nor_4  g16194(new_n18543, new_n18542, new_n18513_1);
nor_4  g16195(new_n18544, new_n18543, new_n18511);
nor_4  g16196(new_n18545, new_n18544, new_n18507);
nor_4  g16197(new_n18546, new_n18545, new_n18503);
nor_4  g16198(new_n18547, new_n18546, new_n18501);
xnor_3 g16199(new_n18548, new_n18547, new_n18499);
nor_4  g16200(new_n18549, new_n18548, new_n18489);
not_3  g16201(new_n18550, new_n18458);
xnor_3 g16202(new_n18551, new_n18488, new_n18550);
not_3  g16203(new_n18552, new_n18548);
nor_4  g16204(new_n18553, new_n18552, new_n18551);
nor_4  g16205(new_n18554, new_n18553, new_n18549);
xnor_3 g16206(new_n18555, new_n18545, new_n18503);
xnor_3 g16207(new_n18556, new_n18486, new_n18462);
nor_4  g16208(new_n18557, new_n18556, new_n18555);
not_3  g16209(new_n18558_1, new_n18557);
xnor_3 g16210(new_n18559, new_n18543, new_n18511);
xnor_3 g16211(new_n18560, new_n18484, new_n18468);
nor_4  g16212(new_n18561, new_n18560, new_n18559);
not_3  g16213(new_n18562, new_n18561);
not_3  g16214(new_n18563, new_n18559);
not_3  g16215(new_n18564, new_n18468);
xnor_3 g16216(new_n18565, new_n18484, new_n18564);
nor_4  g16217(new_n18566, new_n18565, new_n18563);
nor_4  g16218(new_n18567, new_n18566, new_n18561);
xnor_3 g16219(new_n18568, new_n18540, new_n18516);
not_3  g16220(new_n18569, new_n18568);
not_3  g16221(new_n18570, new_n18477);
xnor_3 g16222(new_n18571, new_n18482_1, new_n18570);
nand_4 g16223(new_n18572_1, new_n18571, new_n18569);
xnor_3 g16224(new_n18573, new_n18538, new_n18535);
not_3  g16225(new_n18574_1, new_n18573);
nand_4 g16226(new_n18575, new_n18574_1, new_n16486);
xnor_3 g16227(new_n18576_1, new_n18573, new_n16486);
xnor_3 g16228(new_n18577, new_n18533, new_n18527);
not_3  g16229(new_n18578_1, new_n18577);
nor_4  g16230(new_n18579, new_n18578_1, new_n16508);
xnor_3 g16231(new_n18580, new_n18578_1, new_n16508);
xnor_3 g16232(new_n18581, new_n18531, new_n18530);
not_3  g16233(new_n18582_1, new_n18581);
nand_4 g16234(new_n18583_1, new_n18582_1, new_n16524_1);
xor_3  g16235(new_n18584_1, n23541, new_n11458);
nor_4  g16236(new_n18585, new_n18584_1, new_n16515);
not_3  g16237(new_n18586, new_n18585);
not_3  g16238(new_n18587, new_n18583_1);
nor_4  g16239(new_n18588, new_n18582_1, new_n16524_1);
nor_4  g16240(new_n18589, new_n18588, new_n18587);
nand_4 g16241(new_n18590, new_n18589, new_n18586);
nand_4 g16242(new_n18591, new_n18590, new_n18583_1);
nor_4  g16243(new_n18592, new_n18591, new_n18580);
nor_4  g16244(new_n18593, new_n18592, new_n18579);
nand_4 g16245(new_n18594, new_n18593, new_n18576_1);
nand_4 g16246(new_n18595, new_n18594, new_n18575);
xnor_3 g16247(new_n18596, new_n18571, new_n18568);
nand_4 g16248(new_n18597, new_n18596, new_n18595);
nand_4 g16249(new_n18598, new_n18597, new_n18572_1);
nand_4 g16250(new_n18599, new_n18598, new_n18567);
nand_4 g16251(new_n18600, new_n18599, new_n18562);
not_3  g16252(new_n18601, new_n18555);
not_3  g16253(new_n18602, new_n18462);
xnor_3 g16254(new_n18603, new_n18486, new_n18602);
nor_4  g16255(new_n18604, new_n18603, new_n18601);
nor_4  g16256(new_n18605, new_n18604, new_n18557);
nand_4 g16257(new_n18606, new_n18605, new_n18600);
nand_4 g16258(new_n18607, new_n18606, new_n18558_1);
xnor_3 g16259(n3263, new_n18607, new_n18554);
not_3  g16260(new_n18609, new_n14777);
xor_3  g16261(n3289, new_n14796, new_n18609);
xor_3  g16262(new_n18611, n21832, n5211);
nand_4 g16263(new_n18612, n26913, n12956);
not_3  g16264(new_n18613, new_n18612);
nor_4  g16265(new_n18614, n26913, n12956);
nor_4  g16266(new_n18615, new_n5771, new_n5758);
not_3  g16267(new_n18616, new_n18615);
nor_4  g16268(new_n18617, new_n18616, new_n18614);
nor_4  g16269(new_n18618, new_n18617, new_n18613);
nor_4  g16270(new_n18619, new_n18618, new_n18611);
not_3  g16271(new_n18620, new_n18611);
not_3  g16272(new_n18621, new_n18618);
nor_4  g16273(new_n18622, new_n18621, new_n18620);
nor_4  g16274(new_n18623, new_n18622, new_n18619);
not_3  g16275(new_n18624, new_n18623);
nor_4  g16276(new_n18625, new_n18624, new_n10143);
nor_4  g16277(new_n18626, new_n18623, n18537);
nor_4  g16278(new_n18627, new_n18626, new_n18625);
nor_4  g16279(new_n18628, new_n18614, new_n18613);
xnor_3 g16280(new_n18629, new_n18628, new_n18616);
nand_4 g16281(new_n18630, new_n18629, new_n10148);
not_3  g16282(new_n18631, new_n18629);
nor_4  g16283(new_n18632, new_n18631, n7057);
nor_4  g16284(new_n18633, new_n18629, new_n10148);
nor_4  g16285(new_n18634, new_n18633, new_n18632);
nand_4 g16286(new_n18635_1, new_n5791, new_n5777);
nand_4 g16287(new_n18636, new_n18635_1, new_n5774);
nand_4 g16288(new_n18637, new_n18636, new_n18634);
nand_4 g16289(new_n18638, new_n18637, new_n18630);
xnor_3 g16290(new_n18639, new_n18638, new_n18627);
nor_4  g16291(new_n18640, new_n17406, n21649);
nor_4  g16292(new_n18641, new_n17408, new_n5941);
nor_4  g16293(new_n18642, new_n18641, new_n18640);
nor_4  g16294(new_n18643, new_n11348_1, n18274);
not_3  g16295(new_n18644, new_n18643);
nor_4  g16296(new_n18645, new_n11318, new_n5945);
nor_4  g16297(new_n18646, new_n18645, new_n18643);
nor_4  g16298(new_n18647, new_n11357, n3828);
not_3  g16299(new_n18648, new_n18647);
nand_4 g16300(new_n18649_1, new_n11360, new_n5795);
nand_4 g16301(new_n18650, new_n11363, n21654);
not_3  g16302(new_n18651, new_n18649_1);
nor_4  g16303(new_n18652, new_n11360, new_n5795);
nor_4  g16304(new_n18653_1, new_n18652, new_n18651);
nand_4 g16305(new_n18654, new_n18653_1, new_n18650);
nand_4 g16306(new_n18655, new_n18654, new_n18649_1);
nor_4  g16307(new_n18656, new_n11353, new_n5818);
nor_4  g16308(new_n18657, new_n18656, new_n18647);
nand_4 g16309(new_n18658, new_n18657, new_n18655);
nand_4 g16310(new_n18659, new_n18658, new_n18648);
nand_4 g16311(new_n18660, new_n18659, new_n18646);
nand_4 g16312(new_n18661, new_n18660, new_n18644);
xnor_3 g16313(new_n18662, new_n18661, new_n18642);
nor_4  g16314(new_n18663, new_n18662, new_n18639);
not_3  g16315(new_n18664, new_n18639);
not_3  g16316(new_n18665, new_n18662);
nor_4  g16317(new_n18666, new_n18665, new_n18664);
nor_4  g16318(new_n18667, new_n18666, new_n18663);
not_3  g16319(new_n18668, new_n18667);
xnor_3 g16320(new_n18669, new_n18636, new_n18634);
xnor_3 g16321(new_n18670, new_n18659, new_n18646);
nor_4  g16322(new_n18671, new_n18670, new_n18669);
not_3  g16323(new_n18672, new_n18671);
not_3  g16324(new_n18673, new_n18669);
not_3  g16325(new_n18674, new_n18670);
nor_4  g16326(new_n18675, new_n18674, new_n18673);
nor_4  g16327(new_n18676, new_n18675, new_n18671);
not_3  g16328(new_n18677, new_n18655);
xnor_3 g16329(new_n18678, new_n18657, new_n18677);
nand_4 g16330(new_n18679_1, new_n18678, new_n5837);
xnor_3 g16331(new_n18680, new_n18653_1, new_n18650);
not_3  g16332(new_n18681, new_n18680);
nand_4 g16333(new_n18682, new_n18681, new_n5847);
xor_3  g16334(new_n18683, new_n11364, new_n5803);
nand_4 g16335(new_n18684, new_n18683, new_n5850_1);
xnor_3 g16336(new_n18685, new_n18680, new_n5847);
nand_4 g16337(new_n18686, new_n18685, new_n18684);
nand_4 g16338(new_n18687, new_n18686, new_n18682);
xnor_3 g16339(new_n18688, new_n18678, new_n5792);
nand_4 g16340(new_n18689, new_n18688, new_n18687);
nand_4 g16341(new_n18690_1, new_n18689, new_n18679_1);
nand_4 g16342(new_n18691, new_n18690_1, new_n18676);
nand_4 g16343(new_n18692, new_n18691, new_n18672);
xor_3  g16344(n3301, new_n18692, new_n18668);
xnor_3 g16345(new_n18694, new_n12908, n3030);
not_3  g16346(new_n18695, new_n12898);
nand_4 g16347(new_n18696, new_n18695, n19515);
not_3  g16348(new_n18697, new_n18696);
nor_4  g16349(new_n18698, new_n18695, n19515);
nor_4  g16350(new_n18699, new_n18698, new_n18697);
not_3  g16351(new_n18700, new_n12888);
nor_4  g16352(new_n18701, new_n18700, new_n16488);
not_3  g16353(new_n18702, new_n18701);
nor_4  g16354(new_n18703, new_n12888, n22588);
nor_4  g16355(new_n18704, new_n18703, new_n18701);
nor_4  g16356(new_n18705, new_n12878, n12209);
nor_4  g16357(new_n18706, new_n16223_1, new_n18705);
nand_4 g16358(new_n18707, new_n18706, new_n18704);
nand_4 g16359(new_n18708_1, new_n18707, new_n18702);
nand_4 g16360(new_n18709, new_n18708_1, new_n18699);
nand_4 g16361(new_n18710, new_n18709, new_n18696);
not_3  g16362(new_n18711, new_n18710);
xnor_3 g16363(new_n18712, new_n18711, new_n18694);
xnor_3 g16364(new_n18713, new_n18712, new_n12053);
xnor_3 g16365(new_n18714, new_n18708_1, new_n18699);
nor_4  g16366(new_n18715, new_n18714, new_n12057);
not_3  g16367(new_n18716, new_n18715);
not_3  g16368(new_n18717, new_n18714);
xnor_3 g16369(new_n18718, new_n18717, new_n12057);
not_3  g16370(new_n18719, new_n18707);
nor_4  g16371(new_n18720, new_n18706, new_n18704);
nor_4  g16372(new_n18721_1, new_n18720, new_n18719);
not_3  g16373(new_n18722, new_n18721_1);
nor_4  g16374(new_n18723, new_n18722, new_n12062);
not_3  g16375(new_n18724, new_n18723);
xnor_3 g16376(new_n18725_1, new_n18721_1, new_n12062);
not_3  g16377(new_n18726, new_n16228);
nor_4  g16378(new_n18727, new_n18726, new_n16215_1);
nor_4  g16379(new_n18728, new_n18727, new_n16227);
not_3  g16380(new_n18729, new_n18728);
nand_4 g16381(new_n18730, new_n18729, new_n18725_1);
nand_4 g16382(new_n18731, new_n18730, new_n18724);
nand_4 g16383(new_n18732, new_n18731, new_n18718);
nand_4 g16384(new_n18733, new_n18732, new_n18716);
xor_3  g16385(n3316, new_n18733, new_n18713);
not_3  g16386(new_n18735, new_n16204);
xor_3  g16387(n3332, new_n18735, new_n16183);
nor_4  g16388(new_n18737_1, new_n12871_1, n17458);
xnor_3 g16389(new_n18738, new_n9446, new_n13199_1);
nor_4  g16390(new_n18739, new_n12957, n1222);
xnor_3 g16391(new_n18740, new_n9451_1, new_n8501);
nor_4  g16392(new_n18741, new_n9454, n25240);
nand_4 g16393(new_n18742, new_n12665_1, new_n12644);
not_3  g16394(new_n18743, new_n18742);
nor_4  g16395(new_n18744, new_n18743, new_n18741);
nor_4  g16396(new_n18745_1, new_n18744, new_n18740);
nor_4  g16397(new_n18746, new_n18745_1, new_n18739);
nor_4  g16398(new_n18747, new_n18746, new_n18738);
nor_4  g16399(new_n18748, new_n18747, new_n18737_1);
nand_4 g16400(new_n18749, new_n18748, new_n9524);
nand_4 g16401(new_n18750, new_n15535, n8827);
nand_4 g16402(new_n18751_1, new_n15554, new_n15558_1);
nand_4 g16403(new_n18752, new_n18751_1, new_n18750);
nor_4  g16404(new_n18753, n23166, n11898);
and_4  g16405(new_n18754, new_n15534, new_n15525);
nor_4  g16406(new_n18755, new_n18754, new_n18753);
nand_4 g16407(new_n18756, new_n18755, new_n18752);
xnor_3 g16408(new_n18757, new_n18756, new_n18749);
xnor_3 g16409(new_n18758, new_n18748, new_n9651);
xnor_3 g16410(new_n18759, new_n18755, new_n18752);
nor_4  g16411(new_n18760, new_n18759, new_n18758);
not_3  g16412(new_n18761, new_n18760);
not_3  g16413(new_n18762, new_n18758);
not_3  g16414(new_n18763, new_n18756);
nor_4  g16415(new_n18764, new_n18755, new_n18752);
nor_4  g16416(new_n18765, new_n18764, new_n18763);
nor_4  g16417(new_n18766, new_n18765, new_n18762);
nor_4  g16418(new_n18767, new_n18766, new_n18760);
not_3  g16419(new_n18768, new_n18738);
xnor_3 g16420(new_n18769, new_n18746, new_n18768);
nor_4  g16421(new_n18770, new_n18769, new_n15555_1);
xnor_3 g16422(new_n18771, new_n18769, new_n15555_1);
xnor_3 g16423(new_n18772, new_n18744, new_n18740);
nor_4  g16424(new_n18773, new_n18772, new_n15562);
not_3  g16425(new_n18774, new_n18773);
xnor_3 g16426(new_n18775, new_n18772, new_n15566);
not_3  g16427(new_n18776, new_n12712);
nand_4 g16428(new_n18777, new_n12741, new_n12713);
nand_4 g16429(new_n18778, new_n18777, new_n18776);
nand_4 g16430(new_n18779, new_n18778, new_n18775);
nand_4 g16431(new_n18780_1, new_n18779, new_n18774);
nor_4  g16432(new_n18781, new_n18780_1, new_n18771);
nor_4  g16433(new_n18782_1, new_n18781, new_n18770);
nand_4 g16434(new_n18783, new_n18782_1, new_n18767);
nand_4 g16435(new_n18784, new_n18783, new_n18761);
xnor_3 g16436(n3340, new_n18784, new_n18757);
xor_3  g16437(new_n18786, n13851, new_n12668);
nor_4  g16438(new_n18787, n24937, new_n12692);
not_3  g16439(new_n18788, new_n18787);
xor_3  g16440(new_n18789, n24937, new_n12692);
nor_4  g16441(new_n18790, new_n18066, n5098);
not_3  g16442(new_n18791, new_n18790);
not_3  g16443(new_n18792, n5098);
xor_3  g16444(new_n18793, n26452, new_n18792);
nor_4  g16445(new_n18794, new_n4668, n3030);
not_3  g16446(new_n18795, new_n18794);
xor_3  g16447(new_n18796, n19905, n3030);
not_3  g16448(new_n18797, new_n18796);
not_3  g16449(new_n18798, n19515);
nor_4  g16450(new_n18799, new_n18798, n17035);
nor_4  g16451(new_n18800, new_n16498, new_n16487);
nor_4  g16452(new_n18801, new_n18800, new_n18799);
nand_4 g16453(new_n18802_1, new_n18801, new_n18797);
nand_4 g16454(new_n18803, new_n18802_1, new_n18795);
nand_4 g16455(new_n18804, new_n18803, new_n18793);
nand_4 g16456(new_n18805, new_n18804, new_n18791);
nand_4 g16457(new_n18806, new_n18805, new_n18789);
nand_4 g16458(new_n18807, new_n18806, new_n18788);
xor_3  g16459(new_n18808, new_n18807, new_n18786);
xnor_3 g16460(new_n18809, new_n18808, new_n18551);
xor_3  g16461(new_n18810, new_n18805, new_n18789);
nor_4  g16462(new_n18811, new_n18810, new_n18556);
not_3  g16463(new_n18812, new_n18811);
not_3  g16464(new_n18813, new_n18810);
nor_4  g16465(new_n18814, new_n18813, new_n18603);
nor_4  g16466(new_n18815, new_n18814, new_n18811);
xor_3  g16467(new_n18816, new_n18803, new_n18793);
nor_4  g16468(new_n18817, new_n18816, new_n18560);
not_3  g16469(new_n18818, new_n18817);
not_3  g16470(new_n18819, new_n18816);
nor_4  g16471(new_n18820, new_n18819, new_n18565);
nor_4  g16472(new_n18821, new_n18820, new_n18817);
xor_3  g16473(new_n18822, new_n18801, new_n18796);
nor_4  g16474(new_n18823, new_n18822, new_n18571);
xnor_3 g16475(new_n18824, new_n18822, new_n18571);
nand_4 g16476(new_n18825, new_n16499, new_n16486);
nand_4 g16477(new_n18826, new_n16531, new_n16501);
nand_4 g16478(new_n18827, new_n18826, new_n18825);
nor_4  g16479(new_n18828, new_n18827, new_n18824);
nor_4  g16480(new_n18829, new_n18828, new_n18823);
nand_4 g16481(new_n18830_1, new_n18829, new_n18821);
nand_4 g16482(new_n18831_1, new_n18830_1, new_n18818);
nand_4 g16483(new_n18832, new_n18831_1, new_n18815);
nand_4 g16484(new_n18833, new_n18832, new_n18812);
xor_3  g16485(n3343, new_n18833, new_n18809);
nor_4  g16486(new_n18835, new_n15004_1, n10250);
not_3  g16487(new_n18836, new_n18835);
xnor_3 g16488(new_n18837, new_n14995, new_n10324);
not_3  g16489(new_n18838, new_n18837);
nand_4 g16490(new_n18839, new_n15007, new_n10329);
xor_3  g16491(new_n18840, new_n15007, new_n10329);
not_3  g16492(new_n18841, new_n15012);
nand_4 g16493(new_n18842, new_n18841, new_n10331);
xor_3  g16494(new_n18843_1, new_n18841, new_n10331);
nand_4 g16495(new_n18844, new_n15021, new_n7209);
xor_3  g16496(new_n18845, new_n15021, new_n7209);
nand_4 g16497(new_n18846, new_n15027, new_n14427);
xor_3  g16498(new_n18847, new_n15027, new_n14427);
nor_4  g16499(new_n18848, new_n15034, n21226);
not_3  g16500(new_n18849, new_n18848);
nor_4  g16501(new_n18850, new_n15030, new_n14431);
nor_4  g16502(new_n18851, new_n18850, new_n18848);
nor_4  g16503(new_n18852, new_n15041, n4426);
not_3  g16504(new_n18853, new_n18852);
nor_4  g16505(new_n18854, new_n15040, new_n14435);
nor_4  g16506(new_n18855, new_n18854, new_n18852);
nor_4  g16507(new_n18856, new_n15053_1, n20036);
not_3  g16508(new_n18857, new_n18856);
nor_4  g16509(new_n18858_1, new_n15049, new_n10346);
nor_4  g16510(new_n18859_1, new_n18858_1, new_n18856);
nor_4  g16511(new_n18860, new_n15061, new_n4607);
nor_4  g16512(new_n18861, new_n15057, n9380);
xnor_3 g16513(new_n18862, new_n15061, new_n4607);
nor_4  g16514(new_n18863, new_n18862, new_n18861);
nor_4  g16515(new_n18864_1, new_n18863, new_n18860);
nand_4 g16516(new_n18865_1, new_n18864_1, new_n18859_1);
nand_4 g16517(new_n18866, new_n18865_1, new_n18857);
nand_4 g16518(new_n18867, new_n18866, new_n18855);
nand_4 g16519(new_n18868, new_n18867, new_n18853);
nand_4 g16520(new_n18869, new_n18868, new_n18851);
nand_4 g16521(new_n18870, new_n18869, new_n18849);
nand_4 g16522(new_n18871, new_n18870, new_n18847);
nand_4 g16523(new_n18872, new_n18871, new_n18846);
nand_4 g16524(new_n18873, new_n18872, new_n18845);
nand_4 g16525(new_n18874, new_n18873, new_n18844);
nand_4 g16526(new_n18875, new_n18874, new_n18843_1);
nand_4 g16527(new_n18876, new_n18875, new_n18842);
nand_4 g16528(new_n18877, new_n18876, new_n18840);
nand_4 g16529(new_n18878, new_n18877, new_n18839);
nand_4 g16530(new_n18879, new_n18878, new_n18838);
nand_4 g16531(new_n18880_1, new_n18879, new_n18836);
xnor_3 g16532(new_n18881, new_n18880_1, new_n14868);
nor_4  g16533(new_n18882, new_n18496_1, n19270);
not_3  g16534(new_n18883, new_n18882);
xor_3  g16535(new_n18884, new_n18883, n14704);
nor_4  g16536(new_n18885, new_n18884, n19531);
not_3  g16537(new_n18886_1, new_n18884);
xor_3  g16538(new_n18887_1, new_n18886_1, new_n10379);
not_3  g16539(new_n18888, new_n18887_1);
nor_4  g16540(new_n18889, new_n18497, n18345);
not_3  g16541(new_n18890, new_n18499);
nor_4  g16542(new_n18891, new_n18547, new_n18890);
nor_4  g16543(new_n18892, new_n18891, new_n18889);
nor_4  g16544(new_n18893, new_n18892, new_n18888);
nor_4  g16545(new_n18894, new_n18893, new_n18885);
nor_4  g16546(new_n18895, new_n18883, n14704);
xor_3  g16547(new_n18896, new_n18895, new_n2611);
nor_4  g16548(new_n18897, new_n18896, n20040);
not_3  g16549(new_n18898, n20040);
not_3  g16550(new_n18899, new_n18896);
nor_4  g16551(new_n18900, new_n18899, new_n18898);
nor_4  g16552(new_n18901_1, new_n18900, new_n18897);
xnor_3 g16553(new_n18902, new_n18901_1, new_n18894);
nor_4  g16554(new_n18903, new_n18902, new_n16946);
not_3  g16555(new_n18904, new_n18903);
not_3  g16556(new_n18905, new_n18902);
nor_4  g16557(new_n18906, new_n18905, new_n16944);
not_3  g16558(new_n18907_1, new_n18892);
nor_4  g16559(new_n18908, new_n18907_1, new_n18887_1);
nor_4  g16560(new_n18909, new_n18908, new_n18893);
nor_4  g16561(new_n18910, new_n18909, new_n16928);
xnor_3 g16562(new_n18911, new_n18892, new_n18888);
xnor_3 g16563(new_n18912, new_n18911, new_n16928);
nor_4  g16564(new_n18913, new_n18548, new_n16932);
not_3  g16565(new_n18914, new_n18913);
nor_4  g16566(new_n18915, new_n18552, new_n16930);
nor_4  g16567(new_n18916, new_n18915, new_n18913);
not_3  g16568(new_n18917, new_n7569_1);
nor_4  g16569(new_n18918, new_n18601, new_n18917);
not_3  g16570(new_n18919_1, new_n18918);
nor_4  g16571(new_n18920, new_n18555, new_n7569_1);
nor_4  g16572(new_n18921, new_n18920, new_n18918);
nor_4  g16573(new_n18922, new_n18563, new_n7580);
not_3  g16574(new_n18923, new_n18922);
nor_4  g16575(new_n18924, new_n18569, new_n7584);
not_3  g16576(new_n18925, new_n18924);
nor_4  g16577(new_n18926_1, new_n18568, new_n7586);
nor_4  g16578(new_n18927, new_n18926_1, new_n18924);
nor_4  g16579(new_n18928, new_n18573, new_n7592);
xnor_3 g16580(new_n18929, new_n18573, new_n7592);
nor_4  g16581(new_n18930, new_n18578_1, new_n7595);
not_3  g16582(new_n18931, new_n18930);
nor_4  g16583(new_n18932, new_n18577, new_n7596);
nor_4  g16584(new_n18933, new_n18932, new_n18930);
nor_4  g16585(new_n18934, new_n18581, new_n7606);
not_3  g16586(new_n18935, n4939);
nor_4  g16587(new_n18936, new_n18584_1, new_n18935);
xnor_3 g16588(new_n18937, new_n18581, new_n7606);
nor_4  g16589(new_n18938, new_n18937, new_n18936);
nor_4  g16590(new_n18939, new_n18938, new_n18934);
nand_4 g16591(new_n18940_1, new_n18939, new_n18933);
nand_4 g16592(new_n18941, new_n18940_1, new_n18931);
nor_4  g16593(new_n18942, new_n18941, new_n18929);
nor_4  g16594(new_n18943, new_n18942, new_n18928);
nand_4 g16595(new_n18944, new_n18943, new_n18927);
nand_4 g16596(new_n18945_1, new_n18944, new_n18925);
nor_4  g16597(new_n18946, new_n18559, new_n7576);
nor_4  g16598(new_n18947, new_n18946, new_n18922);
nand_4 g16599(new_n18948, new_n18947, new_n18945_1);
nand_4 g16600(new_n18949, new_n18948, new_n18923);
nand_4 g16601(new_n18950, new_n18949, new_n18921);
nand_4 g16602(new_n18951, new_n18950, new_n18919_1);
nand_4 g16603(new_n18952, new_n18951, new_n18916);
nand_4 g16604(new_n18953, new_n18952, new_n18914);
nand_4 g16605(new_n18954, new_n18953, new_n18912);
not_3  g16606(new_n18955, new_n18954);
nor_4  g16607(new_n18956, new_n18955, new_n18910);
nor_4  g16608(new_n18957, new_n18956, new_n18906);
nor_4  g16609(new_n18958, new_n18957, new_n16974);
nand_4 g16610(new_n18959, new_n18958, new_n18904);
not_3  g16611(new_n18960, new_n18895);
nor_4  g16612(new_n18961, new_n18960, n25365);
nor_4  g16613(new_n18962_1, new_n18900, new_n18894);
nor_4  g16614(new_n18963, new_n18962_1, new_n18897);
nor_4  g16615(new_n18964, new_n18963, new_n18961);
xnor_3 g16616(new_n18965, new_n18964, new_n18959);
not_3  g16617(new_n18966, new_n18965);
nand_4 g16618(new_n18967, new_n18966, new_n18881);
xnor_3 g16619(new_n18968, new_n18878, new_n18837);
nor_4  g16620(new_n18969, new_n18906, new_n18903);
xnor_3 g16621(new_n18970_1, new_n18969, new_n18956);
not_3  g16622(new_n18971, new_n18970_1);
nand_4 g16623(new_n18972, new_n18971, new_n18968);
xnor_3 g16624(new_n18973, new_n18970_1, new_n18968);
not_3  g16625(new_n18974, new_n18840);
xnor_3 g16626(new_n18975, new_n18876, new_n18974);
nor_4  g16627(new_n18976, new_n18953, new_n18912);
nor_4  g16628(new_n18977_1, new_n18976, new_n18955);
not_3  g16629(new_n18978, new_n18977_1);
nand_4 g16630(new_n18979, new_n18978, new_n18975);
xnor_3 g16631(new_n18980, new_n18977_1, new_n18975);
xnor_3 g16632(new_n18981, new_n18874, new_n18843_1);
xnor_3 g16633(new_n18982_1, new_n18951, new_n18916);
not_3  g16634(new_n18983, new_n18982_1);
nor_4  g16635(new_n18984, new_n18983, new_n18981);
not_3  g16636(new_n18985, new_n18984);
not_3  g16637(new_n18986, new_n18981);
nor_4  g16638(new_n18987, new_n18982_1, new_n18986);
nor_4  g16639(new_n18988, new_n18987, new_n18984);
xnor_3 g16640(new_n18989, new_n18872, new_n18845);
not_3  g16641(new_n18990, new_n18989);
xnor_3 g16642(new_n18991, new_n18949, new_n18921);
nand_4 g16643(new_n18992, new_n18991, new_n18990);
xnor_3 g16644(new_n18993, new_n18991, new_n18989);
xnor_3 g16645(new_n18994, new_n18870, new_n18847);
not_3  g16646(new_n18995, new_n18994);
xnor_3 g16647(new_n18996, new_n18947, new_n18945_1);
nand_4 g16648(new_n18997, new_n18996, new_n18995);
xnor_3 g16649(new_n18998, new_n18996, new_n18994);
xnor_3 g16650(new_n18999_1, new_n18868, new_n18851);
not_3  g16651(new_n19000, new_n18999_1);
xnor_3 g16652(new_n19001, new_n18943, new_n18927);
nand_4 g16653(new_n19002, new_n19001, new_n19000);
xnor_3 g16654(new_n19003, new_n19001, new_n18999_1);
not_3  g16655(new_n19004, new_n18855);
xnor_3 g16656(new_n19005_1, new_n18866, new_n19004);
xnor_3 g16657(new_n19006, new_n18941, new_n18929);
not_3  g16658(new_n19007, new_n19006);
nand_4 g16659(new_n19008, new_n19007, new_n19005_1);
xnor_3 g16660(new_n19009, new_n19006, new_n19005_1);
xnor_3 g16661(new_n19010, new_n18864_1, new_n18859_1);
not_3  g16662(new_n19011, new_n19010);
xnor_3 g16663(new_n19012, new_n18939, new_n18933);
nand_4 g16664(new_n19013, new_n19012, new_n19011);
xnor_3 g16665(new_n19014, new_n18937, new_n18936);
not_3  g16666(new_n19015, new_n19014);
not_3  g16667(new_n19016, new_n18861);
xnor_3 g16668(new_n19017, new_n18862, new_n19016);
not_3  g16669(new_n19018, new_n19017);
nor_4  g16670(new_n19019, new_n19018, new_n19015);
nor_4  g16671(new_n19020, new_n18302, n4939);
nor_4  g16672(new_n19021, new_n19020, new_n18936);
not_3  g16673(new_n19022, new_n15057);
xor_3  g16674(new_n19023, new_n19022, n9380);
nand_4 g16675(new_n19024, new_n19023, new_n19021);
xnor_3 g16676(new_n19025, new_n19017, new_n19014);
nor_4  g16677(new_n19026, new_n19025, new_n19024);
nor_4  g16678(new_n19027, new_n19026, new_n19019);
not_3  g16679(new_n19028, new_n19013);
nor_4  g16680(new_n19029, new_n19012, new_n19011);
nor_4  g16681(new_n19030, new_n19029, new_n19028);
nand_4 g16682(new_n19031, new_n19030, new_n19027);
nand_4 g16683(new_n19032, new_n19031, new_n19013);
nand_4 g16684(new_n19033_1, new_n19032, new_n19009);
nand_4 g16685(new_n19034, new_n19033_1, new_n19008);
nand_4 g16686(new_n19035, new_n19034, new_n19003);
nand_4 g16687(new_n19036, new_n19035, new_n19002);
nand_4 g16688(new_n19037, new_n19036, new_n18998);
nand_4 g16689(new_n19038, new_n19037, new_n18997);
nand_4 g16690(new_n19039, new_n19038, new_n18993);
nand_4 g16691(new_n19040, new_n19039, new_n18992);
nand_4 g16692(new_n19041, new_n19040, new_n18988);
nand_4 g16693(new_n19042_1, new_n19041, new_n18985);
nand_4 g16694(new_n19043, new_n19042_1, new_n18980);
nand_4 g16695(new_n19044_1, new_n19043, new_n18979);
nand_4 g16696(new_n19045, new_n19044_1, new_n18973);
nand_4 g16697(new_n19046, new_n19045, new_n18972);
xnor_3 g16698(new_n19047, new_n18965, new_n18881);
nand_4 g16699(new_n19048, new_n19047, new_n19046);
nand_4 g16700(new_n19049, new_n19048, new_n18967);
nor_4  g16701(new_n19050, new_n18880_1, new_n14868);
nor_4  g16702(new_n19051, new_n18964, new_n18959);
xnor_3 g16703(new_n19052, new_n19051, new_n19050);
xnor_3 g16704(n3390, new_n19052, new_n19049);
not_3  g16705(new_n19054, new_n7715);
xor_3  g16706(n3426, new_n7717, new_n19054);
xor_3  g16707(n3451, new_n5397, new_n5394);
not_3  g16708(new_n19057, new_n14677);
xor_3  g16709(n3459, new_n19057, new_n14649);
xnor_3 g16710(new_n19059, n6773, n583);
xor_3  g16711(new_n19060, new_n19059, n21687);
nor_4  g16712(new_n19061, new_n19060, new_n16641);
nand_4 g16713(new_n19062, new_n19059, n21687);
nand_4 g16714(new_n19063, new_n19062, new_n14693);
not_3  g16715(new_n19064, new_n19063);
not_3  g16716(new_n19065, new_n19059);
nor_4  g16717(new_n19066, new_n19065, new_n4521);
nor_4  g16718(new_n19067, new_n19066, new_n19064);
nand_4 g16719(new_n19068, n6773, n583);
nor_4  g16720(new_n19069, n22173, n17090);
nand_4 g16721(new_n19070, n22173, n17090);
not_3  g16722(new_n19071, new_n19070);
nor_4  g16723(new_n19072, new_n19071, new_n19069);
xor_3  g16724(new_n19073, new_n19072, new_n19068);
not_3  g16725(new_n19074, new_n19073);
xnor_3 g16726(new_n19075, new_n19074, new_n19067);
nand_4 g16727(new_n19076, new_n19075, new_n16644);
not_3  g16728(new_n19077, new_n19076);
nor_4  g16729(new_n19078, new_n19075, new_n16644);
nor_4  g16730(new_n19079, new_n19078, new_n19077);
xor_3  g16731(n3502, new_n19079, new_n19061);
xnor_3 g16732(n3516, new_n13067, new_n13023);
not_3  g16733(new_n19082, n18145);
not_3  g16734(new_n19083, n25126);
not_3  g16735(new_n19084, n1689);
nor_4  g16736(new_n19085, n24129, n22274);
nand_4 g16737(new_n19086, new_n19085, new_n19084);
nor_4  g16738(new_n19087, new_n19086, n19608);
nand_4 g16739(new_n19088, new_n19087, new_n19083);
nor_4  g16740(new_n19089, new_n19088, n10712);
xor_3  g16741(new_n19090, new_n19089, new_n19082);
not_3  g16742(new_n19091, new_n19090);
xor_3  g16743(new_n19092, new_n19091, n15761);
xor_3  g16744(new_n19093, new_n19088, n10712);
nor_4  g16745(new_n19094, new_n19093, new_n12333);
not_3  g16746(new_n19095, new_n19094);
not_3  g16747(new_n19096, new_n19093);
xor_3  g16748(new_n19097, new_n19096, n11201);
not_3  g16749(new_n19098, new_n19088);
nor_4  g16750(new_n19099, new_n19087, new_n19083);
nor_4  g16751(new_n19100, new_n19099, new_n19098);
nor_4  g16752(new_n19101, new_n19100, new_n12338);
not_3  g16753(new_n19102, new_n19100);
nor_4  g16754(new_n19103, new_n19102, n18690);
nor_4  g16755(new_n19104, new_n19103, new_n19101);
nand_4 g16756(new_n19105, new_n19086, n19608);
not_3  g16757(new_n19106, new_n19105);
nor_4  g16758(new_n19107_1, new_n19106, new_n19087);
nor_4  g16759(new_n19108, new_n19107_1, new_n12344);
not_3  g16760(new_n19109, new_n19108);
not_3  g16761(new_n19110, new_n19107_1);
nor_4  g16762(new_n19111, new_n19110, n12153);
nor_4  g16763(new_n19112, new_n19111, new_n19108);
not_3  g16764(new_n19113, new_n19086);
nor_4  g16765(new_n19114, new_n19085, new_n19084);
nor_4  g16766(new_n19115, new_n19114, new_n19113);
nor_4  g16767(new_n19116_1, new_n19115, new_n12347);
not_3  g16768(new_n19117, new_n19116_1);
not_3  g16769(new_n19118, new_n19115);
nor_4  g16770(new_n19119, new_n19118, n13044);
nor_4  g16771(new_n19120, new_n19119, new_n19116_1);
xnor_3 g16772(new_n19121, n24129, n22274);
nand_4 g16773(new_n19122, new_n19121, n18745);
not_3  g16774(new_n19123, n24129);
nand_4 g16775(new_n19124, new_n19123, n16167);
not_3  g16776(new_n19125_1, new_n19124);
xnor_3 g16777(new_n19126, new_n19121, n18745);
not_3  g16778(new_n19127, new_n19126);
nand_4 g16779(new_n19128, new_n19127, new_n19125_1);
nand_4 g16780(new_n19129, new_n19128, new_n19122);
nand_4 g16781(new_n19130, new_n19129, new_n19120);
nand_4 g16782(new_n19131, new_n19130, new_n19117);
nand_4 g16783(new_n19132, new_n19131, new_n19112);
nand_4 g16784(new_n19133, new_n19132, new_n19109);
nand_4 g16785(new_n19134, new_n19133, new_n19104);
not_3  g16786(new_n19135, new_n19134);
nor_4  g16787(new_n19136, new_n19135, new_n19101);
not_3  g16788(new_n19137, new_n19136);
nand_4 g16789(new_n19138, new_n19137, new_n19097);
nand_4 g16790(new_n19139, new_n19138, new_n19095);
nand_4 g16791(new_n19140, new_n19139, new_n19092);
not_3  g16792(new_n19141_1, new_n19140);
nor_4  g16793(new_n19142, new_n19139, new_n19092);
nor_4  g16794(new_n19143, new_n19142, new_n19141_1);
xnor_3 g16795(new_n19144_1, new_n19143, new_n8087);
not_3  g16796(new_n19145, new_n19138);
nor_4  g16797(new_n19146, new_n19137, new_n19097);
nor_4  g16798(new_n19147, new_n19146, new_n19145);
nand_4 g16799(new_n19148, new_n19147, new_n8092);
xnor_3 g16800(new_n19149, new_n19147, new_n8095_1);
nor_4  g16801(new_n19150, new_n19133, new_n19104);
nor_4  g16802(new_n19151, new_n19150, new_n19135);
nand_4 g16803(new_n19152, new_n19151, new_n8099);
xnor_3 g16804(new_n19153, new_n19151, new_n8102);
xnor_3 g16805(new_n19154, new_n19131, new_n19112);
nor_4  g16806(new_n19155, new_n19154, new_n8106);
not_3  g16807(new_n19156, new_n19155);
not_3  g16808(new_n19157, new_n19154);
nor_4  g16809(new_n19158, new_n19157, new_n8107);
nor_4  g16810(new_n19159, new_n19158, new_n19155);
xnor_3 g16811(new_n19160, new_n19129, new_n19120);
nand_4 g16812(new_n19161, new_n19160, new_n8119);
not_3  g16813(new_n19162, new_n19161);
xnor_3 g16814(new_n19163_1, new_n19160, new_n8119);
xnor_3 g16815(new_n19164_1, new_n19126, new_n19124);
not_3  g16816(new_n19165, new_n19164_1);
nor_4  g16817(new_n19166, new_n19165, new_n4618);
xor_3  g16818(new_n19167, n24129, n16167);
nand_4 g16819(new_n19168, new_n19167, new_n4625);
xnor_3 g16820(new_n19169, new_n19164_1, new_n4629);
nor_4  g16821(new_n19170, new_n19169, new_n19168);
nor_4  g16822(new_n19171, new_n19170, new_n19166);
nor_4  g16823(new_n19172, new_n19171, new_n19163_1);
nor_4  g16824(new_n19173, new_n19172, new_n19162);
nand_4 g16825(new_n19174_1, new_n19173, new_n19159);
nand_4 g16826(new_n19175, new_n19174_1, new_n19156);
nand_4 g16827(new_n19176_1, new_n19175, new_n19153);
nand_4 g16828(new_n19177, new_n19176_1, new_n19152);
nand_4 g16829(new_n19178, new_n19177, new_n19149);
nand_4 g16830(new_n19179, new_n19178, new_n19148);
xnor_3 g16831(new_n19180, new_n19179, new_n19144_1);
nand_4 g16832(new_n19181, new_n19180, new_n12488);
xnor_3 g16833(new_n19182, new_n19143, new_n8084);
xnor_3 g16834(new_n19183, new_n19179, new_n19182);
nand_4 g16835(new_n19184, new_n19183, new_n12487);
nand_4 g16836(new_n19185, new_n19184, new_n19181);
not_3  g16837(new_n19186, new_n19149);
xnor_3 g16838(new_n19187, new_n19177, new_n19186);
nand_4 g16839(new_n19188, new_n19187, new_n12496);
xnor_3 g16840(new_n19189, new_n19187, new_n12497);
not_3  g16841(new_n19190, new_n19159);
not_3  g16842(new_n19191, new_n19163_1);
not_3  g16843(new_n19192, new_n19166);
not_3  g16844(new_n19193, new_n19168);
nor_4  g16845(new_n19194, new_n19164_1, new_n4629);
nor_4  g16846(new_n19195, new_n19194, new_n19166);
nand_4 g16847(new_n19196_1, new_n19195, new_n19193);
nand_4 g16848(new_n19197, new_n19196_1, new_n19192);
nand_4 g16849(new_n19198, new_n19197, new_n19191);
nand_4 g16850(new_n19199, new_n19198, new_n19161);
nor_4  g16851(new_n19200, new_n19199, new_n19190);
nor_4  g16852(new_n19201, new_n19200, new_n19155);
xnor_3 g16853(new_n19202_1, new_n19201, new_n19153);
nand_4 g16854(new_n19203, new_n19202_1, new_n12509);
xnor_3 g16855(new_n19204, new_n19202_1, new_n12510);
nor_4  g16856(new_n19205, new_n19173, new_n19159);
nor_4  g16857(new_n19206, new_n19205, new_n19200);
nand_4 g16858(new_n19207, new_n19206, new_n12519);
nor_4  g16859(new_n19208, new_n19197, new_n19191);
nor_4  g16860(new_n19209, new_n19208, new_n19172);
not_3  g16861(new_n19210, new_n19209);
nand_4 g16862(new_n19211, new_n19210, new_n12526);
xnor_3 g16863(new_n19212, new_n19209, new_n12526);
not_3  g16864(new_n19213, new_n6802_1);
xnor_3 g16865(new_n19214, new_n19169, new_n19168);
nand_4 g16866(new_n19215, new_n19214, new_n19213);
not_3  g16867(new_n19216, new_n6777);
nor_4  g16868(new_n19217, new_n19167, new_n4625);
nor_4  g16869(new_n19218, new_n19217, new_n19193);
nand_4 g16870(new_n19219, new_n19218, new_n19216);
xnor_3 g16871(new_n19220_1, new_n19214, new_n6802_1);
nand_4 g16872(new_n19221_1, new_n19220_1, new_n19219);
nand_4 g16873(new_n19222, new_n19221_1, new_n19215);
nand_4 g16874(new_n19223_1, new_n19222, new_n19212);
nand_4 g16875(new_n19224_1, new_n19223_1, new_n19211);
xnor_3 g16876(new_n19225, new_n19206, new_n12520);
nand_4 g16877(new_n19226, new_n19225, new_n19224_1);
nand_4 g16878(new_n19227, new_n19226, new_n19207);
nand_4 g16879(new_n19228_1, new_n19227, new_n19204);
nand_4 g16880(new_n19229, new_n19228_1, new_n19203);
nand_4 g16881(new_n19230, new_n19229, new_n19189);
nand_4 g16882(new_n19231, new_n19230, new_n19188);
xor_3  g16883(n3528, new_n19231, new_n19185);
xnor_3 g16884(n3555, new_n10864, new_n10790);
nor_4  g16885(new_n19234_1, new_n2907, new_n2824);
nor_4  g16886(new_n19235, new_n19234_1, new_n2820);
not_3  g16887(new_n19236, new_n19235);
not_3  g16888(new_n19237, new_n2769);
nor_4  g16889(new_n19238, new_n19237, n13951);
not_3  g16890(new_n19239, new_n19238);
nor_4  g16891(new_n19240, new_n12164, new_n19239);
nand_4 g16892(new_n19241, new_n19240, new_n19236);
not_3  g16893(new_n19242, new_n19241);
not_3  g16894(new_n19243, new_n12164);
nor_4  g16895(new_n19244_1, new_n19243, new_n19238);
nand_4 g16896(new_n19245, new_n19244_1, new_n19235);
nand_4 g16897(new_n19246, new_n19245, new_n19241);
nand_4 g16898(new_n19247, new_n19246, new_n17817);
xnor_3 g16899(new_n19248, new_n19246, new_n17816);
nor_4  g16900(new_n19249, new_n19244_1, new_n19240);
xnor_3 g16901(new_n19250, new_n19249, new_n19235);
nand_4 g16902(new_n19251, new_n19250, new_n17820_1);
xnor_3 g16903(new_n19252, new_n19250, new_n17821);
nand_4 g16904(new_n19253, new_n2908, new_n17826);
nand_4 g16905(new_n19254, new_n2981, new_n2909);
nand_4 g16906(new_n19255, new_n19254, new_n19253);
nand_4 g16907(new_n19256, new_n19255, new_n19252);
nand_4 g16908(new_n19257, new_n19256, new_n19251);
nand_4 g16909(new_n19258, new_n19257, new_n19248);
nand_4 g16910(new_n19259, new_n19258, new_n19247);
not_3  g16911(new_n19260, new_n19259);
nor_4  g16912(n3561, new_n19260, new_n19242);
xor_3  g16913(new_n19262, n16439, new_n9083);
nor_4  g16914(new_n19263, new_n9087, n15241);
not_3  g16915(new_n19264, new_n19263);
nand_4 g16916(new_n19265, new_n12768, new_n12743);
nand_4 g16917(new_n19266, new_n19265, new_n19264);
not_3  g16918(new_n19267, new_n19266);
xnor_3 g16919(new_n19268, new_n19267, new_n19262);
xor_3  g16920(new_n19269, new_n11603, new_n9036);
not_3  g16921(new_n19270_1, new_n19269);
nand_4 g16922(new_n19271, new_n11607_1, new_n8849_1);
nand_4 g16923(new_n19272, new_n12783_1, new_n12770);
nand_4 g16924(new_n19273, new_n19272, new_n19271);
xnor_3 g16925(new_n19274, new_n19273, new_n19270_1);
not_3  g16926(new_n19275, new_n19274);
xnor_3 g16927(new_n19276, new_n19275, new_n19268);
not_3  g16928(new_n19277, new_n12769);
not_3  g16929(new_n19278, new_n12784);
nand_4 g16930(new_n19279, new_n19278, new_n19277);
not_3  g16931(new_n19280, new_n12785);
not_3  g16932(new_n19281, new_n12799);
not_3  g16933(new_n19282_1, new_n12800);
not_3  g16934(new_n19283, new_n12829);
nand_4 g16935(new_n19284, new_n19283, new_n19282_1);
nand_4 g16936(new_n19285, new_n19284, new_n19281);
nand_4 g16937(new_n19286, new_n19285, new_n19280);
nand_4 g16938(new_n19287, new_n19286, new_n19279);
xnor_3 g16939(new_n19288, new_n19287, new_n19276);
xnor_3 g16940(new_n19289, new_n19288, new_n6529);
nand_4 g16941(new_n19290, new_n12833, new_n19286);
nor_4  g16942(new_n19291, new_n19290, new_n6531);
nor_4  g16943(new_n19292, new_n12868, new_n12836);
nor_4  g16944(new_n19293, new_n19292, new_n19291);
xor_3  g16945(n3563, new_n19293, new_n19289);
xor_3  g16946(n3617, new_n7181, new_n7180);
xor_3  g16947(new_n19296, n22253, new_n15331);
not_3  g16948(new_n19297, new_n19296);
not_3  g16949(new_n19298, n1255);
nor_4  g16950(new_n19299, n12861, new_n19298);
xor_3  g16951(new_n19300, n12861, new_n19298);
not_3  g16952(new_n19301, n9512);
or_4   g16953(new_n19302, n13333, new_n19301);
xor_3  g16954(new_n19303, n13333, new_n19301);
nand_4 g16955(new_n19304, n16608, new_n8298);
nand_4 g16956(new_n19305, n21735, new_n5229);
nand_4 g16957(new_n19306, new_n5259, new_n5230);
nand_4 g16958(new_n19307, new_n19306, new_n19305);
xor_3  g16959(new_n19308, n16608, new_n8298);
nand_4 g16960(new_n19309, new_n19308, new_n19307);
nand_4 g16961(new_n19310, new_n19309, new_n19304);
nand_4 g16962(new_n19311, new_n19310, new_n19303);
nand_4 g16963(new_n19312, new_n19311, new_n19302);
nand_4 g16964(new_n19313, new_n19312, new_n19300);
not_3  g16965(new_n19314_1, new_n19313);
nor_4  g16966(new_n19315_1, new_n19314_1, new_n19299);
xor_3  g16967(new_n19316, new_n19315_1, new_n19297);
not_3  g16968(new_n19317, new_n19316);
nor_4  g16969(new_n19318, new_n19317, new_n13638);
not_3  g16970(new_n19319, new_n13638);
nor_4  g16971(new_n19320, new_n19316, new_n19319);
nor_4  g16972(new_n19321, new_n19320, new_n19318);
xor_3  g16973(new_n19322, new_n19312, new_n19300);
nor_4  g16974(new_n19323_1, new_n19322, new_n13642);
not_3  g16975(new_n19324, new_n19322);
nor_4  g16976(new_n19325, new_n19324, new_n13646);
nor_4  g16977(new_n19326, new_n19325, new_n19323_1);
not_3  g16978(new_n19327_1, new_n19326);
xor_3  g16979(new_n19328, new_n19310, new_n19303);
nor_4  g16980(new_n19329, new_n19328, new_n13651);
not_3  g16981(new_n19330, new_n19329);
xor_3  g16982(new_n19331, new_n19308, new_n19307);
nand_4 g16983(new_n19332, new_n19331, new_n13661);
not_3  g16984(new_n19333_1, new_n19332);
xnor_3 g16985(new_n19334, new_n19331, new_n13661);
nand_4 g16986(new_n19335, new_n5373, new_n5260);
not_3  g16987(new_n19336, new_n19335);
nor_4  g16988(new_n19337, new_n5415, new_n5374);
nor_4  g16989(new_n19338, new_n19337, new_n19336);
nor_4  g16990(new_n19339, new_n19338, new_n19334);
nor_4  g16991(new_n19340, new_n19339, new_n19333_1);
not_3  g16992(new_n19341, new_n19328);
nor_4  g16993(new_n19342, new_n19341, new_n13656);
nor_4  g16994(new_n19343, new_n19342, new_n19329);
nand_4 g16995(new_n19344, new_n19343, new_n19340);
nand_4 g16996(new_n19345, new_n19344, new_n19330);
not_3  g16997(new_n19346, new_n19345);
nor_4  g16998(new_n19347, new_n19346, new_n19327_1);
nor_4  g16999(new_n19348_1, new_n19347, new_n19323_1);
nand_4 g17000(new_n19349, new_n19348_1, new_n19321);
not_3  g17001(new_n19350, new_n19349);
nor_4  g17002(new_n19351, new_n19348_1, new_n19321);
nor_4  g17003(n3642, new_n19351, new_n19350);
not_3  g17004(new_n19353, n3324);
xor_3  g17005(new_n19354_1, n16544, n4319);
nand_4 g17006(new_n19355, new_n13462, new_n10732);
xor_3  g17007(new_n19356, n23463, n6814);
nor_4  g17008(new_n19357_1, n19701, n13074);
not_3  g17009(new_n19358, new_n19357_1);
xor_3  g17010(new_n19359, n19701, n13074);
nor_4  g17011(new_n19360, n23529, n10739);
not_3  g17012(new_n19361_1, new_n19360);
xor_3  g17013(new_n19362, n23529, n10739);
nor_4  g17014(new_n19363, n24620, n21753);
not_3  g17015(new_n19364, new_n19363);
xor_3  g17016(new_n19365, n24620, n21753);
nor_4  g17017(new_n19366, n21832, n5211);
nor_4  g17018(new_n19367_1, new_n18622, new_n19366);
not_3  g17019(new_n19368, new_n19367_1);
nand_4 g17020(new_n19369, new_n19368, new_n19365);
nand_4 g17021(new_n19370, new_n19369, new_n19364);
nand_4 g17022(new_n19371, new_n19370, new_n19362);
nand_4 g17023(new_n19372, new_n19371, new_n19361_1);
nand_4 g17024(new_n19373, new_n19372, new_n19359);
nand_4 g17025(new_n19374, new_n19373, new_n19358);
nand_4 g17026(new_n19375, new_n19374, new_n19356);
nand_4 g17027(new_n19376, new_n19375, new_n19355);
nor_4  g17028(new_n19377, new_n19376, new_n19354_1);
nand_4 g17029(new_n19378, new_n19376, new_n19354_1);
not_3  g17030(new_n19379, new_n19378);
nor_4  g17031(new_n19380, new_n19379, new_n19377);
not_3  g17032(new_n19381, new_n19380);
nor_4  g17033(new_n19382, new_n19381, new_n19353);
nor_4  g17034(new_n19383, new_n19380, n3324);
nor_4  g17035(new_n19384, new_n19383, new_n19382);
not_3  g17036(new_n19385_1, n17911);
xnor_3 g17037(new_n19386, new_n19374, new_n19356);
nand_4 g17038(new_n19387, new_n19386, new_n19385_1);
xnor_3 g17039(new_n19388, new_n19386, n17911);
not_3  g17040(new_n19389_1, n21997);
xnor_3 g17041(new_n19390, new_n19372, new_n19359);
nand_4 g17042(new_n19391, new_n19390, new_n19389_1);
not_3  g17043(new_n19392, new_n19390);
nor_4  g17044(new_n19393, new_n19392, n21997);
nor_4  g17045(new_n19394, new_n19390, new_n19389_1);
nor_4  g17046(new_n19395, new_n19394, new_n19393);
xnor_3 g17047(new_n19396, new_n19370, new_n19362);
nand_4 g17048(new_n19397, new_n19396, new_n10137);
not_3  g17049(new_n19398, new_n19396);
nor_4  g17050(new_n19399, new_n19398, n25119);
nor_4  g17051(new_n19400, new_n19396, new_n10137);
nor_4  g17052(new_n19401_1, new_n19400, new_n19399);
xnor_3 g17053(new_n19402, new_n19368, new_n19365);
nor_4  g17054(new_n19403, new_n19402, new_n10139);
nand_4 g17055(new_n19404, new_n18624, new_n10143);
nand_4 g17056(new_n19405, new_n18638, new_n18627);
nand_4 g17057(new_n19406, new_n19405, new_n19404);
xnor_3 g17058(new_n19407, new_n19402, new_n10139);
nor_4  g17059(new_n19408, new_n19407, new_n19406);
nor_4  g17060(new_n19409, new_n19408, new_n19403);
nand_4 g17061(new_n19410, new_n19409, new_n19401_1);
nand_4 g17062(new_n19411, new_n19410, new_n19397);
nand_4 g17063(new_n19412, new_n19411, new_n19395);
nand_4 g17064(new_n19413, new_n19412, new_n19391);
nand_4 g17065(new_n19414_1, new_n19413, new_n19388);
nand_4 g17066(new_n19415, new_n19414_1, new_n19387);
xnor_3 g17067(new_n19416, new_n19415, new_n19384);
not_3  g17068(new_n19417, n13419);
not_3  g17069(new_n19418, n5101);
xor_3  g17070(new_n19419, n6659, new_n19418);
not_3  g17071(new_n19420, n23250);
nor_4  g17072(new_n19421, new_n19420, n16507);
not_3  g17073(new_n19422, n16507);
xor_3  g17074(new_n19423, n23250, new_n19422);
not_3  g17075(new_n19424_1, new_n19423);
not_3  g17076(new_n19425, n11455);
or_4   g17077(new_n19426, n22470, new_n19425);
xor_3  g17078(new_n19427, n22470, new_n19425);
nand_4 g17079(new_n19428, new_n3275, n3945);
not_3  g17080(new_n19429, n3945);
xor_3  g17081(new_n19430, n19116, new_n19429);
not_3  g17082(new_n19431, n6861);
nand_4 g17083(new_n19432, new_n19431, n5255);
not_3  g17084(new_n19433, n5255);
xor_3  g17085(new_n19434, n6861, new_n19433);
nor_4  g17086(new_n19435, new_n5941, n19357);
not_3  g17087(new_n19436, new_n19435);
xor_3  g17088(new_n19437, n21649, n19357);
not_3  g17089(new_n19438, new_n19437);
nor_4  g17090(new_n19439, new_n5945, n2328);
not_3  g17091(new_n19440, new_n19439);
nor_4  g17092(new_n19441, new_n5826, new_n5817);
not_3  g17093(new_n19442, n2328);
nor_4  g17094(new_n19443, n18274, new_n19442);
nor_4  g17095(new_n19444, new_n19443, new_n19439);
nand_4 g17096(new_n19445, new_n19444, new_n19441);
nand_4 g17097(new_n19446, new_n19445, new_n19440);
nand_4 g17098(new_n19447, new_n19446, new_n19438);
nand_4 g17099(new_n19448, new_n19447, new_n19436);
nand_4 g17100(new_n19449, new_n19448, new_n19434);
nand_4 g17101(new_n19450_1, new_n19449, new_n19432);
nand_4 g17102(new_n19451, new_n19450_1, new_n19430);
nand_4 g17103(new_n19452, new_n19451, new_n19428);
nand_4 g17104(new_n19453, new_n19452, new_n19427);
nand_4 g17105(new_n19454_1, new_n19453, new_n19426);
not_3  g17106(new_n19455, new_n19454_1);
nor_4  g17107(new_n19456, new_n19455, new_n19424_1);
nor_4  g17108(new_n19457, new_n19456, new_n19421);
not_3  g17109(new_n19458_1, new_n19457);
nor_4  g17110(new_n19459, new_n19458_1, new_n19419);
not_3  g17111(new_n19460, new_n19419);
nor_4  g17112(new_n19461, new_n19457, new_n19460);
nor_4  g17113(new_n19462, new_n19461, new_n19459);
not_3  g17114(new_n19463, new_n19462);
nor_4  g17115(new_n19464, new_n19463, new_n19417);
nor_4  g17116(new_n19465, new_n19462, n13419);
nor_4  g17117(new_n19466, new_n19465, new_n19464);
nor_4  g17118(new_n19467_1, new_n19454_1, new_n19423);
nor_4  g17119(new_n19468, new_n19467_1, new_n19456);
nor_4  g17120(new_n19469, new_n19468, n4967);
not_3  g17121(new_n19470, new_n19469);
not_3  g17122(new_n19471, n4967);
nor_4  g17123(new_n19472_1, new_n19468, new_n19471);
not_3  g17124(new_n19473, new_n19468);
nor_4  g17125(new_n19474, new_n19473, n4967);
nor_4  g17126(new_n19475, new_n19474, new_n19472_1);
not_3  g17127(new_n19476, new_n19475);
xnor_3 g17128(new_n19477_1, new_n19452, new_n19427);
not_3  g17129(new_n19478, new_n19477_1);
nor_4  g17130(new_n19479, new_n19478, n15602);
not_3  g17131(new_n19480, new_n19479);
not_3  g17132(new_n19481, n8694);
xnor_3 g17133(new_n19482, new_n19450_1, new_n19430);
nor_4  g17134(new_n19483, new_n19482, new_n19481);
xnor_3 g17135(new_n19484, new_n19448, new_n19434);
not_3  g17136(new_n19485, new_n19484);
nor_4  g17137(new_n19486, new_n19485, n12380);
not_3  g17138(new_n19487, new_n19486);
not_3  g17139(new_n19488, n12380);
nor_4  g17140(new_n19489, new_n19484, new_n19488);
nor_4  g17141(new_n19490, new_n19489, new_n19486);
xnor_3 g17142(new_n19491, new_n19446, new_n19437);
nor_4  g17143(new_n19492, new_n19491, n8943);
xnor_3 g17144(new_n19493, new_n19491, n8943);
not_3  g17145(new_n19494_1, new_n19444);
xnor_3 g17146(new_n19495, new_n19494_1, new_n19441);
nand_4 g17147(new_n19496_1, new_n19495, n8255);
not_3  g17148(new_n19497, new_n19496_1);
nor_4  g17149(new_n19498, new_n5833_1, new_n5815);
nand_4 g17150(new_n19499, new_n5831, n11184);
not_3  g17151(new_n19500, new_n19499);
nor_4  g17152(new_n19501, new_n19500, new_n19498);
xnor_3 g17153(new_n19502, new_n19495, n8255);
nor_4  g17154(new_n19503, new_n19502, new_n19501);
nor_4  g17155(new_n19504, new_n19503, new_n19497);
not_3  g17156(new_n19505, new_n19504);
nor_4  g17157(new_n19506, new_n19505, new_n19493);
nor_4  g17158(new_n19507, new_n19506, new_n19492);
not_3  g17159(new_n19508, new_n19507);
nand_4 g17160(new_n19509, new_n19508, new_n19490);
nand_4 g17161(new_n19510, new_n19509, new_n19487);
not_3  g17162(new_n19511, new_n19482);
nor_4  g17163(new_n19512, new_n19511, n8694);
nor_4  g17164(new_n19513, new_n19512, new_n19483);
not_3  g17165(new_n19514_1, new_n19513);
nor_4  g17166(new_n19515_1, new_n19514_1, new_n19510);
nor_4  g17167(new_n19516, new_n19515_1, new_n19483);
not_3  g17168(new_n19517, n15602);
xnor_3 g17169(new_n19518, new_n19477_1, new_n19517);
not_3  g17170(new_n19519, new_n19518);
nand_4 g17171(new_n19520, new_n19519, new_n19516);
nand_4 g17172(new_n19521, new_n19520, new_n19480);
nand_4 g17173(new_n19522, new_n19521, new_n19476);
nand_4 g17174(new_n19523_1, new_n19522, new_n19470);
nand_4 g17175(new_n19524, new_n19523_1, new_n19466);
not_3  g17176(new_n19525, new_n19524);
nor_4  g17177(new_n19526, new_n19523_1, new_n19466);
nor_4  g17178(new_n19527, new_n19526, new_n19525);
xnor_3 g17179(new_n19528, new_n19527, new_n19416);
xnor_3 g17180(new_n19529, new_n19413, new_n19388);
not_3  g17181(new_n19530, new_n19529);
xnor_3 g17182(new_n19531_1, new_n19521, new_n19475);
nand_4 g17183(new_n19532, new_n19531_1, new_n19530);
xnor_3 g17184(new_n19533, new_n19531_1, new_n19529);
xnor_3 g17185(new_n19534, new_n19411, new_n19395);
not_3  g17186(new_n19535, new_n19534);
xnor_3 g17187(new_n19536, new_n19518, new_n19516);
nand_4 g17188(new_n19537, new_n19536, new_n19535);
xnor_3 g17189(new_n19538, new_n19536, new_n19534);
xnor_3 g17190(new_n19539_1, new_n19409, new_n19401_1);
not_3  g17191(new_n19540, new_n19539_1);
xnor_3 g17192(new_n19541, new_n19514_1, new_n19510);
nand_4 g17193(new_n19542, new_n19541, new_n19540);
xnor_3 g17194(new_n19543, new_n19541, new_n19539_1);
not_3  g17195(new_n19544, new_n19490);
xnor_3 g17196(new_n19545, new_n19507, new_n19544);
xnor_3 g17197(new_n19546, new_n19407, new_n19406);
not_3  g17198(new_n19547, new_n19546);
nor_4  g17199(new_n19548, new_n19547, new_n19545);
not_3  g17200(new_n19549, new_n19548);
not_3  g17201(new_n19550, new_n19545);
nor_4  g17202(new_n19551, new_n19546, new_n19550);
nor_4  g17203(new_n19552, new_n19551, new_n19548);
not_3  g17204(new_n19553, n8943);
not_3  g17205(new_n19554, new_n19491);
nor_4  g17206(new_n19555, new_n19554, new_n19553);
nor_4  g17207(new_n19556, new_n19555, new_n19492);
nor_4  g17208(new_n19557, new_n19504, new_n19556);
nor_4  g17209(new_n19558, new_n19557, new_n19506);
nand_4 g17210(new_n19559, new_n19558, new_n18664);
xnor_3 g17211(new_n19560, new_n19558, new_n18639);
xnor_3 g17212(new_n19561, new_n19502, new_n19501);
nand_4 g17213(new_n19562, new_n19561, new_n18673);
xnor_3 g17214(new_n19563, new_n19561, new_n18669);
not_3  g17215(new_n19564, new_n5836);
nand_4 g17216(new_n19565, new_n5857, new_n5839);
nand_4 g17217(new_n19566, new_n19565, new_n19564);
nand_4 g17218(new_n19567, new_n19566, new_n19563);
nand_4 g17219(new_n19568, new_n19567, new_n19562);
nand_4 g17220(new_n19569, new_n19568, new_n19560);
nand_4 g17221(new_n19570_1, new_n19569, new_n19559);
nand_4 g17222(new_n19571, new_n19570_1, new_n19552);
nand_4 g17223(new_n19572, new_n19571, new_n19549);
nand_4 g17224(new_n19573, new_n19572, new_n19543);
nand_4 g17225(new_n19574, new_n19573, new_n19542);
nand_4 g17226(new_n19575_1, new_n19574, new_n19538);
nand_4 g17227(new_n19576, new_n19575_1, new_n19537);
nand_4 g17228(new_n19577, new_n19576, new_n19533);
nand_4 g17229(new_n19578, new_n19577, new_n19532);
not_3  g17230(new_n19579, new_n19578);
xor_3  g17231(n3649, new_n19579, new_n19528);
nor_4  g17232(new_n19581, n26625, n14230);
nand_4 g17233(new_n19582, new_n19581, new_n13931);
nor_4  g17234(new_n19583, new_n19582, n11566);
nand_4 g17235(new_n19584_1, new_n19583, new_n13921);
nor_4  g17236(new_n19585, new_n19584_1, n26565);
xor_3  g17237(new_n19586, new_n19585, new_n13723);
xnor_3 g17238(new_n19587, new_n19586, n26191);
not_3  g17239(new_n19588, new_n19584_1);
xor_3  g17240(new_n19589, new_n19588, new_n13915);
nand_4 g17241(new_n19590, new_n19589, new_n13825);
xnor_3 g17242(new_n19591, new_n19589, n26512);
xor_3  g17243(new_n19592, new_n19583, new_n13921);
nand_4 g17244(new_n19593, new_n19592, new_n11441);
xnor_3 g17245(new_n19594, new_n19592, n19575);
not_3  g17246(new_n19595, n15378);
nand_4 g17247(new_n19596, new_n19582, n11566);
not_3  g17248(new_n19597, new_n19596);
nor_4  g17249(new_n19598, new_n19597, new_n19583);
nand_4 g17250(new_n19599, new_n19598, new_n19595);
xnor_3 g17251(new_n19600, new_n19598, n15378);
not_3  g17252(new_n19601, new_n19582);
nor_4  g17253(new_n19602_1, new_n19581, new_n13931);
nor_4  g17254(new_n19603, new_n19602_1, new_n19601);
not_3  g17255(new_n19604, new_n19603);
nor_4  g17256(new_n19605, new_n19604, n17095);
not_3  g17257(new_n19606, new_n19605);
nand_4 g17258(new_n19607, new_n13935, new_n7729);
nand_4 g17259(new_n19608_1, n26625, n14230);
nand_4 g17260(new_n19609, new_n19608_1, new_n19607);
not_3  g17261(new_n19610, new_n19609);
nor_4  g17262(new_n19611, new_n19610, new_n11497);
nor_4  g17263(new_n19612, new_n8491, n14230);
not_3  g17264(new_n19613, new_n19612);
xnor_3 g17265(new_n19614, new_n19609, n22591);
nor_4  g17266(new_n19615, new_n19614, new_n19613);
nor_4  g17267(new_n19616, new_n19615, new_n19611);
nor_4  g17268(new_n19617_1, new_n19603, new_n11442);
nor_4  g17269(new_n19618_1, new_n19617_1, new_n19605);
nand_4 g17270(new_n19619, new_n19618_1, new_n19616);
nand_4 g17271(new_n19620, new_n19619, new_n19606);
nand_4 g17272(new_n19621, new_n19620, new_n19600);
nand_4 g17273(new_n19622, new_n19621, new_n19599);
nand_4 g17274(new_n19623_1, new_n19622, new_n19594);
nand_4 g17275(new_n19624, new_n19623_1, new_n19593);
nand_4 g17276(new_n19625, new_n19624, new_n19591);
nand_4 g17277(new_n19626, new_n19625, new_n19590);
xnor_3 g17278(new_n19627, new_n19626, new_n19587);
xnor_3 g17279(new_n19628, new_n19627, new_n17576);
xnor_3 g17280(new_n19629, new_n19624, new_n19591);
nor_4  g17281(new_n19630, new_n19629, n17302);
not_3  g17282(new_n19631, new_n19630);
not_3  g17283(new_n19632, n17302);
xnor_3 g17284(new_n19633, new_n19629, new_n19632);
xnor_3 g17285(new_n19634, new_n19592, new_n11441);
xnor_3 g17286(new_n19635, new_n19622, new_n19634);
nor_4  g17287(new_n19636, new_n19635, new_n17584);
xnor_3 g17288(new_n19637, new_n19622, new_n19594);
xnor_3 g17289(new_n19638, new_n19637, n2013);
xnor_3 g17290(new_n19639, new_n19620, new_n19600);
not_3  g17291(new_n19640, new_n19639);
nor_4  g17292(new_n19641_1, new_n19640, new_n17603);
nor_4  g17293(new_n19642, new_n19639, n23755);
nor_4  g17294(new_n19643, new_n19642, new_n19641_1);
not_3  g17295(new_n19644, new_n19643);
not_3  g17296(new_n19645, new_n19618_1);
xnor_3 g17297(new_n19646, new_n19645, new_n19616);
nor_4  g17298(new_n19647, new_n19646, new_n17592_1);
not_3  g17299(new_n19648_1, new_n19646);
nor_4  g17300(new_n19649, new_n19648_1, n19163);
nor_4  g17301(new_n19650, new_n19649, new_n19647);
not_3  g17302(new_n19651, new_n19650);
xnor_3 g17303(new_n19652_1, new_n19614, new_n19612);
not_3  g17304(new_n19653, new_n19652_1);
nor_4  g17305(new_n19654, new_n19653, new_n17595);
nor_4  g17306(new_n19655, new_n19652_1, n22358);
xor_3  g17307(new_n19656, n26167, new_n7729);
nand_4 g17308(new_n19657, new_n19656, n9646);
nor_4  g17309(new_n19658, new_n19657, new_n19655);
nor_4  g17310(new_n19659, new_n19658, new_n19654);
nor_4  g17311(new_n19660, new_n19659, new_n19651);
nor_4  g17312(new_n19661, new_n19660, new_n19647);
nor_4  g17313(new_n19662, new_n19661, new_n19644);
nor_4  g17314(new_n19663, new_n19662, new_n19641_1);
nor_4  g17315(new_n19664_1, new_n19663, new_n19638);
nor_4  g17316(new_n19665, new_n19664_1, new_n19636);
nand_4 g17317(new_n19666, new_n19665, new_n19633);
nand_4 g17318(new_n19667, new_n19666, new_n19631);
xnor_3 g17319(new_n19668, new_n19667, new_n19628);
xnor_3 g17320(new_n19669, new_n19668, new_n8143);
xnor_3 g17321(new_n19670, new_n19629, n17302);
not_3  g17322(new_n19671, new_n19636);
nor_4  g17323(new_n19672, new_n19637, n2013);
nor_4  g17324(new_n19673, new_n19672, new_n19636);
not_3  g17325(new_n19674, new_n19663);
nand_4 g17326(new_n19675, new_n19674, new_n19673);
nand_4 g17327(new_n19676, new_n19675, new_n19671);
xnor_3 g17328(new_n19677, new_n19676, new_n19670);
not_3  g17329(new_n19678, new_n19677);
nor_4  g17330(new_n19679, new_n19678, new_n8148_1);
not_3  g17331(new_n19680_1, new_n19679);
nor_4  g17332(new_n19681, new_n19677, new_n8150);
nor_4  g17333(new_n19682, new_n19681, new_n19679);
nor_4  g17334(new_n19683, new_n19674, new_n19673);
nor_4  g17335(new_n19684, new_n19683, new_n19664_1);
nand_4 g17336(new_n19685, new_n19684, new_n8155);
xnor_3 g17337(new_n19686, new_n19684, new_n8152);
not_3  g17338(new_n19687, new_n19661);
nor_4  g17339(new_n19688, new_n19687, new_n19643);
nor_4  g17340(new_n19689, new_n19688, new_n19662);
nand_4 g17341(new_n19690, new_n19689, new_n8160);
xnor_3 g17342(new_n19691, new_n19689, new_n8161);
xnor_3 g17343(new_n19692, new_n19659, new_n19651);
nor_4  g17344(new_n19693, new_n19692, new_n8169);
not_3  g17345(new_n19694, new_n19693);
not_3  g17346(new_n19695, new_n19692);
nor_4  g17347(new_n19696, new_n19695, new_n8168);
nor_4  g17348(new_n19697, new_n19696, new_n19693);
not_3  g17349(new_n19698, new_n19657);
nor_4  g17350(new_n19699, new_n19655, new_n19654);
xnor_3 g17351(new_n19700, new_n19699, new_n19698);
nor_4  g17352(new_n19701_1, new_n19700, new_n8175);
not_3  g17353(new_n19702, new_n19701_1);
not_3  g17354(new_n19703, new_n19656);
xor_3  g17355(new_n19704, new_n19703, n9646);
nand_4 g17356(new_n19705, new_n19704, new_n8177);
not_3  g17357(new_n19706, new_n8175);
not_3  g17358(new_n19707, new_n19700);
nor_4  g17359(new_n19708, new_n19707, new_n19706);
nor_4  g17360(new_n19709, new_n19708, new_n19701_1);
nand_4 g17361(new_n19710, new_n19709, new_n19705);
nand_4 g17362(new_n19711, new_n19710, new_n19702);
nand_4 g17363(new_n19712, new_n19711, new_n19697);
nand_4 g17364(new_n19713, new_n19712, new_n19694);
nand_4 g17365(new_n19714, new_n19713, new_n19691);
nand_4 g17366(new_n19715, new_n19714, new_n19690);
nand_4 g17367(new_n19716, new_n19715, new_n19686);
nand_4 g17368(new_n19717, new_n19716, new_n19685);
nand_4 g17369(new_n19718, new_n19717, new_n19682);
nand_4 g17370(new_n19719, new_n19718, new_n19680_1);
xnor_3 g17371(n3665, new_n19719, new_n19669);
xor_3  g17372(n3679, new_n6782, new_n6779);
nor_4  g17373(new_n19722, n16521, n7139);
nand_4 g17374(new_n19723, new_n19722, new_n3852);
nor_4  g17375(new_n19724, new_n19723, n604);
not_3  g17376(new_n19725, new_n19724);
nor_4  g17377(new_n19726, new_n19725, n4913);
not_3  g17378(new_n19727, new_n19726);
nor_4  g17379(new_n19728, new_n19727, n9172);
not_3  g17380(new_n19729, new_n19728);
nor_4  g17381(new_n19730, new_n19729, n442);
not_3  g17382(new_n19731, new_n19730);
nor_4  g17383(new_n19732, new_n19731, n13719);
xor_3  g17384(new_n19733, new_n19732, new_n3828_1);
not_3  g17385(new_n19734, new_n19733);
xnor_3 g17386(new_n19735, new_n19734, new_n6930);
xor_3  g17387(new_n19736_1, new_n19730, new_n3831);
not_3  g17388(new_n19737, new_n19736_1);
nor_4  g17389(new_n19738, new_n19737, new_n6937);
xnor_3 g17390(new_n19739, new_n19737, new_n6937);
xor_3  g17391(new_n19740, new_n19728, new_n3836);
nor_4  g17392(new_n19741, new_n19740, new_n6947);
not_3  g17393(new_n19742, new_n19741);
not_3  g17394(new_n19743, new_n19740);
nor_4  g17395(new_n19744, new_n19743, new_n6945);
nor_4  g17396(new_n19745, new_n19744, new_n19741);
xor_3  g17397(new_n19746, new_n19726, new_n3840);
nor_4  g17398(new_n19747, new_n19746, new_n6955);
not_3  g17399(new_n19748, new_n19747);
not_3  g17400(new_n19749_1, new_n19746);
nor_4  g17401(new_n19750, new_n19749_1, new_n6952);
nor_4  g17402(new_n19751, new_n19750, new_n19747);
xor_3  g17403(new_n19752, new_n19724, new_n3842_1);
nor_4  g17404(new_n19753, new_n19752, new_n6963);
not_3  g17405(new_n19754, new_n19753);
not_3  g17406(new_n19755, new_n19752);
nor_4  g17407(new_n19756_1, new_n19755, new_n6960);
nor_4  g17408(new_n19757, new_n19756_1, new_n19753);
xor_3  g17409(new_n19758, new_n19723, new_n3846);
not_3  g17410(new_n19759, new_n19758);
nor_4  g17411(new_n19760, new_n19759, new_n6974);
not_3  g17412(new_n19761, new_n19760);
nor_4  g17413(new_n19762, new_n19758, new_n6971_1);
nor_4  g17414(new_n19763, new_n19762, new_n19760);
xor_3  g17415(new_n19764, new_n19722, n16824);
nand_4 g17416(new_n19765, new_n19764, new_n6982);
not_3  g17417(new_n19766, new_n19765);
nor_4  g17418(new_n19767_1, new_n19764, new_n6982);
nor_4  g17419(new_n19768, new_n19767_1, new_n19766);
not_3  g17420(new_n19769, new_n6985_1);
nand_4 g17421(new_n19770_1, new_n19722, new_n19769);
not_3  g17422(new_n19771, new_n19770_1);
nor_4  g17423(new_n19772, new_n19769, n7139);
xnor_3 g17424(new_n19773, new_n19772, n16521);
nor_4  g17425(new_n19774, new_n19773, new_n6993);
nor_4  g17426(new_n19775, new_n19774, new_n19771);
not_3  g17427(new_n19776, new_n19775);
nand_4 g17428(new_n19777, new_n19776, new_n19768);
nand_4 g17429(new_n19778, new_n19777, new_n19765);
nand_4 g17430(new_n19779, new_n19778, new_n19763);
nand_4 g17431(new_n19780_1, new_n19779, new_n19761);
nand_4 g17432(new_n19781, new_n19780_1, new_n19757);
nand_4 g17433(new_n19782, new_n19781, new_n19754);
nand_4 g17434(new_n19783, new_n19782, new_n19751);
nand_4 g17435(new_n19784, new_n19783, new_n19748);
nand_4 g17436(new_n19785, new_n19784, new_n19745);
nand_4 g17437(new_n19786, new_n19785, new_n19742);
nor_4  g17438(new_n19787, new_n19786, new_n19739);
nor_4  g17439(new_n19788, new_n19787, new_n19738);
not_3  g17440(new_n19789_1, new_n19788);
xnor_3 g17441(new_n19790, new_n19789_1, new_n19735);
xnor_3 g17442(new_n19791, new_n7072, n2858);
nor_4  g17443(new_n19792_1, new_n7078, new_n5602);
xnor_3 g17444(new_n19793, new_n7077, new_n5602);
nand_4 g17445(new_n19794, new_n7081, n24327);
nand_4 g17446(new_n19795, new_n10134, new_n10106);
nand_4 g17447(new_n19796, new_n19795, new_n19794);
nand_4 g17448(new_n19797, new_n19796, new_n19793);
not_3  g17449(new_n19798_1, new_n19797);
nor_4  g17450(new_n19799, new_n19798_1, new_n19792_1);
xnor_3 g17451(new_n19800, new_n19799, new_n19791);
xnor_3 g17452(new_n19801, new_n19800, new_n19790);
xnor_3 g17453(new_n19802, new_n19796, new_n19793);
nand_4 g17454(new_n19803_1, new_n19786, new_n19739);
not_3  g17455(new_n19804, new_n19803_1);
nor_4  g17456(new_n19805, new_n19804, new_n19787);
not_3  g17457(new_n19806, new_n19805);
nand_4 g17458(new_n19807, new_n19806, new_n19802);
xnor_3 g17459(new_n19808, new_n19805, new_n19802);
not_3  g17460(new_n19809, new_n19785);
nor_4  g17461(new_n19810, new_n19784, new_n19745);
nor_4  g17462(new_n19811, new_n19810, new_n19809);
nand_4 g17463(new_n19812, new_n19811, new_n10136);
xnor_3 g17464(new_n19813, new_n19811, new_n10135);
not_3  g17465(new_n19814, new_n19783);
nor_4  g17466(new_n19815, new_n19782, new_n19751);
nor_4  g17467(new_n19816, new_n19815, new_n19814);
nand_4 g17468(new_n19817, new_n19816, new_n10173);
xnor_3 g17469(new_n19818, new_n19816, new_n10174);
not_3  g17470(new_n19819, new_n19757);
xnor_3 g17471(new_n19820, new_n19780_1, new_n19819);
nand_4 g17472(new_n19821, new_n19820, new_n10181);
xnor_3 g17473(new_n19822, new_n19820, new_n10182);
xnor_3 g17474(new_n19823, new_n19778, new_n19763);
not_3  g17475(new_n19824, new_n19823);
nand_4 g17476(new_n19825, new_n19824, new_n10188);
not_3  g17477(new_n19826, new_n19825);
nor_4  g17478(new_n19827, new_n19824, new_n10188);
nor_4  g17479(new_n19828, new_n19827, new_n19826);
xnor_3 g17480(new_n19829, new_n19776, new_n19768);
not_3  g17481(new_n19830, new_n19829);
nor_4  g17482(new_n19831, new_n19830, new_n10196);
xnor_3 g17483(new_n19832, new_n19830, new_n10196);
not_3  g17484(new_n19833, new_n10203);
xor_3  g17485(new_n19834, new_n19773, new_n6993);
nand_4 g17486(new_n19835, new_n19834, new_n19833);
xor_3  g17487(new_n19836, new_n6985_1, new_n3858);
nand_4 g17488(new_n19837, new_n19836, new_n10207);
xnor_3 g17489(new_n19838, new_n19834, new_n10203);
nand_4 g17490(new_n19839, new_n19838, new_n19837);
nand_4 g17491(new_n19840, new_n19839, new_n19835);
nor_4  g17492(new_n19841, new_n19840, new_n19832);
nor_4  g17493(new_n19842, new_n19841, new_n19831);
nand_4 g17494(new_n19843, new_n19842, new_n19828);
nand_4 g17495(new_n19844, new_n19843, new_n19825);
nand_4 g17496(new_n19845, new_n19844, new_n19822);
nand_4 g17497(new_n19846, new_n19845, new_n19821);
nand_4 g17498(new_n19847, new_n19846, new_n19818);
nand_4 g17499(new_n19848, new_n19847, new_n19817);
nand_4 g17500(new_n19849, new_n19848, new_n19813);
nand_4 g17501(new_n19850, new_n19849, new_n19812);
nand_4 g17502(new_n19851, new_n19850, new_n19808);
nand_4 g17503(new_n19852, new_n19851, new_n19807);
xor_3  g17504(n3725, new_n19852, new_n19801);
not_3  g17505(new_n19854, new_n18003);
nor_4  g17506(new_n19855, n11220, n3425);
nor_4  g17507(new_n19856, new_n15733, new_n15731);
nor_4  g17508(new_n19857, new_n19856, new_n19855);
nor_4  g17509(new_n19858, n7335, n2160);
not_3  g17510(new_n19859, new_n15724);
nor_4  g17511(new_n19860, new_n15728, new_n19859);
nor_4  g17512(new_n19861, new_n19860, new_n19858);
not_3  g17513(new_n19862, new_n19861);
nor_4  g17514(new_n19863, new_n19862, new_n19857);
not_3  g17515(new_n19864, new_n19857);
nor_4  g17516(new_n19865, new_n19861, new_n19864);
nor_4  g17517(new_n19866, new_n19865, new_n19863);
nor_4  g17518(new_n19867, new_n15734, new_n15729);
not_3  g17519(new_n19868, new_n19867);
not_3  g17520(new_n19869, new_n15735);
nand_4 g17521(new_n19870, new_n15738, new_n19869);
nand_4 g17522(new_n19871, new_n19870, new_n19868);
xnor_3 g17523(new_n19872, new_n19871, new_n19866);
nor_4  g17524(new_n19873_1, new_n19872, new_n19854);
not_3  g17525(new_n19874, new_n19871);
xnor_3 g17526(new_n19875, new_n19874, new_n19866);
nor_4  g17527(new_n19876, new_n19875, new_n18003);
nor_4  g17528(new_n19877, new_n19876, new_n19873_1);
xnor_3 g17529(new_n19878, new_n15738, new_n19869);
nand_4 g17530(new_n19879, new_n18007, new_n19878);
xnor_3 g17531(new_n19880, new_n18009, new_n19878);
nor_4  g17532(new_n19881, new_n18020, new_n6238);
xnor_3 g17533(new_n19882, new_n18020, new_n6238);
xnor_3 g17534(new_n19883, new_n6235, new_n6164);
nor_4  g17535(new_n19884, new_n18024, new_n19883);
not_3  g17536(new_n19885, new_n6253);
nand_4 g17537(new_n19886, new_n18027, new_n19885);
xnor_3 g17538(new_n19887, new_n18027, new_n6253);
not_3  g17539(new_n19888, new_n6259);
nand_4 g17540(new_n19889, new_n17924, new_n19888);
xnor_3 g17541(new_n19890, new_n17924, new_n6259);
nor_4  g17542(new_n19891, new_n6265, new_n4779);
xnor_3 g17543(new_n19892, new_n6265, new_n4779);
nor_4  g17544(new_n19893, new_n6271_1, new_n4788);
not_3  g17545(new_n19894, new_n19893);
nor_4  g17546(new_n19895, new_n6270, new_n4789);
nor_4  g17547(new_n19896, new_n19895, new_n19893);
nor_4  g17548(new_n19897, new_n6279, new_n4795);
xnor_3 g17549(new_n19898, new_n6279, new_n4795);
nor_4  g17550(new_n19899, new_n6288, new_n4799);
nor_4  g17551(new_n19900, new_n6289, new_n4771);
nor_4  g17552(new_n19901, new_n6299, new_n4802);
not_3  g17553(new_n19902, new_n19901);
nor_4  g17554(new_n19903, new_n19902, new_n19900);
nor_4  g17555(new_n19904, new_n19903, new_n19899);
nor_4  g17556(new_n19905_1, new_n19904, new_n19898);
nor_4  g17557(new_n19906, new_n19905_1, new_n19897);
nand_4 g17558(new_n19907, new_n19906, new_n19896);
nand_4 g17559(new_n19908, new_n19907, new_n19894);
nor_4  g17560(new_n19909_1, new_n19908, new_n19892);
nor_4  g17561(new_n19910, new_n19909_1, new_n19891);
nand_4 g17562(new_n19911_1, new_n19910, new_n19890);
nand_4 g17563(new_n19912, new_n19911_1, new_n19889);
nand_4 g17564(new_n19913, new_n19912, new_n19887);
nand_4 g17565(new_n19914, new_n19913, new_n19886);
xnor_3 g17566(new_n19915, new_n18036, new_n6242);
nor_4  g17567(new_n19916_1, new_n19915, new_n19914);
nor_4  g17568(new_n19917, new_n19916_1, new_n19884);
nor_4  g17569(new_n19918, new_n19917, new_n19882);
nor_4  g17570(new_n19919, new_n19918, new_n19881);
nand_4 g17571(new_n19920, new_n19919, new_n19880);
nand_4 g17572(new_n19921, new_n19920, new_n19879);
xnor_3 g17573(n3733, new_n19921, new_n19877);
xnor_3 g17574(new_n19923_1, new_n12925, n24937);
nand_4 g17575(new_n19924, new_n12918, n5098);
nor_4  g17576(new_n19925, new_n12917_1, new_n18792);
nor_4  g17577(new_n19926, new_n12918, n5098);
nor_4  g17578(new_n19927, new_n19926, new_n19925);
not_3  g17579(new_n19928, new_n12908);
nand_4 g17580(new_n19929, new_n19928, n3030);
nand_4 g17581(new_n19930_1, new_n18710, new_n18694);
nand_4 g17582(new_n19931, new_n19930_1, new_n19929);
nand_4 g17583(new_n19932, new_n19931, new_n19927);
nand_4 g17584(new_n19933, new_n19932, new_n19924);
xnor_3 g17585(new_n19934, new_n19933, new_n19923_1);
xnor_3 g17586(new_n19935, new_n19934, new_n12040);
not_3  g17587(new_n19936, new_n19935);
nor_4  g17588(new_n19937, new_n11997, new_n11955);
nor_4  g17589(new_n19938, new_n19937, new_n11999);
xnor_3 g17590(new_n19939, new_n19931, new_n19927);
not_3  g17591(new_n19940, new_n19939);
nor_4  g17592(new_n19941_1, new_n19940, new_n19938);
not_3  g17593(new_n19942, new_n19941_1);
nor_4  g17594(new_n19943, new_n19939, new_n12045);
nor_4  g17595(new_n19944, new_n19943, new_n19941_1);
nor_4  g17596(new_n19945, new_n18712, new_n12053);
not_3  g17597(new_n19946, new_n19945);
not_3  g17598(new_n19947, new_n18712);
nor_4  g17599(new_n19948, new_n19947, new_n12050);
nor_4  g17600(new_n19949, new_n19948, new_n19945);
xnor_3 g17601(new_n19950, new_n18714, new_n12057);
xnor_3 g17602(new_n19951, new_n18722, new_n12062);
nor_4  g17603(new_n19952, new_n18728, new_n19951);
nor_4  g17604(new_n19953, new_n19952, new_n18723);
nor_4  g17605(new_n19954, new_n19953, new_n19950);
nor_4  g17606(new_n19955, new_n19954, new_n18715);
nand_4 g17607(new_n19956, new_n19955, new_n19949);
nand_4 g17608(new_n19957, new_n19956, new_n19946);
nand_4 g17609(new_n19958, new_n19957, new_n19944);
nand_4 g17610(new_n19959, new_n19958, new_n19942);
xor_3  g17611(n3755, new_n19959, new_n19936);
not_3  g17612(new_n19961, new_n10812);
xor_3  g17613(n3758, new_n10855, new_n19961);
not_3  g17614(new_n19963, n655);
not_3  g17615(new_n19964, new_n19089);
nor_4  g17616(new_n19965, new_n19964, n18145);
nand_4 g17617(new_n19966, new_n19965, new_n19963);
nor_4  g17618(new_n19967, new_n19966, n19033);
not_3  g17619(new_n19968_1, new_n19967);
xor_3  g17620(new_n19969, new_n19968_1, n2570);
not_3  g17621(new_n19970, new_n19969);
xor_3  g17622(new_n19971, new_n19970, n14692);
not_3  g17623(new_n19972, new_n19971);
not_3  g17624(new_n19973, n19033);
not_3  g17625(new_n19974, new_n19966);
xor_3  g17626(new_n19975, new_n19974, new_n19973);
nor_4  g17627(new_n19976, new_n19975, new_n12320);
not_3  g17628(new_n19977, new_n19976);
not_3  g17629(new_n19978, new_n19975);
xor_3  g17630(new_n19979, new_n19978, n4100);
not_3  g17631(new_n19980, n21957);
xor_3  g17632(new_n19981, new_n19965, new_n19963);
nor_4  g17633(new_n19982, new_n19981, new_n19980);
not_3  g17634(new_n19983, new_n19982);
not_3  g17635(new_n19984, new_n19981);
xor_3  g17636(new_n19985, new_n19984, n21957);
nor_4  g17637(new_n19986, new_n19090, new_n12328);
nor_4  g17638(new_n19987, new_n19141_1, new_n19986);
not_3  g17639(new_n19988_1, new_n19987);
nand_4 g17640(new_n19989, new_n19988_1, new_n19985);
nand_4 g17641(new_n19990, new_n19989, new_n19983);
nand_4 g17642(new_n19991, new_n19990, new_n19979);
nand_4 g17643(new_n19992, new_n19991, new_n19977);
xnor_3 g17644(new_n19993, new_n19992, new_n19972);
not_3  g17645(new_n19994, new_n19993);
nor_4  g17646(new_n19995, new_n19994, new_n14415);
xnor_3 g17647(new_n19996, new_n19993, new_n14412_1);
not_3  g17648(new_n19997, new_n19979);
xnor_3 g17649(new_n19998, new_n19990, new_n19997);
nand_4 g17650(new_n19999, new_n19998, new_n8074);
not_3  g17651(new_n20000, new_n19999);
xnor_3 g17652(new_n20001, new_n19998, new_n8074);
xnor_3 g17653(new_n20002, new_n19987, new_n19985);
nand_4 g17654(new_n20003, new_n20002, new_n8077);
xnor_3 g17655(new_n20004_1, new_n20002, new_n8078);
nand_4 g17656(new_n20005, new_n19143, new_n8084);
nand_4 g17657(new_n20006, new_n19179, new_n19144_1);
nand_4 g17658(new_n20007, new_n20006, new_n20005);
nand_4 g17659(new_n20008, new_n20007, new_n20004_1);
nand_4 g17660(new_n20009, new_n20008, new_n20003);
not_3  g17661(new_n20010, new_n20009);
nor_4  g17662(new_n20011, new_n20010, new_n20001);
nor_4  g17663(new_n20012, new_n20011, new_n20000);
nor_4  g17664(new_n20013_1, new_n20012, new_n19996);
nor_4  g17665(new_n20014, new_n20013_1, new_n19995);
nor_4  g17666(new_n20015, new_n19968_1, n2570);
nand_4 g17667(new_n20016, new_n19970, n14692);
nand_4 g17668(new_n20017_1, new_n19992, new_n19971);
nand_4 g17669(new_n20018, new_n20017_1, new_n20016);
xnor_3 g17670(new_n20019, new_n20018, new_n20015);
xnor_3 g17671(new_n20020, new_n20019, new_n14468);
xnor_3 g17672(new_n20021, new_n20020, new_n20014);
nor_4  g17673(new_n20022, new_n20021, new_n12459);
xnor_3 g17674(new_n20023, new_n20021, new_n12459);
xnor_3 g17675(new_n20024, new_n20012, new_n19996);
nor_4  g17676(new_n20025, new_n20024, new_n12465);
xnor_3 g17677(new_n20026, new_n20024, new_n12465);
not_3  g17678(new_n20027, new_n20001);
xnor_3 g17679(new_n20028, new_n20009, new_n20027);
not_3  g17680(new_n20029, new_n20028);
nand_4 g17681(new_n20030, new_n20029, new_n12470);
xnor_3 g17682(new_n20031, new_n20028, new_n12470);
xnor_3 g17683(new_n20032, new_n20007, new_n20004_1);
not_3  g17684(new_n20033_1, new_n20032);
nand_4 g17685(new_n20034, new_n20033_1, new_n12476);
xnor_3 g17686(new_n20035, new_n20032, new_n12476);
not_3  g17687(new_n20036_1, new_n19181);
nor_4  g17688(new_n20037, new_n19231, new_n19185);
nor_4  g17689(new_n20038, new_n20037, new_n20036_1);
nand_4 g17690(new_n20039, new_n20038, new_n20035);
nand_4 g17691(new_n20040_1, new_n20039, new_n20034);
nand_4 g17692(new_n20041, new_n20040_1, new_n20031);
nand_4 g17693(new_n20042, new_n20041, new_n20030);
not_3  g17694(new_n20043, new_n20042);
nor_4  g17695(new_n20044, new_n20043, new_n20026);
nor_4  g17696(new_n20045, new_n20044, new_n20025);
nor_4  g17697(new_n20046, new_n20045, new_n20023);
nor_4  g17698(new_n20047, new_n20046, new_n20022);
nand_4 g17699(new_n20048, new_n20019, new_n14468);
not_3  g17700(new_n20049, new_n20015);
nor_4  g17701(new_n20050, new_n20018, new_n20049);
not_3  g17702(new_n20051, new_n20014);
nor_4  g17703(new_n20052, new_n20019, new_n14468);
nor_4  g17704(new_n20053, new_n20052, new_n20051);
nor_4  g17705(new_n20054, new_n20053, new_n20050);
nand_4 g17706(new_n20055, new_n20054, new_n20048);
xnor_3 g17707(n3760, new_n20055, new_n20047);
not_3  g17708(new_n20057, new_n4297);
xor_3  g17709(n3781, new_n4328, new_n20057);
xnor_3 g17710(n3794, new_n16414, new_n16378);
nand_4 g17711(new_n20060, new_n13074_1, new_n5719);
nand_4 g17712(new_n20061_1, new_n20060, new_n5728);
nor_4  g17713(new_n20062, new_n20060, new_n5726);
not_3  g17714(new_n20063, new_n20062);
nand_4 g17715(new_n20064, new_n20063, new_n20061_1);
nor_4  g17716(new_n20065, new_n13073, new_n6985_1);
not_3  g17717(new_n20066, new_n20065);
nand_4 g17718(new_n20067, new_n6993, new_n6985_1);
nand_4 g17719(new_n20068, new_n19769, new_n6907);
nand_4 g17720(new_n20069_1, new_n20068, new_n20067);
nor_4  g17721(new_n20070, new_n20069_1, new_n15810);
nand_4 g17722(new_n20071, new_n20069_1, new_n15810);
not_3  g17723(new_n20072, new_n20071);
nor_4  g17724(new_n20073, new_n20072, new_n20070);
nor_4  g17725(new_n20074, new_n20073, new_n20066);
nand_4 g17726(new_n20075, new_n20073, new_n20066);
not_3  g17727(new_n20076, new_n20075);
nor_4  g17728(new_n20077_1, new_n20076, new_n20074);
xor_3  g17729(n3842, new_n20077_1, new_n20064);
not_3  g17730(new_n20079, new_n10643);
xor_3  g17731(n3850, new_n14790_1, new_n20079);
xor_3  g17732(n3869, new_n17952, new_n4832);
not_3  g17733(new_n20082, n19584);
xor_3  g17734(new_n20083, n21749, n919);
nor_4  g17735(new_n20084, n25316, n7769);
not_3  g17736(new_n20085, new_n20084);
nand_4 g17737(new_n20086_1, n21138, n20385);
nand_4 g17738(new_n20087, n25316, n7769);
not_3  g17739(new_n20088, new_n20087);
nor_4  g17740(new_n20089, new_n20088, new_n20084);
nand_4 g17741(new_n20090, new_n20089, new_n20086_1);
nand_4 g17742(new_n20091, new_n20090, new_n20085);
nor_4  g17743(new_n20092, new_n20091, new_n20083);
nand_4 g17744(new_n20093, new_n20091, new_n20083);
not_3  g17745(new_n20094, new_n20093);
nor_4  g17746(new_n20095, new_n20094, new_n20092);
xnor_3 g17747(new_n20096_1, new_n20095, new_n20082);
not_3  g17748(new_n20097, n5060);
xnor_3 g17749(new_n20098, n21138, n20385);
nand_4 g17750(new_n20099, new_n20098, n15332);
nand_4 g17751(new_n20100, new_n20099, new_n20097);
not_3  g17752(new_n20101, new_n20100);
xor_3  g17753(new_n20102, new_n20089, new_n20086_1);
xor_3  g17754(new_n20103_1, new_n20099, n5060);
nor_4  g17755(new_n20104, new_n20103_1, new_n20102);
nor_4  g17756(new_n20105, new_n20104, new_n20101);
xnor_3 g17757(new_n20106, new_n20105, new_n20096_1);
xnor_3 g17758(new_n20107, new_n20106, new_n19012);
not_3  g17759(new_n20108, new_n20107);
xnor_3 g17760(new_n20109, new_n20103_1, new_n20102);
nand_4 g17761(new_n20110, new_n20109, new_n19015);
xor_3  g17762(new_n20111, new_n20098, n15332);
not_3  g17763(new_n20112, new_n20111);
nand_4 g17764(new_n20113, new_n20112, new_n19021);
xnor_3 g17765(new_n20114, new_n20109, new_n19014);
nand_4 g17766(new_n20115, new_n20114, new_n20113);
nand_4 g17767(new_n20116, new_n20115, new_n20110);
xor_3  g17768(n3871, new_n20116, new_n20108);
xor_3  g17769(n3891, new_n19840, new_n19832);
not_3  g17770(new_n20119, new_n7433);
xor_3  g17771(new_n20120, new_n10324, n2570);
not_3  g17772(new_n20121, new_n20120);
nor_4  g17773(new_n20122, n19033, new_n10329);
xor_3  g17774(new_n20123, n19033, new_n10329);
nand_4 g17775(new_n20124, n6397, new_n19963);
xor_3  g17776(new_n20125, n6397, new_n19963);
nand_4 g17777(new_n20126_1, n19196, new_n19082);
xor_3  g17778(new_n20127, n19196, new_n19082);
not_3  g17779(new_n20128, n10712);
nand_4 g17780(new_n20129, n23586, new_n20128);
xor_3  g17781(new_n20130, n23586, new_n20128);
nor_4  g17782(new_n20131, n25126, new_n14431);
not_3  g17783(new_n20132, new_n20131);
xor_3  g17784(new_n20133, n25126, new_n14431);
nor_4  g17785(new_n20134, n19608, new_n14435);
not_3  g17786(new_n20135, new_n20134);
nor_4  g17787(new_n20136, n20036, new_n19084);
nor_4  g17788(new_n20137, new_n4612, new_n4604);
nor_4  g17789(new_n20138_1, new_n20137, new_n20136);
xor_3  g17790(new_n20139, n19608, new_n14435);
nand_4 g17791(new_n20140, new_n20139, new_n20138_1);
nand_4 g17792(new_n20141, new_n20140, new_n20135);
nand_4 g17793(new_n20142, new_n20141, new_n20133);
nand_4 g17794(new_n20143, new_n20142, new_n20132);
nand_4 g17795(new_n20144, new_n20143, new_n20130);
nand_4 g17796(new_n20145, new_n20144, new_n20129);
nand_4 g17797(new_n20146, new_n20145, new_n20127);
nand_4 g17798(new_n20147, new_n20146, new_n20126_1);
nand_4 g17799(new_n20148, new_n20147, new_n20125);
nand_4 g17800(new_n20149_1, new_n20148, new_n20124);
nand_4 g17801(new_n20150, new_n20149_1, new_n20123);
not_3  g17802(new_n20151_1, new_n20150);
nor_4  g17803(new_n20152, new_n20151_1, new_n20122);
xor_3  g17804(new_n20153, new_n20152, new_n20121);
not_3  g17805(new_n20154, new_n20153);
xnor_3 g17806(new_n20155, new_n20154, new_n14412_1);
not_3  g17807(new_n20156, new_n20155);
xnor_3 g17808(new_n20157, new_n20149_1, new_n20123);
not_3  g17809(new_n20158, new_n20157);
nor_4  g17810(new_n20159, new_n20158, new_n8073);
not_3  g17811(new_n20160, new_n20159);
nor_4  g17812(new_n20161, new_n20157, new_n8074);
nor_4  g17813(new_n20162, new_n20161, new_n20159);
xnor_3 g17814(new_n20163, new_n20147, new_n20125);
nand_4 g17815(new_n20164, new_n20163, new_n8077);
xnor_3 g17816(new_n20165, new_n20163, new_n8078);
xnor_3 g17817(new_n20166, new_n20145, new_n20127);
nand_4 g17818(new_n20167, new_n20166, new_n8084);
xnor_3 g17819(new_n20168, new_n20166, new_n8087);
xnor_3 g17820(new_n20169_1, new_n20143, new_n20130);
nand_4 g17821(new_n20170, new_n20169_1, new_n8092);
xnor_3 g17822(new_n20171, new_n20169_1, new_n8095_1);
xnor_3 g17823(new_n20172, new_n20141, new_n20133);
not_3  g17824(new_n20173, new_n20172);
nor_4  g17825(new_n20174, new_n20173, new_n8102);
not_3  g17826(new_n20175, new_n20174);
nor_4  g17827(new_n20176, new_n20172, new_n8099);
nor_4  g17828(new_n20177, new_n20176, new_n20174);
xnor_3 g17829(new_n20178, new_n20139, new_n20138_1);
not_3  g17830(new_n20179_1, new_n20178);
nor_4  g17831(new_n20180, new_n20179_1, new_n8106);
not_3  g17832(new_n20181, new_n20180);
nor_4  g17833(new_n20182, new_n20178, new_n8107);
nor_4  g17834(new_n20183, new_n20182, new_n20180);
nor_4  g17835(new_n20184, new_n4613, new_n8119);
not_3  g17836(new_n20185, new_n20184);
nand_4 g17837(new_n20186, new_n4638, new_n4635);
nand_4 g17838(new_n20187_1, new_n20186, new_n20185);
nand_4 g17839(new_n20188, new_n20187_1, new_n20183);
nand_4 g17840(new_n20189, new_n20188, new_n20181);
nand_4 g17841(new_n20190, new_n20189, new_n20177);
nand_4 g17842(new_n20191, new_n20190, new_n20175);
nand_4 g17843(new_n20192, new_n20191, new_n20171);
nand_4 g17844(new_n20193, new_n20192, new_n20170);
nand_4 g17845(new_n20194, new_n20193, new_n20168);
nand_4 g17846(new_n20195, new_n20194, new_n20167);
nand_4 g17847(new_n20196, new_n20195, new_n20165);
nand_4 g17848(new_n20197, new_n20196, new_n20164);
nand_4 g17849(new_n20198, new_n20197, new_n20162);
nand_4 g17850(new_n20199, new_n20198, new_n20160);
xnor_3 g17851(new_n20200, new_n20199, new_n20156);
xnor_3 g17852(new_n20201, new_n20200, new_n20119);
not_3  g17853(new_n20202, new_n20198);
nor_4  g17854(new_n20203, new_n20197, new_n20162);
nor_4  g17855(new_n20204, new_n20203, new_n20202);
nand_4 g17856(new_n20205, new_n20204, new_n7439);
xnor_3 g17857(new_n20206, new_n20204, new_n7440);
xnor_3 g17858(new_n20207, new_n20195, new_n20165);
not_3  g17859(new_n20208, new_n20207);
nand_4 g17860(new_n20209, new_n20208, new_n7446);
xnor_3 g17861(new_n20210, new_n20207, new_n7446);
xnor_3 g17862(new_n20211, new_n20166, new_n8084);
xnor_3 g17863(new_n20212, new_n20193, new_n20211);
nand_4 g17864(new_n20213_1, new_n20212, new_n7452);
xnor_3 g17865(new_n20214, new_n20212, new_n7451);
not_3  g17866(new_n20215, new_n20171);
xnor_3 g17867(new_n20216, new_n20191, new_n20215);
nand_4 g17868(new_n20217, new_n20216, new_n7460_1);
not_3  g17869(new_n20218, new_n7460_1);
xnor_3 g17870(new_n20219, new_n20216, new_n20218);
xnor_3 g17871(new_n20220, new_n20189, new_n20177);
not_3  g17872(new_n20221, new_n20220);
nand_4 g17873(new_n20222, new_n20221, new_n7466);
xnor_3 g17874(new_n20223, new_n20220, new_n7466);
xnor_3 g17875(new_n20224, new_n20187_1, new_n20183);
nor_4  g17876(new_n20225, new_n20224, new_n7477_1);
not_3  g17877(new_n20226, new_n20225);
nor_4  g17878(new_n20227, new_n4634, new_n20184);
xnor_3 g17879(new_n20228, new_n20227, new_n20183);
nor_4  g17880(new_n20229, new_n20228, new_n7475_1);
nor_4  g17881(new_n20230, new_n20229, new_n20225);
nand_4 g17882(new_n20231, new_n7484, new_n4640);
nand_4 g17883(new_n20232, new_n4666, new_n4652);
nand_4 g17884(new_n20233, new_n20232, new_n20231);
nand_4 g17885(new_n20234, new_n20233, new_n20230);
nand_4 g17886(new_n20235_1, new_n20234, new_n20226);
nand_4 g17887(new_n20236, new_n20235_1, new_n20223);
nand_4 g17888(new_n20237, new_n20236, new_n20222);
nand_4 g17889(new_n20238, new_n20237, new_n20219);
nand_4 g17890(new_n20239, new_n20238, new_n20217);
nand_4 g17891(new_n20240, new_n20239, new_n20214);
nand_4 g17892(new_n20241, new_n20240, new_n20213_1);
nand_4 g17893(new_n20242, new_n20241, new_n20210);
nand_4 g17894(new_n20243, new_n20242, new_n20209);
nand_4 g17895(new_n20244, new_n20243, new_n20206);
nand_4 g17896(new_n20245, new_n20244, new_n20205);
xnor_3 g17897(n3932, new_n20245, new_n20201);
not_3  g17898(new_n20247, new_n4319_1);
xor_3  g17899(n3934, new_n4322, new_n20247);
xor_3  g17900(n3971, new_n4581, new_n4577);
nor_4  g17901(new_n20250_1, n8581, n5026);
nand_4 g17902(new_n20251, new_n20250_1, new_n7792);
nor_4  g17903(new_n20252, new_n20251, n18157);
nand_4 g17904(new_n20253, new_n20252, new_n12653);
nor_4  g17905(new_n20254, new_n20253, n8067);
nand_4 g17906(new_n20255, new_n20254, new_n8506);
nor_4  g17907(new_n20256, new_n20255, n25240);
xor_3  g17908(new_n20257, new_n20256, new_n8501);
not_3  g17909(new_n20258, new_n20257);
nor_4  g17910(new_n20259_1, new_n20258, new_n10438);
nor_4  g17911(new_n20260, new_n20257, n15077);
nor_4  g17912(new_n20261, new_n20260, new_n20259_1);
xor_3  g17913(new_n20262, new_n20255, n25240);
nor_4  g17914(new_n20263, new_n20262, n3710);
xnor_3 g17915(new_n20264, new_n20262, new_n10445);
not_3  g17916(new_n20265, new_n20264);
xor_3  g17917(new_n20266, new_n20254, n10125);
nor_4  g17918(new_n20267, new_n20266, new_n10454);
not_3  g17919(new_n20268, new_n20267);
xor_3  g17920(new_n20269, new_n20254, new_n8506);
nor_4  g17921(new_n20270, new_n20269, n26318);
not_3  g17922(new_n20271, new_n20270);
nand_4 g17923(new_n20272, new_n20253, n8067);
not_3  g17924(new_n20273, new_n20272);
nor_4  g17925(new_n20274, new_n20273, new_n20254);
nor_4  g17926(new_n20275, new_n20274, n26054);
xnor_3 g17927(new_n20276, new_n20274, new_n12106);
not_3  g17928(new_n20277, new_n20276);
xnor_3 g17929(new_n20278, new_n20252, n20923);
nor_4  g17930(new_n20279_1, new_n20278, n19081);
xnor_3 g17931(new_n20280, new_n20278, new_n10462);
nand_4 g17932(new_n20281, new_n20251, n18157);
not_3  g17933(new_n20282, new_n20281);
nor_4  g17934(new_n20283, new_n20282, new_n20252);
nor_4  g17935(new_n20284, new_n20283, n8309);
not_3  g17936(new_n20285, new_n20284);
xnor_3 g17937(new_n20286, new_n20250_1, n12161);
nor_4  g17938(new_n20287_1, new_n20286, n19144);
not_3  g17939(new_n20288, new_n20287_1);
not_3  g17940(new_n20289, new_n20286);
nor_4  g17941(new_n20290, new_n20289, new_n10474);
nor_4  g17942(new_n20291, new_n20290, new_n20287_1);
xnor_3 g17943(new_n20292, n8581, n5026);
nand_4 g17944(new_n20293, new_n20292, new_n10483);
nand_4 g17945(new_n20294, n13714, n8581);
xnor_3 g17946(new_n20295, new_n20292, n12593);
nand_4 g17947(new_n20296, new_n20295, new_n20294);
nand_4 g17948(new_n20297, new_n20296, new_n20293);
nand_4 g17949(new_n20298, new_n20297, new_n20291);
nand_4 g17950(new_n20299, new_n20298, new_n20288);
not_3  g17951(new_n20300, new_n20283);
nor_4  g17952(new_n20301_1, new_n20300, new_n10490);
nor_4  g17953(new_n20302, new_n20301_1, new_n20284);
nand_4 g17954(new_n20303, new_n20302, new_n20299);
nand_4 g17955(new_n20304, new_n20303, new_n20285);
nand_4 g17956(new_n20305, new_n20304, new_n20280);
not_3  g17957(new_n20306, new_n20305);
nor_4  g17958(new_n20307, new_n20306, new_n20279_1);
nor_4  g17959(new_n20308, new_n20307, new_n20277);
nor_4  g17960(new_n20309, new_n20308, new_n20275);
nand_4 g17961(new_n20310, new_n20309, new_n20271);
nand_4 g17962(new_n20311, new_n20310, new_n20268);
nor_4  g17963(new_n20312, new_n20311, new_n20265);
nor_4  g17964(new_n20313, new_n20312, new_n20263);
xnor_3 g17965(new_n20314, new_n20313, new_n20261);
xnor_3 g17966(new_n20315, new_n20314, n26797);
not_3  g17967(new_n20316, n23913);
xnor_3 g17968(new_n20317, new_n20311, new_n20264);
nor_4  g17969(new_n20318, new_n20317, new_n20316);
xnor_3 g17970(new_n20319, new_n20317, new_n20316);
nor_4  g17971(new_n20320, new_n20270, new_n20267);
xnor_3 g17972(new_n20321, new_n20320, new_n20309);
nor_4  g17973(new_n20322, new_n20321, new_n6434);
xnor_3 g17974(new_n20323, new_n20321, new_n6434);
not_3  g17975(new_n20324, n20429);
xnor_3 g17976(new_n20325, new_n20307, new_n20276);
nor_4  g17977(new_n20326, new_n20325, new_n20324);
xnor_3 g17978(new_n20327, new_n20325, new_n20324);
xnor_3 g17979(new_n20328, new_n20304, new_n20280);
not_3  g17980(new_n20329, new_n20328);
nor_4  g17981(new_n20330_1, new_n20329, new_n6435);
not_3  g17982(new_n20331, new_n20330_1);
nor_4  g17983(new_n20332, new_n20328, n3909);
nor_4  g17984(new_n20333_1, new_n20332, new_n20330_1);
xnor_3 g17985(new_n20334, new_n20302, new_n20299);
not_3  g17986(new_n20335, new_n20334);
nor_4  g17987(new_n20336, new_n20335, new_n9541);
not_3  g17988(new_n20337, new_n20336);
nor_4  g17989(new_n20338, new_n20334, n23974);
nor_4  g17990(new_n20339, new_n20338, new_n20336);
xnor_3 g17991(new_n20340, new_n20297, new_n20291);
not_3  g17992(new_n20341, new_n20340);
nor_4  g17993(new_n20342, new_n20341, new_n6436);
not_3  g17994(new_n20343, new_n20342);
nor_4  g17995(new_n20344, new_n20340, n2146);
nor_4  g17996(new_n20345, new_n20344, new_n20342);
xnor_3 g17997(new_n20346, new_n20295, new_n20294);
not_3  g17998(new_n20347, new_n20346);
nor_4  g17999(new_n20348, new_n20347, new_n9551);
not_3  g18000(new_n20349_1, new_n20348);
xor_3  g18001(new_n20350, n13714, n8581);
not_3  g18002(new_n20351, new_n20350);
nor_4  g18003(new_n20352, new_n20351, new_n9549);
nor_4  g18004(new_n20353, new_n20346, n22173);
nor_4  g18005(new_n20354, new_n20353, new_n20348);
nand_4 g18006(new_n20355_1, new_n20354, new_n20352);
nand_4 g18007(new_n20356, new_n20355_1, new_n20349_1);
nand_4 g18008(new_n20357, new_n20356, new_n20345);
nand_4 g18009(new_n20358, new_n20357, new_n20343);
nand_4 g18010(new_n20359_1, new_n20358, new_n20339);
nand_4 g18011(new_n20360, new_n20359_1, new_n20337);
nand_4 g18012(new_n20361, new_n20360, new_n20333_1);
nand_4 g18013(new_n20362, new_n20361, new_n20331);
not_3  g18014(new_n20363, new_n20362);
nor_4  g18015(new_n20364, new_n20363, new_n20327);
nor_4  g18016(new_n20365, new_n20364, new_n20326);
nor_4  g18017(new_n20366_1, new_n20365, new_n20323);
nor_4  g18018(new_n20367, new_n20366_1, new_n20322);
nor_4  g18019(new_n20368, new_n20367, new_n20319);
nor_4  g18020(new_n20369, new_n20368, new_n20318);
xnor_3 g18021(new_n20370, new_n20369, new_n20315);
xnor_3 g18022(new_n20371, new_n20370, new_n9667);
not_3  g18023(new_n20372, new_n20319);
xnor_3 g18024(new_n20373, new_n20367, new_n20372);
nor_4  g18025(new_n20374, new_n20373, new_n9675);
not_3  g18026(new_n20375, new_n20374);
xnor_3 g18027(new_n20376, new_n20373, new_n9674);
xnor_3 g18028(new_n20377, new_n20321, n22554);
xnor_3 g18029(new_n20378, new_n20365, new_n20377);
nor_4  g18030(new_n20379, new_n20378, new_n9682);
not_3  g18031(new_n20380, new_n20379);
xnor_3 g18032(new_n20381, new_n20378, new_n9686);
xnor_3 g18033(new_n20382, new_n20362, new_n20327);
nor_4  g18034(new_n20383, new_n20382, new_n9690);
not_3  g18035(new_n20384, new_n20383);
not_3  g18036(new_n20385_1, new_n20382);
nor_4  g18037(new_n20386, new_n20385_1, new_n9691);
nor_4  g18038(new_n20387, new_n20386, new_n20383);
xnor_3 g18039(new_n20388_1, new_n20360, new_n20333_1);
nand_4 g18040(new_n20389, new_n20388_1, new_n9697);
not_3  g18041(new_n20390, new_n20388_1);
xnor_3 g18042(new_n20391, new_n20390, new_n9697);
xnor_3 g18043(new_n20392, new_n20358, new_n20339);
nand_4 g18044(new_n20393, new_n20392, new_n9703);
xnor_3 g18045(new_n20394, new_n20392, new_n9702);
xnor_3 g18046(new_n20395, new_n20356, new_n20345);
nand_4 g18047(new_n20396, new_n20395, new_n9709);
xnor_3 g18048(new_n20397, new_n20354, new_n20352);
nand_4 g18049(new_n20398, new_n20397, new_n9722);
xor_3  g18050(new_n20399, new_n20351, new_n9549);
nand_4 g18051(new_n20400, new_n20399, new_n2595);
xor_3  g18052(new_n20401, new_n9502, new_n9497);
xnor_3 g18053(new_n20402_1, new_n20397, new_n20401);
nand_4 g18054(new_n20403_1, new_n20402_1, new_n20400);
nand_4 g18055(new_n20404, new_n20403_1, new_n20398);
xnor_3 g18056(new_n20405, new_n20395, new_n9710);
nand_4 g18057(new_n20406, new_n20405, new_n20404);
nand_4 g18058(new_n20407, new_n20406, new_n20396);
nand_4 g18059(new_n20408, new_n20407, new_n20394);
nand_4 g18060(new_n20409_1, new_n20408, new_n20393);
nand_4 g18061(new_n20410, new_n20409_1, new_n20391);
nand_4 g18062(new_n20411_1, new_n20410, new_n20389);
nand_4 g18063(new_n20412, new_n20411_1, new_n20387);
nand_4 g18064(new_n20413, new_n20412, new_n20384);
nand_4 g18065(new_n20414, new_n20413, new_n20381);
nand_4 g18066(new_n20415, new_n20414, new_n20380);
nand_4 g18067(new_n20416, new_n20415, new_n20376);
nand_4 g18068(new_n20417, new_n20416, new_n20375);
not_3  g18069(new_n20418, new_n20417);
xor_3  g18070(n3983, new_n20418, new_n20371);
xor_3  g18071(new_n20420, n13714, n583);
nor_4  g18072(new_n20421, new_n20420, n6611);
nand_4 g18073(new_n20422, new_n20420, n6611);
not_3  g18074(new_n20423, new_n20422);
nor_4  g18075(new_n20424_1, new_n20423, new_n20421);
nor_4  g18076(new_n20425, new_n20424_1, new_n7842);
nand_4 g18077(new_n20426, n13714, n583);
not_3  g18078(new_n20427, new_n20426);
xnor_3 g18079(new_n20428, n22173, n12593);
xor_3  g18080(new_n20429_1, new_n20428, new_n20427);
xnor_3 g18081(new_n20430, new_n20429_1, new_n6479);
nor_4  g18082(new_n20431, new_n20430, new_n20423);
xor_3  g18083(new_n20432, new_n20428, new_n20426);
nor_4  g18084(new_n20433, new_n20432, n27188);
nor_4  g18085(new_n20434, new_n20429_1, new_n6479);
nor_4  g18086(new_n20435, new_n20434, new_n20433);
nor_4  g18087(new_n20436_1, new_n20435, new_n20422);
nor_4  g18088(new_n20437, new_n20436_1, new_n20431);
xnor_3 g18089(new_n20438, new_n20437, new_n20425);
xor_3  g18090(n4000, new_n20438, new_n7837);
xor_3  g18091(new_n20440, n26823, new_n8803_1);
nand_4 g18092(new_n20441_1, new_n8807, n4812);
xor_3  g18093(new_n20442, n19228, new_n15864);
nand_4 g18094(new_n20443, n24278, new_n8811);
xor_3  g18095(new_n20444, n24278, new_n8811);
nand_4 g18096(new_n20445_1, n24618, new_n8815);
nand_4 g18097(new_n20446, new_n3314, n8052);
nand_4 g18098(new_n20447, n10158, new_n13536);
nand_4 g18099(new_n20448, new_n13537, new_n13535);
nand_4 g18100(new_n20449, new_n20448, new_n20447);
not_3  g18101(new_n20450_1, new_n20449);
nand_4 g18102(new_n20451, new_n20450_1, new_n20446);
nand_4 g18103(new_n20452, new_n20451, new_n20445_1);
nand_4 g18104(new_n20453, new_n20452, new_n20444);
nand_4 g18105(new_n20454, new_n20453, new_n20443);
nand_4 g18106(new_n20455_1, new_n20454, new_n20442);
nand_4 g18107(new_n20456, new_n20455_1, new_n20441_1);
xor_3  g18108(new_n20457, new_n20456, new_n20440);
xnor_3 g18109(new_n20458, new_n20457, new_n8737);
not_3  g18110(new_n20459, new_n20458);
xor_3  g18111(new_n20460, new_n20454, new_n20442);
not_3  g18112(new_n20461, new_n20460);
nand_4 g18113(new_n20462, new_n20461, new_n8743);
xnor_3 g18114(new_n20463, new_n20460, new_n8743);
not_3  g18115(new_n20464, new_n20444);
xor_3  g18116(new_n20465, new_n20452, new_n20464);
nand_4 g18117(new_n20466, new_n20465, new_n8747);
nand_4 g18118(new_n20467, new_n20446, new_n20445_1);
xor_3  g18119(new_n20468, new_n20467, new_n20450_1);
nand_4 g18120(new_n20469, new_n20468, new_n8751);
not_3  g18121(new_n20470_1, new_n20468);
xnor_3 g18122(new_n20471, new_n20470_1, new_n8751);
not_3  g18123(new_n20472, new_n13534);
not_3  g18124(new_n20473, new_n13539);
nor_4  g18125(new_n20474, new_n20473, new_n20472);
nor_4  g18126(new_n20475, new_n13540, new_n8765);
nor_4  g18127(new_n20476, new_n20475, new_n20474);
nand_4 g18128(new_n20477, new_n20476, new_n20471);
nand_4 g18129(new_n20478_1, new_n20477, new_n20469);
xnor_3 g18130(new_n20479, new_n20465, new_n8746);
nand_4 g18131(new_n20480, new_n20479, new_n20478_1);
nand_4 g18132(new_n20481, new_n20480, new_n20466);
nand_4 g18133(new_n20482, new_n20481, new_n20463);
nand_4 g18134(new_n20483, new_n20482, new_n20462);
xor_3  g18135(n4010, new_n20483, new_n20459);
xor_3  g18136(new_n20485, n11220, new_n14210);
not_3  g18137(new_n20486, new_n20485);
not_3  g18138(new_n20487, n10763);
nor_4  g18139(new_n20488, n22379, new_n20487);
xor_3  g18140(new_n20489_1, n22379, new_n20487);
nor_4  g18141(new_n20490_1, new_n14261, n1662);
not_3  g18142(new_n20491, new_n20490_1);
xor_3  g18143(new_n20492, n7437, new_n2987);
nor_4  g18144(new_n20493, new_n3037, n12875);
not_3  g18145(new_n20494, new_n20493);
not_3  g18146(new_n20495_1, n7099);
nor_4  g18147(new_n20496, new_n20495_1, n2035);
not_3  g18148(new_n20497, new_n20496);
nand_4 g18149(new_n20498, new_n17913, new_n17889_1);
nand_4 g18150(new_n20499, new_n20498, new_n20497);
xor_3  g18151(new_n20500, n20700, new_n2989);
nand_4 g18152(new_n20501, new_n20500, new_n20499);
nand_4 g18153(new_n20502, new_n20501, new_n20494);
nand_4 g18154(new_n20503, new_n20502, new_n20492);
nand_4 g18155(new_n20504, new_n20503, new_n20491);
nand_4 g18156(new_n20505, new_n20504, new_n20489_1);
not_3  g18157(new_n20506, new_n20505);
nor_4  g18158(new_n20507, new_n20506, new_n20488);
xor_3  g18159(new_n20508, new_n20507, new_n20486);
xnor_3 g18160(new_n20509, new_n20508, new_n18093);
not_3  g18161(new_n20510, new_n20509);
xnor_3 g18162(new_n20511, new_n20504, new_n20489_1);
nand_4 g18163(new_n20512, new_n20511, new_n18104);
xnor_3 g18164(new_n20513, new_n20511, new_n18103);
not_3  g18165(new_n20514, new_n20492);
xor_3  g18166(new_n20515_1, new_n20502, new_n20514);
nand_4 g18167(new_n20516, new_n20515_1, new_n18113);
not_3  g18168(new_n20517, new_n20500);
xor_3  g18169(new_n20518, new_n20517, new_n20499);
nor_4  g18170(new_n20519, new_n20518, new_n18126);
xnor_3 g18171(new_n20520, new_n20518, new_n18126);
nor_4  g18172(new_n20521, new_n17930, new_n17914);
nor_4  g18173(new_n20522, new_n17961, new_n17931_1);
nor_4  g18174(new_n20523, new_n20522, new_n20521);
nor_4  g18175(new_n20524, new_n20523, new_n20520);
nor_4  g18176(new_n20525, new_n20524, new_n20519);
xnor_3 g18177(new_n20526, new_n20515_1, new_n18109);
nand_4 g18178(new_n20527, new_n20526, new_n20525);
nand_4 g18179(new_n20528, new_n20527, new_n20516);
nand_4 g18180(new_n20529, new_n20528, new_n20513);
nand_4 g18181(new_n20530, new_n20529, new_n20512);
xnor_3 g18182(n4014, new_n20530, new_n20510);
not_3  g18183(new_n20532, new_n14348);
xor_3  g18184(new_n20533_1, new_n17178, n18496);
nor_4  g18185(new_n20534, new_n17183, n26224);
xor_3  g18186(new_n20535, new_n17185, n26224);
nor_4  g18187(new_n20536, new_n4082, n19327);
nor_4  g18188(new_n20537, new_n4133, new_n4084);
nor_4  g18189(new_n20538, new_n20537, new_n20536);
nor_4  g18190(new_n20539, new_n20538, new_n20535);
nor_4  g18191(new_n20540, new_n20539, new_n20534);
xnor_3 g18192(new_n20541, new_n20540, new_n20533_1);
nor_4  g18193(new_n20542, new_n20541, n647);
not_3  g18194(new_n20543, new_n20541);
nor_4  g18195(new_n20544, new_n20543, new_n8656_1);
nor_4  g18196(new_n20545, new_n20544, new_n20542);
xnor_3 g18197(new_n20546, new_n20538, new_n20535);
not_3  g18198(new_n20547, new_n20546);
nor_4  g18199(new_n20548, new_n20547, new_n8659);
xnor_3 g18200(new_n20549, new_n20546, n20409);
not_3  g18201(new_n20550, new_n4134_1);
nor_4  g18202(new_n20551, new_n20550, new_n5472_1);
nor_4  g18203(new_n20552, new_n4183, new_n4135);
nor_4  g18204(new_n20553, new_n20552, new_n20551);
nor_4  g18205(new_n20554, new_n20553, new_n20549);
nor_4  g18206(new_n20555, new_n20554, new_n20548);
not_3  g18207(new_n20556, new_n20555);
xnor_3 g18208(new_n20557, new_n20556, new_n20545);
xnor_3 g18209(new_n20558, new_n20557, new_n20532);
not_3  g18210(new_n20559, new_n20549);
not_3  g18211(new_n20560, new_n20551);
not_3  g18212(new_n20561, new_n20552);
nand_4 g18213(new_n20562, new_n20561, new_n20560);
nor_4  g18214(new_n20563, new_n20562, new_n20559);
nor_4  g18215(new_n20564, new_n20563, new_n20554);
nor_4  g18216(new_n20565, new_n20564, new_n14354);
xnor_3 g18217(new_n20566, new_n20564, new_n14354);
not_3  g18218(new_n20567, new_n4184);
nor_4  g18219(new_n20568, new_n4282, new_n20567);
not_3  g18220(new_n20569, new_n4331);
nor_4  g18221(new_n20570, new_n20569, new_n4289);
nor_4  g18222(new_n20571, new_n20570, new_n4284);
nor_4  g18223(new_n20572, new_n20571, new_n20568);
nor_4  g18224(new_n20573, new_n20572, new_n20566);
nor_4  g18225(new_n20574, new_n20573, new_n20565);
xnor_3 g18226(n4071, new_n20574, new_n20558);
not_3  g18227(new_n20576, new_n15600);
xor_3  g18228(n4088, new_n20576, new_n15591);
not_3  g18229(new_n20578, new_n15742);
nor_4  g18230(new_n20579, new_n20578, n7593);
not_3  g18231(new_n20580, new_n20579);
not_3  g18232(new_n20581, new_n15746);
not_3  g18233(new_n20582_1, new_n15745);
nand_4 g18234(new_n20583, new_n15755, new_n20582_1);
nand_4 g18235(new_n20584, new_n20583, new_n20581);
nand_4 g18236(new_n20585, new_n20584, new_n20580);
not_3  g18237(new_n20586, new_n19865);
not_3  g18238(new_n20587, new_n19863);
nand_4 g18239(new_n20588, new_n19874, new_n20587);
nand_4 g18240(new_n20589, new_n20588, new_n20586);
nor_4  g18241(new_n20590_1, new_n20589, new_n20585);
not_3  g18242(new_n20591, new_n20585);
nor_4  g18243(new_n20592, new_n20591, new_n19875);
nor_4  g18244(new_n20593, new_n20585, new_n19872);
nor_4  g18245(new_n20594, new_n15756, new_n19878);
not_3  g18246(new_n20595, new_n20594);
nand_4 g18247(new_n20596, new_n15762_1, new_n20595);
nor_4  g18248(new_n20597, new_n20596, new_n20593);
nor_4  g18249(new_n20598, new_n20597, new_n20592);
nor_4  g18250(new_n20599, new_n20598, new_n20590_1);
not_3  g18251(new_n20600, new_n20589);
nor_4  g18252(new_n20601, new_n20600, new_n20591);
nor_4  g18253(new_n20602_1, new_n20601, new_n20597);
nor_4  g18254(n4089, new_n20602_1, new_n20599);
not_3  g18255(new_n20604_1, n3228);
nand_4 g18256(new_n20605, new_n14587, new_n7937_1);
xor_3  g18257(new_n20606, new_n20605, n2289);
not_3  g18258(new_n20607, new_n20606);
nor_4  g18259(new_n20608, new_n20607, new_n20604_1);
nor_4  g18260(new_n20609_1, new_n20606, n3228);
nor_4  g18261(new_n20610, new_n20609_1, new_n20608);
nand_4 g18262(new_n20611, new_n14588, n5302);
xor_3  g18263(new_n20612, new_n14587, n1112);
nand_4 g18264(new_n20613, new_n20612, new_n3274);
not_3  g18265(new_n20614, n25738);
not_3  g18266(new_n20615, new_n14595);
nor_4  g18267(new_n20616, new_n20615, new_n20614);
not_3  g18268(new_n20617, new_n20616);
nor_4  g18269(new_n20618, new_n14595, n25738);
not_3  g18270(new_n20619, new_n20618);
nor_4  g18271(new_n20620, new_n10232, n21471);
nor_4  g18272(new_n20621, new_n10262_1, new_n10233);
nor_4  g18273(new_n20622, new_n20621, new_n20620);
nand_4 g18274(new_n20623_1, new_n20622, new_n20619);
nand_4 g18275(new_n20624, new_n20623_1, new_n20617);
nand_4 g18276(new_n20625, new_n20624, new_n20613);
nand_4 g18277(new_n20626, new_n20625, new_n20611);
xnor_3 g18278(new_n20627, new_n20626, new_n20610);
xnor_3 g18279(new_n20628, new_n20627, new_n8045);
not_3  g18280(new_n20629_1, new_n20628);
nand_4 g18281(new_n20630, new_n20613, new_n20611);
xnor_3 g18282(new_n20631, new_n20630, new_n20624);
nor_4  g18283(new_n20632, new_n20631, n1293);
not_3  g18284(new_n20633, new_n20632);
nor_4  g18285(new_n20634, new_n20612, new_n3274);
nor_4  g18286(new_n20635, new_n14588, n5302);
nor_4  g18287(new_n20636, new_n20635, new_n20634);
xnor_3 g18288(new_n20637, new_n20636, new_n20624);
nor_4  g18289(new_n20638, new_n20637, new_n10335);
nor_4  g18290(new_n20639, new_n20638, new_n20632);
nor_4  g18291(new_n20640, new_n20618, new_n20616);
xnor_3 g18292(new_n20641, new_n20640, new_n20622);
nor_4  g18293(new_n20642, new_n20641, new_n10337);
not_3  g18294(new_n20643, new_n20642);
not_3  g18295(new_n20644, new_n10267);
nand_4 g18296(new_n20645, new_n10294, new_n10268);
nand_4 g18297(new_n20646, new_n20645, new_n20644);
not_3  g18298(new_n20647, new_n20641);
nor_4  g18299(new_n20648, new_n20647, n19042);
nor_4  g18300(new_n20649, new_n20648, new_n20642);
nand_4 g18301(new_n20650, new_n20649, new_n20646);
nand_4 g18302(new_n20651, new_n20650, new_n20643);
not_3  g18303(new_n20652, new_n20651);
nand_4 g18304(new_n20653, new_n20652, new_n20639);
nand_4 g18305(new_n20654, new_n20653, new_n20633);
nor_4  g18306(new_n20655, new_n20654, new_n20629_1);
xnor_3 g18307(new_n20656, new_n20631, n1293);
nor_4  g18308(new_n20657, new_n20651, new_n20656);
nor_4  g18309(new_n20658_1, new_n20657, new_n20632);
nor_4  g18310(new_n20659, new_n20658_1, new_n20628);
nor_4  g18311(new_n20660, new_n20659, new_n20655);
xnor_3 g18312(new_n20661_1, new_n8917, new_n6330_1);
nand_4 g18313(new_n20662, new_n8923, n23200);
nor_4  g18314(new_n20663, new_n2483, new_n8081);
nor_4  g18315(new_n20664, new_n8923, n23200);
nor_4  g18316(new_n20665, new_n20664, new_n20663);
nand_4 g18317(new_n20666, new_n2494, n17959);
xnor_3 g18318(new_n20667, new_n2494, new_n6335);
nand_4 g18319(new_n20668, new_n2497, n7566);
nand_4 g18320(new_n20669, new_n7869, new_n7855);
nand_4 g18321(new_n20670, new_n20669, new_n20668);
nand_4 g18322(new_n20671, new_n20670, new_n20667);
nand_4 g18323(new_n20672, new_n20671, new_n20666);
nand_4 g18324(new_n20673_1, new_n20672, new_n20665);
nand_4 g18325(new_n20674, new_n20673_1, new_n20662);
xnor_3 g18326(new_n20675, new_n20674, new_n20661_1);
not_3  g18327(new_n20676, new_n20675);
xnor_3 g18328(new_n20677, new_n20676, new_n20660);
not_3  g18329(new_n20678_1, new_n20677);
xnor_3 g18330(new_n20679, new_n20651, new_n20656);
not_3  g18331(new_n20680_1, new_n20679);
not_3  g18332(new_n20681, new_n20672);
xnor_3 g18333(new_n20682, new_n20681, new_n20665);
not_3  g18334(new_n20683, new_n20682);
nand_4 g18335(new_n20684, new_n20683, new_n20680_1);
not_3  g18336(new_n20685_1, new_n20684);
xnor_3 g18337(new_n20686, new_n20682, new_n20679);
xnor_3 g18338(new_n20687, new_n20670, new_n20667);
xnor_3 g18339(new_n20688, new_n20649, new_n20646);
nand_4 g18340(new_n20689, new_n20688, new_n20687);
not_3  g18341(new_n20690, new_n20689);
nand_4 g18342(new_n20691_1, new_n10295_1, new_n7870);
not_3  g18343(new_n20692, new_n20691_1);
nor_4  g18344(new_n20693, new_n10322, new_n10296);
nor_4  g18345(new_n20694, new_n20693, new_n20692);
xnor_3 g18346(new_n20695, new_n20688, new_n20687);
nor_4  g18347(new_n20696_1, new_n20695, new_n20694);
nor_4  g18348(new_n20697, new_n20696_1, new_n20690);
nor_4  g18349(new_n20698, new_n20697, new_n20686);
nor_4  g18350(new_n20699, new_n20698, new_n20685_1);
xor_3  g18351(n4103, new_n20699, new_n20678_1);
nor_4  g18352(new_n20701, new_n18003, new_n15425);
nor_4  g18353(new_n20702, new_n19854, new_n15424_1);
nor_4  g18354(new_n20703, new_n20702, new_n20701);
not_3  g18355(new_n20704_1, new_n20703);
nand_4 g18356(new_n20705_1, new_n18007, new_n15338);
nand_4 g18357(new_n20706, new_n18020, new_n15347);
xnor_3 g18358(new_n20707, new_n18012, new_n15347);
nand_4 g18359(new_n20708, new_n18024, new_n15356);
xnor_3 g18360(new_n20709_1, new_n18036, new_n15356);
nor_4  g18361(new_n20710, new_n18119, new_n15362);
not_3  g18362(new_n20711, new_n20710);
not_3  g18363(new_n20712, new_n15362);
nor_4  g18364(new_n20713_1, new_n18027, new_n20712);
nor_4  g18365(new_n20714, new_n20713_1, new_n20710);
not_3  g18366(new_n20715, new_n15368);
nand_4 g18367(new_n20716, new_n17986, new_n17917);
xnor_3 g18368(new_n20717, new_n17923, new_n20716);
nor_4  g18369(new_n20718, new_n20717, new_n20715);
not_3  g18370(new_n20719, new_n20718);
nor_4  g18371(new_n20720, new_n15374, new_n4783);
not_3  g18372(new_n20721, new_n20720);
nor_4  g18373(new_n20722_1, new_n15376, new_n4779);
nor_4  g18374(new_n20723_1, new_n20722_1, new_n20720);
nor_4  g18375(new_n20724, new_n15380, new_n4789);
xnor_3 g18376(new_n20725, new_n15379, new_n4788);
nor_4  g18377(new_n20726, new_n15386, new_n4796);
not_3  g18378(new_n20727, new_n20726);
nor_4  g18379(new_n20728, new_n15389, new_n4795);
nor_4  g18380(new_n20729, new_n20728, new_n20726);
nor_4  g18381(new_n20730, new_n15392, new_n4798);
not_3  g18382(new_n20731, new_n20730);
not_3  g18383(new_n20732, new_n4802);
nand_4 g18384(new_n20733, new_n15394, new_n20732);
nor_4  g18385(new_n20734, new_n15397, new_n4799);
nor_4  g18386(new_n20735, new_n20734, new_n20730);
nand_4 g18387(new_n20736, new_n20735, new_n20733);
nand_4 g18388(new_n20737, new_n20736, new_n20731);
nand_4 g18389(new_n20738, new_n20737, new_n20729);
nand_4 g18390(new_n20739, new_n20738, new_n20727);
nor_4  g18391(new_n20740, new_n20739, new_n20725);
nor_4  g18392(new_n20741, new_n20740, new_n20724);
nand_4 g18393(new_n20742, new_n20741, new_n20723_1);
nand_4 g18394(new_n20743, new_n20742, new_n20721);
nor_4  g18395(new_n20744, new_n17924, new_n15368);
nor_4  g18396(new_n20745, new_n20744, new_n20718);
nand_4 g18397(new_n20746, new_n20745, new_n20743);
nand_4 g18398(new_n20747, new_n20746, new_n20719);
nand_4 g18399(new_n20748_1, new_n20747, new_n20714);
nand_4 g18400(new_n20749, new_n20748_1, new_n20711);
nand_4 g18401(new_n20750, new_n20749, new_n20709_1);
nand_4 g18402(new_n20751, new_n20750, new_n20708);
nand_4 g18403(new_n20752, new_n20751, new_n20707);
nand_4 g18404(new_n20753, new_n20752, new_n20706);
not_3  g18405(new_n20754, new_n20705_1);
nor_4  g18406(new_n20755, new_n18007, new_n15338);
nor_4  g18407(new_n20756, new_n20755, new_n20754);
nand_4 g18408(new_n20757, new_n20756, new_n20753);
nand_4 g18409(new_n20758, new_n20757, new_n20705_1);
nor_4  g18410(new_n20759, new_n20758, new_n20704_1);
nor_4  g18411(new_n20760, new_n20759, new_n20701);
not_3  g18412(new_n20761_1, new_n20760);
nor_4  g18413(new_n20762, new_n6876, new_n16695);
not_3  g18414(new_n20763, new_n20762);
nor_4  g18415(new_n20764, new_n6875, n6456);
nor_4  g18416(new_n20765, new_n6928, n4085);
xor_3  g18417(new_n20766, new_n6929, new_n16702);
not_3  g18418(new_n20767, new_n20766);
nor_4  g18419(new_n20768, new_n6936, n26725);
xor_3  g18420(new_n20769, new_n6940, new_n16709);
not_3  g18421(new_n20770, new_n20769);
nor_4  g18422(new_n20771, new_n6943, n11980);
xnor_3 g18423(new_n20772, new_n6943, n11980);
nor_4  g18424(new_n20773, new_n6954, n3253);
nor_4  g18425(new_n20774_1, new_n6951, new_n6888);
nor_4  g18426(new_n20775, new_n20774_1, new_n20773);
not_3  g18427(new_n20776, new_n20775);
nor_4  g18428(new_n20777, new_n6962, n7759);
xor_3  g18429(new_n20778, new_n6962, n7759);
nand_4 g18430(new_n20779, new_n6970, new_n15793_1);
nand_4 g18431(new_n20780, new_n6981, new_n15801);
xor_3  g18432(new_n20781, new_n6980, n7949);
nand_4 g18433(new_n20782, new_n6996, new_n15819);
nand_4 g18434(new_n20783, n20658, n14575);
xor_3  g18435(new_n20784, new_n6996, new_n15819);
nand_4 g18436(new_n20785, new_n20784, new_n20783);
nand_4 g18437(new_n20786, new_n20785, new_n20782);
nand_4 g18438(new_n20787, new_n20786, new_n20781);
nand_4 g18439(new_n20788_1, new_n20787, new_n20780);
xor_3  g18440(new_n20789, new_n6969, n12562);
nand_4 g18441(new_n20790, new_n20789, new_n20788_1);
nand_4 g18442(new_n20791, new_n20790, new_n20779);
nand_4 g18443(new_n20792, new_n20791, new_n20778);
not_3  g18444(new_n20793, new_n20792);
nor_4  g18445(new_n20794_1, new_n20793, new_n20777);
nor_4  g18446(new_n20795_1, new_n20794_1, new_n20776);
nor_4  g18447(new_n20796, new_n20795_1, new_n20773);
nor_4  g18448(new_n20797, new_n20796, new_n20772);
nor_4  g18449(new_n20798, new_n20797, new_n20771);
nor_4  g18450(new_n20799, new_n20798, new_n20770);
nor_4  g18451(new_n20800, new_n20799, new_n20768);
nor_4  g18452(new_n20801, new_n20800, new_n20767);
nor_4  g18453(new_n20802, new_n20801, new_n20765);
not_3  g18454(new_n20803_1, new_n20802);
nor_4  g18455(new_n20804, new_n20803_1, new_n20764);
nor_4  g18456(new_n20805, new_n20804, new_n16750);
nand_4 g18457(new_n20806, new_n20805, new_n20763);
not_3  g18458(new_n20807, new_n20806);
nand_4 g18459(new_n20808, new_n20807, new_n20761_1);
xnor_3 g18460(new_n20809, new_n20758, new_n20703);
nor_4  g18461(new_n20810, new_n20809, new_n20807);
not_3  g18462(new_n20811, new_n20810);
xnor_3 g18463(new_n20812, new_n20758, new_n20704_1);
nor_4  g18464(new_n20813, new_n20812, new_n20806);
nor_4  g18465(new_n20814, new_n20813, new_n20810);
xnor_3 g18466(new_n20815, new_n18007, new_n15338);
xnor_3 g18467(new_n20816, new_n20815, new_n20753);
nor_4  g18468(new_n20817, new_n20764, new_n20762);
xnor_3 g18469(new_n20818, new_n20817, new_n20802);
nand_4 g18470(new_n20819, new_n20818, new_n20816);
xnor_3 g18471(new_n20820, new_n20756, new_n20753);
xnor_3 g18472(new_n20821, new_n20818, new_n20820);
not_3  g18473(new_n20822, new_n20800);
nor_4  g18474(new_n20823, new_n20822, new_n20766);
nor_4  g18475(new_n20824, new_n20823, new_n20801);
xnor_3 g18476(new_n20825, new_n20751, new_n20707);
not_3  g18477(new_n20826_1, new_n20825);
nand_4 g18478(new_n20827, new_n20826_1, new_n20824);
xnor_3 g18479(new_n20828, new_n20825, new_n20824);
not_3  g18480(new_n20829, new_n20798);
nor_4  g18481(new_n20830, new_n20829, new_n20769);
nor_4  g18482(new_n20831, new_n20830, new_n20799);
xnor_3 g18483(new_n20832, new_n20749, new_n20709_1);
not_3  g18484(new_n20833, new_n20832);
nand_4 g18485(new_n20834, new_n20833, new_n20831);
xnor_3 g18486(new_n20835, new_n20832, new_n20831);
xor_3  g18487(new_n20836, new_n20796, new_n20772);
xnor_3 g18488(new_n20837, new_n20747, new_n20714);
not_3  g18489(new_n20838, new_n20837);
nand_4 g18490(new_n20839, new_n20838, new_n20836);
xnor_3 g18491(new_n20840, new_n20837, new_n20836);
xor_3  g18492(new_n20841, new_n20794_1, new_n20776);
xnor_3 g18493(new_n20842, new_n20745, new_n20743);
not_3  g18494(new_n20843, new_n20842);
nand_4 g18495(new_n20844, new_n20843, new_n20841);
xnor_3 g18496(new_n20845, new_n20842, new_n20841);
nor_4  g18497(new_n20846, new_n20791, new_n20778);
nor_4  g18498(new_n20847, new_n20846, new_n20793);
xnor_3 g18499(new_n20848, new_n20741, new_n20723_1);
not_3  g18500(new_n20849, new_n20848);
nand_4 g18501(new_n20850, new_n20849, new_n20847);
xnor_3 g18502(new_n20851, new_n20848, new_n20847);
xnor_3 g18503(new_n20852, new_n20739, new_n20725);
xnor_3 g18504(new_n20853, new_n20789, new_n20788_1);
not_3  g18505(new_n20854, new_n20853);
nand_4 g18506(new_n20855, new_n20854, new_n20852);
not_3  g18507(new_n20856, new_n20855);
nor_4  g18508(new_n20857, new_n20854, new_n20852);
nor_4  g18509(new_n20858, new_n20857, new_n20856);
not_3  g18510(new_n20859, new_n20781);
xnor_3 g18511(new_n20860, new_n20786, new_n20859);
not_3  g18512(new_n20861, new_n20729);
xnor_3 g18513(new_n20862, new_n20737, new_n20861);
nor_4  g18514(new_n20863, new_n20862, new_n20860);
xnor_3 g18515(new_n20864, new_n20862, new_n20860);
xnor_3 g18516(new_n20865, new_n20735, new_n20733);
nor_4  g18517(new_n20866, new_n20865, new_n20784);
not_3  g18518(new_n20867, new_n20866);
not_3  g18519(new_n20868, new_n20784);
xor_3  g18520(new_n20869_1, new_n20868, new_n20783);
nand_4 g18521(new_n20870, new_n20869_1, new_n20865);
xor_3  g18522(new_n20871, n20658, n14575);
xor_3  g18523(new_n20872, new_n15395, new_n4802);
nand_4 g18524(new_n20873, new_n20872, new_n20871);
nand_4 g18525(new_n20874, new_n20873, new_n20870);
nand_4 g18526(new_n20875, new_n20874, new_n20867);
nor_4  g18527(new_n20876, new_n20875, new_n20864);
nor_4  g18528(new_n20877, new_n20876, new_n20863);
nand_4 g18529(new_n20878, new_n20877, new_n20858);
nand_4 g18530(new_n20879_1, new_n20878, new_n20855);
nand_4 g18531(new_n20880, new_n20879_1, new_n20851);
nand_4 g18532(new_n20881, new_n20880, new_n20850);
nand_4 g18533(new_n20882, new_n20881, new_n20845);
nand_4 g18534(new_n20883, new_n20882, new_n20844);
nand_4 g18535(new_n20884, new_n20883, new_n20840);
nand_4 g18536(new_n20885, new_n20884, new_n20839);
nand_4 g18537(new_n20886, new_n20885, new_n20835);
nand_4 g18538(new_n20887, new_n20886, new_n20834);
nand_4 g18539(new_n20888, new_n20887, new_n20828);
nand_4 g18540(new_n20889, new_n20888, new_n20827);
nand_4 g18541(new_n20890, new_n20889, new_n20821);
nand_4 g18542(new_n20891, new_n20890, new_n20819);
nand_4 g18543(new_n20892, new_n20891, new_n20814);
nand_4 g18544(new_n20893, new_n20892, new_n20811);
nand_4 g18545(new_n20894, new_n20893, new_n20808);
nand_4 g18546(new_n20895, new_n20806, new_n20760);
nand_4 g18547(new_n20896, new_n20895, new_n20892);
nand_4 g18548(new_n20897, new_n20896, new_n20894);
not_3  g18549(n4123, new_n20897);
nor_4  g18550(new_n20899, new_n16094, new_n9348);
nor_4  g18551(new_n20900, new_n16093, new_n9349);
nor_4  g18552(new_n20901, new_n20900, new_n20899);
nor_4  g18553(new_n20902, new_n16104, new_n9356);
not_3  g18554(new_n20903, new_n20902);
nor_4  g18555(new_n20904, new_n16103, new_n9357);
nor_4  g18556(new_n20905, new_n20904, new_n20902);
not_3  g18557(new_n20906, new_n9377);
nor_4  g18558(new_n20907, new_n16113, new_n20906);
not_3  g18559(new_n20908, new_n20907);
not_3  g18560(new_n20909, new_n16113);
nor_4  g18561(new_n20910, new_n20909, new_n9377);
nor_4  g18562(new_n20911, new_n20910, new_n20907);
nor_4  g18563(new_n20912, new_n16125, new_n9365);
not_3  g18564(new_n20913, new_n11716);
nand_4 g18565(new_n20914, new_n20913, new_n9367);
xnor_3 g18566(new_n20915_1, new_n16125, new_n9365);
nor_4  g18567(new_n20916, new_n20915_1, new_n20914);
nor_4  g18568(new_n20917, new_n20916, new_n20912);
nand_4 g18569(new_n20918, new_n20917, new_n20911);
nand_4 g18570(new_n20919, new_n20918, new_n20908);
nand_4 g18571(new_n20920, new_n20919, new_n20905);
nand_4 g18572(new_n20921, new_n20920, new_n20903);
not_3  g18573(new_n20922, new_n20921);
xor_3  g18574(n4134, new_n20922, new_n20901);
xnor_3 g18575(n4146, new_n10862, new_n10794);
nor_4  g18576(new_n20925, new_n18717, new_n17287);
nor_4  g18577(new_n20926, new_n18714, new_n17288);
nor_4  g18578(new_n20927, new_n20926, new_n20925);
nor_4  g18579(new_n20928, new_n18721_1, new_n17300);
xnor_3 g18580(new_n20929_1, new_n18722, new_n17299);
nor_4  g18581(new_n20930, new_n17303, new_n16224);
not_3  g18582(new_n20931, new_n20930);
nor_4  g18583(new_n20932, new_n17307, new_n16213);
xor_3  g18584(new_n20933, new_n17303, new_n16224);
nand_4 g18585(new_n20934, new_n20933, new_n20932);
nand_4 g18586(new_n20935_1, new_n20934, new_n20931);
nor_4  g18587(new_n20936_1, new_n20935_1, new_n20929_1);
nor_4  g18588(new_n20937, new_n20936_1, new_n20928);
not_3  g18589(new_n20938, new_n20937);
xor_3  g18590(n4150, new_n20938, new_n20927);
not_3  g18591(new_n20940, new_n15118_1);
xor_3  g18592(n4151, new_n15119, new_n20940);
nor_4  g18593(new_n20942, new_n15514, new_n15453);
xnor_3 g18594(n4152, new_n20942, new_n15446);
xnor_3 g18595(n4153, new_n7191, new_n7143);
not_3  g18596(new_n20945, n25972);
nor_4  g18597(new_n20946_1, new_n20945, n10250);
nor_4  g18598(new_n20947, new_n10373, new_n10326_1);
nor_4  g18599(new_n20948, new_n20947, new_n20946_1);
not_3  g18600(new_n20949, new_n20948);
nor_4  g18601(new_n20950, new_n20949, new_n14752);
nor_4  g18602(new_n20951, new_n20948, new_n14750);
nor_4  g18603(new_n20952, new_n20951, new_n20950);
nand_4 g18604(new_n20953, new_n20949, new_n14760);
nand_4 g18605(new_n20954, new_n20948, new_n14757);
nor_4  g18606(new_n20955, new_n10584, new_n10375);
nor_4  g18607(new_n20956, new_n10663, new_n20955);
nand_4 g18608(new_n20957, new_n20956, new_n20954);
nand_4 g18609(new_n20958, new_n20957, new_n20953);
xnor_3 g18610(n4165, new_n20958, new_n20952);
xnor_3 g18611(n4172, new_n13893, new_n13857);
xor_3  g18612(n4173, new_n13685, new_n5403_1);
not_3  g18613(new_n20962, new_n7696);
xor_3  g18614(n4176, new_n7723, new_n20962);
not_3  g18615(new_n20964, new_n10843);
xor_3  g18616(n4186, new_n10846, new_n20964);
not_3  g18617(new_n20966, new_n20387);
xor_3  g18618(n4204, new_n20411_1, new_n20966);
not_3  g18619(new_n20968, new_n13771);
not_3  g18620(new_n20969, new_n13741);
nor_4  g18621(new_n20970, new_n20969, new_n6377);
nor_4  g18622(new_n20971, new_n13741, n13494);
nor_4  g18623(new_n20972, new_n20971, new_n20970);
not_3  g18624(new_n20973, new_n7979);
nand_4 g18625(new_n20974, new_n8042_1, new_n7981);
nand_4 g18626(new_n20975, new_n20974, new_n20973);
nand_4 g18627(new_n20976, new_n20975, new_n20972);
not_3  g18628(new_n20977, new_n20976);
nor_4  g18629(new_n20978, new_n20977, new_n20970);
nor_4  g18630(new_n20979, new_n20978, new_n20968);
nand_4 g18631(new_n20980, new_n19585, new_n13723);
nor_4  g18632(new_n20981, new_n20980, n19652);
xor_3  g18633(new_n20982, new_n20981, new_n13903);
not_3  g18634(new_n20983, new_n20982);
nor_4  g18635(new_n20984, new_n20983, n17037);
xor_3  g18636(new_n20985, new_n20983, new_n13804);
xor_3  g18637(new_n20986_1, new_n20980, new_n13907);
nand_4 g18638(new_n20987, new_n20986_1, n5386);
not_3  g18639(new_n20988, new_n19586);
nor_4  g18640(new_n20989, new_n20988, n26191);
nand_4 g18641(new_n20990, new_n19626, new_n19587);
not_3  g18642(new_n20991, new_n20990);
nor_4  g18643(new_n20992, new_n20991, new_n20989);
xnor_3 g18644(new_n20993, new_n20986_1, new_n13812);
nand_4 g18645(new_n20994, new_n20993, new_n20992);
nand_4 g18646(new_n20995, new_n20994, new_n20987);
nor_4  g18647(new_n20996, new_n20995, new_n20985);
nor_4  g18648(new_n20997, new_n20996, new_n20984);
not_3  g18649(new_n20998, new_n20981);
nor_4  g18650(new_n20999, new_n20998, n3984);
xor_3  g18651(new_n21000, new_n20999, new_n13897);
nor_4  g18652(new_n21001, new_n21000, new_n13795);
not_3  g18653(new_n21002, new_n21000);
nor_4  g18654(new_n21003, new_n21002, n7569);
nor_4  g18655(new_n21004, new_n21003, new_n21001);
xnor_3 g18656(new_n21005, new_n21004, new_n20997);
nor_4  g18657(new_n21006, new_n21005, new_n17620);
not_3  g18658(new_n21007, new_n21006);
not_3  g18659(new_n21008_1, new_n21005);
nor_4  g18660(new_n21009, new_n21008_1, n25586);
nor_4  g18661(new_n21010, new_n21009, new_n21006);
not_3  g18662(new_n21011, n25751);
not_3  g18663(new_n21012, new_n20985);
xnor_3 g18664(new_n21013, new_n20995, new_n21012);
nor_4  g18665(new_n21014, new_n21013, new_n21011);
not_3  g18666(new_n21015, new_n21014);
xnor_3 g18667(new_n21016, new_n21013, new_n21011);
not_3  g18668(new_n21017_1, new_n21016);
xnor_3 g18669(new_n21018, new_n20993, new_n20992);
nand_4 g18670(new_n21019, new_n21018, new_n17572);
not_3  g18671(new_n21020, new_n21019);
xnor_3 g18672(new_n21021, new_n21018, new_n17572);
nor_4  g18673(new_n21022, new_n19627, n7917);
xnor_3 g18674(new_n21023, new_n19627, n7917);
nor_4  g18675(new_n21024, new_n19676, new_n19670);
nor_4  g18676(new_n21025, new_n21024, new_n19630);
nor_4  g18677(new_n21026, new_n21025, new_n21023);
nor_4  g18678(new_n21027, new_n21026, new_n21022);
nor_4  g18679(new_n21028, new_n21027, new_n21021);
nor_4  g18680(new_n21029, new_n21028, new_n21020);
nand_4 g18681(new_n21030, new_n21029, new_n21017_1);
nand_4 g18682(new_n21031, new_n21030, new_n21015);
nand_4 g18683(new_n21032, new_n21031, new_n21010);
nand_4 g18684(new_n21033, new_n21032, new_n21007);
not_3  g18685(new_n21034_1, new_n20999);
nor_4  g18686(new_n21035, new_n21034_1, n4514);
nor_4  g18687(new_n21036, new_n21001, new_n20997);
and_4  g18688(new_n21037, new_n21036, new_n21035);
not_3  g18689(new_n21038, new_n21037);
nor_4  g18690(new_n21039, new_n21038, new_n21033);
not_3  g18691(new_n21040, new_n21035);
xnor_3 g18692(new_n21041, new_n21036, new_n21040);
nor_4  g18693(new_n21042, new_n21041, new_n21003);
nand_4 g18694(new_n21043, new_n21042, new_n21033);
nor_4  g18695(new_n21044, new_n21043, new_n21037);
nor_4  g18696(new_n21045, new_n21044, new_n21039);
nor_4  g18697(new_n21046_1, new_n21045, new_n20979);
xnor_3 g18698(new_n21047, new_n21042, new_n21033);
xnor_3 g18699(new_n21048, new_n20978, new_n20968);
not_3  g18700(new_n21049, new_n21048);
nor_4  g18701(new_n21050, new_n21049, new_n21047);
not_3  g18702(new_n21051, new_n21050);
xnor_3 g18703(new_n21052, new_n21048, new_n21047);
not_3  g18704(new_n21053, new_n21021);
not_3  g18705(new_n21054, new_n21022);
nand_4 g18706(new_n21055, new_n19667, new_n19628);
nand_4 g18707(new_n21056, new_n21055, new_n21054);
nand_4 g18708(new_n21057, new_n21056, new_n21053);
nand_4 g18709(new_n21058, new_n21057, new_n21019);
nor_4  g18710(new_n21059, new_n21058, new_n21016);
nor_4  g18711(new_n21060, new_n21059, new_n21014);
xnor_3 g18712(new_n21061, new_n21060, new_n21010);
nor_4  g18713(new_n21062_1, new_n20975, new_n20972);
nor_4  g18714(new_n21063, new_n21062_1, new_n20977);
not_3  g18715(new_n21064, new_n21063);
nand_4 g18716(new_n21065, new_n21064, new_n21061);
not_3  g18717(new_n21066, new_n21065);
nor_4  g18718(new_n21067, new_n21064, new_n21061);
nor_4  g18719(new_n21068, new_n21067, new_n21066);
xnor_3 g18720(new_n21069, new_n21058, new_n21017_1);
nand_4 g18721(new_n21070, new_n21069, new_n8043);
not_3  g18722(new_n21071, new_n21070);
nor_4  g18723(new_n21072, new_n21069, new_n8043);
nor_4  g18724(new_n21073, new_n21072, new_n21071);
nor_4  g18725(new_n21074, new_n21056, new_n21053);
nor_4  g18726(new_n21075, new_n21074, new_n21028);
not_3  g18727(new_n21076, new_n21075);
nand_4 g18728(new_n21077, new_n21076, new_n8137);
nand_4 g18729(new_n21078_1, new_n19668, new_n8142);
nand_4 g18730(new_n21079, new_n19719, new_n19669);
nand_4 g18731(new_n21080, new_n21079, new_n21078_1);
xnor_3 g18732(new_n21081, new_n21075, new_n8137);
nand_4 g18733(new_n21082, new_n21081, new_n21080);
nand_4 g18734(new_n21083, new_n21082, new_n21077);
nand_4 g18735(new_n21084, new_n21083, new_n21073);
nand_4 g18736(new_n21085, new_n21084, new_n21070);
nand_4 g18737(new_n21086, new_n21085, new_n21068);
nand_4 g18738(new_n21087, new_n21086, new_n21065);
nand_4 g18739(new_n21088, new_n21087, new_n21052);
nand_4 g18740(new_n21089, new_n21088, new_n21051);
nor_4  g18741(new_n21090, new_n21089, new_n21046_1);
not_3  g18742(new_n21091, new_n21039);
nand_4 g18743(new_n21092, new_n21045, new_n20979);
nand_4 g18744(new_n21093_1, new_n21092, new_n21091);
nor_4  g18745(n4205, new_n21093_1, new_n21090);
nand_4 g18746(new_n21095_1, new_n15992, new_n5606);
xor_3  g18747(new_n21096, new_n21095_1, n2659);
not_3  g18748(new_n21097, new_n21096);
xor_3  g18749(new_n21098, new_n21097, n18444);
xor_3  g18750(new_n21099, new_n15992, new_n5606);
nor_4  g18751(new_n21100, new_n21099, n24638);
xnor_3 g18752(new_n21101, new_n21099, n24638);
nor_4  g18753(new_n21102, new_n16032, new_n16000);
nor_4  g18754(new_n21103, new_n21102, new_n15998);
nor_4  g18755(new_n21104, new_n21103, new_n21101);
nor_4  g18756(new_n21105, new_n21104, new_n21100);
not_3  g18757(new_n21106, new_n21105);
xnor_3 g18758(new_n21107, new_n21106, new_n21098);
xnor_3 g18759(new_n21108, new_n21107, new_n9151);
xnor_3 g18760(new_n21109, new_n21103, new_n21101);
nand_4 g18761(new_n21110, new_n21109, new_n9161);
not_3  g18762(new_n21111, new_n21110);
nor_4  g18763(new_n21112, new_n21109, new_n9161);
nor_4  g18764(new_n21113, new_n21112, new_n21111);
nor_4  g18765(new_n21114, new_n16033, new_n9179);
nor_4  g18766(new_n21115, new_n16062_1, new_n21114);
nand_4 g18767(new_n21116, new_n21115, new_n21113);
nand_4 g18768(new_n21117, new_n21116, new_n21110);
nand_4 g18769(new_n21118, new_n21117, new_n21108);
not_3  g18770(new_n21119, new_n21118);
nor_4  g18771(new_n21120, new_n21117, new_n21108);
nor_4  g18772(new_n21121, new_n21120, new_n21119);
xor_3  g18773(new_n21122, n21997, new_n9840);
nand_4 g18774(new_n21123_1, new_n10137, n23923);
xor_3  g18775(new_n21124, n25119, new_n8258);
nand_4 g18776(new_n21125, new_n10139, n329);
nand_4 g18777(new_n21126, new_n16086, new_n16067);
nand_4 g18778(new_n21127, new_n21126, new_n21125);
nand_4 g18779(new_n21128, new_n21127, new_n21124);
nand_4 g18780(new_n21129, new_n21128, new_n21123_1);
xor_3  g18781(new_n21130, new_n21129, new_n21122);
xnor_3 g18782(new_n21131, new_n21130, new_n21121);
xor_3  g18783(new_n21132, new_n21127, new_n21124);
xnor_3 g18784(new_n21133, new_n21115, new_n21113);
not_3  g18785(new_n21134_1, new_n21133);
nand_4 g18786(new_n21135, new_n21134_1, new_n21132);
not_3  g18787(new_n21136, new_n21135);
xnor_3 g18788(new_n21137, new_n21134_1, new_n21132);
nor_4  g18789(new_n21138_1, new_n16087, new_n16066);
not_3  g18790(new_n21139, new_n21138_1);
not_3  g18791(new_n21140, new_n16087);
nor_4  g18792(new_n21141, new_n21140, new_n16065);
nor_4  g18793(new_n21142, new_n21138_1, new_n21141);
nand_4 g18794(new_n21143, new_n16136, new_n21142);
nand_4 g18795(new_n21144, new_n21143, new_n21139);
nor_4  g18796(new_n21145, new_n21144, new_n21137);
nor_4  g18797(new_n21146, new_n21145, new_n21136);
xor_3  g18798(n4215, new_n21146, new_n21131);
not_3  g18799(new_n21148, n3740);
nand_4 g18800(new_n21149, new_n17342, new_n9080);
not_3  g18801(new_n21150, new_n21149);
xor_3  g18802(new_n21151, new_n21150, new_n9076);
not_3  g18803(new_n21152, new_n21151);
nor_4  g18804(new_n21153, new_n21152, new_n21148);
nor_4  g18805(new_n21154_1, new_n21151, n3740);
nor_4  g18806(new_n21155, new_n21154_1, new_n21153);
nor_4  g18807(new_n21156, new_n17380, new_n17346);
nor_4  g18808(new_n21157_1, new_n21156, new_n17345);
xnor_3 g18809(new_n21158, new_n21157_1, new_n21155);
not_3  g18810(new_n21159, new_n21158);
not_3  g18811(new_n21160, n22626);
nor_4  g18812(new_n21161, new_n11598, n27089);
xor_3  g18813(new_n21162, new_n21161, new_n4853);
not_3  g18814(new_n21163, new_n21162);
nor_4  g18815(new_n21164, new_n21163, new_n21160);
nor_4  g18816(new_n21165, new_n21162, n22626);
nor_4  g18817(new_n21166, new_n21165, new_n21164);
not_3  g18818(new_n21167, n14440);
nand_4 g18819(new_n21168_1, new_n11600, new_n21167);
xor_3  g18820(new_n21169, new_n11600, new_n21167);
nand_4 g18821(new_n21170, new_n11603, new_n9036);
nand_4 g18822(new_n21171, new_n19273, new_n19269);
nand_4 g18823(new_n21172, new_n21171, new_n21170);
nand_4 g18824(new_n21173_1, new_n21172, new_n21169);
nand_4 g18825(new_n21174, new_n21173_1, new_n21168_1);
xnor_3 g18826(new_n21175, new_n21174, new_n21166);
xnor_3 g18827(new_n21176_1, new_n21175, new_n21159);
not_3  g18828(new_n21177, new_n21169);
xnor_3 g18829(new_n21178, new_n21172, new_n21177);
nor_4  g18830(new_n21179, new_n21178, new_n17382);
nand_4 g18831(new_n21180, new_n19274, new_n17389);
xnor_3 g18832(new_n21181, new_n19274, new_n17389);
not_3  g18833(new_n21182_1, new_n21181);
nand_4 g18834(new_n21183, new_n17395, new_n12784);
xnor_3 g18835(new_n21184, new_n17395, new_n12784);
not_3  g18836(new_n21185, new_n21184);
xnor_3 g18837(new_n21186, new_n12781, new_n12775);
nor_4  g18838(new_n21187, new_n17399, new_n21186);
not_3  g18839(new_n21188, new_n21187);
xnor_3 g18840(new_n21189, new_n17399, new_n21186);
nand_4 g18841(new_n21190, new_n17406, new_n12808);
xnor_3 g18842(new_n21191, new_n17406, new_n12807);
not_3  g18843(new_n21192, new_n11346);
nand_4 g18844(new_n21193_1, new_n11372, new_n11351);
nand_4 g18845(new_n21194, new_n21193_1, new_n21192);
nand_4 g18846(new_n21195, new_n21194, new_n21191);
nand_4 g18847(new_n21196, new_n21195, new_n21190);
nor_4  g18848(new_n21197, new_n21196, new_n21189);
not_3  g18849(new_n21198, new_n21197);
nand_4 g18850(new_n21199, new_n21198, new_n21188);
nand_4 g18851(new_n21200, new_n21199, new_n21185);
nand_4 g18852(new_n21201, new_n21200, new_n21183);
nand_4 g18853(new_n21202, new_n21201, new_n21182_1);
nand_4 g18854(new_n21203_1, new_n21202, new_n21180);
xnor_3 g18855(new_n21204, new_n21172, new_n21169);
nor_4  g18856(new_n21205, new_n21204, new_n17381);
nor_4  g18857(new_n21206, new_n21205, new_n21179);
not_3  g18858(new_n21207, new_n21206);
nor_4  g18859(new_n21208, new_n21207, new_n21203_1);
nor_4  g18860(new_n21209, new_n21208, new_n21179);
xnor_3 g18861(new_n21210, new_n21209, new_n21176_1);
not_3  g18862(new_n21211, n23166);
nor_4  g18863(new_n21212, new_n18307, n10611);
not_3  g18864(new_n21213, new_n21212);
nor_4  g18865(new_n21214, new_n21213, n3164);
not_3  g18866(new_n21215, new_n21214);
nor_4  g18867(new_n21216, new_n21215, n11356);
nand_4 g18868(new_n21217, new_n21216, new_n10893);
nor_4  g18869(new_n21218, new_n21217, n6381);
not_3  g18870(new_n21219, new_n21218);
nor_4  g18871(new_n21220, new_n21219, n10577);
xor_3  g18872(new_n21221, new_n21220, new_n21211);
not_3  g18873(new_n21222_1, new_n21221);
nor_4  g18874(new_n21223, new_n21222_1, new_n9258);
nor_4  g18875(new_n21224, new_n21221, n9554);
nor_4  g18876(new_n21225_1, new_n21224, new_n21223);
xor_3  g18877(new_n21226_1, new_n21218, new_n10886);
nor_4  g18878(new_n21227, new_n21226_1, n26408);
not_3  g18879(new_n21228, n26408);
not_3  g18880(new_n21229, new_n21226_1);
xor_3  g18881(new_n21230, new_n21229, new_n21228);
not_3  g18882(new_n21231, n18227);
xor_3  g18883(new_n21232, new_n21217, n6381);
not_3  g18884(new_n21233, new_n21232);
nand_4 g18885(new_n21234, new_n21233, new_n21231);
xor_3  g18886(new_n21235, new_n21233, new_n21231);
xor_3  g18887(new_n21236, new_n21216, new_n10893);
not_3  g18888(new_n21237, new_n21236);
nand_4 g18889(new_n21238_1, new_n21237, new_n5471);
xor_3  g18890(new_n21239, new_n21237, new_n5471);
not_3  g18891(new_n21240, n11630);
xor_3  g18892(new_n21241, new_n21215, n11356);
not_3  g18893(new_n21242, new_n21241);
nand_4 g18894(new_n21243, new_n21242, new_n21240);
xor_3  g18895(new_n21244, new_n21212, new_n10898);
nor_4  g18896(new_n21245, new_n21244, n13453);
not_3  g18897(new_n21246, new_n21245);
not_3  g18898(new_n21247, new_n21244);
xor_3  g18899(new_n21248, new_n21247, new_n9246_1);
nor_4  g18900(new_n21249, new_n18325, new_n18311_1);
nor_4  g18901(new_n21250, new_n21249, new_n18310_1);
nand_4 g18902(new_n21251, new_n21250, new_n21248);
nand_4 g18903(new_n21252, new_n21251, new_n21246);
xor_3  g18904(new_n21253, new_n21242, new_n21240);
nand_4 g18905(new_n21254_1, new_n21253, new_n21252);
nand_4 g18906(new_n21255, new_n21254_1, new_n21243);
nand_4 g18907(new_n21256, new_n21255, new_n21239);
nand_4 g18908(new_n21257, new_n21256, new_n21238_1);
nand_4 g18909(new_n21258, new_n21257, new_n21235);
nand_4 g18910(new_n21259, new_n21258, new_n21234);
nand_4 g18911(new_n21260, new_n21259, new_n21230);
not_3  g18912(new_n21261, new_n21260);
nor_4  g18913(new_n21262, new_n21261, new_n21227);
xnor_3 g18914(new_n21263, new_n21262, new_n21225_1);
not_3  g18915(new_n21264, new_n21263);
xnor_3 g18916(new_n21265, new_n21264, new_n21210);
xnor_3 g18917(new_n21266, new_n21259, new_n21230);
not_3  g18918(new_n21267, new_n21266);
xnor_3 g18919(new_n21268, new_n21207, new_n21203_1);
nand_4 g18920(new_n21269, new_n21268, new_n21267);
xnor_3 g18921(new_n21270, new_n21268, new_n21267);
not_3  g18922(new_n21271, new_n21270);
xnor_3 g18923(new_n21272, new_n21257, new_n21235);
not_3  g18924(new_n21273, new_n21272);
xnor_3 g18925(new_n21274, new_n21201, new_n21181);
nand_4 g18926(new_n21275, new_n21274, new_n21273);
xnor_3 g18927(new_n21276_1, new_n21274, new_n21272);
not_3  g18928(new_n21277, new_n21239);
xnor_3 g18929(new_n21278, new_n21255, new_n21277);
xnor_3 g18930(new_n21279, new_n21199, new_n21184);
nand_4 g18931(new_n21280, new_n21279, new_n21278);
not_3  g18932(new_n21281, new_n21279);
xnor_3 g18933(new_n21282, new_n21281, new_n21278);
xnor_3 g18934(new_n21283, new_n21196, new_n21189);
xnor_3 g18935(new_n21284, new_n21253, new_n21252);
nor_4  g18936(new_n21285, new_n21284, new_n21283);
not_3  g18937(new_n21286, new_n21285);
not_3  g18938(new_n21287_1, new_n21283);
not_3  g18939(new_n21288, new_n21284);
nor_4  g18940(new_n21289, new_n21288, new_n21287_1);
nor_4  g18941(new_n21290, new_n21289, new_n21285);
not_3  g18942(new_n21291, new_n21248);
xnor_3 g18943(new_n21292, new_n21250, new_n21291);
xnor_3 g18944(new_n21293, new_n21194, new_n21191);
nand_4 g18945(new_n21294, new_n21293, new_n21292);
not_3  g18946(new_n21295, new_n21293);
xnor_3 g18947(new_n21296, new_n21295, new_n21292);
not_3  g18948(new_n21297, new_n11373);
nor_4  g18949(new_n21298_1, new_n18326, new_n21297);
not_3  g18950(new_n21299, new_n21298_1);
not_3  g18951(new_n21300, new_n18326);
nor_4  g18952(new_n21301, new_n21300, new_n11373);
nor_4  g18953(new_n21302_1, new_n21301, new_n21298_1);
nor_4  g18954(new_n21303, new_n18328, new_n11397);
xnor_3 g18955(new_n21304, new_n18328, new_n11397);
nor_4  g18956(new_n21305, new_n18335, new_n11408);
not_3  g18957(new_n21306, new_n18338);
nor_4  g18958(new_n21307, new_n21306, new_n11401);
not_3  g18959(new_n21308, new_n21307);
xnor_3 g18960(new_n21309, new_n18335, new_n11408);
nor_4  g18961(new_n21310, new_n21309, new_n21308);
nor_4  g18962(new_n21311, new_n21310, new_n21305);
nor_4  g18963(new_n21312, new_n21311, new_n21304);
nor_4  g18964(new_n21313, new_n21312, new_n21303);
nand_4 g18965(new_n21314, new_n21313, new_n21302_1);
nand_4 g18966(new_n21315, new_n21314, new_n21299);
nand_4 g18967(new_n21316, new_n21315, new_n21296);
nand_4 g18968(new_n21317_1, new_n21316, new_n21294);
nand_4 g18969(new_n21318, new_n21317_1, new_n21290);
nand_4 g18970(new_n21319, new_n21318, new_n21286);
nand_4 g18971(new_n21320, new_n21319, new_n21282);
nand_4 g18972(new_n21321, new_n21320, new_n21280);
nand_4 g18973(new_n21322, new_n21321, new_n21276_1);
nand_4 g18974(new_n21323, new_n21322, new_n21275);
nand_4 g18975(new_n21324, new_n21323, new_n21271);
nand_4 g18976(new_n21325, new_n21324, new_n21269);
nor_4  g18977(new_n21326, new_n21325, new_n21265);
not_3  g18978(new_n21327, new_n21265);
not_3  g18979(new_n21328, new_n21325);
nor_4  g18980(new_n21329, new_n21328, new_n21327);
nor_4  g18981(n4221, new_n21329, new_n21326);
xnor_3 g18982(new_n21331, new_n12688, new_n21231);
not_3  g18983(new_n21332, new_n21331);
nand_4 g18984(new_n21333, new_n12690, n7377);
xnor_3 g18985(new_n21334, new_n12690, new_n5471);
nand_4 g18986(new_n21335, new_n12694, n11630);
nand_4 g18987(new_n21336, new_n12697, n13453);
nand_4 g18988(new_n21337, new_n15652_1, new_n15646);
nand_4 g18989(new_n21338, new_n21337, new_n21336);
xnor_3 g18990(new_n21339, new_n12694, new_n21240);
nand_4 g18991(new_n21340, new_n21339, new_n21338);
nand_4 g18992(new_n21341, new_n21340, new_n21335);
nand_4 g18993(new_n21342, new_n21341, new_n21334);
nand_4 g18994(new_n21343, new_n21342, new_n21333);
xnor_3 g18995(new_n21344, new_n21343, new_n21332);
xnor_3 g18996(new_n21345, new_n21344, new_n19802);
not_3  g18997(new_n21346, new_n21334);
xnor_3 g18998(new_n21347, new_n21341, new_n21346);
nand_4 g18999(new_n21348, new_n21347, new_n10136);
xnor_3 g19000(new_n21349_1, new_n21347, new_n10135);
not_3  g19001(new_n21350, new_n21339);
xnor_3 g19002(new_n21351, new_n21350, new_n21338);
nand_4 g19003(new_n21352, new_n21351, new_n10173);
not_3  g19004(new_n21353, new_n21352);
nor_4  g19005(new_n21354, new_n21351, new_n10173);
nor_4  g19006(new_n21355, new_n21354, new_n21353);
nand_4 g19007(new_n21356, new_n15654, new_n10181);
not_3  g19008(new_n21357, new_n21356);
nor_4  g19009(new_n21358, new_n15654, new_n10181);
nor_4  g19010(new_n21359, new_n21358, new_n21357);
nand_4 g19011(new_n21360, new_n10188, new_n7777);
not_3  g19012(new_n21361, new_n21360);
nor_4  g19013(new_n21362, new_n10188, new_n7777);
nor_4  g19014(new_n21363, new_n21362, new_n21361);
nand_4 g19015(new_n21364, new_n10196, new_n7830_1);
not_3  g19016(new_n21365_1, new_n21364);
nor_4  g19017(new_n21366, new_n10196, new_n7830_1);
nor_4  g19018(new_n21367_1, new_n21366, new_n21365_1);
not_3  g19019(new_n21368, new_n7835);
nor_4  g19020(new_n21369, new_n10203, new_n21368);
not_3  g19021(new_n21370, new_n21369);
nor_4  g19022(new_n21371, new_n10207, new_n7841_1);
nor_4  g19023(new_n21372, new_n19833, new_n7835);
nor_4  g19024(new_n21373, new_n21372, new_n21369);
nand_4 g19025(new_n21374, new_n21373, new_n21371);
nand_4 g19026(new_n21375, new_n21374, new_n21370);
nand_4 g19027(new_n21376, new_n21375, new_n21367_1);
nand_4 g19028(new_n21377, new_n21376, new_n21364);
nand_4 g19029(new_n21378, new_n21377, new_n21363);
nand_4 g19030(new_n21379, new_n21378, new_n21360);
nand_4 g19031(new_n21380, new_n21379, new_n21359);
nand_4 g19032(new_n21381, new_n21380, new_n21356);
nand_4 g19033(new_n21382, new_n21381, new_n21355);
nand_4 g19034(new_n21383, new_n21382, new_n21352);
nand_4 g19035(new_n21384, new_n21383, new_n21349_1);
nand_4 g19036(new_n21385, new_n21384, new_n21348);
xor_3  g19037(n4224, new_n21385, new_n21345);
xor_3  g19038(n4231, new_n12859, new_n12858);
not_3  g19039(new_n21388, new_n14345_1);
nor_4  g19040(new_n21389, new_n17171, new_n15250);
nor_4  g19041(new_n21390, new_n17169, n9934);
nor_4  g19042(new_n21391, new_n21390, new_n21389);
nor_4  g19043(new_n21392, new_n17176, n18496);
nor_4  g19044(new_n21393, new_n20540, new_n20533_1);
nor_4  g19045(new_n21394, new_n21393, new_n21392);
xnor_3 g19046(new_n21395, new_n21394, new_n21391);
not_3  g19047(new_n21396_1, new_n21395);
nor_4  g19048(new_n21397, new_n21396_1, n2979);
nor_4  g19049(new_n21398_1, new_n21395, new_n6863_1);
nor_4  g19050(new_n21399_1, new_n21398_1, new_n21397);
not_3  g19051(new_n21400, new_n21399_1);
not_3  g19052(new_n21401, new_n20545);
nor_4  g19053(new_n21402, new_n20555, new_n21401);
nor_4  g19054(new_n21403, new_n21402, new_n20544);
xnor_3 g19055(new_n21404_1, new_n21403, new_n21400);
xnor_3 g19056(new_n21405, new_n21404_1, new_n21388);
not_3  g19057(new_n21406, new_n20557);
nor_4  g19058(new_n21407, new_n21406, new_n14348);
nor_4  g19059(new_n21408, new_n20574, new_n20558);
nor_4  g19060(new_n21409, new_n21408, new_n21407);
xnor_3 g19061(n4266, new_n21409, new_n21405);
not_3  g19062(new_n21411, new_n8156);
xor_3  g19063(n4340, new_n8190, new_n21411);
xnor_3 g19064(new_n21413, new_n20067, new_n6982);
xnor_3 g19065(new_n21414, new_n21413, new_n15798);
nand_4 g19066(new_n21415, new_n20075, new_n20071);
xnor_3 g19067(new_n21416, new_n21415, new_n21414);
not_3  g19068(new_n21417, new_n21416);
xnor_3 g19069(new_n21418, new_n21417, new_n5712);
nor_4  g19070(new_n21419, new_n20077_1, new_n20064);
nor_4  g19071(new_n21420, new_n21419, new_n20062);
xor_3  g19072(n4374, new_n21420, new_n21418);
xnor_3 g19073(n4401, new_n13454, new_n13389);
not_3  g19074(new_n21423, new_n15717);
xor_3  g19075(n4424, new_n15720, new_n21423);
not_3  g19076(new_n21425, n1881);
nor_4  g19077(new_n21426, new_n12952, new_n21425);
xnor_3 g19078(new_n21427, new_n12951, n1881);
nor_4  g19079(new_n21428, new_n12943, n5834);
not_3  g19080(new_n21429, new_n21428);
not_3  g19081(new_n21430, n5834);
xnor_3 g19082(new_n21431, new_n12942_1, new_n21430);
not_3  g19083(new_n21432, new_n21431);
not_3  g19084(new_n21433, n13851);
nor_4  g19085(new_n21434, new_n12935, new_n21433);
nor_4  g19086(new_n21435, new_n12936, n13851);
nor_4  g19087(new_n21436, new_n21435, new_n21434);
nand_4 g19088(new_n21437, new_n12924, n24937);
nand_4 g19089(new_n21438, new_n19933, new_n19923_1);
nand_4 g19090(new_n21439, new_n21438, new_n21437);
nand_4 g19091(new_n21440, new_n21439, new_n21436);
not_3  g19092(new_n21441, new_n21440);
nor_4  g19093(new_n21442, new_n21441, new_n21434);
nand_4 g19094(new_n21443, new_n21442, new_n21432);
nand_4 g19095(new_n21444, new_n21443, new_n21429);
nor_4  g19096(new_n21445, new_n21444, new_n21427);
nor_4  g19097(new_n21446_1, new_n21445, new_n21426);
nor_4  g19098(new_n21447, n8827, n4306);
nor_4  g19099(new_n21448, new_n12950, new_n12946);
nor_4  g19100(new_n21449, new_n21448, new_n21447);
not_3  g19101(new_n21450, new_n21449);
nor_4  g19102(new_n21451, new_n21450, new_n21446_1);
not_3  g19103(new_n21452, new_n21446_1);
nor_4  g19104(new_n21453, new_n21449, new_n21452);
nor_4  g19105(new_n21454, new_n21453, new_n21451);
nor_4  g19106(new_n21455, new_n21454, new_n12020);
not_3  g19107(new_n21456, new_n21454);
nor_4  g19108(new_n21457, new_n21456, new_n12018);
nor_4  g19109(new_n21458, new_n21457, new_n21455);
not_3  g19110(new_n21459, new_n21427);
not_3  g19111(new_n21460, new_n21444);
nor_4  g19112(new_n21461, new_n21460, new_n21459);
nor_4  g19113(new_n21462, new_n21461, new_n21445);
not_3  g19114(new_n21463, new_n21462);
nor_4  g19115(new_n21464, new_n21463, new_n12025);
not_3  g19116(new_n21465, new_n21464);
nor_4  g19117(new_n21466, new_n21462, new_n12024);
nor_4  g19118(new_n21467, new_n21466, new_n21464);
not_3  g19119(new_n21468, new_n21443);
nor_4  g19120(new_n21469, new_n21442, new_n21432);
nor_4  g19121(new_n21470, new_n21469, new_n21468);
nor_4  g19122(new_n21471_1, new_n21470, new_n12029);
not_3  g19123(new_n21472_1, new_n21471_1);
xnor_3 g19124(new_n21473, new_n21439, new_n21436);
nand_4 g19125(new_n21474, new_n21473, new_n12035);
xnor_3 g19126(new_n21475, new_n21473, new_n12035);
not_3  g19127(new_n21476, new_n21475);
nand_4 g19128(new_n21477, new_n19934, new_n12040);
nand_4 g19129(new_n21478, new_n19959, new_n19936);
nand_4 g19130(new_n21479, new_n21478, new_n21477);
nand_4 g19131(new_n21480, new_n21479, new_n21476);
nand_4 g19132(new_n21481, new_n21480, new_n21474);
not_3  g19133(new_n21482, new_n21481);
not_3  g19134(new_n21483, new_n21470);
nor_4  g19135(new_n21484, new_n21483, new_n12031);
nor_4  g19136(new_n21485, new_n21484, new_n21471_1);
nand_4 g19137(new_n21486, new_n21485, new_n21482);
nand_4 g19138(new_n21487, new_n21486, new_n21472_1);
nand_4 g19139(new_n21488, new_n21487, new_n21467);
nand_4 g19140(new_n21489_1, new_n21488, new_n21465);
xnor_3 g19141(n4432, new_n21489_1, new_n21458);
not_3  g19142(new_n21491, new_n17959_1);
xor_3  g19143(n4441, new_n21491, new_n17958);
nor_4  g19144(new_n21493, n27120, n23065);
nand_4 g19145(new_n21494, new_n21493, new_n10272);
nor_4  g19146(new_n21495, new_n21494, n25370);
not_3  g19147(new_n21496, new_n21495);
nor_4  g19148(new_n21497, new_n21496, n19472);
not_3  g19149(new_n21498, new_n21497);
nor_4  g19150(new_n21499, new_n21498, n19042);
not_3  g19151(new_n21500, new_n21499);
nor_4  g19152(new_n21501, new_n21500, n1293);
xor_3  g19153(new_n21502, new_n21501, new_n8045);
not_3  g19154(new_n21503, new_n21502);
nor_4  g19155(new_n21504, new_n21503, new_n20627);
not_3  g19156(new_n21505, new_n20627);
nor_4  g19157(new_n21506, new_n21502, new_n21505);
nor_4  g19158(new_n21507, new_n21506, new_n21504);
xor_3  g19159(new_n21508, new_n21499, new_n10335);
nor_4  g19160(new_n21509, new_n21508, new_n20631);
xnor_3 g19161(new_n21510, new_n21508, new_n20631);
xor_3  g19162(new_n21511, new_n21497, new_n10337);
nor_4  g19163(new_n21512, new_n21511, new_n20647);
xor_3  g19164(new_n21513, new_n21495, new_n10265);
nor_4  g19165(new_n21514, new_n21513, new_n10263);
not_3  g19166(new_n21515, new_n21513);
nor_4  g19167(new_n21516, new_n21515, new_n10266);
nor_4  g19168(new_n21517, new_n21516, new_n21514);
not_3  g19169(new_n21518, new_n21517);
xor_3  g19170(new_n21519, new_n21494, n25370);
not_3  g19171(new_n21520, new_n21519);
nor_4  g19172(new_n21521, new_n21520, new_n10269);
not_3  g19173(new_n21522, new_n21521);
nor_4  g19174(new_n21523, new_n21519, new_n10270);
nor_4  g19175(new_n21524, new_n21523, new_n21521);
not_3  g19176(new_n21525_1, new_n10273);
xor_3  g19177(new_n21526, new_n21493, new_n10272);
nor_4  g19178(new_n21527, new_n21526, new_n21525_1);
xnor_3 g19179(new_n21528, new_n21526, new_n21525_1);
xor_3  g19180(new_n21529, n27120, n23065);
nor_4  g19181(new_n21530, new_n21529, new_n10281);
nor_4  g19182(new_n21531, new_n21530, new_n10285);
nor_4  g19183(new_n21532, new_n21531, new_n21528);
nor_4  g19184(new_n21533, new_n21532, new_n21527);
nand_4 g19185(new_n21534, new_n21533, new_n21524);
nand_4 g19186(new_n21535, new_n21534, new_n21522);
nor_4  g19187(new_n21536, new_n21535, new_n21518);
nor_4  g19188(new_n21537, new_n21536, new_n21514);
not_3  g19189(new_n21538_1, new_n21511);
nor_4  g19190(new_n21539, new_n21538_1, new_n20641);
nor_4  g19191(new_n21540, new_n21539, new_n21512);
not_3  g19192(new_n21541, new_n21540);
nor_4  g19193(new_n21542, new_n21541, new_n21537);
nor_4  g19194(new_n21543, new_n21542, new_n21512);
nor_4  g19195(new_n21544, new_n21543, new_n21510);
nor_4  g19196(new_n21545, new_n21544, new_n21509);
xnor_3 g19197(new_n21546, new_n21545, new_n21507);
nor_4  g19198(new_n21547, new_n14550, n26318);
xor_3  g19199(new_n21548, new_n21547, n3710);
xnor_3 g19200(new_n21549_1, new_n21548, new_n6159);
not_3  g19201(new_n21550, new_n14551);
nand_4 g19202(new_n21551, new_n21550, new_n6167);
nand_4 g19203(new_n21552, new_n14585, new_n14552);
nand_4 g19204(new_n21553, new_n21552, new_n21551);
nor_4  g19205(new_n21554, new_n21553, new_n21549_1);
nand_4 g19206(new_n21555, new_n21553, new_n21549_1);
not_3  g19207(new_n21556, new_n21555);
nor_4  g19208(new_n21557, new_n21556, new_n21554);
xnor_3 g19209(new_n21558, new_n21557, new_n21546);
not_3  g19210(new_n21559, new_n21510);
not_3  g19211(new_n21560, new_n21512);
not_3  g19212(new_n21561, new_n21514);
not_3  g19213(new_n21562, new_n21536);
nand_4 g19214(new_n21563, new_n21562, new_n21561);
nand_4 g19215(new_n21564, new_n21540, new_n21563);
nand_4 g19216(new_n21565, new_n21564, new_n21560);
nor_4  g19217(new_n21566, new_n21565, new_n21559);
nor_4  g19218(new_n21567, new_n21566, new_n21544);
nand_4 g19219(new_n21568, new_n21567, new_n14627);
xnor_3 g19220(new_n21569, new_n21567, new_n14586);
xnor_3 g19221(new_n21570, new_n21540, new_n21563);
nor_4  g19222(new_n21571, new_n21570, new_n14632);
not_3  g19223(new_n21572, new_n21571);
not_3  g19224(new_n21573, new_n21570);
nor_4  g19225(new_n21574, new_n21573, new_n14633_1);
nor_4  g19226(new_n21575, new_n21574, new_n21571);
not_3  g19227(new_n21576, new_n21535);
nor_4  g19228(new_n21577, new_n21576, new_n21517);
nor_4  g19229(new_n21578, new_n21577, new_n21536);
nor_4  g19230(new_n21579, new_n21578, new_n14637);
xnor_3 g19231(new_n21580, new_n21533, new_n21524);
nand_4 g19232(new_n21581, new_n21580, new_n14643);
xnor_3 g19233(new_n21582, new_n21580, new_n14642);
not_3  g19234(new_n21583, new_n21528);
not_3  g19235(new_n21584, new_n21531);
nor_4  g19236(new_n21585, new_n21584, new_n21583);
nor_4  g19237(new_n21586, new_n21585, new_n21532);
nor_4  g19238(new_n21587, new_n21586, new_n14655);
not_3  g19239(new_n21588, new_n21586);
nor_4  g19240(new_n21589, new_n21588, new_n14650);
xnor_3 g19241(new_n21590, new_n21529, new_n10286);
nand_4 g19242(new_n21591, new_n21590, new_n14671);
nand_4 g19243(new_n21592, new_n14669, new_n10309);
not_3  g19244(new_n21593, new_n21591);
nor_4  g19245(new_n21594, new_n21590, new_n14671);
nor_4  g19246(new_n21595, new_n21594, new_n21593);
nand_4 g19247(new_n21596, new_n21595, new_n21592);
nand_4 g19248(new_n21597, new_n21596, new_n21591);
nor_4  g19249(new_n21598, new_n21597, new_n21589);
nor_4  g19250(new_n21599_1, new_n21598, new_n21587);
nand_4 g19251(new_n21600, new_n21599_1, new_n21582);
nand_4 g19252(new_n21601, new_n21600, new_n21581);
xnor_3 g19253(new_n21602, new_n21578, new_n14637);
nor_4  g19254(new_n21603, new_n21602, new_n21601);
nor_4  g19255(new_n21604, new_n21603, new_n21579);
nand_4 g19256(new_n21605, new_n21604, new_n21575);
nand_4 g19257(new_n21606, new_n21605, new_n21572);
nand_4 g19258(new_n21607, new_n21606, new_n21569);
nand_4 g19259(new_n21608, new_n21607, new_n21568);
xnor_3 g19260(n4451, new_n21608, new_n21558);
not_3  g19261(new_n21610, n6659);
xor_3  g19262(new_n21611, n25494, new_n21610);
not_3  g19263(new_n21612, new_n21611);
nor_4  g19264(new_n21613, new_n19420, n10117);
xor_3  g19265(new_n21614, new_n19420, n10117);
nand_4 g19266(new_n21615_1, new_n13566, n11455);
xor_3  g19267(new_n21616, n13460, new_n19425);
nand_4 g19268(new_n21617, new_n13569, n3945);
xor_3  g19269(new_n21618, n6104, new_n19429);
nand_4 g19270(new_n21619, n5255, new_n3693);
nand_4 g19271(new_n21620, new_n5963, new_n5940);
nand_4 g19272(new_n21621, new_n21620, new_n21619);
nand_4 g19273(new_n21622, new_n21621, new_n21618);
nand_4 g19274(new_n21623, new_n21622, new_n21617);
nand_4 g19275(new_n21624, new_n21623, new_n21616);
nand_4 g19276(new_n21625, new_n21624, new_n21615_1);
nand_4 g19277(new_n21626, new_n21625, new_n21614);
not_3  g19278(new_n21627, new_n21626);
nor_4  g19279(new_n21628_1, new_n21627, new_n21613);
xor_3  g19280(new_n21629, new_n21628_1, new_n21612);
nor_4  g19281(new_n21630, new_n21629, new_n15942);
not_3  g19282(new_n21631, new_n21629);
nor_4  g19283(new_n21632, new_n21631, new_n15941);
nor_4  g19284(new_n21633, new_n21632, new_n21630);
xor_3  g19285(new_n21634, new_n21625, new_n21614);
nor_4  g19286(new_n21635, new_n21634, new_n15949);
not_3  g19287(new_n21636, new_n21634);
nor_4  g19288(new_n21637_1, new_n21636, new_n15950);
nor_4  g19289(new_n21638, new_n21637_1, new_n21635);
not_3  g19290(new_n21639, new_n21638);
xor_3  g19291(new_n21640, new_n21623, new_n21616);
nor_4  g19292(new_n21641, new_n21640, new_n15955);
xnor_3 g19293(new_n21642, new_n21640, new_n15955);
xor_3  g19294(new_n21643, new_n21621, new_n21618);
not_3  g19295(new_n21644, new_n21643);
nor_4  g19296(new_n21645_1, new_n21644, new_n15962);
not_3  g19297(new_n21646, new_n21645_1);
nor_4  g19298(new_n21647, new_n21643, new_n15961);
nor_4  g19299(new_n21648, new_n21647, new_n21645_1);
not_3  g19300(new_n21649_1, new_n5964_1);
nor_4  g19301(new_n21650, new_n21649_1, new_n15967_1);
not_3  g19302(new_n21651, new_n21650);
not_3  g19303(new_n21652, new_n5965);
nor_4  g19304(new_n21653, new_n14401, new_n5970);
nor_4  g19305(new_n21654_1, new_n21653, new_n5968);
nand_4 g19306(new_n21655, new_n21654_1, new_n21652);
nand_4 g19307(new_n21656, new_n21655, new_n21651);
nand_4 g19308(new_n21657, new_n21656, new_n21648);
nand_4 g19309(new_n21658, new_n21657, new_n21646);
nor_4  g19310(new_n21659, new_n21658, new_n21642);
nor_4  g19311(new_n21660, new_n21659, new_n21641);
nor_4  g19312(new_n21661, new_n21660, new_n21639);
nor_4  g19313(new_n21662, new_n21661, new_n21635);
nand_4 g19314(new_n21663, new_n21662, new_n21633);
not_3  g19315(new_n21664, new_n21663);
nor_4  g19316(new_n21665_1, new_n21662, new_n21633);
nor_4  g19317(n4476, new_n21665_1, new_n21664);
not_3  g19318(new_n21667, new_n4433);
nor_4  g19319(new_n21668, new_n21667, n12398);
not_3  g19320(new_n21669, new_n21668);
nor_4  g19321(new_n21670, new_n21669, n21317);
not_3  g19322(new_n21671, new_n21670);
nor_4  g19323(new_n21672, new_n21671, n18452);
not_3  g19324(new_n21673, new_n21672);
nor_4  g19325(new_n21674_1, new_n21673, n13137);
not_3  g19326(new_n21675, new_n21674_1);
nor_4  g19327(new_n21676, new_n21675, n1831);
xnor_3 g19328(new_n21677, new_n21676, new_n7293);
xor_3  g19329(new_n21678, new_n21674_1, new_n16881);
not_3  g19330(new_n21679, new_n21678);
nand_4 g19331(new_n21680_1, new_n21679, new_n7310);
xor_3  g19332(new_n21681, new_n21672, new_n16885_1);
nor_4  g19333(new_n21682, new_n21681, new_n7313_1);
not_3  g19334(new_n21683, new_n21682);
not_3  g19335(new_n21684, new_n7288);
nor_4  g19336(new_n21685_1, new_n21684, new_n7268_1);
nor_4  g19337(new_n21686, new_n21685_1, new_n7289);
not_3  g19338(new_n21687_1, new_n21681);
nor_4  g19339(new_n21688, new_n21687_1, new_n21686);
nor_4  g19340(new_n21689, new_n21688, new_n21682);
xor_3  g19341(new_n21690, new_n21670, new_n16889);
nor_4  g19342(new_n21691, new_n21690, new_n7317);
not_3  g19343(new_n21692, new_n21691);
not_3  g19344(new_n21693, new_n21690);
nor_4  g19345(new_n21694, new_n21693, new_n7323);
nor_4  g19346(new_n21695, new_n21694, new_n21691);
xor_3  g19347(new_n21696, new_n21668, new_n7210);
not_3  g19348(new_n21697, new_n21696);
nor_4  g19349(new_n21698, new_n21697, new_n7327);
xnor_3 g19350(new_n21699, new_n21697, new_n7327);
xnor_3 g19351(new_n21700, new_n4490, new_n4435);
nor_4  g19352(new_n21701, new_n4544, new_n4543);
nor_4  g19353(new_n21702, new_n21701, new_n4498);
nor_4  g19354(new_n21703, new_n21702, new_n21700);
nor_4  g19355(new_n21704, new_n21703, new_n4491);
nor_4  g19356(new_n21705, new_n21704, new_n21699);
nor_4  g19357(new_n21706, new_n21705, new_n21698);
nand_4 g19358(new_n21707, new_n21706, new_n21695);
nand_4 g19359(new_n21708, new_n21707, new_n21692);
nand_4 g19360(new_n21709, new_n21708, new_n21689);
nand_4 g19361(new_n21710, new_n21709, new_n21683);
not_3  g19362(new_n21711, new_n21680_1);
nor_4  g19363(new_n21712, new_n21679, new_n7310);
nor_4  g19364(new_n21713, new_n21712, new_n21711);
nand_4 g19365(new_n21714, new_n21713, new_n21710);
nand_4 g19366(new_n21715, new_n21714, new_n21680_1);
xnor_3 g19367(new_n21716, new_n21715, new_n21677);
xnor_3 g19368(new_n21717_1, new_n21716, new_n14072);
xnor_3 g19369(new_n21718, new_n21681, new_n7313_1);
xnor_3 g19370(new_n21719_1, new_n21690, new_n7317);
not_3  g19371(new_n21720, new_n21698);
xnor_3 g19372(new_n21721, new_n21696, new_n7327);
not_3  g19373(new_n21722, new_n4491);
nand_4 g19374(new_n21723, new_n4540, new_n4494);
nand_4 g19375(new_n21724, new_n21723, new_n21722);
nand_4 g19376(new_n21725, new_n21724, new_n21721);
nand_4 g19377(new_n21726, new_n21725, new_n21720);
nor_4  g19378(new_n21727, new_n21726, new_n21719_1);
nor_4  g19379(new_n21728, new_n21727, new_n21691);
nor_4  g19380(new_n21729, new_n21728, new_n21718);
nor_4  g19381(new_n21730, new_n21729, new_n21682);
xnor_3 g19382(new_n21731, new_n21679, new_n7310);
xnor_3 g19383(new_n21732, new_n21731, new_n21730);
nor_4  g19384(new_n21733, new_n21732, new_n14077);
xnor_3 g19385(new_n21734, new_n21732, new_n14077);
xnor_3 g19386(new_n21735_1, new_n21728, new_n21718);
nor_4  g19387(new_n21736, new_n21735_1, new_n14085);
xnor_3 g19388(new_n21737, new_n21735_1, new_n14085);
xnor_3 g19389(new_n21738, new_n21726, new_n21695);
nand_4 g19390(new_n21739, new_n21738, new_n14092);
xnor_3 g19391(new_n21740, new_n21738, new_n14091);
xnor_3 g19392(new_n21741, new_n21724, new_n21721);
nand_4 g19393(new_n21742, new_n21741, new_n14098);
xnor_3 g19394(new_n21743, new_n21741, new_n14097);
nand_4 g19395(new_n21744, new_n4541, new_n14110);
nand_4 g19396(new_n21745, new_n4589, new_n4542);
nand_4 g19397(new_n21746, new_n21745, new_n21744);
nand_4 g19398(new_n21747, new_n21746, new_n21743);
nand_4 g19399(new_n21748, new_n21747, new_n21742);
nand_4 g19400(new_n21749_1, new_n21748, new_n21740);
nand_4 g19401(new_n21750_1, new_n21749_1, new_n21739);
not_3  g19402(new_n21751, new_n21750_1);
nor_4  g19403(new_n21752, new_n21751, new_n21737);
nor_4  g19404(new_n21753_1, new_n21752, new_n21736);
nor_4  g19405(new_n21754, new_n21753_1, new_n21734);
nor_4  g19406(new_n21755, new_n21754, new_n21733);
xnor_3 g19407(n4478, new_n21755, new_n21717_1);
xnor_3 g19408(n4529, new_n15075, new_n15028);
xnor_3 g19409(n4552, new_n7193, new_n7138);
not_3  g19410(new_n21759, new_n7152);
xor_3  g19411(n4595, new_n7189, new_n21759);
xnor_3 g19412(n4624, new_n17323, new_n17274);
nor_4  g19413(new_n21762, new_n21095_1, n2659);
xor_3  g19414(new_n21763, new_n21762, new_n17338);
nor_4  g19415(new_n21764, new_n21763, n14899);
not_3  g19416(new_n21765_1, new_n21763);
xor_3  g19417(new_n21766, new_n21765_1, n14899);
nor_4  g19418(new_n21767, new_n21096, n18444);
nor_4  g19419(new_n21768, new_n21105, new_n21098);
nor_4  g19420(new_n21769, new_n21768, new_n21767);
nor_4  g19421(new_n21770, new_n21769, new_n21766);
nor_4  g19422(new_n21771, new_n21770, new_n21764);
not_3  g19423(new_n21772, new_n21762);
nor_4  g19424(new_n21773, new_n21772, n2858);
xor_3  g19425(new_n21774, new_n21773, new_n21148);
nor_4  g19426(new_n21775, new_n21774, n3506);
not_3  g19427(new_n21776, new_n21774);
nor_4  g19428(new_n21777, new_n21776, new_n9753_1);
nor_4  g19429(new_n21778, new_n21777, new_n21775);
xnor_3 g19430(new_n21779_1, new_n21778, new_n21771);
not_3  g19431(new_n21780, new_n21779_1);
nand_4 g19432(new_n21781, new_n21780, new_n9132);
xnor_3 g19433(new_n21782, new_n21779_1, new_n9132);
not_3  g19434(new_n21783, new_n21769);
xnor_3 g19435(new_n21784_1, new_n21783, new_n21766);
not_3  g19436(new_n21785, new_n21784_1);
nand_4 g19437(new_n21786, new_n21785, new_n9141);
xnor_3 g19438(new_n21787, new_n21784_1, new_n9141);
not_3  g19439(new_n21788, new_n21107);
nand_4 g19440(new_n21789, new_n21788, new_n9151);
nand_4 g19441(new_n21790, new_n21118, new_n21789);
nand_4 g19442(new_n21791, new_n21790, new_n21787);
nand_4 g19443(new_n21792, new_n21791, new_n21786);
nand_4 g19444(new_n21793, new_n21792, new_n21782);
nand_4 g19445(new_n21794, new_n21793, new_n21781);
not_3  g19446(new_n21795, new_n21775);
nand_4 g19447(new_n21796, new_n21795, new_n21771);
not_3  g19448(new_n21797, new_n21773);
nor_4  g19449(new_n21798, new_n21797, n3740);
nor_4  g19450(new_n21799, new_n21777, new_n21798);
nand_4 g19451(new_n21800_1, new_n21799, new_n21796);
not_3  g19452(new_n21801, new_n21800_1);
xnor_3 g19453(new_n21802, new_n21801, new_n21794);
nand_4 g19454(new_n21803, new_n21802, new_n9075);
not_3  g19455(new_n21804, new_n9075);
xnor_3 g19456(new_n21805, new_n21800_1, new_n21794);
nand_4 g19457(new_n21806, new_n21805, new_n21804);
nand_4 g19458(new_n21807, new_n21806, new_n21803);
xnor_3 g19459(new_n21808, new_n21807, new_n9313);
not_3  g19460(new_n21809, new_n21793);
nor_4  g19461(new_n21810, new_n21792, new_n21782);
nor_4  g19462(new_n21811, new_n21810, new_n21809);
not_3  g19463(new_n21812, new_n21811);
nand_4 g19464(new_n21813, new_n21812, new_n9318_1);
xnor_3 g19465(new_n21814, new_n21790, new_n21787);
not_3  g19466(new_n21815, new_n21814);
nor_4  g19467(new_n21816, new_n21815, new_n9324);
not_3  g19468(new_n21817, new_n21816);
nor_4  g19469(new_n21818, new_n21814, new_n9325);
nor_4  g19470(new_n21819, new_n21818, new_n21816);
not_3  g19471(new_n21820_1, new_n21121);
nand_4 g19472(new_n21821, new_n21820_1, new_n9331);
xnor_3 g19473(new_n21822, new_n21121, new_n9331);
nor_4  g19474(new_n21823, new_n21134_1, new_n9340);
not_3  g19475(new_n21824, new_n21823);
nor_4  g19476(new_n21825, new_n21133, new_n9338);
nor_4  g19477(new_n21826, new_n21825, new_n21823);
nor_4  g19478(new_n21827, new_n16065, new_n9344_1);
not_3  g19479(new_n21828, new_n20899);
nand_4 g19480(new_n21829, new_n20921, new_n20901);
nand_4 g19481(new_n21830, new_n21829, new_n21828);
xnor_3 g19482(new_n21831, new_n16065, new_n9344_1);
nor_4  g19483(new_n21832_1, new_n21831, new_n21830);
nor_4  g19484(new_n21833, new_n21832_1, new_n21827);
nand_4 g19485(new_n21834, new_n21833, new_n21826);
nand_4 g19486(new_n21835, new_n21834, new_n21824);
nand_4 g19487(new_n21836, new_n21835, new_n21822);
nand_4 g19488(new_n21837, new_n21836, new_n21821);
nand_4 g19489(new_n21838, new_n21837, new_n21819);
nand_4 g19490(new_n21839_1, new_n21838, new_n21817);
xnor_3 g19491(new_n21840, new_n21811, new_n9318_1);
nand_4 g19492(new_n21841, new_n21840, new_n21839_1);
nand_4 g19493(new_n21842, new_n21841, new_n21813);
nor_4  g19494(new_n21843, new_n21842, new_n21808);
nor_4  g19495(new_n21844, new_n21807, new_n9313);
nor_4  g19496(new_n21845, new_n21805, new_n21804);
nor_4  g19497(new_n21846, new_n21802, new_n9075);
nor_4  g19498(new_n21847, new_n21846, new_n21845);
nor_4  g19499(new_n21848, new_n21847, new_n16536);
nor_4  g19500(new_n21849, new_n21848, new_n21844);
not_3  g19501(new_n21850, new_n21842);
nor_4  g19502(new_n21851, new_n21850, new_n21849);
nor_4  g19503(n4646, new_n21851, new_n21843);
xnor_3 g19504(n4674, new_n17332, new_n17250_1);
xor_3  g19505(new_n21854, n7057, n3480);
nor_4  g19506(new_n21855, new_n9050, n8381);
nor_4  g19507(new_n21856, n16722, new_n5757);
nor_4  g19508(new_n21857, n20235, new_n9053);
nor_4  g19509(new_n21858, new_n5778, n11486);
nand_4 g19510(new_n21859, n13781, new_n10209);
nor_4  g19511(new_n21860, new_n21859, new_n21858);
nor_4  g19512(new_n21861, new_n21860, new_n21857);
nor_4  g19513(new_n21862, new_n21861, new_n21856);
nor_4  g19514(new_n21863, new_n21862, new_n21855);
xor_3  g19515(new_n21864, new_n21863, new_n21854);
xnor_3 g19516(new_n21865, new_n21864, new_n3216);
nor_4  g19517(new_n21866, new_n21856, new_n21855);
xor_3  g19518(new_n21867, new_n21866, new_n21861);
nor_4  g19519(new_n21868, new_n21867, new_n3224);
not_3  g19520(new_n21869, new_n21868);
xnor_3 g19521(new_n21870, new_n21867, new_n3224);
not_3  g19522(new_n21871, new_n21870);
xor_3  g19523(new_n21872, n13781, new_n10209);
nor_4  g19524(new_n21873, new_n21872, new_n3237);
nor_4  g19525(new_n21874_1, new_n21873, new_n3244_1);
not_3  g19526(new_n21875, new_n21874_1);
not_3  g19527(new_n21876, new_n21873);
nor_4  g19528(new_n21877, new_n21876, new_n3245);
nor_4  g19529(new_n21878, new_n21877, new_n21874_1);
not_3  g19530(new_n21879, new_n21859);
nor_4  g19531(new_n21880, new_n21858, new_n21857);
xor_3  g19532(new_n21881, new_n21880, new_n21879);
nand_4 g19533(new_n21882, new_n21881, new_n21878);
nand_4 g19534(new_n21883, new_n21882, new_n21875);
nand_4 g19535(new_n21884, new_n21883, new_n21871);
nand_4 g19536(new_n21885, new_n21884, new_n21869);
xor_3  g19537(n4693, new_n21885, new_n21865);
xor_3  g19538(n4731, new_n12861_1, new_n12852);
nor_4  g19539(new_n21888, new_n7068, new_n7022);
nor_4  g19540(new_n21889, new_n7125, new_n7069);
nor_4  g19541(new_n21890, new_n21889, new_n21888);
nor_4  g19542(new_n21891, n21784, n3582);
not_3  g19543(new_n21892, new_n7023);
nor_4  g19544(new_n21893, new_n7067, new_n21892);
nor_4  g19545(new_n21894, new_n21893, new_n21891);
not_3  g19546(new_n21895, new_n21894);
nor_4  g19547(new_n21896, new_n21895, new_n21890);
nor_4  g19548(new_n21897, new_n21896, new_n18756);
not_3  g19549(new_n21898_1, new_n21896);
nor_4  g19550(new_n21899, new_n21898_1, new_n18763);
nor_4  g19551(new_n21900, new_n21899, new_n21897);
xnor_3 g19552(new_n21901, new_n21895, new_n21890);
not_3  g19553(new_n21902, new_n21901);
nor_4  g19554(new_n21903, new_n21902, new_n18759);
not_3  g19555(new_n21904, new_n21903);
nor_4  g19556(new_n21905_1, new_n21901, new_n18765);
nor_4  g19557(new_n21906, new_n21905_1, new_n21903);
not_3  g19558(new_n21907, new_n15560);
nand_4 g19559(new_n21908, new_n15614_1, new_n15561);
nand_4 g19560(new_n21909, new_n21908, new_n21907);
nand_4 g19561(new_n21910, new_n21909, new_n21906);
nand_4 g19562(new_n21911, new_n21910, new_n21904);
xnor_3 g19563(n4745, new_n21911, new_n21900);
xor_3  g19564(new_n21913, new_n7355, new_n6353);
xor_3  g19565(n4747, new_n21913, new_n11690);
not_3  g19566(new_n21915_1, new_n6696);
xor_3  g19567(n4766, new_n6699, new_n21915_1);
not_3  g19568(new_n21917, new_n16622);
xor_3  g19569(n4770, new_n16651, new_n21917);
xor_3  g19570(n4777, new_n20112, new_n19021);
xor_3  g19571(new_n21920, n17959, new_n19431);
not_3  g19572(new_n21921, n19357);
nor_4  g19573(new_n21922, new_n21921, n7566);
xor_3  g19574(new_n21923, n19357, new_n6339_1);
not_3  g19575(new_n21924, new_n21923);
nor_4  g19576(new_n21925, n7731, new_n19442);
xor_3  g19577(new_n21926, n7731, n2328);
nor_4  g19578(new_n21927, n15053, new_n6348);
nor_4  g19579(new_n21928, new_n5816, n12341);
nor_4  g19580(new_n21929, n25471, new_n6351);
nor_4  g19581(new_n21930, new_n3291, n20986);
nand_4 g19582(new_n21931, new_n5793, n12384);
nor_4  g19583(new_n21932, new_n21931, new_n21930);
nor_4  g19584(new_n21933, new_n21932, new_n21929);
nor_4  g19585(new_n21934_1, new_n21933, new_n21928);
nor_4  g19586(new_n21935, new_n21934_1, new_n21927);
not_3  g19587(new_n21936, new_n21935);
nor_4  g19588(new_n21937, new_n21936, new_n21926);
nor_4  g19589(new_n21938, new_n21937, new_n21925);
nor_4  g19590(new_n21939, new_n21938, new_n21924);
nor_4  g19591(new_n21940, new_n21939, new_n21922);
not_3  g19592(new_n21941, new_n21940);
xor_3  g19593(new_n21942, new_n21941, new_n21920);
nor_4  g19594(new_n21943_1, n20077, n6794);
nand_4 g19595(new_n21944, new_n21943_1, new_n6401);
nor_4  g19596(new_n21945, new_n21944, n8745);
nand_4 g19597(new_n21946, new_n21945, new_n6391);
xor_3  g19598(new_n21947, new_n21946, n22660);
not_3  g19599(new_n21948, new_n21947);
xor_3  g19600(new_n21949, new_n21948, new_n10744);
not_3  g19601(new_n21950, new_n21946);
nor_4  g19602(new_n21951, new_n21945, new_n6391);
nor_4  g19603(new_n21952, new_n21951, new_n21950);
nor_4  g19604(new_n21953, new_n21952, new_n6463);
not_3  g19605(new_n21954, new_n21952);
nor_4  g19606(new_n21955, new_n21954, n15884);
nor_4  g19607(new_n21956, new_n21955, new_n21953);
nand_4 g19608(new_n21957_1, new_n21944, n8745);
not_3  g19609(new_n21958, new_n21957_1);
nor_4  g19610(new_n21959, new_n21958, new_n21945);
nor_4  g19611(new_n21960_1, new_n21959, new_n6488);
not_3  g19612(new_n21961, new_n21960_1);
not_3  g19613(new_n21962, new_n21959);
nor_4  g19614(new_n21963, new_n21962, n6356);
nor_4  g19615(new_n21964, new_n21963, new_n21960_1);
not_3  g19616(new_n21965, new_n21944);
nor_4  g19617(new_n21966, new_n21943_1, new_n6401);
nor_4  g19618(new_n21967, new_n21966, new_n21965);
nor_4  g19619(new_n21968, new_n21967, new_n6475);
not_3  g19620(new_n21969, new_n21968);
not_3  g19621(new_n21970, new_n21967);
nor_4  g19622(new_n21971, new_n21970, n27104);
nor_4  g19623(new_n21972, new_n21971, new_n21968);
not_3  g19624(new_n21973, new_n21943_1);
nand_4 g19625(new_n21974, new_n21973, new_n8019);
nand_4 g19626(new_n21975, new_n21974, n27188);
nor_4  g19627(new_n21976_1, n6794, new_n10762);
xnor_3 g19628(new_n21977, new_n21974, new_n6479);
nand_4 g19629(new_n21978, new_n21977, new_n21976_1);
nand_4 g19630(new_n21979, new_n21978, new_n21975);
nand_4 g19631(new_n21980, new_n21979, new_n21972);
nand_4 g19632(new_n21981_1, new_n21980, new_n21969);
nand_4 g19633(new_n21982, new_n21981_1, new_n21964);
nand_4 g19634(new_n21983, new_n21982, new_n21961);
nand_4 g19635(new_n21984, new_n21983, new_n21956);
not_3  g19636(new_n21985, new_n21984);
nor_4  g19637(new_n21986_1, new_n21985, new_n21953);
nor_4  g19638(new_n21987, new_n21986_1, new_n21949);
xor_3  g19639(new_n21988, new_n21948, n11580);
not_3  g19640(new_n21989, new_n21986_1);
nor_4  g19641(new_n21990, new_n21989, new_n21988);
nor_4  g19642(new_n21991, new_n21990, new_n21987);
xnor_3 g19643(new_n21992, new_n21991, new_n19402);
xnor_3 g19644(new_n21993_1, new_n21983, new_n21956);
nand_4 g19645(new_n21994, new_n21993_1, new_n18624);
xnor_3 g19646(new_n21995, new_n21981_1, new_n21964);
nor_4  g19647(new_n21996, new_n21995, new_n18629);
xnor_3 g19648(new_n21997_1, new_n21995, new_n18629);
xnor_3 g19649(new_n21998, new_n21979, new_n21972);
nand_4 g19650(new_n21999, new_n21998, new_n5773);
xnor_3 g19651(new_n22000, new_n21998, new_n5772);
xnor_3 g19652(new_n22001, new_n21977, new_n21976_1);
nand_4 g19653(new_n22002, new_n22001, new_n5845);
xor_3  g19654(new_n22003, n6794, new_n10762);
nor_4  g19655(new_n22004, new_n22003, new_n5779);
xnor_3 g19656(new_n22005, new_n22001, new_n5788);
nand_4 g19657(new_n22006, new_n22005, new_n22004);
nand_4 g19658(new_n22007, new_n22006, new_n22002);
nand_4 g19659(new_n22008, new_n22007, new_n22000);
nand_4 g19660(new_n22009, new_n22008, new_n21999);
nor_4  g19661(new_n22010, new_n22009, new_n21997_1);
nor_4  g19662(new_n22011, new_n22010, new_n21996);
xnor_3 g19663(new_n22012, new_n21993_1, new_n18623);
nand_4 g19664(new_n22013, new_n22012, new_n22011);
nand_4 g19665(new_n22014, new_n22013, new_n21994);
xnor_3 g19666(new_n22015, new_n22014, new_n21992);
not_3  g19667(new_n22016_1, new_n22015);
xnor_3 g19668(new_n22017, new_n22016_1, new_n21942);
xor_3  g19669(new_n22018, new_n21938, new_n21923);
xnor_3 g19670(new_n22019, new_n22012, new_n22011);
nand_4 g19671(new_n22020, new_n22019, new_n22018);
xnor_3 g19672(new_n22021, new_n22019, new_n22018);
not_3  g19673(new_n22022, new_n22021);
xnor_3 g19674(new_n22023, new_n22009, new_n21997_1);
xor_3  g19675(new_n22024, new_n21936, new_n21926);
nor_4  g19676(new_n22025, new_n22024, new_n22023);
not_3  g19677(new_n22026, new_n22025);
xnor_3 g19678(new_n22027_1, new_n22024, new_n22023);
not_3  g19679(new_n22028, new_n22027_1);
not_3  g19680(new_n22029, new_n22000);
xnor_3 g19681(new_n22030, new_n22007, new_n22029);
nor_4  g19682(new_n22031, new_n21928, new_n21927);
xor_3  g19683(new_n22032, new_n22031, new_n21933);
nor_4  g19684(new_n22033, new_n22032, new_n22030);
not_3  g19685(new_n22034, new_n22033);
not_3  g19686(new_n22035, new_n22030);
not_3  g19687(new_n22036, new_n22032);
nor_4  g19688(new_n22037, new_n22036, new_n22035);
nor_4  g19689(new_n22038, new_n22037, new_n22033);
xnor_3 g19690(new_n22039, new_n22003, new_n5779);
xor_3  g19691(new_n22040, n16502, new_n7881);
nor_4  g19692(new_n22041, new_n22040, new_n22039);
nor_4  g19693(new_n22042, new_n21930, new_n21929);
xor_3  g19694(new_n22043_1, new_n22042, new_n21931);
nor_4  g19695(new_n22044, new_n22043_1, new_n22041);
not_3  g19696(new_n22045, new_n22005);
xnor_3 g19697(new_n22046, new_n22045, new_n22004);
xnor_3 g19698(new_n22047, new_n22043_1, new_n22041);
nor_4  g19699(new_n22048, new_n22047, new_n22046);
nor_4  g19700(new_n22049, new_n22048, new_n22044);
not_3  g19701(new_n22050_1, new_n22049);
nand_4 g19702(new_n22051, new_n22050_1, new_n22038);
nand_4 g19703(new_n22052, new_n22051, new_n22034);
nand_4 g19704(new_n22053, new_n22052, new_n22028);
nand_4 g19705(new_n22054, new_n22053, new_n22026);
nand_4 g19706(new_n22055, new_n22054, new_n22022);
nand_4 g19707(new_n22056, new_n22055, new_n22020);
xor_3  g19708(n4785, new_n22056, new_n22017);
xnor_3 g19709(n4804, new_n17039, new_n17001);
not_3  g19710(new_n22059, new_n19032);
xor_3  g19711(n4810, new_n22059, new_n19009);
nor_4  g19712(new_n22061, new_n21211, n18105);
nor_4  g19713(new_n22062, new_n10930, new_n10885);
nor_4  g19714(new_n22063_1, new_n22062, new_n22061);
not_3  g19715(new_n22064, new_n22063_1);
nand_4 g19716(new_n22065, new_n12953, new_n9446);
nand_4 g19717(new_n22066, new_n13006, new_n12954);
nand_4 g19718(new_n22067, new_n22066, new_n22065);
not_3  g19719(new_n22068_1, new_n12944);
nor_4  g19720(new_n22069, new_n12951, new_n22068_1);
not_3  g19721(new_n22070, new_n22069);
nand_4 g19722(new_n22071, new_n21449, new_n22070);
nand_4 g19723(new_n22072_1, new_n22069, new_n21447);
nand_4 g19724(new_n22073, new_n22072_1, new_n22071);
not_3  g19725(new_n22074, new_n22073);
nor_4  g19726(new_n22075, new_n22074, new_n9524);
nor_4  g19727(new_n22076_1, new_n22073, new_n9651);
nor_4  g19728(new_n22077, new_n22076_1, new_n22075);
xnor_3 g19729(new_n22078, new_n22077, new_n22067);
nor_4  g19730(new_n22079, new_n22078, new_n22064);
not_3  g19731(new_n22080, new_n22079);
xnor_3 g19732(new_n22081, new_n22078, new_n22063_1);
not_3  g19733(new_n22082, new_n13008);
nand_4 g19734(new_n22083, new_n13071, new_n13011);
nand_4 g19735(new_n22084, new_n22083, new_n22082);
nand_4 g19736(new_n22085, new_n22084, new_n22081);
nand_4 g19737(new_n22086, new_n22085, new_n22080);
not_3  g19738(new_n22087, new_n22086);
not_3  g19739(new_n22088, new_n22075);
not_3  g19740(new_n22089, new_n22076_1);
nand_4 g19741(new_n22090_1, new_n22089, new_n22067);
nand_4 g19742(new_n22091, new_n22090_1, new_n22088);
nand_4 g19743(new_n22092, new_n22091, new_n22072_1);
nand_4 g19744(n4814, new_n22092, new_n22087);
not_3  g19745(new_n22094, new_n19838);
xor_3  g19746(n4850, new_n22094, new_n19837);
xnor_3 g19747(n4891, new_n20883, new_n20840);
xnor_3 g19748(n4925, new_n21087, new_n21052);
not_3  g19749(new_n22098, new_n19844);
xor_3  g19750(n4947, new_n22098, new_n19822);
xor_3  g19751(n4952, new_n11279, new_n11277);
xor_3  g19752(new_n22101, n25068, new_n11820);
not_3  g19753(new_n22102, new_n22101);
nor_4  g19754(new_n22103, n22879, new_n9474);
not_3  g19755(new_n22104, new_n22103);
xor_3  g19756(new_n22105, n22879, new_n9474);
nor_4  g19757(new_n22106, new_n9485, n2117);
not_3  g19758(new_n22107_1, new_n22106);
xor_3  g19759(new_n22108, n22631, new_n11830);
nor_4  g19760(new_n22109, n16743, new_n11854);
nor_4  g19761(new_n22110, new_n9488, n5882);
nor_4  g19762(new_n22111, n15258, new_n11847);
nor_4  g19763(new_n22112, new_n11842_1, n4588);
not_3  g19764(new_n22113_1, new_n22112);
nor_4  g19765(new_n22114, new_n9492, n11775);
nor_4  g19766(new_n22115, new_n22114, new_n22113_1);
nor_4  g19767(new_n22116, new_n22115, new_n22111);
nor_4  g19768(new_n22117, new_n22116, new_n22110);
nor_4  g19769(new_n22118, new_n22117, new_n22109);
nand_4 g19770(new_n22119, new_n22118, new_n22108);
nand_4 g19771(new_n22120, new_n22119, new_n22107_1);
nand_4 g19772(new_n22121, new_n22120, new_n22105);
nand_4 g19773(new_n22122, new_n22121, new_n22104);
xnor_3 g19774(new_n22123, new_n22122, new_n22102);
nand_4 g19775(new_n22124_1, new_n22123, new_n18559);
not_3  g19776(new_n22125, new_n22124_1);
nor_4  g19777(new_n22126_1, new_n22123, new_n18559);
nor_4  g19778(new_n22127, new_n22126_1, new_n22125);
not_3  g19779(new_n22128, new_n22105);
xnor_3 g19780(new_n22129, new_n22120, new_n22128);
nor_4  g19781(new_n22130_1, new_n22129, new_n18568);
xnor_3 g19782(new_n22131, new_n22129, new_n18568);
not_3  g19783(new_n22132, new_n22118);
xnor_3 g19784(new_n22133, new_n22132, new_n22108);
nor_4  g19785(new_n22134, new_n22133, new_n18573);
xnor_3 g19786(new_n22135, new_n22133, new_n18573);
not_3  g19787(new_n22136, new_n22116);
not_3  g19788(new_n22137, new_n22109);
not_3  g19789(new_n22138, new_n22110);
nand_4 g19790(new_n22139, new_n22138, new_n22137);
xnor_3 g19791(new_n22140, new_n22139, new_n22136);
nor_4  g19792(new_n22141, new_n22140, new_n18578_1);
not_3  g19793(new_n22142, new_n22141);
not_3  g19794(new_n22143, new_n22140);
nor_4  g19795(new_n22144_1, new_n22143, new_n18577);
nor_4  g19796(new_n22145, new_n22144_1, new_n22141);
nor_4  g19797(new_n22146, new_n22114, new_n22111);
xnor_3 g19798(new_n22147, new_n22146, new_n22113_1);
nor_4  g19799(new_n22148, new_n22147, new_n18582_1);
not_3  g19800(new_n22149, new_n22148);
nand_4 g19801(new_n22150_1, new_n18303, new_n18302);
not_3  g19802(new_n22151, new_n22150_1);
not_3  g19803(new_n22152, new_n22147);
nor_4  g19804(new_n22153, new_n22152, new_n18581);
nor_4  g19805(new_n22154, new_n22153, new_n22148);
nand_4 g19806(new_n22155, new_n22154, new_n22151);
nand_4 g19807(new_n22156, new_n22155, new_n22149);
nand_4 g19808(new_n22157_1, new_n22156, new_n22145);
nand_4 g19809(new_n22158, new_n22157_1, new_n22142);
nor_4  g19810(new_n22159, new_n22158, new_n22135);
nor_4  g19811(new_n22160, new_n22159, new_n22134);
nor_4  g19812(new_n22161, new_n22160, new_n22131);
nor_4  g19813(new_n22162, new_n22161, new_n22130_1);
xnor_3 g19814(new_n22163, new_n22162, new_n22127);
xnor_3 g19815(new_n22164, new_n22163, new_n18464);
not_3  g19816(new_n22165, new_n22164);
not_3  g19817(new_n22166, new_n22131);
not_3  g19818(new_n22167, new_n22160);
nor_4  g19819(new_n22168, new_n22167, new_n22166);
nor_4  g19820(new_n22169, new_n22168, new_n22161);
nand_4 g19821(new_n22170, new_n22169, new_n18475);
xnor_3 g19822(new_n22171, new_n22169, new_n18471);
not_3  g19823(new_n22172, new_n22135);
not_3  g19824(new_n22173_1, new_n22158);
nor_4  g19825(new_n22174, new_n22173_1, new_n22172);
nor_4  g19826(new_n22175, new_n22174, new_n22159);
nand_4 g19827(new_n22176, new_n22175, new_n16450);
xnor_3 g19828(new_n22177, new_n22175, new_n16452);
not_3  g19829(new_n22178, new_n22157_1);
nor_4  g19830(new_n22179, new_n22156, new_n22145);
nor_4  g19831(new_n22180, new_n22179, new_n22178);
nor_4  g19832(new_n22181, new_n22180, new_n16461);
not_3  g19833(new_n22182, new_n22181);
not_3  g19834(new_n22183, new_n22180);
nor_4  g19835(new_n22184, new_n22183, new_n16462);
nor_4  g19836(new_n22185, new_n22184, new_n22181);
nor_4  g19837(new_n22186, new_n18304_1, new_n11983);
nor_4  g19838(new_n22187, new_n22186, new_n16481_1);
not_3  g19839(new_n22188, new_n22187);
not_3  g19840(new_n22189, new_n22186);
nor_4  g19841(new_n22190, new_n22189, new_n16505);
nor_4  g19842(new_n22191, new_n22190, new_n22187);
not_3  g19843(new_n22192, new_n22154);
xnor_3 g19844(new_n22193, new_n22192, new_n22150_1);
nand_4 g19845(new_n22194, new_n22193, new_n22191);
nand_4 g19846(new_n22195, new_n22194, new_n22188);
nand_4 g19847(new_n22196, new_n22195, new_n22185);
nand_4 g19848(new_n22197, new_n22196, new_n22182);
nand_4 g19849(new_n22198_1, new_n22197, new_n22177);
nand_4 g19850(new_n22199, new_n22198_1, new_n22176);
nand_4 g19851(new_n22200, new_n22199, new_n22171);
nand_4 g19852(new_n22201_1, new_n22200, new_n22170);
xor_3  g19853(n4966, new_n22201_1, new_n22165);
xor_3  g19854(n4972, new_n21485, new_n21481);
nor_4  g19855(new_n22204, new_n8903, n23895);
xnor_3 g19856(new_n22205, new_n8903, new_n6319);
not_3  g19857(new_n22206, new_n22205);
xnor_3 g19858(new_n22207, new_n8892, new_n8883);
nor_4  g19859(new_n22208, new_n22207, new_n6324);
not_3  g19860(new_n22209, new_n22208);
nor_4  g19861(new_n22210, new_n8911_1, n17351);
nor_4  g19862(new_n22211, new_n22210, new_n22208);
nand_4 g19863(new_n22212, new_n8918, n11736);
nor_4  g19864(new_n22213_1, new_n8918, n11736);
nor_4  g19865(new_n22214, new_n8917, new_n6330_1);
nor_4  g19866(new_n22215, new_n22214, new_n22213_1);
nand_4 g19867(new_n22216, new_n20674, new_n22215);
nand_4 g19868(new_n22217, new_n22216, new_n22212);
nand_4 g19869(new_n22218, new_n22217, new_n22211);
nand_4 g19870(new_n22219, new_n22218, new_n22209);
nor_4  g19871(new_n22220, new_n22219, new_n22206);
nor_4  g19872(new_n22221, new_n22220, new_n22204);
nand_4 g19873(new_n22222, new_n22221, new_n8898);
nor_4  g19874(new_n22223, new_n20605, n2289);
not_3  g19875(new_n22224, new_n22223);
nor_4  g19876(new_n22225, new_n22224, n23697);
xor_3  g19877(new_n22226, new_n22225, new_n8789);
nor_4  g19878(new_n22227, new_n22226, n7593);
not_3  g19879(new_n22228, new_n22226);
nor_4  g19880(new_n22229, new_n22228, new_n15741);
nor_4  g19881(new_n22230, new_n22229, new_n22227);
not_3  g19882(new_n22231, n337);
xor_3  g19883(new_n22232, new_n22224, n23697);
not_3  g19884(new_n22233, new_n22232);
nor_4  g19885(new_n22234, new_n22233, new_n22231);
nor_4  g19886(new_n22235, new_n22232, n337);
not_3  g19887(new_n22236, new_n22235);
not_3  g19888(new_n22237, new_n20608);
not_3  g19889(new_n22238, new_n20609_1);
nand_4 g19890(new_n22239, new_n20626, new_n22238);
nand_4 g19891(new_n22240, new_n22239, new_n22237);
nand_4 g19892(new_n22241, new_n22240, new_n22236);
not_3  g19893(new_n22242, new_n22241);
nor_4  g19894(new_n22243, new_n22242, new_n22234);
xnor_3 g19895(new_n22244, new_n22243, new_n22230);
nor_4  g19896(new_n22245, new_n22244, n25972);
not_3  g19897(new_n22246, new_n22245);
xnor_3 g19898(new_n22247, new_n22244, n25972);
not_3  g19899(new_n22248, new_n22247);
nor_4  g19900(new_n22249, new_n22235, new_n22234);
xnor_3 g19901(new_n22250, new_n22249, new_n22240);
nand_4 g19902(new_n22251, new_n22250, new_n10327_1);
nand_4 g19903(new_n22252, new_n20627, new_n8045);
nand_4 g19904(new_n22253_1, new_n20654, new_n20629_1);
nand_4 g19905(new_n22254, new_n22253_1, new_n22252);
not_3  g19906(new_n22255, new_n22251);
nor_4  g19907(new_n22256, new_n22250, new_n10327_1);
nor_4  g19908(new_n22257, new_n22256, new_n22255);
nand_4 g19909(new_n22258, new_n22257, new_n22254);
nand_4 g19910(new_n22259, new_n22258, new_n22251);
nand_4 g19911(new_n22260, new_n22259, new_n22248);
nand_4 g19912(new_n22261, new_n22260, new_n22246);
nor_4  g19913(new_n22262, new_n22243, new_n22227);
not_3  g19914(new_n22263, new_n22225);
nor_4  g19915(new_n22264, new_n22263, n2978);
nor_4  g19916(new_n22265, new_n22229, new_n22264);
not_3  g19917(new_n22266, new_n22265);
nor_4  g19918(new_n22267, new_n22266, new_n22262);
not_3  g19919(new_n22268, new_n22267);
nor_4  g19920(new_n22269, new_n22268, new_n22261);
not_3  g19921(new_n22270_1, new_n22222);
nor_4  g19922(new_n22271, new_n22221, new_n8898);
nor_4  g19923(new_n22272, new_n22271, new_n22270_1);
not_3  g19924(new_n22273, new_n22272);
xnor_3 g19925(new_n22274_1, new_n22267, new_n22261);
not_3  g19926(new_n22275, new_n22274_1);
nand_4 g19927(new_n22276, new_n22275, new_n22273);
not_3  g19928(new_n22277, new_n22276);
xnor_3 g19929(new_n22278, new_n22274_1, new_n22272);
xnor_3 g19930(new_n22279, new_n22219, new_n22205);
xnor_3 g19931(new_n22280, new_n22259, new_n22247);
nor_4  g19932(new_n22281, new_n22280, new_n22279);
not_3  g19933(new_n22282, new_n22281);
not_3  g19934(new_n22283_1, new_n22279);
not_3  g19935(new_n22284, new_n22280);
nor_4  g19936(new_n22285, new_n22284, new_n22283_1);
nor_4  g19937(new_n22286, new_n22285, new_n22281);
xnor_3 g19938(new_n22287, new_n22217, new_n22211);
not_3  g19939(new_n22288, new_n22252);
nor_4  g19940(new_n22289, new_n20659, new_n22288);
xnor_3 g19941(new_n22290_1, new_n22257, new_n22289);
nor_4  g19942(new_n22291, new_n22290_1, new_n22287);
not_3  g19943(new_n22292, new_n22291);
nand_4 g19944(new_n22293, new_n20676, new_n20660);
not_3  g19945(new_n22294, new_n22293);
nor_4  g19946(new_n22295, new_n20699, new_n20677);
nor_4  g19947(new_n22296, new_n22295, new_n22294);
not_3  g19948(new_n22297, new_n22287);
xnor_3 g19949(new_n22298, new_n22257, new_n22254);
nor_4  g19950(new_n22299, new_n22298, new_n22297);
nor_4  g19951(new_n22300, new_n22299, new_n22291);
nand_4 g19952(new_n22301, new_n22300, new_n22296);
nand_4 g19953(new_n22302, new_n22301, new_n22292);
nand_4 g19954(new_n22303, new_n22302, new_n22286);
nand_4 g19955(new_n22304, new_n22303, new_n22282);
nor_4  g19956(new_n22305, new_n22304, new_n22278);
nor_4  g19957(new_n22306, new_n22305, new_n22277);
xnor_3 g19958(new_n22307, new_n22306, new_n22269);
xnor_3 g19959(n5011, new_n22307, new_n22222);
not_3  g19960(new_n22309_1, n11220);
nor_4  g19961(new_n22310, new_n22309_1, n2944);
xor_3  g19962(new_n22311_1, n11220, new_n13250);
not_3  g19963(new_n22312, new_n22311_1);
not_3  g19964(new_n22313, n22379);
nor_4  g19965(new_n22314, new_n22313, n767);
nand_4 g19966(new_n22315, new_n3031, new_n2984);
not_3  g19967(new_n22316, new_n22315);
nor_4  g19968(new_n22317_1, new_n22316, new_n22314);
nor_4  g19969(new_n22318, new_n22317_1, new_n22312);
nor_4  g19970(new_n22319, new_n22318, new_n22310);
not_3  g19971(new_n22320, new_n22319);
nand_4 g19972(new_n22321, n16544, n2160);
nor_4  g19973(new_n22322, n16544, n2160);
not_3  g19974(new_n22323, new_n22322);
nor_4  g19975(new_n22324, n10763, n6814);
not_3  g19976(new_n22325, new_n3033);
nor_4  g19977(new_n22326, new_n3073, new_n22325);
nor_4  g19978(new_n22327, new_n22326, new_n22324);
nand_4 g19979(new_n22328, new_n22327, new_n22323);
nand_4 g19980(new_n22329, new_n22328, new_n22321);
not_3  g19981(new_n22330, new_n22329);
nor_4  g19982(new_n22331, new_n22330, new_n18388);
xor_3  g19983(new_n22332_1, new_n22329, new_n18388);
not_3  g19984(new_n22333, new_n22321);
nor_4  g19985(new_n22334, new_n22322, new_n22333);
xnor_3 g19986(new_n22335_1, new_n22334, new_n22327);
nor_4  g19987(new_n22336, new_n22335_1, new_n18353);
xnor_3 g19988(new_n22337, new_n22335_1, new_n18350_1);
not_3  g19989(new_n22338, new_n22337);
nor_4  g19990(new_n22339, new_n3119, new_n3074);
nor_4  g19991(new_n22340, new_n3186, new_n3120);
nor_4  g19992(new_n22341_1, new_n22340, new_n22339);
nor_4  g19993(new_n22342, new_n22341_1, new_n22338);
nor_4  g19994(new_n22343, new_n22342, new_n22336);
nor_4  g19995(new_n22344, new_n22343, new_n22332_1);
nor_4  g19996(new_n22345, new_n22344, new_n22331);
nor_4  g19997(new_n22346, new_n22345, new_n22320);
xnor_3 g19998(new_n22347, new_n22343, new_n22332_1);
not_3  g19999(new_n22348, new_n22347);
nor_4  g20000(new_n22349, new_n22348, new_n22319);
nor_4  g20001(new_n22350, new_n22347, new_n22320);
xor_3  g20002(new_n22351, new_n22317_1, new_n22312);
xnor_3 g20003(new_n22352, new_n22341_1, new_n22338);
not_3  g20004(new_n22353_1, new_n22352);
nor_4  g20005(new_n22354, new_n22353_1, new_n22351);
xnor_3 g20006(new_n22355, new_n22353_1, new_n22351);
not_3  g20007(new_n22356, new_n3187);
nor_4  g20008(new_n22357, new_n22356, new_n3032);
not_3  g20009(new_n22358_1, new_n3188);
nor_4  g20010(new_n22359_1, new_n3263_1, new_n22358_1);
nor_4  g20011(new_n22360, new_n22359_1, new_n22357);
nor_4  g20012(new_n22361, new_n22360, new_n22355);
nor_4  g20013(new_n22362, new_n22361, new_n22354);
nor_4  g20014(new_n22363, new_n22362, new_n22350);
nor_4  g20015(new_n22364, new_n22363, new_n22349);
nor_4  g20016(new_n22365, new_n22364, new_n22346);
not_3  g20017(new_n22366, new_n22345);
nor_4  g20018(new_n22367, new_n22366, new_n22319);
nor_4  g20019(new_n22368, new_n22367, new_n22363);
nor_4  g20020(n5020, new_n22368, new_n22365);
nor_4  g20021(new_n22370, n13781, n11486);
not_3  g20022(new_n22371, new_n22370);
nor_4  g20023(new_n22372, new_n22371, n16722);
not_3  g20024(new_n22373, new_n22372);
nor_4  g20025(new_n22374, new_n22373, n3480);
xor_3  g20026(new_n22375, new_n22374, new_n9045);
xnor_3 g20027(new_n22376, new_n22375, new_n3139);
xor_3  g20028(new_n22377, new_n22372, new_n2426);
nor_4  g20029(new_n22378, new_n22377, new_n3145);
xnor_3 g20030(new_n22379_1, new_n22377, new_n3145);
xor_3  g20031(new_n22380, new_n22370, new_n9050);
nor_4  g20032(new_n22381, new_n22380, new_n3155);
xnor_3 g20033(new_n22382, new_n22380, new_n3155);
not_3  g20034(new_n22383, new_n6752);
nor_4  g20035(new_n22384, new_n22370, new_n22383);
nor_4  g20036(new_n22385, new_n22384, new_n3162);
nand_4 g20037(new_n22386, new_n3166, new_n2390);
xnor_3 g20038(new_n22387, new_n22384, new_n3162);
nor_4  g20039(new_n22388, new_n22387, new_n22386);
nor_4  g20040(new_n22389, new_n22388, new_n22385);
nor_4  g20041(new_n22390, new_n22389, new_n22382);
nor_4  g20042(new_n22391, new_n22390, new_n22381);
nor_4  g20043(new_n22392, new_n22391, new_n22379_1);
nor_4  g20044(new_n22393, new_n22392, new_n22378);
xnor_3 g20045(new_n22394, new_n22393, new_n22376);
xnor_3 g20046(new_n22395, new_n22394, new_n8152);
not_3  g20047(new_n22396, new_n22395);
xnor_3 g20048(new_n22397, new_n22391, new_n22379_1);
not_3  g20049(new_n22398, new_n22397);
nand_4 g20050(new_n22399, new_n22398, new_n8160);
xnor_3 g20051(new_n22400, new_n22397, new_n8160);
xnor_3 g20052(new_n22401, new_n22389, new_n22382);
not_3  g20053(new_n22402, new_n22401);
nand_4 g20054(new_n22403, new_n22402, new_n8168);
not_3  g20055(new_n22404, new_n22386);
not_3  g20056(new_n22405, new_n22387);
nor_4  g20057(new_n22406, new_n22405, new_n22404);
nor_4  g20058(new_n22407, new_n22406, new_n22388);
nand_4 g20059(new_n22408, new_n22407, new_n19706);
xor_3  g20060(new_n22409, new_n3167, new_n2390);
nand_4 g20061(new_n22410, new_n22409, new_n8177);
xnor_3 g20062(new_n22411, new_n22407, new_n8175);
nand_4 g20063(new_n22412, new_n22411, new_n22410);
nand_4 g20064(new_n22413, new_n22412, new_n22408);
xnor_3 g20065(new_n22414, new_n22401, new_n8168);
nand_4 g20066(new_n22415, new_n22414, new_n22413);
nand_4 g20067(new_n22416, new_n22415, new_n22403);
nand_4 g20068(new_n22417, new_n22416, new_n22400);
nand_4 g20069(new_n22418, new_n22417, new_n22399);
xor_3  g20070(n5024, new_n22418, new_n22396);
not_3  g20071(new_n22420, new_n4014_1);
xor_3  g20072(n5046, new_n4064, new_n22420);
xor_3  g20073(n5062, new_n6855, new_n4169);
xnor_3 g20074(n5064, new_n15128_1, new_n15101);
nand_4 g20075(new_n22424, n12495, n11479);
not_3  g20076(new_n22425, new_n22424);
nor_4  g20077(new_n22426, n12495, n11479);
nor_4  g20078(new_n22427, new_n22426, new_n22425);
xor_3  g20079(new_n22428, new_n22427, new_n2392);
xor_3  g20080(new_n22429, n9251, new_n9869);
nor_4  g20081(new_n22430, new_n22429, new_n22428);
nor_4  g20082(new_n22431, new_n2374_1, n7428);
xor_3  g20083(new_n22432, n20138, new_n8273);
xnor_3 g20084(new_n22433_1, new_n22432, new_n22431);
nand_4 g20085(new_n22434, new_n22433_1, new_n22430);
not_3  g20086(new_n22435, new_n22434);
nor_4  g20087(new_n22436, new_n22433_1, new_n22430);
nor_4  g20088(new_n22437, new_n22436, new_n22435);
nor_4  g20089(new_n22438, new_n22427, new_n2392);
xnor_3 g20090(new_n22439, n20235, n8259);
xnor_3 g20091(new_n22440, new_n22439, new_n22424);
xnor_3 g20092(new_n22441, new_n22440, new_n2396);
xor_3  g20093(new_n22442_1, new_n22441, new_n22438);
xor_3  g20094(n5082, new_n22442_1, new_n22437);
xor_3  g20095(n5120, new_n16640_1, new_n16637);
not_3  g20096(new_n22445, new_n18129);
xor_3  g20097(n5158, new_n18139, new_n22445);
not_3  g20098(new_n22447, new_n19842);
xor_3  g20099(n5168, new_n22447, new_n19828);
not_3  g20100(new_n22449, new_n19416);
xnor_3 g20101(new_n22450, new_n21158, n6659);
nor_4  g20102(new_n22451, new_n17381, n23250);
xnor_3 g20103(new_n22452, new_n17381, n23250);
nor_4  g20104(new_n22453, new_n17388, n11455);
xnor_3 g20105(new_n22454, new_n17388, n11455);
nor_4  g20106(new_n22455, new_n17393, n3945);
xnor_3 g20107(new_n22456, new_n17393, n3945);
nand_4 g20108(new_n22457, new_n17399, n5255);
not_3  g20109(new_n22458, new_n22457);
nor_4  g20110(new_n22459, new_n17399, n5255);
nor_4  g20111(new_n22460, new_n22459, new_n22458);
not_3  g20112(new_n22461, new_n18640);
nand_4 g20113(new_n22462, new_n18661, new_n18642);
nand_4 g20114(new_n22463, new_n22462, new_n22461);
not_3  g20115(new_n22464, new_n22463);
nand_4 g20116(new_n22465, new_n22464, new_n22460);
nand_4 g20117(new_n22466, new_n22465, new_n22457);
nor_4  g20118(new_n22467_1, new_n22466, new_n22456);
nor_4  g20119(new_n22468, new_n22467_1, new_n22455);
nor_4  g20120(new_n22469, new_n22468, new_n22454);
nor_4  g20121(new_n22470_1, new_n22469, new_n22453);
nor_4  g20122(new_n22471, new_n22470_1, new_n22452);
nor_4  g20123(new_n22472, new_n22471, new_n22451);
not_3  g20124(new_n22473, new_n22472);
xnor_3 g20125(new_n22474, new_n22473, new_n22450);
nand_4 g20126(new_n22475, new_n22474, new_n22449);
not_3  g20127(new_n22476, new_n22475);
nor_4  g20128(new_n22477, new_n22474, new_n22449);
nor_4  g20129(new_n22478, new_n22477, new_n22476);
not_3  g20130(new_n22479, new_n22470_1);
xnor_3 g20131(new_n22480, new_n22479, new_n22452);
nand_4 g20132(new_n22481, new_n22480, new_n19530);
not_3  g20133(new_n22482, new_n22481);
nor_4  g20134(new_n22483, new_n22480, new_n19530);
nor_4  g20135(new_n22484_1, new_n22483, new_n22482);
not_3  g20136(new_n22485, new_n22468);
xnor_3 g20137(new_n22486, new_n22485, new_n22454);
nand_4 g20138(new_n22487, new_n22486, new_n19535);
not_3  g20139(new_n22488, new_n22487);
nor_4  g20140(new_n22489_1, new_n22486, new_n19535);
nor_4  g20141(new_n22490, new_n22489_1, new_n22488);
xnor_3 g20142(new_n22491, new_n22466, new_n22456);
nor_4  g20143(new_n22492_1, new_n22491, new_n19539_1);
not_3  g20144(new_n22493, new_n22492_1);
not_3  g20145(new_n22494_1, new_n22491);
nor_4  g20146(new_n22495, new_n22494_1, new_n19540);
nor_4  g20147(new_n22496, new_n22495, new_n22492_1);
xnor_3 g20148(new_n22497, new_n22464, new_n22460);
not_3  g20149(new_n22498, new_n22497);
nor_4  g20150(new_n22499, new_n22498, new_n19547);
not_3  g20151(new_n22500, new_n22499);
nor_4  g20152(new_n22501, new_n22497, new_n19546);
nor_4  g20153(new_n22502, new_n22501, new_n22499);
not_3  g20154(new_n22503, new_n18663);
nand_4 g20155(new_n22504, new_n18692, new_n18667);
nand_4 g20156(new_n22505, new_n22504, new_n22503);
nand_4 g20157(new_n22506, new_n22505, new_n22502);
nand_4 g20158(new_n22507, new_n22506, new_n22500);
nand_4 g20159(new_n22508, new_n22507, new_n22496);
nand_4 g20160(new_n22509, new_n22508, new_n22493);
nand_4 g20161(new_n22510, new_n22509, new_n22490);
nand_4 g20162(new_n22511, new_n22510, new_n22487);
nand_4 g20163(new_n22512, new_n22511, new_n22484_1);
nand_4 g20164(new_n22513, new_n22512, new_n22481);
xnor_3 g20165(n5184, new_n22513, new_n22478);
not_3  g20166(new_n22515, new_n5135);
nor_4  g20167(new_n22516, new_n5137, new_n5136);
nor_4  g20168(new_n22517, new_n22516, new_n5135);
not_3  g20169(new_n22518, new_n5142);
not_3  g20170(new_n22519, new_n5144);
not_3  g20171(new_n22520, new_n5147);
not_3  g20172(new_n22521, new_n5156);
nand_4 g20173(new_n22522, new_n5219, new_n22521);
nand_4 g20174(new_n22523, new_n22522, new_n5149);
nand_4 g20175(new_n22524, new_n22523, new_n22520);
nand_4 g20176(new_n22525, new_n22524, new_n22519);
nand_4 g20177(new_n22526, new_n22525, new_n22518);
nand_4 g20178(new_n22527, new_n22526, new_n22517);
nand_4 g20179(new_n22528, new_n22527, new_n22515);
nand_4 g20180(new_n22529, new_n22528, new_n5128_1);
nand_4 g20181(new_n22530, new_n5227, new_n5130);
nand_4 g20182(n5228, new_n22530, new_n22529);
nor_4  g20183(new_n22532, n25494, new_n9766);
not_3  g20184(new_n22533_1, new_n13563);
nor_4  g20185(new_n22534, new_n13581, new_n22533_1);
nor_4  g20186(new_n22535, new_n22534, new_n22532);
xnor_3 g20187(new_n22536, new_n22535, new_n8486);
nor_4  g20188(new_n22537, new_n13583, new_n8389);
not_3  g20189(new_n22538, new_n22537);
nor_4  g20190(new_n22539, new_n8394, new_n8315);
nor_4  g20191(new_n22540, new_n22539, new_n8311);
nor_4  g20192(new_n22541, new_n8387, new_n22540);
nor_4  g20193(new_n22542, new_n8388, new_n8374);
nor_4  g20194(new_n22543, new_n22542, new_n22541);
nor_4  g20195(new_n22544, new_n13582, new_n22543);
nor_4  g20196(new_n22545, new_n22544, new_n22537);
nand_4 g20197(new_n22546, new_n13606, new_n8398);
nand_4 g20198(new_n22547, new_n15130, new_n15099);
nand_4 g20199(new_n22548, new_n22547, new_n22546);
nand_4 g20200(new_n22549, new_n22548, new_n22545);
nand_4 g20201(new_n22550, new_n22549, new_n22538);
xnor_3 g20202(n5256, new_n22550, new_n22536);
xor_3  g20203(n5265, new_n7847, new_n7834_1);
xnor_3 g20204(n5273, new_n20885, new_n20835);
xor_3  g20205(new_n22554_1, n20946, new_n8796);
nand_4 g20206(new_n22555, n7751, new_n7937_1);
xor_3  g20207(new_n22556, n7751, new_n7937_1);
nand_4 g20208(new_n22557, n26823, new_n8803_1);
nand_4 g20209(new_n22558, new_n20456, new_n20440);
nand_4 g20210(new_n22559, new_n22558, new_n22557);
nand_4 g20211(new_n22560, new_n22559, new_n22556);
nand_4 g20212(new_n22561, new_n22560, new_n22555);
xor_3  g20213(new_n22562, new_n22561, new_n22554_1);
xnor_3 g20214(new_n22563, new_n22562, new_n8721_1);
not_3  g20215(new_n22564, new_n22556);
xor_3  g20216(new_n22565, new_n22559, new_n22564);
nand_4 g20217(new_n22566, new_n22565, new_n8731);
xnor_3 g20218(new_n22567, new_n22565, new_n8730);
not_3  g20219(new_n22568, new_n20457);
nand_4 g20220(new_n22569, new_n22568, new_n8737);
nand_4 g20221(new_n22570, new_n20483, new_n20458);
nand_4 g20222(new_n22571, new_n22570, new_n22569);
nand_4 g20223(new_n22572, new_n22571, new_n22567);
nand_4 g20224(new_n22573, new_n22572, new_n22566);
xnor_3 g20225(n5274, new_n22573, new_n22563);
nor_4  g20226(new_n22575, n25316, n20385);
nand_4 g20227(new_n22576, new_n22575, new_n14842);
nor_4  g20228(new_n22577, new_n22576, n3918);
xor_3  g20229(new_n22578, new_n22577, n6513);
xnor_3 g20230(new_n22579, new_n22578, new_n10539);
xor_3  g20231(new_n22580, new_n22576, new_n14840);
nand_4 g20232(new_n22581, new_n22580, new_n10541);
xor_3  g20233(new_n22582, new_n22575, new_n14842);
not_3  g20234(new_n22583, new_n22582);
nand_4 g20235(new_n22584_1, new_n22583, new_n10552);
xnor_3 g20236(new_n22585, new_n22582, new_n10552);
xor_3  g20237(new_n22586, n25316, n20385);
nand_4 g20238(new_n22587, new_n22586, new_n10565);
not_3  g20239(new_n22588_1, new_n22587);
not_3  g20240(new_n22589_1, new_n10670);
xnor_3 g20241(new_n22590, new_n22586, new_n10565);
nor_4  g20242(new_n22591_1, new_n22590, new_n22589_1);
nor_4  g20243(new_n22592, new_n22591_1, new_n22588_1);
nand_4 g20244(new_n22593, new_n22592, new_n22585);
nand_4 g20245(new_n22594, new_n22593, new_n22584_1);
xnor_3 g20246(new_n22595, new_n22580, new_n10542);
nand_4 g20247(new_n22596, new_n22595, new_n22594);
nand_4 g20248(new_n22597_1, new_n22596, new_n22581);
xnor_3 g20249(new_n22598, new_n22597_1, new_n22579);
xor_3  g20250(new_n22599, new_n20173, new_n10265);
nor_4  g20251(new_n22600, new_n20179_1, new_n10291);
not_3  g20252(new_n22601, new_n22600);
xor_3  g20253(new_n22602, new_n20179_1, new_n10291);
nand_4 g20254(new_n22603, new_n4614, n24786);
xor_3  g20255(new_n22604, new_n4614, n24786);
not_3  g20256(new_n22605, n27120);
nor_4  g20257(new_n22606, new_n4621, new_n22605);
not_3  g20258(new_n22607, new_n22606);
not_3  g20259(new_n22608, n23065);
nand_4 g20260(new_n22609, new_n4626, new_n22608);
nor_4  g20261(new_n22610, new_n4622, n27120);
nor_4  g20262(new_n22611, new_n22610, new_n22606);
nand_4 g20263(new_n22612, new_n22611, new_n22609);
nand_4 g20264(new_n22613, new_n22612, new_n22607);
nand_4 g20265(new_n22614, new_n22613, new_n22604);
nand_4 g20266(new_n22615, new_n22614, new_n22603);
nand_4 g20267(new_n22616, new_n22615, new_n22602);
nand_4 g20268(new_n22617, new_n22616, new_n22601);
xnor_3 g20269(new_n22618, new_n22617, new_n22599);
xnor_3 g20270(new_n22619_1, new_n22618, new_n22598);
not_3  g20271(new_n22620_1, new_n22619_1);
xnor_3 g20272(new_n22621, new_n22615, new_n22602);
xnor_3 g20273(new_n22622, new_n22595, new_n22594);
not_3  g20274(new_n22623_1, new_n22622);
nand_4 g20275(new_n22624, new_n22623_1, new_n22621);
xnor_3 g20276(new_n22625, new_n22622, new_n22621);
xnor_3 g20277(new_n22626_1, new_n22613, new_n22604);
xnor_3 g20278(new_n22627, new_n22592, new_n22585);
not_3  g20279(new_n22628, new_n22627);
nand_4 g20280(new_n22629, new_n22628, new_n22626_1);
xnor_3 g20281(new_n22630, new_n22627, new_n22626_1);
not_3  g20282(new_n22631_1, new_n22590);
nor_4  g20283(new_n22632, new_n22631_1, new_n10670);
nor_4  g20284(new_n22633, new_n22632, new_n22591_1);
xnor_3 g20285(new_n22634, new_n22611, new_n22609);
not_3  g20286(new_n22635, new_n22634);
nor_4  g20287(new_n22636, new_n22635, new_n22633);
not_3  g20288(new_n22637, new_n22636);
xnor_3 g20289(new_n22638, new_n4626, new_n22608);
not_3  g20290(new_n22639, new_n22638);
nor_4  g20291(new_n22640, new_n22639, new_n10672);
not_3  g20292(new_n22641, new_n22640);
not_3  g20293(new_n22642, new_n22633);
nor_4  g20294(new_n22643, new_n22634, new_n22642);
nor_4  g20295(new_n22644, new_n22643, new_n22636);
nand_4 g20296(new_n22645, new_n22644, new_n22641);
nand_4 g20297(new_n22646, new_n22645, new_n22637);
nand_4 g20298(new_n22647, new_n22646, new_n22630);
nand_4 g20299(new_n22648, new_n22647, new_n22629);
nand_4 g20300(new_n22649, new_n22648, new_n22625);
nand_4 g20301(new_n22650, new_n22649, new_n22624);
xor_3  g20302(n5300, new_n22650, new_n22620_1);
not_3  g20303(new_n22652, new_n8471);
nor_4  g20304(new_n22653, new_n8475, new_n22652);
nor_4  g20305(new_n22654, new_n8480_1, new_n22653);
nor_4  g20306(new_n22655, new_n22654, new_n22535);
not_3  g20307(new_n22656, new_n22535);
not_3  g20308(new_n22657, new_n22654);
nor_4  g20309(new_n22658, new_n22657, new_n22656);
nor_4  g20310(new_n22659, new_n22658, new_n22655);
not_3  g20311(new_n22660_1, new_n22659);
nand_4 g20312(new_n22661, new_n22656, new_n8486);
nand_4 g20313(new_n22662, new_n22550, new_n22536);
nand_4 g20314(new_n22663, new_n22662, new_n22661);
nor_4  g20315(new_n22664, new_n22663, new_n22660_1);
nor_4  g20316(n5325, new_n22664, new_n22655);
xor_3  g20317(new_n22666, n25120, n17458);
not_3  g20318(new_n22667, n8363);
nand_4 g20319(new_n22668, new_n22667, new_n8501);
xor_3  g20320(new_n22669, n8363, n1222);
nand_4 g20321(new_n22670, new_n8503, new_n9083);
xor_3  g20322(new_n22671, n25240, n14680);
nand_4 g20323(new_n22672, new_n9087, new_n8506);
xor_3  g20324(new_n22673, n17250, n10125);
nand_4 g20325(new_n22674, n23160, n8067);
not_3  g20326(new_n22675, new_n22674);
nor_4  g20327(new_n22676, n23160, n8067);
nor_4  g20328(new_n22677, n20923, n16524);
not_3  g20329(new_n22678, new_n22677);
not_3  g20330(new_n22679, new_n15657);
nand_4 g20331(new_n22680, new_n7789, new_n7778);
nand_4 g20332(new_n22681, new_n22680, new_n22679);
nand_4 g20333(new_n22682, new_n22681, new_n15655);
nand_4 g20334(new_n22683, new_n22682, new_n22678);
nor_4  g20335(new_n22684, new_n22683, new_n22676);
nor_4  g20336(new_n22685, new_n22684, new_n22675);
nand_4 g20337(new_n22686, new_n22685, new_n22673);
nand_4 g20338(new_n22687, new_n22686, new_n22672);
nand_4 g20339(new_n22688, new_n22687, new_n22671);
nand_4 g20340(new_n22689, new_n22688, new_n22670);
nand_4 g20341(new_n22690, new_n22689, new_n22669);
nand_4 g20342(new_n22691, new_n22690, new_n22668);
not_3  g20343(new_n22692, new_n22691);
xor_3  g20344(new_n22693, new_n22692, new_n22666);
not_3  g20345(new_n22694, new_n22693);
nand_4 g20346(new_n22695, new_n22694, new_n4907);
xnor_3 g20347(new_n22696, new_n22693, new_n4907);
xnor_3 g20348(new_n22697_1, new_n22689, new_n22669);
nor_4  g20349(new_n22698, new_n22697_1, n11481);
not_3  g20350(new_n22699, new_n22698);
not_3  g20351(new_n22700, n11481);
xnor_3 g20352(new_n22701, new_n22697_1, new_n22700);
not_3  g20353(new_n22702, n16439);
xnor_3 g20354(new_n22703, new_n22687, new_n22671);
not_3  g20355(new_n22704, new_n22703);
nand_4 g20356(new_n22705, new_n22704, new_n22702);
xnor_3 g20357(new_n22706, new_n22703, new_n22702);
xnor_3 g20358(new_n22707, new_n22685, new_n22673);
nor_4  g20359(new_n22708, new_n22707, n15241);
not_3  g20360(new_n22709, new_n22708);
xnor_3 g20361(new_n22710, new_n22707, new_n4922);
nor_4  g20362(new_n22711, new_n22676, new_n22675);
not_3  g20363(new_n22712, new_n22711);
xnor_3 g20364(new_n22713, new_n22712, new_n22683);
nand_4 g20365(new_n22714_1, new_n22713, new_n12765);
xnor_3 g20366(new_n22715, new_n22713, n7678);
not_3  g20367(new_n22716, new_n15660);
nand_4 g20368(new_n22717, new_n15665, new_n15663);
nand_4 g20369(new_n22718, new_n22717, new_n22716);
nand_4 g20370(new_n22719, new_n22718, new_n22715);
nand_4 g20371(new_n22720, new_n22719, new_n22714_1);
nand_4 g20372(new_n22721, new_n22720, new_n22710);
nand_4 g20373(new_n22722, new_n22721, new_n22709);
nand_4 g20374(new_n22723, new_n22722, new_n22706);
nand_4 g20375(new_n22724, new_n22723, new_n22705);
nand_4 g20376(new_n22725, new_n22724, new_n22701);
nand_4 g20377(new_n22726, new_n22725, new_n22699);
nand_4 g20378(new_n22727, new_n22726, new_n22696);
nand_4 g20379(new_n22728, new_n22727, new_n22695);
nor_4  g20380(new_n22729, n25120, n17458);
not_3  g20381(new_n22730, new_n22666);
nor_4  g20382(new_n22731, new_n22692, new_n22730);
nor_4  g20383(new_n22732, new_n22731, new_n22729);
not_3  g20384(new_n22733, new_n22732);
nor_4  g20385(new_n22734, new_n22733, new_n22728);
not_3  g20386(new_n22735, new_n22734);
xor_3  g20387(new_n22736, n12702, n12507);
nand_4 g20388(new_n22737, new_n6433, new_n10438);
xor_3  g20389(new_n22738, n26797, n15077);
nor_4  g20390(new_n22739, n23913, n3710);
not_3  g20391(new_n22740, new_n22739);
xor_3  g20392(new_n22741, n23913, n3710);
nor_4  g20393(new_n22742, n26318, n22554);
not_3  g20394(new_n22743, new_n22742);
xor_3  g20395(new_n22744, n26318, n22554);
nor_4  g20396(new_n22745, n26054, n20429);
not_3  g20397(new_n22746, new_n22745);
xor_3  g20398(new_n22747, n26054, n20429);
nor_4  g20399(new_n22748, n19081, n3909);
not_3  g20400(new_n22749, new_n22748);
xor_3  g20401(new_n22750, n19081, n3909);
nor_4  g20402(new_n22751, n23974, n8309);
not_3  g20403(new_n22752, new_n22751);
xor_3  g20404(new_n22753, n23974, n8309);
nand_4 g20405(new_n22754, n19144, n2146);
not_3  g20406(new_n22755, new_n22754);
nor_4  g20407(new_n22756, n19144, n2146);
nor_4  g20408(new_n22757, n22173, n12593);
nor_4  g20409(new_n22758, new_n20428, new_n20427);
nor_4  g20410(new_n22759, new_n22758, new_n22757);
not_3  g20411(new_n22760, new_n22759);
nor_4  g20412(new_n22761_1, new_n22760, new_n22756);
nor_4  g20413(new_n22762, new_n22761_1, new_n22755);
nand_4 g20414(new_n22763, new_n22762, new_n22753);
nand_4 g20415(new_n22764_1, new_n22763, new_n22752);
nand_4 g20416(new_n22765, new_n22764_1, new_n22750);
nand_4 g20417(new_n22766, new_n22765, new_n22749);
nand_4 g20418(new_n22767, new_n22766, new_n22747);
nand_4 g20419(new_n22768, new_n22767, new_n22746);
nand_4 g20420(new_n22769, new_n22768, new_n22744);
nand_4 g20421(new_n22770, new_n22769, new_n22743);
nand_4 g20422(new_n22771, new_n22770, new_n22741);
nand_4 g20423(new_n22772, new_n22771, new_n22740);
nand_4 g20424(new_n22773, new_n22772, new_n22738);
nand_4 g20425(new_n22774, new_n22773, new_n22737);
not_3  g20426(new_n22775, new_n22774);
xor_3  g20427(new_n22776, new_n22775, new_n22736);
not_3  g20428(new_n22777, new_n22776);
nand_4 g20429(new_n22778, new_n22777, new_n6510);
xnor_3 g20430(new_n22779_1, new_n22776, new_n6510);
xnor_3 g20431(new_n22780, new_n22772, new_n22738);
nor_4  g20432(new_n22781, new_n22780, n10201);
not_3  g20433(new_n22782, new_n22781);
not_3  g20434(new_n22783, n10201);
not_3  g20435(new_n22784, new_n22780);
xor_3  g20436(new_n22785, new_n22784, new_n22783);
xnor_3 g20437(new_n22786, new_n22770, new_n22741);
nor_4  g20438(new_n22787_1, new_n22786, n10593);
not_3  g20439(new_n22788, new_n22787_1);
not_3  g20440(new_n22789, new_n22786);
xor_3  g20441(new_n22790, new_n22789, new_n10735);
xnor_3 g20442(new_n22791, new_n22768, new_n22744);
nor_4  g20443(new_n22792, new_n22791, n18290);
not_3  g20444(new_n22793_1, new_n22792);
not_3  g20445(new_n22794, new_n22747);
xnor_3 g20446(new_n22795, new_n22766, new_n22794);
nand_4 g20447(new_n22796, new_n22795, new_n10744);
xnor_3 g20448(new_n22797, new_n22795, n11580);
not_3  g20449(new_n22798, new_n22750);
xnor_3 g20450(new_n22799, new_n22764_1, new_n22798);
nand_4 g20451(new_n22800, new_n22799, new_n6463);
xnor_3 g20452(new_n22801, new_n22799, n15884);
not_3  g20453(new_n22802, new_n22753);
xnor_3 g20454(new_n22803, new_n22762, new_n22802);
nand_4 g20455(new_n22804, new_n22803, new_n6488);
nor_4  g20456(new_n22805, new_n22756, new_n22755);
xor_3  g20457(new_n22806, new_n22805, new_n22760);
nor_4  g20458(new_n22807, new_n22806, new_n6475);
xor_3  g20459(new_n22808, new_n22805, new_n22759);
xnor_3 g20460(new_n22809, new_n22808, n27104);
not_3  g20461(new_n22810, new_n20433);
nand_4 g20462(new_n22811, new_n20435, new_n20422);
nand_4 g20463(new_n22812, new_n22811, new_n22810);
nor_4  g20464(new_n22813, new_n22812, new_n22809);
nor_4  g20465(new_n22814, new_n22813, new_n22807);
xor_3  g20466(new_n22815, new_n22803, new_n6488);
nand_4 g20467(new_n22816, new_n22815, new_n22814);
nand_4 g20468(new_n22817, new_n22816, new_n22804);
nand_4 g20469(new_n22818, new_n22817, new_n22801);
nand_4 g20470(new_n22819_1, new_n22818, new_n22800);
nand_4 g20471(new_n22820, new_n22819_1, new_n22797);
nand_4 g20472(new_n22821, new_n22820, new_n22796);
not_3  g20473(new_n22822, new_n22791);
xor_3  g20474(new_n22823, new_n22822, new_n10738);
nand_4 g20475(new_n22824, new_n22823, new_n22821);
nand_4 g20476(new_n22825, new_n22824, new_n22793_1);
nand_4 g20477(new_n22826, new_n22825, new_n22790);
nand_4 g20478(new_n22827, new_n22826, new_n22788);
nand_4 g20479(new_n22828, new_n22827, new_n22785);
nand_4 g20480(new_n22829, new_n22828, new_n22782);
nand_4 g20481(new_n22830, new_n22829, new_n22779_1);
nand_4 g20482(new_n22831, new_n22830, new_n22778);
nor_4  g20483(new_n22832, n12702, n12507);
not_3  g20484(new_n22833, new_n22736);
nor_4  g20485(new_n22834, new_n22775, new_n22833);
nor_4  g20486(new_n22835, new_n22834, new_n22832);
not_3  g20487(new_n22836, new_n22835);
nor_4  g20488(new_n22837, new_n22836, new_n22831);
nor_4  g20489(new_n22838, new_n22837, new_n22735);
not_3  g20490(new_n22839, new_n22837);
nor_4  g20491(new_n22840, new_n22839, new_n22734);
nor_4  g20492(new_n22841, new_n22840, new_n22838);
xnor_3 g20493(new_n22842, new_n22733, new_n22728);
not_3  g20494(new_n22843_1, new_n22842);
xnor_3 g20495(new_n22844, new_n22836, new_n22831);
nand_4 g20496(new_n22845, new_n22844, new_n22843_1);
xnor_3 g20497(new_n22846, new_n22844, new_n22842);
xnor_3 g20498(new_n22847, new_n22726, new_n22696);
not_3  g20499(new_n22848, new_n22829);
xnor_3 g20500(new_n22849, new_n22848, new_n22779_1);
nand_4 g20501(new_n22850, new_n22849, new_n22847);
not_3  g20502(new_n22851, new_n22725);
nor_4  g20503(new_n22852, new_n22851, new_n22698);
xnor_3 g20504(new_n22853, new_n22852, new_n22696);
xnor_3 g20505(new_n22854, new_n22849, new_n22853);
xnor_3 g20506(new_n22855, new_n22724, new_n22701);
not_3  g20507(new_n22856, new_n22785);
xnor_3 g20508(new_n22857, new_n22827, new_n22856);
nand_4 g20509(new_n22858_1, new_n22857, new_n22855);
nor_4  g20510(new_n22859, new_n22724, new_n22701);
nor_4  g20511(new_n22860, new_n22859, new_n22851);
xnor_3 g20512(new_n22861, new_n22857, new_n22860);
xnor_3 g20513(new_n22862, new_n22722, new_n22706);
xor_3  g20514(new_n22863, new_n22789, n10593);
xnor_3 g20515(new_n22864, new_n22825, new_n22863);
nand_4 g20516(new_n22865, new_n22864, new_n22862);
xor_3  g20517(new_n22866, new_n22704, n16439);
xnor_3 g20518(new_n22867, new_n22722, new_n22866);
xnor_3 g20519(new_n22868, new_n22864, new_n22867);
xnor_3 g20520(new_n22869, new_n22720, new_n22710);
xor_3  g20521(new_n22870_1, new_n22822, n18290);
xnor_3 g20522(new_n22871_1, new_n22870_1, new_n22821);
nand_4 g20523(new_n22872, new_n22871_1, new_n22869);
xnor_3 g20524(new_n22873, new_n22707, n15241);
xnor_3 g20525(new_n22874, new_n22720, new_n22873);
xnor_3 g20526(new_n22875, new_n22871_1, new_n22874);
not_3  g20527(new_n22876, new_n22797);
xnor_3 g20528(new_n22877, new_n22819_1, new_n22876);
xnor_3 g20529(new_n22878, new_n22718, new_n22715);
nand_4 g20530(new_n22879_1, new_n22878, new_n22877);
not_3  g20531(new_n22880, new_n22715);
xnor_3 g20532(new_n22881, new_n22718, new_n22880);
xnor_3 g20533(new_n22882, new_n22881, new_n22877);
not_3  g20534(new_n22883, new_n22801);
xnor_3 g20535(new_n22884, new_n22817, new_n22883);
nand_4 g20536(new_n22885, new_n22884, new_n15666);
nor_4  g20537(new_n22886, new_n15675, new_n7803);
xnor_3 g20538(new_n22887, new_n22886, new_n15663);
xnor_3 g20539(new_n22888, new_n22884, new_n22887);
xor_3  g20540(new_n22889, new_n22803, n6356);
xnor_3 g20541(new_n22890, new_n22889, new_n22814);
nand_4 g20542(new_n22891_1, new_n22890, new_n7825);
xnor_3 g20543(new_n22892, new_n22812, new_n22809);
nand_4 g20544(new_n22893, new_n22892, new_n7831);
not_3  g20545(new_n22894, new_n22893);
nor_4  g20546(new_n22895, new_n22892, new_n7831);
nor_4  g20547(new_n22896, new_n22895, new_n22894);
nor_4  g20548(new_n22897_1, new_n20437, new_n20425);
nor_4  g20549(new_n22898, new_n20438, new_n7837);
nor_4  g20550(new_n22899, new_n22898, new_n22897_1);
nand_4 g20551(new_n22900, new_n22899, new_n22896);
nand_4 g20552(new_n22901, new_n22900, new_n22893);
xnor_3 g20553(new_n22902, new_n22890, new_n15677);
nand_4 g20554(new_n22903_1, new_n22902, new_n22901);
nand_4 g20555(new_n22904, new_n22903_1, new_n22891_1);
nand_4 g20556(new_n22905, new_n22904, new_n22888);
nand_4 g20557(new_n22906, new_n22905, new_n22885);
nand_4 g20558(new_n22907_1, new_n22906, new_n22882);
nand_4 g20559(new_n22908, new_n22907_1, new_n22879_1);
nand_4 g20560(new_n22909, new_n22908, new_n22875);
nand_4 g20561(new_n22910_1, new_n22909, new_n22872);
nand_4 g20562(new_n22911, new_n22910_1, new_n22868);
nand_4 g20563(new_n22912, new_n22911, new_n22865);
nand_4 g20564(new_n22913, new_n22912, new_n22861);
nand_4 g20565(new_n22914_1, new_n22913, new_n22858_1);
nand_4 g20566(new_n22915, new_n22914_1, new_n22854);
nand_4 g20567(new_n22916, new_n22915, new_n22850);
nand_4 g20568(new_n22917, new_n22916, new_n22846);
nand_4 g20569(new_n22918_1, new_n22917, new_n22845);
xnor_3 g20570(n5351, new_n22918_1, new_n22841);
nor_4  g20571(n5353, new_n20055, new_n20047);
nor_4  g20572(new_n22921, new_n14253, n2160);
not_3  g20573(new_n22922, new_n22921);
nand_4 g20574(new_n22923, new_n14311, new_n14254);
nand_4 g20575(new_n22924, new_n22923, new_n22922);
nor_4  g20576(new_n22925, n9934, n2272);
nor_4  g20577(new_n22926, new_n14252, new_n14212);
nor_4  g20578(new_n22927, new_n22926, new_n22925);
nor_4  g20579(new_n22928, new_n22927, new_n22924);
not_3  g20580(new_n22929, new_n14319);
nor_4  g20581(new_n22930, new_n22929, n21784);
nor_4  g20582(new_n22931, new_n22930, new_n8567);
not_3  g20583(new_n22932, new_n22931);
nor_4  g20584(new_n22933, new_n14320, new_n8573);
not_3  g20585(new_n22934, new_n14344);
nor_4  g20586(new_n22935, new_n22934, new_n14321);
nor_4  g20587(new_n22936, new_n22935, new_n22933);
nor_4  g20588(new_n22937, new_n22936, new_n22932);
not_3  g20589(new_n22938, new_n22937);
xnor_3 g20590(new_n22939_1, new_n22938, new_n22928);
xnor_3 g20591(new_n22940, new_n22927, new_n22924);
xor_3  g20592(new_n22941, new_n22930, new_n8567);
xnor_3 g20593(new_n22942, new_n22941, new_n22936);
nor_4  g20594(new_n22943, new_n22942, new_n22940);
not_3  g20595(new_n22944, new_n22943);
xnor_3 g20596(new_n22945, new_n22942, new_n22940);
not_3  g20597(new_n22946, new_n22945);
nor_4  g20598(new_n22947, new_n14345_1, new_n14312);
not_3  g20599(new_n22948, new_n22947);
not_3  g20600(new_n22949, new_n14346);
not_3  g20601(new_n22950, new_n14349);
xnor_3 g20602(new_n22951, new_n14309, new_n14260);
nor_4  g20603(new_n22952, new_n20532, new_n22951);
nor_4  g20604(new_n22953, new_n22952, new_n14349);
nand_4 g20605(new_n22954, new_n14396, new_n22953);
nand_4 g20606(new_n22955, new_n22954, new_n22950);
nand_4 g20607(new_n22956, new_n22955, new_n22949);
nand_4 g20608(new_n22957, new_n22956, new_n22948);
nand_4 g20609(new_n22958, new_n22957, new_n22946);
nand_4 g20610(new_n22959, new_n22958, new_n22944);
xnor_3 g20611(n5399, new_n22959, new_n22939_1);
nor_4  g20612(new_n22961, new_n21403, new_n21400);
nor_4  g20613(new_n22962, new_n22961, new_n21398_1);
nor_4  g20614(new_n22963, new_n21394, new_n21389);
nor_4  g20615(new_n22964, new_n22963, new_n21390);
nor_4  g20616(new_n22965, new_n22964, new_n17234);
not_3  g20617(new_n22966, new_n22965);
nor_4  g20618(new_n22967, new_n22966, new_n22962);
xnor_3 g20619(new_n22968, new_n22967, new_n22937);
xnor_3 g20620(new_n22969, new_n22965, new_n22962);
nor_4  g20621(new_n22970, new_n22969, new_n22942);
not_3  g20622(new_n22971, new_n21404_1);
nor_4  g20623(new_n22972, new_n22971, new_n14345_1);
nor_4  g20624(new_n22973, new_n21409, new_n21405);
nor_4  g20625(new_n22974, new_n22973, new_n22972);
xnor_3 g20626(new_n22975, new_n22969, new_n22942);
nor_4  g20627(new_n22976, new_n22975, new_n22974);
nor_4  g20628(new_n22977, new_n22976, new_n22970);
xnor_3 g20629(n5403, new_n22977, new_n22968);
not_3  g20630(new_n22979, new_n18998);
xor_3  g20631(n5430, new_n19036, new_n22979);
not_3  g20632(new_n22981, new_n17755);
nor_4  g20633(new_n22982, new_n22981, new_n17749_1);
nand_4 g20634(new_n22983, new_n17756, new_n17740);
nand_4 g20635(new_n22984, new_n22983, new_n17743);
nor_4  g20636(new_n22985, new_n22984, new_n12368);
not_3  g20637(new_n22986, new_n22985);
nor_4  g20638(n5439, new_n22986, new_n22982);
not_3  g20639(new_n22988, new_n14775);
xor_3  g20640(n5472, new_n14798, new_n22988);
xnor_3 g20641(n5485, new_n9990, new_n9942_1);
xnor_3 g20642(n5524, new_n22304, new_n22278);
nor_4  g20643(new_n22992, new_n20067, new_n6982);
not_3  g20644(new_n22993, new_n22992);
nor_4  g20645(new_n22994, new_n22993, new_n6971_1);
nand_4 g20646(new_n22995, new_n22994, new_n6963);
not_3  g20647(new_n22996, new_n22995);
nand_4 g20648(new_n22997, new_n22996, new_n6955);
nor_4  g20649(new_n22998_1, new_n22997, new_n6945);
not_3  g20650(new_n22999, new_n22998_1);
nor_4  g20651(new_n23000, new_n22999, new_n6937);
not_3  g20652(new_n23001, new_n23000);
nor_4  g20653(new_n23002, new_n23001, new_n6930);
not_3  g20654(new_n23003, new_n23002);
nor_4  g20655(new_n23004, new_n23003, new_n6925);
nor_4  g20656(new_n23005, new_n23002, new_n16281);
nor_4  g20657(new_n23006_1, new_n23005, new_n23004);
nor_4  g20658(new_n23007_1, new_n23006_1, new_n16692);
xnor_3 g20659(new_n23008, new_n23006_1, new_n16692);
nor_4  g20660(new_n23009_1, new_n23000, new_n6933);
nor_4  g20661(new_n23010, new_n23009_1, new_n23002);
nor_4  g20662(new_n23011, new_n23010, new_n16699);
xnor_3 g20663(new_n23012, new_n23010, new_n16699);
nor_4  g20664(new_n23013, new_n22998_1, new_n6938);
nor_4  g20665(new_n23014_1, new_n23013, new_n23000);
nor_4  g20666(new_n23015, new_n23014_1, new_n16706);
xnor_3 g20667(new_n23016, new_n23014_1, new_n16706);
xnor_3 g20668(new_n23017, new_n22997, new_n6945);
not_3  g20669(new_n23018, new_n23017);
nor_4  g20670(new_n23019, new_n23018, new_n16713);
xnor_3 g20671(new_n23020, new_n23017, new_n16713);
not_3  g20672(new_n23021, new_n16718);
xnor_3 g20673(new_n23022, new_n22995, new_n6952);
nand_4 g20674(new_n23023, new_n23022, new_n23021);
xnor_3 g20675(new_n23024, new_n23022, new_n16718);
xnor_3 g20676(new_n23025, new_n22994, new_n6963);
nand_4 g20677(new_n23026, new_n23025, new_n16730);
xnor_3 g20678(new_n23027, new_n23025, new_n16732);
nor_4  g20679(new_n23028, new_n22992, new_n6974);
nor_4  g20680(new_n23029, new_n23028, new_n22994);
not_3  g20681(new_n23030, new_n23029);
nand_4 g20682(new_n23031, new_n21413, new_n15802);
nand_4 g20683(new_n23032, new_n21415, new_n21414);
nand_4 g20684(new_n23033, new_n23032, new_n23031);
nand_4 g20685(new_n23034, new_n23033, new_n23030);
xnor_3 g20686(new_n23035_1, new_n23033, new_n23029);
nand_4 g20687(new_n23036, new_n23035_1, new_n15790);
nand_4 g20688(new_n23037, new_n23036, new_n23034);
nand_4 g20689(new_n23038, new_n23037, new_n23027);
nand_4 g20690(new_n23039_1, new_n23038, new_n23026);
nand_4 g20691(new_n23040, new_n23039_1, new_n23024);
nand_4 g20692(new_n23041, new_n23040, new_n23023);
nand_4 g20693(new_n23042, new_n23041, new_n23020);
not_3  g20694(new_n23043, new_n23042);
nor_4  g20695(new_n23044, new_n23043, new_n23019);
nor_4  g20696(new_n23045, new_n23044, new_n23016);
nor_4  g20697(new_n23046, new_n23045, new_n23015);
nor_4  g20698(new_n23047_1, new_n23046, new_n23012);
nor_4  g20699(new_n23048, new_n23047_1, new_n23011);
nor_4  g20700(new_n23049, new_n23048, new_n23008);
nor_4  g20701(new_n23050, new_n23049, new_n23007_1);
not_3  g20702(new_n23051, new_n23004);
nand_4 g20703(new_n23052, new_n23051, new_n16277);
nand_4 g20704(new_n23053, new_n23004, new_n16275_1);
nand_4 g20705(new_n23054, new_n23053, new_n23052);
nand_4 g20706(new_n23055, new_n23054, new_n16752);
not_3  g20707(new_n23056, new_n16752);
not_3  g20708(new_n23057, new_n23054);
nand_4 g20709(new_n23058_1, new_n23057, new_n23056);
nand_4 g20710(new_n23059, new_n23058_1, new_n23055);
xnor_3 g20711(new_n23060, new_n23059, new_n23050);
nor_4  g20712(new_n23061, new_n23060, new_n5462);
xnor_3 g20713(new_n23062, new_n23060, new_n5462);
xnor_3 g20714(new_n23063, new_n23048, new_n23008);
nor_4  g20715(new_n23064, new_n23063, new_n5660);
xnor_3 g20716(new_n23065_1, new_n23063, new_n5660);
xnor_3 g20717(new_n23066_1, new_n23046, new_n23012);
nor_4  g20718(new_n23067_1, new_n23066_1, new_n5666);
xnor_3 g20719(new_n23068_1, new_n23066_1, new_n5666);
xnor_3 g20720(new_n23069, new_n23044, new_n23016);
nor_4  g20721(new_n23070, new_n23069, new_n5676);
xnor_3 g20722(new_n23071, new_n23069, new_n5676);
nor_4  g20723(new_n23072, new_n23041, new_n23020);
nor_4  g20724(new_n23073, new_n23072, new_n23043);
nand_4 g20725(new_n23074, new_n23073, new_n5680_1);
xnor_3 g20726(new_n23075, new_n23073, new_n5679);
not_3  g20727(new_n23076, new_n23024);
xnor_3 g20728(new_n23077, new_n23039_1, new_n23076);
nand_4 g20729(new_n23078, new_n23077, new_n5687_1);
xnor_3 g20730(new_n23079, new_n23077, new_n5686);
not_3  g20731(new_n23080, new_n23027);
xnor_3 g20732(new_n23081, new_n23037, new_n23080);
nand_4 g20733(new_n23082, new_n23081, new_n5694);
xnor_3 g20734(new_n23083, new_n23081, new_n5693);
xnor_3 g20735(new_n23084, new_n23035_1, new_n15791);
nand_4 g20736(new_n23085, new_n23084, new_n5701);
not_3  g20737(new_n23086, new_n23084);
xnor_3 g20738(new_n23087, new_n23086, new_n5701);
nor_4  g20739(new_n23088, new_n21417, new_n5712);
nor_4  g20740(new_n23089, new_n21420, new_n21418);
nor_4  g20741(new_n23090, new_n23089, new_n23088);
nand_4 g20742(new_n23091, new_n23090, new_n23087);
nand_4 g20743(new_n23092, new_n23091, new_n23085);
nand_4 g20744(new_n23093, new_n23092, new_n23083);
nand_4 g20745(new_n23094, new_n23093, new_n23082);
nand_4 g20746(new_n23095, new_n23094, new_n23079);
nand_4 g20747(new_n23096, new_n23095, new_n23078);
nand_4 g20748(new_n23097, new_n23096, new_n23075);
nand_4 g20749(new_n23098, new_n23097, new_n23074);
not_3  g20750(new_n23099, new_n23098);
nor_4  g20751(new_n23100, new_n23099, new_n23071);
nor_4  g20752(new_n23101, new_n23100, new_n23070);
nor_4  g20753(new_n23102, new_n23101, new_n23068_1);
nor_4  g20754(new_n23103, new_n23102, new_n23067_1);
nor_4  g20755(new_n23104, new_n23103, new_n23065_1);
nor_4  g20756(new_n23105, new_n23104, new_n23064);
nor_4  g20757(new_n23106, new_n23105, new_n23062);
nor_4  g20758(new_n23107, new_n23106, new_n23061);
not_3  g20759(new_n23108, new_n23050);
nand_4 g20760(new_n23109, new_n23058_1, new_n23108);
nand_4 g20761(new_n23110, new_n23109, new_n23055);
nand_4 g20762(new_n23111, new_n23110, new_n23053);
xnor_3 g20763(n5564, new_n23111, new_n23107);
not_3  g20764(new_n23113, new_n8171);
xor_3  g20765(n5593, new_n8186, new_n23113);
xnor_3 g20766(new_n23115, new_n21473, new_n17265);
not_3  g20767(new_n23116, new_n19934);
nand_4 g20768(new_n23117, new_n23116, new_n17272);
xnor_3 g20769(new_n23118, new_n19934, new_n17272);
nand_4 g20770(new_n23119, new_n19940, new_n17277);
xnor_3 g20771(new_n23120_1, new_n19939, new_n17277);
nor_4  g20772(new_n23121, new_n19947, new_n17284);
not_3  g20773(new_n23122, new_n23121);
nor_4  g20774(new_n23123, new_n18712, new_n17282);
nor_4  g20775(new_n23124, new_n23123, new_n23121);
not_3  g20776(new_n23125, new_n20926);
nand_4 g20777(new_n23126, new_n20937, new_n20927);
nand_4 g20778(new_n23127, new_n23126, new_n23125);
nand_4 g20779(new_n23128, new_n23127, new_n23124);
nand_4 g20780(new_n23129, new_n23128, new_n23122);
nand_4 g20781(new_n23130, new_n23129, new_n23120_1);
nand_4 g20782(new_n23131, new_n23130, new_n23119);
nand_4 g20783(new_n23132, new_n23131, new_n23118);
nand_4 g20784(new_n23133, new_n23132, new_n23117);
xnor_3 g20785(n5603, new_n23133, new_n23115);
xor_3  g20786(new_n23135, n17911, new_n21167);
nor_4  g20787(new_n23136, new_n19389_1, n1654);
not_3  g20788(new_n23137, new_n23136);
xor_3  g20789(new_n23138, n21997, new_n9036);
nor_4  g20790(new_n23139, new_n10137, n13783);
not_3  g20791(new_n23140, new_n23139);
xor_3  g20792(new_n23141, n25119, new_n8849_1);
nor_4  g20793(new_n23142, n26660, new_n10139);
not_3  g20794(new_n23143, new_n23142);
xor_3  g20795(new_n23144, n26660, new_n10139);
nor_4  g20796(new_n23145, new_n10143, n3018);
not_3  g20797(new_n23146_1, new_n23145);
nor_4  g20798(new_n23147, n18537, new_n9045);
not_3  g20799(new_n23148, new_n23147);
nor_4  g20800(new_n23149, n7057, new_n2426);
nor_4  g20801(new_n23150, new_n21863, new_n21854);
nor_4  g20802(new_n23151, new_n23150, new_n23149);
nand_4 g20803(new_n23152, new_n23151, new_n23148);
nand_4 g20804(new_n23153, new_n23152, new_n23146_1);
nand_4 g20805(new_n23154, new_n23153, new_n23144);
nand_4 g20806(new_n23155, new_n23154, new_n23143);
nand_4 g20807(new_n23156, new_n23155, new_n23141);
nand_4 g20808(new_n23157, new_n23156, new_n23140);
nand_4 g20809(new_n23158, new_n23157, new_n23138);
nand_4 g20810(new_n23159, new_n23158, new_n23137);
not_3  g20811(new_n23160_1, new_n23159);
xor_3  g20812(new_n23161, new_n23160_1, new_n23135);
nor_4  g20813(new_n23162, new_n23161, new_n3187);
not_3  g20814(new_n23163, new_n23161);
nor_4  g20815(new_n23164, new_n23163, new_n22356);
nor_4  g20816(new_n23165, new_n23164, new_n23162);
xor_3  g20817(new_n23166_1, new_n23157, new_n23138);
nor_4  g20818(new_n23167, new_n23166_1, new_n3192);
xnor_3 g20819(new_n23168, new_n23166_1, new_n3192);
not_3  g20820(new_n23169, new_n23141);
xor_3  g20821(new_n23170, new_n23155, new_n23169);
nand_4 g20822(new_n23171, new_n23170, new_n3200);
not_3  g20823(new_n23172, new_n23171);
xnor_3 g20824(new_n23173, new_n23170, new_n3200);
xor_3  g20825(new_n23174, new_n23153, new_n23144);
nor_4  g20826(new_n23175, new_n23174, new_n3206);
xnor_3 g20827(new_n23176, new_n23174, new_n3206);
nor_4  g20828(new_n23177, new_n23147, new_n23145);
xor_3  g20829(new_n23178, new_n23177, new_n23151);
nand_4 g20830(new_n23179, new_n23178, new_n3211);
nor_4  g20831(new_n23180, new_n21864, new_n3216);
nor_4  g20832(new_n23181, new_n21885, new_n21865);
nor_4  g20833(new_n23182, new_n23181, new_n23180);
not_3  g20834(new_n23183, new_n23182);
xnor_3 g20835(new_n23184, new_n23178, new_n3211);
not_3  g20836(new_n23185, new_n23184);
nand_4 g20837(new_n23186, new_n23185, new_n23183);
nand_4 g20838(new_n23187, new_n23186, new_n23179);
nor_4  g20839(new_n23188, new_n23187, new_n23176);
nor_4  g20840(new_n23189, new_n23188, new_n23175);
nor_4  g20841(new_n23190, new_n23189, new_n23173);
nor_4  g20842(new_n23191, new_n23190, new_n23172);
nor_4  g20843(new_n23192, new_n23191, new_n23168);
nor_4  g20844(new_n23193, new_n23192, new_n23167);
xor_3  g20845(n5609, new_n23193, new_n23165);
not_3  g20846(new_n23195, new_n16176);
xor_3  g20847(n5634, new_n16206_1, new_n23195);
nor_4  g20848(new_n23197, new_n3330, n2978);
xor_3  g20849(new_n23198, n3425, new_n8789);
nor_4  g20850(new_n23199, n23697, new_n3464);
not_3  g20851(new_n23200_1, new_n23199);
xor_3  g20852(new_n23201, n23697, new_n3464);
nand_4 g20853(new_n23202, n20946, new_n8796);
nand_4 g20854(new_n23203, new_n22561, new_n22554_1);
nand_4 g20855(new_n23204, new_n23203, new_n23202);
nand_4 g20856(new_n23205, new_n23204, new_n23201);
nand_4 g20857(new_n23206, new_n23205, new_n23200_1);
and_4  g20858(new_n23207, new_n23206, new_n23198);
nor_4  g20859(new_n23208, new_n23207, new_n23197);
nor_4  g20860(new_n23209, new_n23208, new_n8651);
xor_3  g20861(new_n23210, new_n23206, new_n23198);
nor_4  g20862(new_n23211, new_n23210, new_n8711);
xnor_3 g20863(new_n23212, new_n23210, new_n8711);
xor_3  g20864(new_n23213, new_n23204, new_n23201);
nor_4  g20865(new_n23214, new_n23213, new_n8714);
xnor_3 g20866(new_n23215, new_n23213, new_n8714);
nor_4  g20867(new_n23216, new_n22562, new_n8722);
nand_4 g20868(new_n23217, new_n22573, new_n22563);
not_3  g20869(new_n23218, new_n23217);
nor_4  g20870(new_n23219, new_n23218, new_n23216);
nor_4  g20871(new_n23220, new_n23219, new_n23215);
nor_4  g20872(new_n23221, new_n23220, new_n23214);
nor_4  g20873(new_n23222, new_n23221, new_n23212);
nor_4  g20874(new_n23223, new_n23222, new_n23211);
xnor_3 g20875(new_n23224, new_n23208, new_n8651);
nor_4  g20876(new_n23225, new_n23224, new_n23223);
nor_4  g20877(new_n23226, new_n23225, new_n23209);
not_3  g20878(new_n23227, new_n23208);
and_4  g20879(new_n23228, new_n8567, new_n8546);
not_3  g20880(new_n23229, new_n8568);
not_3  g20881(new_n23230, new_n8650);
nor_4  g20882(new_n23231, new_n23230, new_n23229);
nor_4  g20883(new_n23232, new_n23231, new_n23228);
not_3  g20884(new_n23233, new_n23232);
nor_4  g20885(new_n23234, new_n23233, new_n23227);
nor_4  g20886(new_n23235, new_n23232, new_n23208);
nor_4  g20887(new_n23236, new_n23235, new_n23234);
xnor_3 g20888(n5643, new_n23236, new_n23226);
xor_3  g20889(new_n23238_1, n18035, new_n21430);
nor_4  g20890(new_n23239, n13851, new_n12668);
not_3  g20891(new_n23240, new_n23239);
nand_4 g20892(new_n23241, new_n18807, new_n18786);
nand_4 g20893(new_n23242, new_n23241, new_n23240);
xor_3  g20894(new_n23243, new_n23242, new_n23238_1);
xnor_3 g20895(new_n23244, new_n23243, new_n18227_1);
not_3  g20896(new_n23245, new_n18808);
nand_4 g20897(new_n23246, new_n23245, new_n18259);
xnor_3 g20898(new_n23247_1, new_n18808, new_n18259);
nand_4 g20899(new_n23248_1, new_n18813, new_n18265);
xnor_3 g20900(new_n23249, new_n18810, new_n18265);
nand_4 g20901(new_n23250_1, new_n18819, new_n18271);
xnor_3 g20902(new_n23251, new_n18816, new_n18271);
nand_4 g20903(new_n23252, new_n18822, new_n18275);
nand_4 g20904(new_n23253, new_n16838, new_n16499);
xnor_3 g20905(new_n23254, new_n16838, new_n16500);
nand_4 g20906(new_n23255, new_n16856, new_n16511);
not_3  g20907(new_n23256, new_n16511);
xnor_3 g20908(new_n23257, new_n16856, new_n23256);
not_3  g20909(new_n23258, new_n16520);
nor_4  g20910(new_n23259, new_n16863, new_n16513);
nor_4  g20911(new_n23260, new_n23259, new_n23258);
not_3  g20912(new_n23261, new_n23260);
not_3  g20913(new_n23262, new_n23259);
nor_4  g20914(new_n23263, new_n23262, new_n16520);
nor_4  g20915(new_n23264, new_n23263, new_n23260);
nand_4 g20916(new_n23265, new_n23264, new_n16870);
nand_4 g20917(new_n23266, new_n23265, new_n23261);
nand_4 g20918(new_n23267, new_n23266, new_n23257);
nand_4 g20919(new_n23268, new_n23267, new_n23255);
nand_4 g20920(new_n23269, new_n23268, new_n23254);
nand_4 g20921(new_n23270_1, new_n23269, new_n23253);
xnor_3 g20922(new_n23271, new_n18822, new_n18274_1);
nand_4 g20923(new_n23272_1, new_n23271, new_n23270_1);
nand_4 g20924(new_n23273, new_n23272_1, new_n23252);
nand_4 g20925(new_n23274, new_n23273, new_n23251);
nand_4 g20926(new_n23275, new_n23274, new_n23250_1);
nand_4 g20927(new_n23276, new_n23275, new_n23249);
nand_4 g20928(new_n23277, new_n23276, new_n23248_1);
nand_4 g20929(new_n23278, new_n23277, new_n23247_1);
nand_4 g20930(new_n23279, new_n23278, new_n23246);
xor_3  g20931(n5680, new_n23279, new_n23244);
not_3  g20932(new_n23281, new_n17864);
xor_3  g20933(n5687, new_n17867, new_n23281);
not_3  g20934(new_n23283, new_n19212);
xor_3  g20935(n5700, new_n19222, new_n23283);
not_3  g20936(new_n23285, new_n12571);
nor_4  g20937(new_n23286, new_n12637, new_n23285);
nor_4  g20938(new_n23287, new_n12638, new_n12571);
nor_4  g20939(n5732, new_n23287, new_n23286);
nor_4  g20940(new_n23289_1, n23775, n8381);
nand_4 g20941(new_n23290, n23775, n8381);
not_3  g20942(new_n23291, new_n23290);
nor_4  g20943(new_n23292, new_n23291, new_n23289_1);
nor_4  g20944(new_n23293, n20235, n8259);
nor_4  g20945(new_n23294, new_n22439, new_n22425);
nor_4  g20946(new_n23295, new_n23294, new_n23293);
xnor_3 g20947(new_n23296, new_n23295, new_n23292);
xnor_3 g20948(new_n23297, new_n23296, new_n2409_1);
nor_4  g20949(new_n23298, new_n22440, new_n2396);
nor_4  g20950(new_n23299, new_n22441, new_n22438);
nor_4  g20951(new_n23300, new_n23299, new_n23298);
xnor_3 g20952(new_n23301, new_n23300, new_n23297);
xor_3  g20953(new_n23302, n8869, new_n2366);
nand_4 g20954(new_n23303, n20138, new_n8273);
nand_4 g20955(new_n23304_1, new_n22432, new_n22431);
nand_4 g20956(new_n23305_1, new_n23304_1, new_n23303);
xnor_3 g20957(new_n23306, new_n23305_1, new_n23302);
xnor_3 g20958(new_n23307, new_n23306, new_n23301);
not_3  g20959(new_n23308, new_n23307);
nand_4 g20960(new_n23309, new_n22442_1, new_n22437);
nand_4 g20961(new_n23310, new_n23309, new_n22434);
xor_3  g20962(n5742, new_n23310, new_n23308);
not_3  g20963(new_n23312, new_n16526);
xor_3  g20964(n5765, new_n16529, new_n23312);
xnor_3 g20965(n5776, new_n15077_1, new_n15022);
not_3  g20966(new_n23315, new_n2975);
xor_3  g20967(n5782, new_n23315, new_n2929_1);
xor_3  g20968(new_n23317, n18901, n1163);
nor_4  g20969(new_n23318, n18537, n4376);
not_3  g20970(new_n23319, new_n23318);
xor_3  g20971(new_n23320, n18537, n4376);
nor_4  g20972(new_n23321, n14570, n7057);
not_3  g20973(new_n23322, new_n23321);
xor_3  g20974(new_n23323, n14570, n7057);
not_3  g20975(new_n23324, new_n23289_1);
not_3  g20976(new_n23325, new_n23295);
nand_4 g20977(new_n23326, new_n23325, new_n23292);
nand_4 g20978(new_n23327, new_n23326, new_n23324);
nand_4 g20979(new_n23328, new_n23327, new_n23323);
nand_4 g20980(new_n23329, new_n23328, new_n23322);
nand_4 g20981(new_n23330, new_n23329, new_n23320);
nand_4 g20982(new_n23331, new_n23330, new_n23319);
nor_4  g20983(new_n23332, new_n23331, new_n23317);
nand_4 g20984(new_n23333_1, new_n23331, new_n23317);
not_3  g20985(new_n23334, new_n23333_1);
nor_4  g20986(new_n23335, new_n23334, new_n23332);
xnor_3 g20987(new_n23336, new_n23335, new_n2439);
not_3  g20988(new_n23337, new_n23336);
xnor_3 g20989(new_n23338, new_n23329, new_n23320);
nor_4  g20990(new_n23339, new_n23338, new_n2432);
not_3  g20991(new_n23340, new_n23328);
nor_4  g20992(new_n23341_1, new_n23327, new_n23323);
nor_4  g20993(new_n23342_1, new_n23341_1, new_n23340);
nand_4 g20994(new_n23343, new_n23296, new_n2410);
nand_4 g20995(new_n23344, new_n23300, new_n23297);
nand_4 g20996(new_n23345, new_n23344, new_n23343);
nand_4 g20997(new_n23346, new_n23345, new_n23342_1);
not_3  g20998(new_n23347, new_n23346);
nor_4  g20999(new_n23348, new_n23345, new_n23342_1);
nor_4  g21000(new_n23349, new_n23348, new_n23347);
nand_4 g21001(new_n23350, new_n23349, new_n2417);
nand_4 g21002(new_n23351, new_n23350, new_n23346);
not_3  g21003(new_n23352, new_n23351);
xnor_3 g21004(new_n23353, new_n23338, new_n2432);
nor_4  g21005(new_n23354, new_n23353, new_n23352);
nor_4  g21006(new_n23355_1, new_n23354, new_n23339);
xnor_3 g21007(new_n23356, new_n23355_1, new_n23337);
xor_3  g21008(new_n23357, n23068, new_n20495_1);
nor_4  g21009(new_n23358, n19514, new_n17891);
xor_3  g21010(new_n23359, n19514, new_n17891);
not_3  g21011(new_n23360, new_n23359);
nor_4  g21012(new_n23361, n10053, new_n14280);
xor_3  g21013(new_n23362, n10053, n1118);
nor_4  g21014(new_n23363, n25974, new_n4199);
nor_4  g21015(new_n23364, new_n14285, n8399);
nor_4  g21016(new_n23365, new_n4203, n1630);
nor_4  g21017(new_n23366, n9507, new_n14287);
nor_4  g21018(new_n23367, new_n8820, n1451);
not_3  g21019(new_n23368, new_n23367);
nor_4  g21020(new_n23369_1, new_n23368, new_n23366);
nor_4  g21021(new_n23370, new_n23369_1, new_n23365);
nor_4  g21022(new_n23371_1, new_n23370, new_n23364);
nor_4  g21023(new_n23372, new_n23371_1, new_n23363);
not_3  g21024(new_n23373, new_n23372);
nor_4  g21025(new_n23374, new_n23373, new_n23362);
nor_4  g21026(new_n23375, new_n23374, new_n23361);
nor_4  g21027(new_n23376, new_n23375, new_n23360);
nor_4  g21028(new_n23377, new_n23376, new_n23358);
not_3  g21029(new_n23378, new_n23377);
xor_3  g21030(new_n23379, new_n23378, new_n23357);
not_3  g21031(new_n23380, new_n23379);
nor_4  g21032(new_n23381, new_n23380, new_n23356);
not_3  g21033(new_n23382, new_n23356);
nor_4  g21034(new_n23383, new_n23379, new_n23382);
nor_4  g21035(new_n23384, new_n23383, new_n23381);
not_3  g21036(new_n23385, new_n23384);
xor_3  g21037(new_n23386, new_n23375, new_n23359);
not_3  g21038(new_n23387, new_n23353);
nor_4  g21039(new_n23388, new_n23387, new_n23351);
nor_4  g21040(new_n23389, new_n23388, new_n23354);
nor_4  g21041(new_n23390, new_n23389, new_n23386);
xnor_3 g21042(new_n23391, new_n23349, new_n2417);
not_3  g21043(new_n23392, new_n23391);
xor_3  g21044(new_n23393, new_n23372, new_n23362);
nand_4 g21045(new_n23394, new_n23393, new_n23392);
xnor_3 g21046(new_n23395, new_n23393, new_n23391);
xor_3  g21047(new_n23396, n25974, n8399);
xor_3  g21048(new_n23397, new_n23396, new_n23370);
not_3  g21049(new_n23398, new_n23397);
nor_4  g21050(new_n23399, new_n23398, new_n23301);
not_3  g21051(new_n23400, new_n23399);
xor_3  g21052(new_n23401_1, new_n23398, new_n23301);
xor_3  g21053(new_n23402, n26979, new_n17944);
nor_4  g21054(new_n23403, new_n23402, new_n22428);
nor_4  g21055(new_n23404, new_n23366, new_n23365);
xor_3  g21056(new_n23405, new_n23404, new_n23367);
not_3  g21057(new_n23406, new_n23405);
nor_4  g21058(new_n23407, new_n23406, new_n23403);
not_3  g21059(new_n23408, new_n23407);
not_3  g21060(new_n23409, new_n22442_1);
not_3  g21061(new_n23410, new_n23403);
nor_4  g21062(new_n23411, new_n23405, new_n23410);
nor_4  g21063(new_n23412, new_n23411, new_n23407);
nand_4 g21064(new_n23413, new_n23412, new_n23409);
nand_4 g21065(new_n23414_1, new_n23413, new_n23408);
nand_4 g21066(new_n23415, new_n23414_1, new_n23401_1);
nand_4 g21067(new_n23416, new_n23415, new_n23400);
nand_4 g21068(new_n23417, new_n23416, new_n23395);
nand_4 g21069(new_n23418, new_n23417, new_n23394);
xnor_3 g21070(new_n23419, new_n23389, new_n23386);
nor_4  g21071(new_n23420, new_n23419, new_n23418);
nor_4  g21072(new_n23421, new_n23420, new_n23390);
xor_3  g21073(n5833, new_n23421, new_n23385);
not_3  g21074(new_n23423, new_n15037);
xor_3  g21075(n5840, new_n15073, new_n23423);
xor_3  g21076(n5841, new_n23185, new_n23183);
not_3  g21077(new_n23426, new_n15634);
xor_3  g21078(n5850, new_n23426, new_n15633);
not_3  g21079(new_n23428, new_n23254);
xor_3  g21080(n5903, new_n23268, new_n23428);
xnor_3 g21081(new_n23430_1, new_n20169_1, new_n10337);
nor_4  g21082(new_n23431, new_n20173, new_n10265);
not_3  g21083(new_n23432, new_n23431);
nand_4 g21084(new_n23433_1, new_n22617, new_n22599);
nand_4 g21085(new_n23434_1, new_n23433_1, new_n23432);
xnor_3 g21086(new_n23435, new_n23434_1, new_n23430_1);
not_3  g21087(new_n23436, new_n22577);
nor_4  g21088(new_n23437, new_n23436, n6513);
xor_3  g21089(new_n23438, new_n23437, new_n14831);
not_3  g21090(new_n23439, new_n23438);
xor_3  g21091(new_n23440, new_n23439, new_n10533);
nand_4 g21092(new_n23441, new_n22578, new_n10535);
nand_4 g21093(new_n23442, new_n22597_1, new_n22579);
nand_4 g21094(new_n23443, new_n23442, new_n23441);
xnor_3 g21095(new_n23444, new_n23443, new_n23440);
nor_4  g21096(new_n23445, new_n23444, new_n23435);
not_3  g21097(new_n23446, new_n23430_1);
xnor_3 g21098(new_n23447, new_n23434_1, new_n23446);
not_3  g21099(new_n23448, new_n23444);
nor_4  g21100(new_n23449, new_n23448, new_n23447);
nor_4  g21101(new_n23450_1, new_n23449, new_n23445);
not_3  g21102(new_n23451, new_n23450_1);
not_3  g21103(new_n23452, new_n22598);
nand_4 g21104(new_n23453, new_n22618, new_n23452);
nand_4 g21105(new_n23454, new_n22650, new_n22619_1);
nand_4 g21106(new_n23455, new_n23454, new_n23453);
xor_3  g21107(n5904, new_n23455, new_n23451);
xor_3  g21108(new_n23457, n27089, new_n10732);
not_3  g21109(new_n23458, n11841);
nand_4 g21110(new_n23459, n19701, new_n23458);
xor_3  g21111(new_n23460, n19701, new_n23458);
nor_4  g21112(new_n23461, new_n3038, n10710);
not_3  g21113(new_n23462, new_n23461);
xor_3  g21114(new_n23463_1, n23529, new_n3080);
nor_4  g21115(new_n23464, new_n10741, n20929);
not_3  g21116(new_n23465, new_n23464);
xor_3  g21117(new_n23466, n24620, new_n11610);
nor_4  g21118(new_n23467, n8006, new_n10746);
xor_3  g21119(new_n23468, n8006, new_n10746);
not_3  g21120(new_n23469, new_n23468);
nor_4  g21121(new_n23470, n25074, new_n10750);
xor_3  g21122(new_n23471_1, n25074, n12956);
nor_4  g21123(new_n23472, n18295, new_n4879);
nor_4  g21124(new_n23473, new_n10756_1, n16396);
nor_4  g21125(new_n23474, new_n4883, n6502);
nor_4  g21126(new_n23475, n9399, new_n11146);
nor_4  g21127(new_n23476, n15780, new_n4885);
not_3  g21128(new_n23477, new_n23476);
nor_4  g21129(new_n23478, new_n23477, new_n23475);
nor_4  g21130(new_n23479, new_n23478, new_n23474);
nor_4  g21131(new_n23480_1, new_n23479, new_n23473);
nor_4  g21132(new_n23481, new_n23480_1, new_n23472);
not_3  g21133(new_n23482, new_n23481);
nor_4  g21134(new_n23483, new_n23482, new_n23471_1);
nor_4  g21135(new_n23484, new_n23483, new_n23470);
nor_4  g21136(new_n23485, new_n23484, new_n23469);
nor_4  g21137(new_n23486, new_n23485, new_n23467);
not_3  g21138(new_n23487, new_n23486);
nand_4 g21139(new_n23488, new_n23487, new_n23466);
nand_4 g21140(new_n23489, new_n23488, new_n23465);
nand_4 g21141(new_n23490, new_n23489, new_n23463_1);
nand_4 g21142(new_n23491, new_n23490, new_n23462);
nand_4 g21143(new_n23492, new_n23491, new_n23460);
nand_4 g21144(new_n23493_1, new_n23492, new_n23459);
xor_3  g21145(new_n23494, new_n23493_1, new_n23457);
not_3  g21146(new_n23495, new_n23494);
xnor_3 g21147(new_n23496, new_n23495, new_n12240);
xnor_3 g21148(new_n23497, new_n23491, new_n23460);
nand_4 g21149(new_n23498, new_n23497, new_n12246);
xnor_3 g21150(new_n23499, new_n23497, new_n12245);
not_3  g21151(new_n23500, new_n23463_1);
xor_3  g21152(new_n23501, new_n23489, new_n23500);
nand_4 g21153(new_n23502, new_n23501, new_n12252);
xnor_3 g21154(new_n23503, new_n23501, new_n12251);
xor_3  g21155(new_n23504, new_n23487, new_n23466);
not_3  g21156(new_n23505, new_n23504);
nand_4 g21157(new_n23506, new_n23505, new_n12258);
xor_3  g21158(new_n23507, new_n23484, new_n23469);
not_3  g21159(new_n23508, new_n23507);
nand_4 g21160(new_n23509, new_n23508, new_n12262);
xnor_3 g21161(new_n23510, new_n23507, new_n12262);
xor_3  g21162(new_n23511, new_n23482, new_n23471_1);
not_3  g21163(new_n23512, new_n23511);
nand_4 g21164(new_n23513_1, new_n23512, new_n12265);
not_3  g21165(new_n23514, new_n23479);
nor_4  g21166(new_n23515, new_n23473, new_n23472);
xor_3  g21167(new_n23516, new_n23515, new_n23514);
not_3  g21168(new_n23517, new_n23516);
nor_4  g21169(new_n23518, new_n23517, new_n12269);
not_3  g21170(new_n23519, new_n23518);
nor_4  g21171(new_n23520, new_n23516, new_n12276);
nor_4  g21172(new_n23521, new_n23520, new_n23518);
xor_3  g21173(new_n23522, n15780, new_n4885);
nor_4  g21174(new_n23523, new_n23522, new_n12280);
not_3  g21175(new_n23524, new_n23523);
nor_4  g21176(new_n23525, new_n23475, new_n23474);
xor_3  g21177(new_n23526, new_n23525, new_n23476);
nor_4  g21178(new_n23527, new_n23526, new_n23524);
not_3  g21179(new_n23528, new_n23526);
xor_3  g21180(new_n23529_1, new_n23528, new_n23524);
nor_4  g21181(new_n23530, new_n23529_1, new_n12289);
nor_4  g21182(new_n23531, new_n23530, new_n23527);
nand_4 g21183(new_n23532, new_n23531, new_n23521);
nand_4 g21184(new_n23533, new_n23532, new_n23519);
not_3  g21185(new_n23534, new_n23513_1);
nor_4  g21186(new_n23535, new_n23512, new_n12265);
nor_4  g21187(new_n23536, new_n23535, new_n23534);
nand_4 g21188(new_n23537, new_n23536, new_n23533);
nand_4 g21189(new_n23538, new_n23537, new_n23513_1);
nand_4 g21190(new_n23539, new_n23538, new_n23510);
nand_4 g21191(new_n23540, new_n23539, new_n23509);
xnor_3 g21192(new_n23541_1, new_n23504, new_n12258);
nand_4 g21193(new_n23542, new_n23541_1, new_n23540);
nand_4 g21194(new_n23543, new_n23542, new_n23506);
nand_4 g21195(new_n23544, new_n23543, new_n23503);
nand_4 g21196(new_n23545, new_n23544, new_n23502);
nand_4 g21197(new_n23546_1, new_n23545, new_n23499);
nand_4 g21198(new_n23547, new_n23546_1, new_n23498);
xnor_3 g21199(n5911, new_n23547, new_n23496);
xor_3  g21200(n5936, new_n14378, new_n4318);
xnor_3 g21201(n5943, new_n12083, new_n12042);
xnor_3 g21202(n5964, new_n17321, new_n17279);
not_3  g21203(new_n23552, new_n3466);
not_3  g21204(new_n23553, new_n5829);
nand_4 g21205(new_n23554, new_n5828, n11184);
not_3  g21206(new_n23555, new_n5812);
nand_4 g21207(new_n23556, new_n5811, n23146);
nor_4  g21208(new_n23557, new_n5805, n17968);
nand_4 g21209(new_n23558, new_n23557, new_n23556);
nand_4 g21210(new_n23559, new_n23558, new_n23555);
nand_4 g21211(new_n23560, new_n23559, new_n23554);
nand_4 g21212(new_n23561, new_n23560, new_n23553);
nand_4 g21213(new_n23562, new_n23561, new_n19502);
not_3  g21214(new_n23563, n8255);
not_3  g21215(new_n23564, new_n19495);
not_3  g21216(new_n23565, new_n23557);
nor_4  g21217(new_n23566, new_n23565, new_n5809);
nor_4  g21218(new_n23567, new_n23566, new_n5812);
nor_4  g21219(new_n23568, new_n23567, new_n5832);
nor_4  g21220(new_n23569, new_n23568, new_n5829);
nand_4 g21221(new_n23570, new_n23569, new_n23564);
nand_4 g21222(new_n23571, new_n23570, new_n23563);
nand_4 g21223(new_n23572, new_n23571, new_n23562);
nor_4  g21224(new_n23573, new_n23572, new_n19491);
xnor_3 g21225(new_n23574, new_n19495, new_n23563);
nor_4  g21226(new_n23575, new_n23569, new_n23574);
nor_4  g21227(new_n23576, new_n23561, new_n19495);
nor_4  g21228(new_n23577, new_n23576, n8255);
nor_4  g21229(new_n23578, new_n23577, new_n23575);
nor_4  g21230(new_n23579, new_n23578, new_n19556);
nor_4  g21231(new_n23580, new_n23579, new_n19553);
nor_4  g21232(new_n23581, new_n23580, new_n23573);
nor_4  g21233(new_n23582, new_n23581, new_n19485);
not_3  g21234(new_n23583, new_n23573);
nand_4 g21235(new_n23584, new_n23572, new_n19493);
nand_4 g21236(new_n23585_1, new_n23584, n8943);
nand_4 g21237(new_n23586_1, new_n23585_1, new_n23583);
nor_4  g21238(new_n23587, new_n23586_1, new_n19490);
nor_4  g21239(new_n23588_1, new_n23587, new_n19488);
nor_4  g21240(new_n23589, new_n23588_1, new_n23582);
nor_4  g21241(new_n23590, new_n23589, new_n19511);
not_3  g21242(new_n23591, new_n23582);
nand_4 g21243(new_n23592, new_n23581, new_n19544);
nand_4 g21244(new_n23593, new_n23592, n12380);
nand_4 g21245(new_n23594, new_n23593, new_n23591);
nor_4  g21246(new_n23595, new_n23594, new_n19513);
nor_4  g21247(new_n23596, new_n23595, new_n19481);
nor_4  g21248(new_n23597, new_n23596, new_n23590);
nor_4  g21249(new_n23598, new_n23597, new_n19478);
not_3  g21250(new_n23599, new_n23590);
nand_4 g21251(new_n23600, new_n23589, new_n19514_1);
nand_4 g21252(new_n23601, new_n23600, n8694);
nand_4 g21253(new_n23602, new_n23601, new_n23599);
nor_4  g21254(new_n23603, new_n23602, new_n19519);
nor_4  g21255(new_n23604, new_n23603, new_n19517);
nor_4  g21256(new_n23605, new_n23604, new_n23598);
xnor_3 g21257(new_n23606, new_n23605, new_n19476);
xnor_3 g21258(new_n23607, new_n23606, new_n23552);
xnor_3 g21259(new_n23608, new_n23602, new_n19519);
nor_4  g21260(new_n23609, new_n23608, new_n3471);
not_3  g21261(new_n23610, new_n23609);
not_3  g21262(new_n23611, new_n3471);
not_3  g21263(new_n23612, new_n23608);
nor_4  g21264(new_n23613, new_n23612, new_n23611);
nor_4  g21265(new_n23614, new_n23613, new_n23609);
xnor_3 g21266(new_n23615, new_n23589, new_n19514_1);
nor_4  g21267(new_n23616, new_n23615, new_n3479);
not_3  g21268(new_n23617, new_n23615);
nor_4  g21269(new_n23618, new_n23617, new_n3478);
nor_4  g21270(new_n23619_1, new_n23618, new_n23616);
not_3  g21271(new_n23620, new_n23619_1);
xnor_3 g21272(new_n23621, new_n23586_1, new_n19490);
nor_4  g21273(new_n23622, new_n23621, new_n3485);
xnor_3 g21274(new_n23623, new_n23621, new_n3485);
xnor_3 g21275(new_n23624_1, new_n23572, new_n19493);
nor_4  g21276(new_n23625, new_n23624_1, new_n3490);
xnor_3 g21277(new_n23626, new_n23624_1, new_n3490);
nor_4  g21278(new_n23627, new_n23561, new_n19502);
nor_4  g21279(new_n23628_1, new_n23627, new_n23575);
not_3  g21280(new_n23629, new_n23628_1);
nor_4  g21281(new_n23630, new_n23629, new_n3494);
xnor_3 g21282(new_n23631, new_n23629, new_n3494);
xnor_3 g21283(new_n23632, new_n23559, new_n5833_1);
nor_4  g21284(new_n23633, new_n23632, new_n3503);
xnor_3 g21285(new_n23634, new_n23632, new_n3503);
nor_4  g21286(new_n23635, new_n23565, new_n5813);
nor_4  g21287(new_n23636, new_n23557, new_n5841_1);
nor_4  g21288(new_n23637_1, new_n23636, new_n23635);
nor_4  g21289(new_n23638, new_n23637_1, new_n3515);
nor_4  g21290(new_n23639, new_n15768, new_n3510);
xnor_3 g21291(new_n23640, new_n23637_1, new_n3515);
nor_4  g21292(new_n23641, new_n23640, new_n23639);
nor_4  g21293(new_n23642, new_n23641, new_n23638);
nor_4  g21294(new_n23643, new_n23642, new_n23634);
nor_4  g21295(new_n23644, new_n23643, new_n23633);
nor_4  g21296(new_n23645, new_n23644, new_n23631);
nor_4  g21297(new_n23646, new_n23645, new_n23630);
nor_4  g21298(new_n23647, new_n23646, new_n23626);
nor_4  g21299(new_n23648, new_n23647, new_n23625);
nor_4  g21300(new_n23649, new_n23648, new_n23623);
nor_4  g21301(new_n23650, new_n23649, new_n23622);
nor_4  g21302(new_n23651, new_n23650, new_n23620);
nor_4  g21303(new_n23652, new_n23651, new_n23616);
not_3  g21304(new_n23653, new_n23652);
nand_4 g21305(new_n23654, new_n23653, new_n23614);
nand_4 g21306(new_n23655, new_n23654, new_n23610);
xor_3  g21307(n5980, new_n23655, new_n23607);
xnor_3 g21308(n6012, new_n13528, new_n13500_1);
nor_4  g21309(new_n23658, new_n12228_1, n16544);
nor_4  g21310(new_n23659, new_n12166, new_n10728);
nor_4  g21311(new_n23660, new_n23659, new_n23658);
not_3  g21312(new_n23661, new_n23660);
nor_4  g21313(new_n23662, new_n12172, n6814);
nor_4  g21314(new_n23663_1, new_n12170, new_n10732);
nor_4  g21315(new_n23664, new_n23663_1, new_n23662);
not_3  g21316(new_n23665, new_n23664);
nor_4  g21317(new_n23666, new_n12176, n19701);
not_3  g21318(new_n23667, n19701);
xnor_3 g21319(new_n23668, new_n12176, new_n23667);
nand_4 g21320(new_n23669_1, new_n12218, new_n3038);
nand_4 g21321(new_n23670, new_n11165, new_n11113);
nand_4 g21322(new_n23671, new_n23670, new_n23669_1);
nand_4 g21323(new_n23672, new_n23671, new_n23668);
not_3  g21324(new_n23673, new_n23672);
nor_4  g21325(new_n23674, new_n23673, new_n23666);
nor_4  g21326(new_n23675, new_n23674, new_n23665);
nor_4  g21327(new_n23676, new_n23675, new_n23662);
nor_4  g21328(new_n23677, new_n23676, new_n23661);
nor_4  g21329(new_n23678, new_n23677, new_n23658);
nand_4 g21330(new_n23679, new_n23678, new_n12161_1);
nor_4  g21331(new_n23680, new_n17104_1, n3582);
xnor_3 g21332(new_n23681, new_n17104_1, n3582);
nor_4  g21333(new_n23682, new_n17107, n2145);
xnor_3 g21334(new_n23683, new_n17107, n2145);
nor_4  g21335(new_n23684_1, new_n17113, n5031);
xnor_3 g21336(new_n23685, new_n17112, new_n9085);
not_3  g21337(new_n23686, new_n11199);
nand_4 g21338(new_n23687, new_n11241, new_n11201_1);
nand_4 g21339(new_n23688, new_n23687, new_n23686);
nor_4  g21340(new_n23689, new_n23688, new_n23685);
nor_4  g21341(new_n23690_1, new_n23689, new_n23684_1);
nor_4  g21342(new_n23691, new_n23690_1, new_n23683);
nor_4  g21343(new_n23692, new_n23691, new_n23682);
nor_4  g21344(new_n23693, new_n23692, new_n23681);
nor_4  g21345(new_n23694, new_n23693, new_n23680);
nand_4 g21346(new_n23695, new_n23694, new_n17162);
xnor_3 g21347(new_n23696, new_n23695, new_n23679);
xnor_3 g21348(new_n23697_1, new_n23678, new_n12161_1);
xnor_3 g21349(new_n23698, new_n23694, new_n17162);
not_3  g21350(new_n23699, new_n23698);
nand_4 g21351(new_n23700, new_n23699, new_n23697_1);
xnor_3 g21352(new_n23701, new_n23698, new_n23697_1);
xnor_3 g21353(new_n23702, new_n23676, new_n23660);
xnor_3 g21354(new_n23703, new_n23692, new_n23681);
nand_4 g21355(new_n23704, new_n23703, new_n23702);
not_3  g21356(new_n23705, new_n23703);
xnor_3 g21357(new_n23706, new_n23705, new_n23702);
xnor_3 g21358(new_n23707, new_n23674, new_n23664);
xnor_3 g21359(new_n23708, new_n23690_1, new_n23683);
nand_4 g21360(new_n23709, new_n23708, new_n23707);
not_3  g21361(new_n23710, new_n23708);
xnor_3 g21362(new_n23711, new_n23710, new_n23707);
xnor_3 g21363(new_n23712, new_n23671, new_n23668);
not_3  g21364(new_n23713, new_n23712);
nand_4 g21365(new_n23714_1, new_n23688, new_n23685);
not_3  g21366(new_n23715, new_n23714_1);
nor_4  g21367(new_n23716, new_n23715, new_n23689);
not_3  g21368(new_n23717_1, new_n23716);
nand_4 g21369(new_n23718, new_n23717_1, new_n23713);
xnor_3 g21370(new_n23719_1, new_n23717_1, new_n23712);
not_3  g21371(new_n23720, new_n11166);
nand_4 g21372(new_n23721, new_n11243, new_n23720);
nand_4 g21373(new_n23722, new_n11293, new_n11244);
nand_4 g21374(new_n23723, new_n23722, new_n23721);
nand_4 g21375(new_n23724, new_n23723, new_n23719_1);
nand_4 g21376(new_n23725, new_n23724, new_n23718);
nand_4 g21377(new_n23726, new_n23725, new_n23711);
nand_4 g21378(new_n23727, new_n23726, new_n23709);
nand_4 g21379(new_n23728, new_n23727, new_n23706);
nand_4 g21380(new_n23729, new_n23728, new_n23704);
nand_4 g21381(new_n23730, new_n23729, new_n23701);
nand_4 g21382(new_n23731, new_n23730, new_n23700);
xnor_3 g21383(n6022, new_n23731, new_n23696);
not_3  g21384(new_n23733, new_n23251);
xor_3  g21385(n6031, new_n23273, new_n23733);
nand_4 g21386(new_n23735, new_n20256, new_n8501);
xor_3  g21387(new_n23736, new_n23735, n17458);
nor_4  g21388(new_n23737, new_n23736, n12507);
not_3  g21389(new_n23738, new_n23736);
nor_4  g21390(new_n23739, new_n23738, new_n10423);
nor_4  g21391(new_n23740, new_n23739, new_n23737);
not_3  g21392(new_n23741, new_n20259_1);
not_3  g21393(new_n23742, new_n20260);
nand_4 g21394(new_n23743, new_n20313, new_n23742);
nand_4 g21395(new_n23744, new_n23743, new_n23741);
xnor_3 g21396(new_n23745, new_n23744, new_n23740);
not_3  g21397(new_n23746, new_n23745);
nor_4  g21398(new_n23747, new_n23746, n12702);
nor_4  g21399(new_n23748_1, new_n23745, new_n6505);
nor_4  g21400(new_n23749, new_n23748_1, new_n23747);
nand_4 g21401(new_n23750, new_n20314, new_n6433);
nand_4 g21402(new_n23751, new_n20369, new_n20315);
nand_4 g21403(new_n23752, new_n23751, new_n23750);
xnor_3 g21404(new_n23753, new_n23752, new_n23749);
xnor_3 g21405(new_n23754, new_n23753, new_n9660);
not_3  g21406(new_n23755_1, new_n20370);
nand_4 g21407(new_n23756, new_n23755_1, new_n9667);
nand_4 g21408(new_n23757, new_n20417, new_n20371);
nand_4 g21409(new_n23758, new_n23757, new_n23756);
xnor_3 g21410(n6044, new_n23758, new_n23754);
nand_4 g21411(new_n23760, new_n10931, new_n10883);
xnor_3 g21412(new_n23761, new_n12870_1, new_n10883);
nand_4 g21413(new_n23762, new_n11022, new_n23761);
nand_4 g21414(new_n23763, new_n23762, new_n23760);
not_3  g21415(new_n23764, new_n10882);
nor_4  g21416(new_n23765, new_n23764, n4306);
or_4   g21417(new_n23766, new_n22063_1, new_n23765);
nor_4  g21418(new_n23767, new_n23766, new_n23763);
xor_3  g21419(new_n23768, new_n22063_1, new_n23765);
xnor_3 g21420(new_n23769, new_n23768, new_n23763);
nor_4  g21421(new_n23770, new_n23769, new_n5132);
xnor_3 g21422(new_n23771, new_n23769, new_n5132);
nor_4  g21423(new_n23772, new_n11023_1, new_n5141);
nor_4  g21424(new_n23773, new_n11079, new_n11024);
nor_4  g21425(new_n23774, new_n23773, new_n23772);
nor_4  g21426(new_n23775_1, new_n23774, new_n23771);
nor_4  g21427(new_n23776, new_n23775_1, new_n23770);
nor_4  g21428(new_n23777, new_n23776, new_n23767);
nand_4 g21429(new_n23778, new_n23767, new_n4984);
nand_4 g21430(new_n23779, new_n23776, new_n5129);
nand_4 g21431(new_n23780, new_n23779, new_n23778);
nor_4  g21432(n6046, new_n23780, new_n23777);
xor_3  g21433(new_n23782, n17077, new_n14261);
nand_4 g21434(new_n23783, new_n3081, n20700);
xor_3  g21435(new_n23784, n26510, new_n3037);
nor_4  g21436(new_n23785, n23068, new_n20495_1);
not_3  g21437(new_n23786, new_n23785);
nand_4 g21438(new_n23787, new_n23378, new_n23357);
nand_4 g21439(new_n23788, new_n23787, new_n23786);
nand_4 g21440(new_n23789, new_n23788, new_n23784);
nand_4 g21441(new_n23790, new_n23789, new_n23783);
xor_3  g21442(new_n23791, new_n23790, new_n23782);
not_3  g21443(new_n23792, new_n23791);
xor_3  g21444(new_n23793, n21997, n18483);
nand_4 g21445(new_n23794, n25119, n21934);
not_3  g21446(new_n23795, new_n23794);
nor_4  g21447(new_n23796, n25119, n21934);
nor_4  g21448(new_n23797, n18901, n1163);
not_3  g21449(new_n23798, new_n23797);
nand_4 g21450(new_n23799, new_n23333_1, new_n23798);
nor_4  g21451(new_n23800, new_n23799, new_n23796);
nor_4  g21452(new_n23801, new_n23800, new_n23795);
xnor_3 g21453(new_n23802, new_n23801, new_n23793);
not_3  g21454(new_n23803, new_n23802);
nor_4  g21455(new_n23804, new_n23803, new_n8853);
not_3  g21456(new_n23805, new_n8853);
nor_4  g21457(new_n23806, new_n23802, new_n23805);
nor_4  g21458(new_n23807, new_n23806, new_n23804);
not_3  g21459(new_n23808, new_n2448);
nor_4  g21460(new_n23809, new_n23796, new_n23795);
xnor_3 g21461(new_n23810, new_n23809, new_n23799);
not_3  g21462(new_n23811, new_n23810);
nor_4  g21463(new_n23812, new_n23811, new_n23808);
not_3  g21464(new_n23813, new_n23812);
nor_4  g21465(new_n23814, new_n23335, new_n2439);
not_3  g21466(new_n23815, new_n23814);
nand_4 g21467(new_n23816, new_n23355_1, new_n23337);
nand_4 g21468(new_n23817, new_n23816, new_n23815);
xnor_3 g21469(new_n23818, new_n23810, new_n2448);
not_3  g21470(new_n23819, new_n23818);
nand_4 g21471(new_n23820, new_n23819, new_n23817);
nand_4 g21472(new_n23821, new_n23820, new_n23813);
xnor_3 g21473(new_n23822, new_n23821, new_n23807);
nor_4  g21474(new_n23823, new_n23822, new_n23792);
not_3  g21475(new_n23824, new_n23822);
nor_4  g21476(new_n23825, new_n23824, new_n23791);
nor_4  g21477(new_n23826, new_n23825, new_n23823);
xnor_3 g21478(new_n23827, new_n23788, new_n23784);
xnor_3 g21479(new_n23828, new_n23818, new_n23817);
not_3  g21480(new_n23829, new_n23828);
nand_4 g21481(new_n23830, new_n23829, new_n23827);
not_3  g21482(new_n23831_1, new_n23383);
nand_4 g21483(new_n23832, new_n23421, new_n23384);
nand_4 g21484(new_n23833, new_n23832, new_n23831_1);
xnor_3 g21485(new_n23834, new_n23828, new_n23827);
nand_4 g21486(new_n23835, new_n23834, new_n23833);
nand_4 g21487(new_n23836, new_n23835, new_n23830);
xnor_3 g21488(n6084, new_n23836, new_n23826);
xor_3  g21489(n6160, new_n23529_1, new_n12289);
not_3  g21490(new_n23839, new_n23533);
xor_3  g21491(n6171, new_n23536, new_n23839);
or_4   g21492(new_n23841, n22359, new_n11919);
nand_4 g21493(new_n23842_1, new_n18455, new_n11920);
nand_4 g21494(new_n23843, new_n23842_1, new_n23841);
xnor_3 g21495(new_n23844, new_n23843, new_n11926_1);
not_3  g21496(new_n23845, new_n23844);
xor_3  g21497(new_n23846, n26264, new_n11806);
nand_4 g21498(new_n23847, new_n11813, n7841);
xor_3  g21499(new_n23848, n22918, new_n9457);
nand_4 g21500(new_n23849_1, new_n11815, n16812);
xor_3  g21501(new_n23850, n25923, new_n9460_1);
nand_4 g21502(new_n23851, n25068, new_n11820);
nand_4 g21503(new_n23852, new_n22122, new_n22101);
nand_4 g21504(new_n23853, new_n23852, new_n23851);
nand_4 g21505(new_n23854, new_n23853, new_n23850);
nand_4 g21506(new_n23855, new_n23854, new_n23849_1);
nand_4 g21507(new_n23856_1, new_n23855, new_n23848);
nand_4 g21508(new_n23857, new_n23856_1, new_n23847);
xnor_3 g21509(new_n23858, new_n23857, new_n23846);
nor_4  g21510(new_n23859, new_n23858, new_n18909);
not_3  g21511(new_n23860, new_n23858);
nor_4  g21512(new_n23861, new_n23860, new_n18911);
nor_4  g21513(new_n23862, new_n23861, new_n23859);
not_3  g21514(new_n23863, new_n23848);
xnor_3 g21515(new_n23864, new_n23855, new_n23863);
nor_4  g21516(new_n23865, new_n23864, new_n18552);
xnor_3 g21517(new_n23866, new_n23864, new_n18548);
not_3  g21518(new_n23867, new_n23866);
xnor_3 g21519(new_n23868, new_n23853, new_n23850);
not_3  g21520(new_n23869, new_n23868);
nand_4 g21521(new_n23870, new_n23869, new_n18555);
xnor_3 g21522(new_n23871, new_n23869, new_n18555);
not_3  g21523(new_n23872, new_n23871);
nand_4 g21524(new_n23873, new_n22162, new_n22127);
nand_4 g21525(new_n23874, new_n23873, new_n22124_1);
nand_4 g21526(new_n23875, new_n23874, new_n23872);
nand_4 g21527(new_n23876, new_n23875, new_n23870);
nor_4  g21528(new_n23877, new_n23876, new_n23867);
nor_4  g21529(new_n23878, new_n23877, new_n23865);
nand_4 g21530(new_n23879, new_n23878, new_n23862);
not_3  g21531(new_n23880, new_n23879);
nor_4  g21532(new_n23881, new_n23878, new_n23862);
nor_4  g21533(new_n23882, new_n23881, new_n23880);
xnor_3 g21534(new_n23883_1, new_n23882, new_n23845);
not_3  g21535(new_n23884, new_n23876);
nor_4  g21536(new_n23885, new_n23884, new_n23866);
nor_4  g21537(new_n23886, new_n23885, new_n23877);
nand_4 g21538(new_n23887, new_n23886, new_n18457);
xnor_3 g21539(new_n23888_1, new_n23886, new_n18456);
not_3  g21540(new_n23889, new_n23875);
nor_4  g21541(new_n23890, new_n23874, new_n23872);
nor_4  g21542(new_n23891, new_n23890, new_n23889);
not_3  g21543(new_n23892, new_n23891);
nand_4 g21544(new_n23893, new_n23892, new_n18460);
xnor_3 g21545(new_n23894, new_n23891, new_n18460);
nand_4 g21546(new_n23895_1, new_n22163, new_n18463);
nand_4 g21547(new_n23896, new_n22201_1, new_n22164);
nand_4 g21548(new_n23897, new_n23896, new_n23895_1);
nand_4 g21549(new_n23898, new_n23897, new_n23894);
nand_4 g21550(new_n23899_1, new_n23898, new_n23893);
nand_4 g21551(new_n23900, new_n23899_1, new_n23888_1);
nand_4 g21552(new_n23901, new_n23900, new_n23887);
xor_3  g21553(n6183, new_n23901, new_n23883_1);
xor_3  g21554(new_n23903_1, n14702, new_n10893);
not_3  g21555(new_n23904, new_n23903_1);
nor_4  g21556(new_n23905, new_n10896, n2999);
not_3  g21557(new_n23906, new_n23905);
xor_3  g21558(new_n23907, n11356, new_n10958);
nor_4  g21559(new_n23908, new_n10898, n2547);
not_3  g21560(new_n23909, new_n23908);
xor_3  g21561(new_n23910, n3164, n2547);
not_3  g21562(new_n23911, new_n23910);
nor_4  g21563(new_n23912_1, n10611, new_n10980);
nor_4  g21564(new_n23913_1, new_n17062, new_n17046);
nor_4  g21565(new_n23914, new_n23913_1, new_n23912_1);
nand_4 g21566(new_n23915, new_n23914, new_n23911);
nand_4 g21567(new_n23916, new_n23915, new_n23909);
nand_4 g21568(new_n23917, new_n23916, new_n23907);
nand_4 g21569(new_n23918, new_n23917, new_n23906);
xor_3  g21570(new_n23919, new_n23918, new_n23904);
xnor_3 g21571(new_n23920, new_n23919, new_n10804);
xor_3  g21572(new_n23921, new_n23916, new_n23907);
not_3  g21573(new_n23922, new_n23921);
nand_4 g21574(new_n23923_1, new_n23922, new_n10810);
xnor_3 g21575(new_n23924_1, new_n23921, new_n10810);
xor_3  g21576(new_n23925, new_n23914, new_n23911);
not_3  g21577(new_n23926, new_n23925);
nand_4 g21578(new_n23927, new_n23926, new_n10816);
xnor_3 g21579(new_n23928, new_n23925, new_n10816);
nand_4 g21580(new_n23929, new_n17063, new_n10820);
nand_4 g21581(new_n23930, new_n17085, new_n17064);
nand_4 g21582(new_n23931, new_n23930, new_n23929);
nand_4 g21583(new_n23932, new_n23931, new_n23928);
nand_4 g21584(new_n23933, new_n23932, new_n23927);
nand_4 g21585(new_n23934, new_n23933, new_n23924_1);
nand_4 g21586(new_n23935_1, new_n23934, new_n23923_1);
xor_3  g21587(n6189, new_n23935_1, new_n23920);
xor_3  g21588(new_n23937, n20036, n15167);
nor_4  g21589(new_n23938, new_n7602, n11192);
nor_4  g21590(new_n23939, n21095, new_n4607);
nand_4 g21591(new_n23940, new_n4609, n8656);
nor_4  g21592(new_n23941, new_n23940, new_n23939);
nor_4  g21593(new_n23942_1, new_n23941, new_n23938);
xor_3  g21594(new_n23943, new_n23942_1, new_n23937);
xnor_3 g21595(new_n23944, new_n23943, new_n22180);
xor_3  g21596(new_n23945, n9380, new_n14848);
nor_4  g21597(new_n23946, new_n23945, new_n18304_1);
nor_4  g21598(new_n23947, new_n23939, new_n23938);
xor_3  g21599(new_n23948, new_n23947, new_n23940);
nor_4  g21600(new_n23949, new_n23948, new_n23946);
not_3  g21601(new_n23950, new_n23949);
not_3  g21602(new_n23951, new_n23946);
not_3  g21603(new_n23952, new_n23948);
xor_3  g21604(new_n23953, new_n23952, new_n23951);
nand_4 g21605(new_n23954_1, new_n23953, new_n22193);
nand_4 g21606(new_n23955, new_n23954_1, new_n23950);
not_3  g21607(new_n23956, new_n23955);
xor_3  g21608(n6223, new_n23956, new_n23944);
not_3  g21609(new_n23958_1, new_n17083);
xor_3  g21610(n6233, new_n23958_1, new_n17071);
xnor_3 g21611(n6245, new_n22957, new_n22946);
not_3  g21612(new_n23961, new_n12293);
xor_3  g21613(n6248, new_n23961, new_n12278);
xor_3  g21614(new_n23963, n21839, new_n10728);
not_3  g21615(new_n23964, new_n23963);
nor_4  g21616(new_n23965, n27089, new_n10732);
nand_4 g21617(new_n23966, new_n23493_1, new_n23457);
not_3  g21618(new_n23967, new_n23966);
nor_4  g21619(new_n23968, new_n23967, new_n23965);
xor_3  g21620(new_n23969, new_n23968, new_n23964);
xnor_3 g21621(new_n23970, new_n23969, new_n12236);
nor_4  g21622(new_n23971, new_n23494, new_n12240);
nand_4 g21623(new_n23972, new_n23547, new_n23496);
not_3  g21624(new_n23973, new_n23972);
nor_4  g21625(new_n23974_1, new_n23973, new_n23971);
xnor_3 g21626(n6256, new_n23974_1, new_n23970);
xnor_3 g21627(n6271, new_n18141, new_n18115);
nor_4  g21628(new_n23977, new_n11929, n13549);
nor_4  g21629(new_n23978, new_n11925, n8405);
nand_4 g21630(new_n23979, new_n23843, new_n11926_1);
not_3  g21631(new_n23980, new_n23979);
nor_4  g21632(new_n23981, new_n23980, new_n23978);
nor_4  g21633(new_n23982, new_n23981, new_n11931);
nor_4  g21634(new_n23983, new_n23982, new_n23977);
nor_4  g21635(new_n23984, n13951, new_n13250);
not_3  g21636(new_n23985, new_n23984);
xor_3  g21637(new_n23986_1, n13951, new_n13250);
nor_4  g21638(new_n23987, n22793, new_n2983);
not_3  g21639(new_n23988, new_n23987);
nand_4 g21640(new_n23989, new_n18187, new_n18163);
nand_4 g21641(new_n23990, new_n23989, new_n23988);
nand_4 g21642(new_n23991, new_n23990, new_n23986_1);
nand_4 g21643(new_n23992, new_n23991, new_n23985);
not_3  g21644(new_n23993, new_n23992);
nand_4 g21645(new_n23994, new_n23993, new_n23983);
xnor_3 g21646(new_n23995, new_n23990, new_n23986_1);
not_3  g21647(new_n23996, new_n23995);
xor_3  g21648(new_n23997, new_n23981, new_n11931);
nor_4  g21649(new_n23998, new_n23997, new_n23996);
not_3  g21650(new_n23999, new_n23998);
not_3  g21651(new_n24000, new_n23997);
nor_4  g21652(new_n24001, new_n24000, new_n23995);
nor_4  g21653(new_n24002_1, new_n24001, new_n23998);
nor_4  g21654(new_n24003, new_n23844, new_n18188);
not_3  g21655(new_n24004_1, new_n18188);
nor_4  g21656(new_n24005, new_n23845, new_n24004_1);
nor_4  g21657(new_n24006, new_n24005, new_n24003);
not_3  g21658(new_n24007, new_n24006);
nand_4 g21659(new_n24008, new_n18457, new_n18191);
nand_4 g21660(new_n24009, new_n18488, new_n18550);
nand_4 g21661(new_n24010, new_n24009, new_n24008);
nor_4  g21662(new_n24011, new_n24010, new_n24007);
nor_4  g21663(new_n24012, new_n24011, new_n24003);
nand_4 g21664(new_n24013, new_n24012, new_n24002_1);
nand_4 g21665(new_n24014, new_n24013, new_n23999);
not_3  g21666(new_n24015, new_n23983);
xnor_3 g21667(new_n24016, new_n23992, new_n24015);
not_3  g21668(new_n24017, new_n24016);
nand_4 g21669(new_n24018, new_n24017, new_n24014);
nand_4 g21670(new_n24019, new_n24018, new_n23994);
not_3  g21671(new_n24020, new_n24019);
nor_4  g21672(new_n24021, new_n15557, n1881);
xor_3  g21673(new_n24022, n8827, new_n21425);
not_3  g21674(new_n24023, new_n24022);
nor_4  g21675(new_n24024, new_n15538, n5834);
not_3  g21676(new_n24025, new_n24024);
nand_4 g21677(new_n24026, new_n23242, new_n23238_1);
nand_4 g21678(new_n24027, new_n24026, new_n24025);
not_3  g21679(new_n24028, new_n24027);
nor_4  g21680(new_n24029, new_n24028, new_n24023);
nor_4  g21681(new_n24030, new_n24029, new_n24021);
not_3  g21682(new_n24031, new_n24030);
nor_4  g21683(new_n24032_1, new_n24031, new_n24020);
nor_4  g21684(new_n24033, new_n24030, new_n24019);
nor_4  g21685(new_n24034, new_n24033, new_n24032_1);
xnor_3 g21686(new_n24035, new_n24017, new_n24014);
nor_4  g21687(new_n24036, new_n24035, new_n24030);
not_3  g21688(new_n24037, new_n24036);
xnor_3 g21689(new_n24038, new_n24016, new_n24014);
nor_4  g21690(new_n24039_1, new_n24038, new_n24031);
nor_4  g21691(new_n24040, new_n24039_1, new_n24036);
xor_3  g21692(new_n24041, new_n24028, new_n24023);
not_3  g21693(new_n24042, new_n24041);
xnor_3 g21694(new_n24043, new_n23997, new_n23996);
xnor_3 g21695(new_n24044, new_n24012, new_n24043);
nor_4  g21696(new_n24045, new_n24044, new_n24042);
xnor_3 g21697(new_n24046, new_n24010, new_n24006);
nor_4  g21698(new_n24047, new_n24046, new_n23243);
not_3  g21699(new_n24048_1, new_n24047);
not_3  g21700(new_n24049, new_n23243);
xnor_3 g21701(new_n24050, new_n24010, new_n24007);
nor_4  g21702(new_n24051, new_n24050, new_n24049);
nor_4  g21703(new_n24052_1, new_n24051, new_n24047);
nor_4  g21704(new_n24053, new_n23245, new_n18489);
nor_4  g21705(new_n24054, new_n18833, new_n18809);
nor_4  g21706(new_n24055, new_n24054, new_n24053);
nand_4 g21707(new_n24056, new_n24055, new_n24052_1);
nand_4 g21708(new_n24057, new_n24056, new_n24048_1);
xnor_3 g21709(new_n24058, new_n24044, new_n24042);
nor_4  g21710(new_n24059, new_n24058, new_n24057);
nor_4  g21711(new_n24060, new_n24059, new_n24045);
nand_4 g21712(new_n24061, new_n24060, new_n24040);
nand_4 g21713(new_n24062, new_n24061, new_n24037);
xnor_3 g21714(n6276, new_n24062, new_n24034);
not_3  g21715(new_n24064, new_n22902);
xor_3  g21716(n6308, new_n24064, new_n22901);
xnor_3 g21717(n6311, new_n20528, new_n20513);
xnor_3 g21718(n6323, new_n20237, new_n20219);
nor_4  g21719(new_n24068, new_n6925, new_n6876);
not_3  g21720(new_n24069, new_n24068);
nand_4 g21721(new_n24070, new_n7018, new_n24069);
not_3  g21722(new_n24071, new_n24070);
not_3  g21723(new_n24072, new_n16750);
nor_4  g21724(new_n24073, new_n16277, new_n24072);
not_3  g21725(new_n24074, new_n24073);
nor_4  g21726(new_n24075, new_n24074, new_n24071);
nor_4  g21727(new_n24076, new_n16278, new_n16750);
not_3  g21728(new_n24077, new_n24076);
nor_4  g21729(new_n24078, new_n24077, new_n24070);
nor_4  g21730(new_n24079, new_n24078, new_n24075);
nor_4  g21731(new_n24080, new_n24079, new_n21896);
xnor_3 g21732(new_n24081, new_n24079, new_n21896);
nand_4 g21733(new_n24082, new_n24077, new_n24074);
xnor_3 g21734(new_n24083, new_n24082, new_n24070);
not_3  g21735(new_n24084, new_n24083);
nor_4  g21736(new_n24085_1, new_n24084, new_n21902);
xnor_3 g21737(new_n24086, new_n24083, new_n21901);
nor_4  g21738(new_n24087, new_n7126, new_n7021);
nor_4  g21739(new_n24088, new_n7198, new_n7127);
nor_4  g21740(new_n24089, new_n24088, new_n24087);
nor_4  g21741(new_n24090, new_n24089, new_n24086);
nor_4  g21742(new_n24091, new_n24090, new_n24085_1);
nor_4  g21743(new_n24092_1, new_n24091, new_n24081);
nor_4  g21744(new_n24093_1, new_n24092_1, new_n24080);
nor_4  g21745(n6330, new_n24093_1, new_n24075);
xnor_3 g21746(n6339, new_n10222, new_n10177);
not_3  g21747(new_n24096_1, new_n17037_1);
xor_3  g21748(n6354, new_n24096_1, new_n17009);
not_3  g21749(new_n24098, n7335);
not_3  g21750(new_n24099, new_n3331);
nor_4  g21751(new_n24100, new_n24099, new_n24098);
not_3  g21752(new_n24101, new_n24100);
nor_4  g21753(new_n24102, new_n3331, n7335);
nor_4  g21754(new_n24103, new_n3465, n5696);
not_3  g21755(new_n24104, new_n24103);
xor_3  g21756(new_n24105_1, new_n3468_1, n5696);
not_3  g21757(new_n24106, new_n24105_1);
nor_4  g21758(new_n24107, new_n3470, n13367);
not_3  g21759(new_n24108, new_n24107);
xor_3  g21760(new_n24109, new_n3473, new_n3336);
nor_4  g21761(new_n24110, new_n3476, n932);
not_3  g21762(new_n24111, new_n24110);
not_3  g21763(new_n24112, new_n3476);
xor_3  g21764(new_n24113, new_n24112, new_n6117);
nor_4  g21765(new_n24114, new_n3484, n6691);
not_3  g21766(new_n24115, new_n24114);
xor_3  g21767(new_n24116, new_n3484, n6691);
nor_4  g21768(new_n24117, new_n3489, n3260);
not_3  g21769(new_n24118, new_n24117);
xor_3  g21770(new_n24119_1, new_n3489, n3260);
nor_4  g21771(new_n24120, new_n3493, n20489);
not_3  g21772(new_n24121, new_n24120);
not_3  g21773(new_n24122, n2355);
not_3  g21774(new_n24123, new_n3498);
nand_4 g21775(new_n24124, new_n24123, new_n24122);
xor_3  g21776(new_n24125, new_n24123, new_n24122);
nor_4  g21777(new_n24126, new_n3518, n11121);
not_3  g21778(new_n24127, new_n24126);
nand_4 g21779(new_n24128, n16217, n12315);
xor_3  g21780(new_n24129_1, new_n3518, n11121);
nand_4 g21781(new_n24130, new_n24129_1, new_n24128);
nand_4 g21782(new_n24131, new_n24130, new_n24127);
nand_4 g21783(new_n24132, new_n24131, new_n24125);
nand_4 g21784(new_n24133_1, new_n24132, new_n24124);
not_3  g21785(new_n24134, n20489);
xor_3  g21786(new_n24135, new_n3496, new_n24134);
nand_4 g21787(new_n24136, new_n24135, new_n24133_1);
nand_4 g21788(new_n24137, new_n24136, new_n24121);
nand_4 g21789(new_n24138, new_n24137, new_n24119_1);
nand_4 g21790(new_n24139, new_n24138, new_n24118);
nand_4 g21791(new_n24140, new_n24139, new_n24116);
nand_4 g21792(new_n24141_1, new_n24140, new_n24115);
nand_4 g21793(new_n24142, new_n24141_1, new_n24113);
nand_4 g21794(new_n24143, new_n24142, new_n24111);
nand_4 g21795(new_n24144, new_n24143, new_n24109);
nand_4 g21796(new_n24145_1, new_n24144, new_n24108);
nand_4 g21797(new_n24146_1, new_n24145_1, new_n24106);
nand_4 g21798(new_n24147, new_n24146_1, new_n24104);
nor_4  g21799(new_n24148, new_n24147, new_n24102);
nor_4  g21800(new_n24149, new_n24148, new_n3329);
nand_4 g21801(new_n24150_1, new_n24149, new_n24101);
not_3  g21802(new_n24151, new_n24150_1);
nand_4 g21803(new_n24152, new_n24151, new_n20761_1);
nor_4  g21804(new_n24153, new_n24151, new_n20809);
not_3  g21805(new_n24154, new_n24153);
nor_4  g21806(new_n24155_1, new_n24150_1, new_n20812);
nor_4  g21807(new_n24156, new_n24155_1, new_n24153);
nor_4  g21808(new_n24157, new_n24102, new_n24100);
xnor_3 g21809(new_n24158, new_n24157, new_n24147);
nor_4  g21810(new_n24159, new_n24158, new_n20820);
not_3  g21811(new_n24160_1, new_n24159);
not_3  g21812(new_n24161, new_n24158);
nor_4  g21813(new_n24162, new_n24161, new_n20816);
nor_4  g21814(new_n24163, new_n24162, new_n24159);
xnor_3 g21815(new_n24164, new_n24145_1, new_n24105_1);
nand_4 g21816(new_n24165, new_n24164, new_n20826_1);
xnor_3 g21817(new_n24166, new_n24164, new_n20825);
not_3  g21818(new_n24167_1, new_n24109);
xnor_3 g21819(new_n24168, new_n24143, new_n24167_1);
nand_4 g21820(new_n24169, new_n24168, new_n20833);
xnor_3 g21821(new_n24170_1, new_n24168, new_n20832);
not_3  g21822(new_n24171, new_n24113);
xnor_3 g21823(new_n24172_1, new_n24141_1, new_n24171);
nand_4 g21824(new_n24173, new_n24172_1, new_n20838);
xnor_3 g21825(new_n24174, new_n24172_1, new_n20837);
not_3  g21826(new_n24175, new_n24116);
xnor_3 g21827(new_n24176, new_n24139, new_n24175);
nand_4 g21828(new_n24177_1, new_n24176, new_n20843);
xnor_3 g21829(new_n24178, new_n24176, new_n20842);
not_3  g21830(new_n24179, new_n24138);
nor_4  g21831(new_n24180, new_n24137, new_n24119_1);
nor_4  g21832(new_n24181, new_n24180, new_n24179);
nand_4 g21833(new_n24182, new_n24181, new_n20849);
xnor_3 g21834(new_n24183, new_n24181, new_n20848);
xnor_3 g21835(new_n24184, new_n24135, new_n24133_1);
not_3  g21836(new_n24185, new_n24184);
nand_4 g21837(new_n24186, new_n24185, new_n20852);
xnor_3 g21838(new_n24187, new_n24184, new_n20852);
not_3  g21839(new_n24188, new_n24131);
xnor_3 g21840(new_n24189, new_n24188, new_n24125);
nor_4  g21841(new_n24190, new_n24189, new_n20862);
xnor_3 g21842(new_n24191, new_n24189, new_n20862);
nor_4  g21843(new_n24192, new_n24129_1, new_n20865);
not_3  g21844(new_n24193, new_n24192);
not_3  g21845(new_n24194, new_n24129_1);
xor_3  g21846(new_n24195, new_n24194, new_n24128);
nand_4 g21847(new_n24196_1, new_n24195, new_n20865);
xor_3  g21848(new_n24197, n16217, n12315);
nand_4 g21849(new_n24198, new_n24197, new_n20872);
nand_4 g21850(new_n24199, new_n24198, new_n24196_1);
nand_4 g21851(new_n24200, new_n24199, new_n24193);
nor_4  g21852(new_n24201, new_n24200, new_n24191);
nor_4  g21853(new_n24202, new_n24201, new_n24190);
nand_4 g21854(new_n24203, new_n24202, new_n24187);
nand_4 g21855(new_n24204, new_n24203, new_n24186);
nand_4 g21856(new_n24205, new_n24204, new_n24183);
nand_4 g21857(new_n24206, new_n24205, new_n24182);
nand_4 g21858(new_n24207, new_n24206, new_n24178);
nand_4 g21859(new_n24208, new_n24207, new_n24177_1);
nand_4 g21860(new_n24209, new_n24208, new_n24174);
nand_4 g21861(new_n24210, new_n24209, new_n24173);
nand_4 g21862(new_n24211, new_n24210, new_n24170_1);
nand_4 g21863(new_n24212, new_n24211, new_n24169);
nand_4 g21864(new_n24213, new_n24212, new_n24166);
nand_4 g21865(new_n24214, new_n24213, new_n24165);
nand_4 g21866(new_n24215, new_n24214, new_n24163);
nand_4 g21867(new_n24216, new_n24215, new_n24160_1);
nand_4 g21868(new_n24217, new_n24216, new_n24156);
nand_4 g21869(new_n24218, new_n24217, new_n24154);
nand_4 g21870(new_n24219, new_n24218, new_n24152);
nand_4 g21871(new_n24220, new_n24150_1, new_n20760);
nand_4 g21872(new_n24221, new_n24220, new_n24217);
nand_4 g21873(new_n24222, new_n24221, new_n24219);
not_3  g21874(n6375, new_n24222);
not_3  g21875(new_n24224, new_n23079);
xor_3  g21876(n6383, new_n23094, new_n24224);
not_3  g21877(new_n24226, new_n17558);
xor_3  g21878(n6407, new_n24226, new_n17506);
not_3  g21879(new_n24228_1, new_n10211);
xor_3  g21880(n6431, new_n10214, new_n24228_1);
xnor_3 g21881(n6437, new_n20038, new_n20035);
not_3  g21882(new_n24231, new_n4661);
xor_3  g21883(n6457, new_n4664, new_n24231);
xnor_3 g21884(n6465, new_n14804, new_n14767);
not_3  g21885(new_n24234, new_n21153);
nor_4  g21886(new_n24235, new_n21149, n3582);
nor_4  g21887(new_n24236, new_n21157_1, new_n21154_1);
nor_4  g21888(new_n24237, new_n24236, new_n24235);
nand_4 g21889(new_n24238, new_n24237, new_n24234);
not_3  g21890(new_n24239, new_n24238);
nor_4  g21891(new_n24240, new_n24239, new_n9924);
not_3  g21892(new_n24241, new_n9924);
nor_4  g21893(new_n24242, new_n24238, new_n24241);
nor_4  g21894(new_n24243, new_n24242, new_n24240);
nor_4  g21895(new_n24244, new_n21159, new_n3742);
not_3  g21896(new_n24245, new_n24244);
nor_4  g21897(new_n24246, new_n17443, new_n17386);
nor_4  g21898(new_n24247, new_n24246, new_n17384);
nor_4  g21899(new_n24248, new_n21158, new_n3744);
nor_4  g21900(new_n24249, new_n24248, new_n24244);
nand_4 g21901(new_n24250, new_n24249, new_n24247);
nand_4 g21902(new_n24251, new_n24250, new_n24245);
xnor_3 g21903(new_n24252, new_n24251, new_n24243);
not_3  g21904(new_n24253, new_n3894);
nor_4  g21905(new_n24254, new_n24253, new_n3825);
nor_4  g21906(new_n24255, new_n3893, n9259);
not_3  g21907(new_n24256, new_n24255);
nand_4 g21908(new_n24257, new_n24253, new_n3825);
nand_4 g21909(new_n24258_1, new_n17481, new_n17446);
nand_4 g21910(new_n24259, new_n24258_1, new_n17445);
nand_4 g21911(new_n24260_1, new_n24259, new_n24257);
nand_4 g21912(new_n24261, new_n24260_1, new_n24256);
nor_4  g21913(new_n24262, new_n24261, new_n24254);
not_3  g21914(new_n24263, new_n24262);
nor_4  g21915(new_n24264, new_n24263, new_n24252);
nand_4 g21916(new_n24265, new_n24263, new_n24252);
not_3  g21917(new_n24266, new_n24265);
nor_4  g21918(new_n24267, new_n24266, new_n24264);
not_3  g21919(new_n24268, new_n24250);
nor_4  g21920(new_n24269, new_n24249, new_n24247);
nor_4  g21921(new_n24270, new_n24269, new_n24268);
xor_3  g21922(new_n24271, new_n24253, new_n3825);
not_3  g21923(new_n24272, new_n24271);
xnor_3 g21924(new_n24273, new_n24272, new_n24259);
nor_4  g21925(new_n24274, new_n24273, new_n24270);
xnor_3 g21926(new_n24275, new_n24249, new_n24247);
not_3  g21927(new_n24276, new_n24273);
xnor_3 g21928(new_n24277, new_n24276, new_n24275);
nor_4  g21929(new_n24278_1, new_n17482, new_n17444);
nor_4  g21930(new_n24279, new_n17562, new_n17483);
nor_4  g21931(new_n24280, new_n24279, new_n24278_1);
nor_4  g21932(new_n24281, new_n24280, new_n24277);
nor_4  g21933(new_n24282, new_n24281, new_n24274);
not_3  g21934(new_n24283, new_n24282);
xnor_3 g21935(n6470, new_n24283, new_n24267);
xnor_3 g21936(n6476, new_n13891, new_n13864);
not_3  g21937(new_n24286, new_n22507);
xor_3  g21938(n6506, new_n24286, new_n22496);
not_3  g21939(new_n24288, new_n11228);
nor_4  g21940(new_n24289_1, new_n24288, new_n11226);
not_3  g21941(new_n24290, new_n24289_1);
nor_4  g21942(new_n24291, new_n24290, new_n17139);
nand_4 g21943(new_n24292, new_n24291, new_n11214);
not_3  g21944(new_n24293, new_n24292);
nand_4 g21945(new_n24294, new_n24293, new_n11209);
nor_4  g21946(new_n24295, new_n24294, new_n11202);
not_3  g21947(new_n24296, new_n24295);
nor_4  g21948(new_n24297_1, new_n24296, new_n11197);
not_3  g21949(new_n24298, new_n24297_1);
nor_4  g21950(new_n24299, new_n24298, new_n17113);
not_3  g21951(new_n24300, new_n24299);
nor_4  g21952(new_n24301, new_n24300, new_n17107);
nor_4  g21953(new_n24302, new_n24299, new_n17108);
nor_4  g21954(new_n24303, new_n24302, new_n24301);
xnor_3 g21955(new_n24304, new_n24303, new_n12172);
xnor_3 g21956(new_n24305, new_n24297_1, new_n17112);
nand_4 g21957(new_n24306, new_n24305, new_n12179_1);
xnor_3 g21958(new_n24307_1, new_n24305, new_n12176);
xnor_3 g21959(new_n24308, new_n24296, new_n11197);
nand_4 g21960(new_n24309, new_n24308, new_n12218);
xnor_3 g21961(new_n24310, new_n24308, new_n11112);
xnor_3 g21962(new_n24311, new_n24294, new_n11202);
nand_4 g21963(new_n24312, new_n24311, new_n11115);
xnor_3 g21964(new_n24313, new_n24311, new_n11117);
xnor_3 g21965(new_n24314, new_n24292, new_n11208);
nand_4 g21966(new_n24315, new_n24314, new_n11130);
xnor_3 g21967(new_n24316, new_n24314, new_n11131);
xnor_3 g21968(new_n24317, new_n24291, new_n11214);
nand_4 g21969(new_n24318, new_n24317, new_n11136);
xnor_3 g21970(new_n24319_1, new_n24289_1, new_n11220_1);
nand_4 g21971(new_n24320, new_n24319_1, new_n11142);
not_3  g21972(new_n24321, new_n24320);
xnor_3 g21973(new_n24322, new_n24319_1, new_n11142);
nor_4  g21974(new_n24323_1, new_n11228, new_n11150);
nor_4  g21975(new_n24324, new_n24323_1, new_n11153);
nor_4  g21976(new_n24325, new_n11228, new_n11185);
nor_4  g21977(new_n24326, new_n24325, new_n24289_1);
not_3  g21978(new_n24327_1, new_n24323_1);
nor_4  g21979(new_n24328, new_n24327_1, new_n11123);
nor_4  g21980(new_n24329, new_n24328, new_n24324);
not_3  g21981(new_n24330, new_n24329);
nor_4  g21982(new_n24331, new_n24330, new_n24326);
nor_4  g21983(new_n24332, new_n24331, new_n24324);
nor_4  g21984(new_n24333, new_n24332, new_n24322);
nor_4  g21985(new_n24334, new_n24333, new_n24321);
not_3  g21986(new_n24335, new_n24334);
xnor_3 g21987(new_n24336, new_n24317, new_n11137);
nand_4 g21988(new_n24337, new_n24336, new_n24335);
nand_4 g21989(new_n24338, new_n24337, new_n24318);
nand_4 g21990(new_n24339, new_n24338, new_n24316);
nand_4 g21991(new_n24340, new_n24339, new_n24315);
nand_4 g21992(new_n24341, new_n24340, new_n24313);
nand_4 g21993(new_n24342_1, new_n24341, new_n24312);
nand_4 g21994(new_n24343, new_n24342_1, new_n24310);
nand_4 g21995(new_n24344, new_n24343, new_n24309);
nand_4 g21996(new_n24345_1, new_n24344, new_n24307_1);
nand_4 g21997(new_n24346, new_n24345_1, new_n24306);
xnor_3 g21998(new_n24347_1, new_n24346, new_n24304);
xnor_3 g21999(new_n24348, new_n24347_1, new_n20314);
not_3  g22000(new_n24349, new_n24344);
xnor_3 g22001(new_n24350, new_n24349, new_n24307_1);
nand_4 g22002(new_n24351, new_n24350, new_n20317);
not_3  g22003(new_n24352, new_n20317);
xnor_3 g22004(new_n24353, new_n24350, new_n24352);
xnor_3 g22005(new_n24354, new_n24342_1, new_n24310);
not_3  g22006(new_n24355, new_n24354);
nand_4 g22007(new_n24356, new_n24355, new_n20321);
xnor_3 g22008(new_n24357, new_n24354, new_n20321);
xnor_3 g22009(new_n24358, new_n24311, new_n11115);
xnor_3 g22010(new_n24359, new_n24340, new_n24358);
nand_4 g22011(new_n24360, new_n24359, new_n20325);
not_3  g22012(new_n24361, new_n24360);
nor_4  g22013(new_n24362, new_n24359, new_n20325);
nor_4  g22014(new_n24363, new_n24362, new_n24361);
not_3  g22015(new_n24364, new_n24316);
xnor_3 g22016(new_n24365, new_n24338, new_n24364);
nor_4  g22017(new_n24366, new_n24365, new_n20329);
xnor_3 g22018(new_n24367, new_n24336, new_n24335);
not_3  g22019(new_n24368, new_n24367);
nor_4  g22020(new_n24369, new_n24368, new_n20335);
xnor_3 g22021(new_n24370, new_n24367, new_n20334);
xnor_3 g22022(new_n24371, new_n24332, new_n24322);
not_3  g22023(new_n24372, new_n24371);
nor_4  g22024(new_n24373_1, new_n24372, new_n20341);
xnor_3 g22025(new_n24374_1, new_n24371, new_n20340);
not_3  g22026(new_n24375, new_n24326);
nor_4  g22027(new_n24376, new_n24329, new_n24375);
nor_4  g22028(new_n24377, new_n24376, new_n24331);
nor_4  g22029(new_n24378, new_n24377, new_n20347);
xor_3  g22030(new_n24379, new_n11228, new_n11150);
not_3  g22031(new_n24380, new_n24379);
nor_4  g22032(new_n24381, new_n24380, new_n20351);
not_3  g22033(new_n24382, new_n24381);
xnor_3 g22034(new_n24383, new_n24377, new_n20347);
nor_4  g22035(new_n24384, new_n24383, new_n24382);
nor_4  g22036(new_n24385, new_n24384, new_n24378);
nor_4  g22037(new_n24386, new_n24385, new_n24374_1);
nor_4  g22038(new_n24387, new_n24386, new_n24373_1);
nor_4  g22039(new_n24388, new_n24387, new_n24370);
nor_4  g22040(new_n24389, new_n24388, new_n24369);
xnor_3 g22041(new_n24390, new_n24365, new_n20329);
nor_4  g22042(new_n24391, new_n24390, new_n24389);
nor_4  g22043(new_n24392, new_n24391, new_n24366);
nand_4 g22044(new_n24393, new_n24392, new_n24363);
nand_4 g22045(new_n24394, new_n24393, new_n24360);
nand_4 g22046(new_n24395, new_n24394, new_n24357);
nand_4 g22047(new_n24396, new_n24395, new_n24356);
nand_4 g22048(new_n24397, new_n24396, new_n24353);
nand_4 g22049(new_n24398, new_n24397, new_n24351);
xor_3  g22050(n6514, new_n24398, new_n24348);
nand_4 g22051(new_n24400, new_n13849, new_n13734);
nand_4 g22052(new_n24401, new_n13895, new_n13850_1);
nand_4 g22053(new_n24402, new_n24401, new_n24400);
xor_3  g22054(new_n24403, new_n13787, new_n13773);
nor_4  g22055(new_n24404, new_n24403, new_n13847);
xor_3  g22056(new_n24405, new_n13788, new_n13773);
nor_4  g22057(new_n24406_1, new_n13848, new_n13791);
not_3  g22058(new_n24407, new_n24406_1);
nor_4  g22059(new_n24408, new_n24407, new_n24405);
nor_4  g22060(new_n24409, new_n24408, new_n24404);
xnor_3 g22061(n6542, new_n24409, new_n24402);
not_3  g22062(new_n24411, new_n18676);
xor_3  g22063(n6558, new_n18690_1, new_n24411);
not_3  g22064(new_n24413, new_n21881);
xor_3  g22065(n6560, new_n24413, new_n21878);
nand_4 g22066(new_n24415_1, new_n7343, n10405);
not_3  g22067(new_n24416, new_n24415_1);
nor_4  g22068(new_n24417, new_n7343, n10405);
nor_4  g22069(new_n24418, new_n24417, new_n24416);
nor_4  g22070(new_n24419, new_n7346_1, new_n6346);
not_3  g22071(new_n24420, new_n24419);
xor_3  g22072(new_n24421_1, new_n7346_1, new_n6346);
nor_4  g22073(new_n24422, new_n7357, n17090);
nor_4  g22074(new_n24423, new_n7355, new_n6353);
xor_3  g22075(new_n24424, new_n7357, new_n4477);
nor_4  g22076(new_n24425, new_n24424, new_n24423);
nor_4  g22077(new_n24426, new_n24425, new_n24422);
nand_4 g22078(new_n24427, new_n24426, new_n24421_1);
nand_4 g22079(new_n24428, new_n24427, new_n24420);
xnor_3 g22080(new_n24429, new_n24428, new_n24418);
xnor_3 g22081(new_n24430, new_n24429, new_n11678);
not_3  g22082(new_n24431_1, new_n24430);
xnor_3 g22083(new_n24432, new_n24426, new_n24421_1);
nand_4 g22084(new_n24433, new_n24432, new_n11681);
not_3  g22085(new_n24434, new_n24433);
nor_4  g22086(new_n24435, new_n24432, new_n11681);
nor_4  g22087(new_n24436, new_n24435, new_n24434);
not_3  g22088(new_n24437, new_n24423);
not_3  g22089(new_n24438, new_n24424);
nor_4  g22090(new_n24439, new_n24438, new_n24437);
nor_4  g22091(new_n24440, new_n24439, new_n24425);
nand_4 g22092(new_n24441, new_n24440, new_n11688);
nor_4  g22093(new_n24442, new_n21913, new_n11691);
not_3  g22094(new_n24443, new_n24441);
nor_4  g22095(new_n24444, new_n24440, new_n11688);
nor_4  g22096(new_n24445, new_n24444, new_n24443);
nand_4 g22097(new_n24446, new_n24445, new_n24442);
nand_4 g22098(new_n24447, new_n24446, new_n24441);
nand_4 g22099(new_n24448, new_n24447, new_n24436);
nand_4 g22100(new_n24449, new_n24448, new_n24433);
xor_3  g22101(n6567, new_n24449, new_n24431_1);
not_3  g22102(new_n24451, new_n16547);
nor_4  g22103(new_n24452, new_n24451, n8324);
not_3  g22104(new_n24453, new_n24452);
nor_4  g22105(new_n24454, new_n24453, n1279);
not_3  g22106(new_n24455, new_n24454);
nor_4  g22107(new_n24456, new_n24455, n9445);
not_3  g22108(new_n24457, new_n24456);
nor_4  g22109(new_n24458, new_n24457, n19454);
xor_3  g22110(new_n24459, new_n24458, new_n9573);
not_3  g22111(new_n24460, new_n24459);
nor_4  g22112(new_n24461, new_n24460, new_n5038);
nor_4  g22113(new_n24462, new_n24459, new_n5043);
nor_4  g22114(new_n24463, new_n24462, new_n24461);
xor_3  g22115(new_n24464, new_n24456, new_n9578);
nor_4  g22116(new_n24465, new_n24464, new_n5048);
xnor_3 g22117(new_n24466, new_n24464, new_n5048);
xor_3  g22118(new_n24467, new_n24454, new_n9583);
nor_4  g22119(new_n24468, new_n24467, new_n5057);
xnor_3 g22120(new_n24469, new_n24467, new_n5057);
xor_3  g22121(new_n24470, new_n24452, n1279);
nand_4 g22122(new_n24471, new_n24470, new_n5067);
xnor_3 g22123(new_n24472_1, new_n24470, new_n5062_1);
not_3  g22124(new_n24473, new_n16551);
nand_4 g22125(new_n24474, new_n16584_1, new_n16552);
nand_4 g22126(new_n24475, new_n24474, new_n24473);
nand_4 g22127(new_n24476_1, new_n24475, new_n24472_1);
nand_4 g22128(new_n24477, new_n24476_1, new_n24471);
not_3  g22129(new_n24478, new_n24477);
nor_4  g22130(new_n24479, new_n24478, new_n24469);
nor_4  g22131(new_n24480, new_n24479, new_n24468);
nor_4  g22132(new_n24481, new_n24480, new_n24466);
nor_4  g22133(new_n24482, new_n24481, new_n24465);
nand_4 g22134(new_n24483_1, new_n24482, new_n24463);
not_3  g22135(new_n24484, new_n24483_1);
nor_4  g22136(new_n24485_1, new_n24482, new_n24463);
nor_4  g22137(new_n24486, new_n24485_1, new_n24484);
xnor_3 g22138(new_n24487, new_n9574, n23272);
nand_4 g22139(new_n24488, new_n9579, new_n22700);
xor_3  g22140(new_n24489, new_n9581, n11481);
nand_4 g22141(new_n24490, new_n9584, new_n22702);
xor_3  g22142(new_n24491, new_n9586, n16439);
nand_4 g22143(new_n24492, new_n9589, new_n4922);
nor_4  g22144(new_n24493, new_n9593, new_n12765);
nor_4  g22145(new_n24494, new_n16607, new_n16586);
nor_4  g22146(new_n24495, new_n24494, new_n24493);
xnor_3 g22147(new_n24496, new_n9589, n15241);
nand_4 g22148(new_n24497, new_n24496, new_n24495);
nand_4 g22149(new_n24498, new_n24497, new_n24492);
nand_4 g22150(new_n24499, new_n24498, new_n24491);
nand_4 g22151(new_n24500, new_n24499, new_n24490);
nand_4 g22152(new_n24501_1, new_n24500, new_n24489);
nand_4 g22153(new_n24502, new_n24501_1, new_n24488);
nor_4  g22154(new_n24503, new_n24502, new_n24487);
not_3  g22155(new_n24504, new_n24487);
not_3  g22156(new_n24505, new_n24502);
nor_4  g22157(new_n24506, new_n24505, new_n24504);
nor_4  g22158(new_n24507, new_n24506, new_n24503);
xnor_3 g22159(new_n24508, new_n24507, new_n24486);
xnor_3 g22160(new_n24509, new_n24480, new_n24466);
xnor_3 g22161(new_n24510, new_n24500, new_n24489);
nor_4  g22162(new_n24511, new_n24510, new_n24509);
xnor_3 g22163(new_n24512_1, new_n24510, new_n24509);
not_3  g22164(new_n24513, new_n24469);
nor_4  g22165(new_n24514, new_n24477, new_n24513);
nor_4  g22166(new_n24515, new_n24514, new_n24479);
not_3  g22167(new_n24516, new_n24515);
xnor_3 g22168(new_n24517, new_n24498, new_n24491);
nor_4  g22169(new_n24518, new_n24517, new_n24516);
xnor_3 g22170(new_n24519, new_n24517, new_n24515);
xnor_3 g22171(new_n24520, new_n24475, new_n24472_1);
not_3  g22172(new_n24521, new_n24520);
not_3  g22173(new_n24522, new_n24496);
xnor_3 g22174(new_n24523, new_n24522, new_n24495);
nand_4 g22175(new_n24524, new_n24523, new_n24521);
xnor_3 g22176(new_n24525, new_n24523, new_n24520);
not_3  g22177(new_n24526, new_n16585);
nand_4 g22178(new_n24527, new_n16608_1, new_n24526);
nand_4 g22179(new_n24528, new_n16655, new_n16609);
nand_4 g22180(new_n24529, new_n24528, new_n24527);
nand_4 g22181(new_n24530, new_n24529, new_n24525);
nand_4 g22182(new_n24531, new_n24530, new_n24524);
nand_4 g22183(new_n24532, new_n24531, new_n24519);
not_3  g22184(new_n24533, new_n24532);
nor_4  g22185(new_n24534, new_n24533, new_n24518);
nor_4  g22186(new_n24535, new_n24534, new_n24512_1);
nor_4  g22187(new_n24536, new_n24535, new_n24511);
xnor_3 g22188(n6576, new_n24536, new_n24508);
not_3  g22189(new_n24538, new_n20865);
xor_3  g22190(new_n24539, new_n24195, new_n24538);
xor_3  g22191(n6587, new_n24539, new_n24198);
xnor_3 g22192(n6612, new_n22914_1, new_n22854);
nor_4  g22193(new_n24542, new_n21221, new_n12952);
xnor_3 g22194(new_n24543, new_n21222_1, new_n12951);
nor_4  g22195(new_n24544, new_n21226_1, new_n12942_1);
xnor_3 g22196(new_n24545, new_n21226_1, new_n12942_1);
nor_4  g22197(new_n24546, new_n21232, new_n12935);
xnor_3 g22198(new_n24547, new_n21233, new_n12935);
nand_4 g22199(new_n24548, new_n21237, new_n12924);
nor_4  g22200(new_n24549, new_n21236, new_n12925);
nor_4  g22201(new_n24550, new_n21237, new_n12924);
nor_4  g22202(new_n24551, new_n24550, new_n24549);
nand_4 g22203(new_n24552, new_n21242, new_n12918);
nor_4  g22204(new_n24553, new_n21241, new_n12917_1);
nor_4  g22205(new_n24554, new_n21242, new_n12918);
nor_4  g22206(new_n24555, new_n24554, new_n24553);
nand_4 g22207(new_n24556, new_n21247, new_n19928);
nor_4  g22208(new_n24557, new_n21244, new_n12908);
nor_4  g22209(new_n24558_1, new_n21247, new_n19928);
nor_4  g22210(new_n24559, new_n24558_1, new_n24557);
nor_4  g22211(new_n24560, new_n18308, new_n12898);
not_3  g22212(new_n24561, new_n24560);
xnor_3 g22213(new_n24562, new_n18308, new_n12898);
not_3  g22214(new_n24563, new_n24562);
nor_4  g22215(new_n24564, new_n18313, new_n12888);
nor_4  g22216(new_n24565, new_n12979, n18);
not_3  g22217(new_n24566, new_n24565);
nor_4  g22218(new_n24567, new_n24566, n15490);
nor_4  g22219(new_n24568, new_n24565, new_n18316);
nor_4  g22220(new_n24569, new_n24568, new_n24567);
not_3  g22221(new_n24570, new_n24569);
nor_4  g22222(new_n24571, new_n24570, new_n12877);
nor_4  g22223(new_n24572, new_n24571, new_n24567);
not_3  g22224(new_n24573, new_n24572);
xnor_3 g22225(new_n24574, new_n18313, new_n12888);
nor_4  g22226(new_n24575, new_n24574, new_n24573);
nor_4  g22227(new_n24576_1, new_n24575, new_n24564);
nand_4 g22228(new_n24577, new_n24576_1, new_n24563);
nand_4 g22229(new_n24578, new_n24577, new_n24561);
nand_4 g22230(new_n24579_1, new_n24578, new_n24559);
nand_4 g22231(new_n24580, new_n24579_1, new_n24556);
nand_4 g22232(new_n24581, new_n24580, new_n24555);
nand_4 g22233(new_n24582, new_n24581, new_n24552);
nand_4 g22234(new_n24583, new_n24582, new_n24551);
nand_4 g22235(new_n24584, new_n24583, new_n24548);
nand_4 g22236(new_n24585, new_n24584, new_n24547);
not_3  g22237(new_n24586, new_n24585);
nor_4  g22238(new_n24587, new_n24586, new_n24546);
nor_4  g22239(new_n24588, new_n24587, new_n24545);
nor_4  g22240(new_n24589, new_n24588, new_n24544);
nor_4  g22241(new_n24590, new_n24589, new_n24543);
nor_4  g22242(new_n24591, new_n24590, new_n24542);
not_3  g22243(new_n24592, new_n21220);
nor_4  g22244(new_n24593, new_n24592, n23166);
not_3  g22245(new_n24594, new_n24593);
nor_4  g22246(new_n24595, new_n21449, new_n24594);
and_4  g22247(new_n24596, new_n24595, new_n24591);
nor_4  g22248(new_n24597, new_n21450, new_n24593);
not_3  g22249(new_n24598, new_n24597);
nor_4  g22250(new_n24599, new_n24598, new_n24591);
nor_4  g22251(new_n24600, new_n24599, new_n24596);
not_3  g22252(new_n24601, new_n23695);
nor_4  g22253(new_n24602_1, new_n24597, new_n24595);
not_3  g22254(new_n24603, new_n24602_1);
xnor_3 g22255(new_n24604_1, new_n24603, new_n24591);
nand_4 g22256(new_n24605, new_n24604_1, new_n23698);
not_3  g22257(new_n24606, new_n24605);
xnor_3 g22258(new_n24607, new_n24604_1, new_n23698);
xnor_3 g22259(new_n24608, new_n24589, new_n24543);
nor_4  g22260(new_n24609, new_n24608, new_n23703);
xnor_3 g22261(new_n24610, new_n24608, new_n23703);
xnor_3 g22262(new_n24611, new_n24587, new_n24545);
nor_4  g22263(new_n24612, new_n24611, new_n23708);
xnor_3 g22264(new_n24613, new_n24611, new_n23708);
xnor_3 g22265(new_n24614, new_n24584, new_n24547);
not_3  g22266(new_n24615, new_n24614);
nand_4 g22267(new_n24616, new_n24615, new_n23716);
xnor_3 g22268(new_n24617, new_n24614, new_n23716);
xnor_3 g22269(new_n24618_1, new_n24582, new_n24551);
not_3  g22270(new_n24619, new_n24618_1);
nand_4 g22271(new_n24620_1, new_n24619, new_n11242);
xnor_3 g22272(new_n24621, new_n24618_1, new_n11242);
xnor_3 g22273(new_n24622, new_n24580, new_n24555);
not_3  g22274(new_n24623, new_n24622);
nand_4 g22275(new_n24624, new_n24623, new_n11247);
xnor_3 g22276(new_n24625, new_n24622, new_n11247);
not_3  g22277(new_n24626_1, new_n24559);
xnor_3 g22278(new_n24627, new_n24578, new_n24626_1);
nand_4 g22279(new_n24628, new_n24627, new_n11253);
xnor_3 g22280(new_n24629_1, new_n24627, new_n11254);
not_3  g22281(new_n24630, new_n11261_1);
xnor_3 g22282(new_n24631, new_n24576_1, new_n24562);
nand_4 g22283(new_n24632, new_n24631, new_n24630);
not_3  g22284(new_n24633, new_n24632);
nor_4  g22285(new_n24634, new_n24631, new_n24630);
nor_4  g22286(new_n24635, new_n24634, new_n24633);
xnor_3 g22287(new_n24636_1, new_n24574, new_n24572);
not_3  g22288(new_n24637, new_n24636_1);
nand_4 g22289(new_n24638_1, new_n24637, new_n11268);
not_3  g22290(new_n24639, new_n24638_1);
nor_4  g22291(new_n24640, new_n24637, new_n11268);
nor_4  g22292(new_n24641, new_n24640, new_n24639);
nor_4  g22293(new_n24642, new_n24569, new_n12878);
nor_4  g22294(new_n24643, new_n24642, new_n24571);
not_3  g22295(new_n24644, new_n24643);
nor_4  g22296(new_n24645, new_n24644, new_n11274);
not_3  g22297(new_n24646, new_n24645);
xor_3  g22298(new_n24647, new_n12875_1, new_n10912);
not_3  g22299(new_n24648, new_n24647);
nand_4 g22300(new_n24649, new_n24648, new_n11277);
not_3  g22301(new_n24650, new_n11274);
nor_4  g22302(new_n24651, new_n24643, new_n24650);
nor_4  g22303(new_n24652, new_n24651, new_n24645);
nand_4 g22304(new_n24653, new_n24652, new_n24649);
nand_4 g22305(new_n24654, new_n24653, new_n24646);
nand_4 g22306(new_n24655, new_n24654, new_n24641);
nand_4 g22307(new_n24656, new_n24655, new_n24638_1);
nand_4 g22308(new_n24657, new_n24656, new_n24635);
nand_4 g22309(new_n24658, new_n24657, new_n24632);
nand_4 g22310(new_n24659, new_n24658, new_n24629_1);
nand_4 g22311(new_n24660, new_n24659, new_n24628);
nand_4 g22312(new_n24661, new_n24660, new_n24625);
nand_4 g22313(new_n24662, new_n24661, new_n24624);
nand_4 g22314(new_n24663, new_n24662, new_n24621);
nand_4 g22315(new_n24664, new_n24663, new_n24620_1);
nand_4 g22316(new_n24665, new_n24664, new_n24617);
nand_4 g22317(new_n24666, new_n24665, new_n24616);
not_3  g22318(new_n24667, new_n24666);
nor_4  g22319(new_n24668, new_n24667, new_n24613);
nor_4  g22320(new_n24669, new_n24668, new_n24612);
nor_4  g22321(new_n24670, new_n24669, new_n24610);
nor_4  g22322(new_n24671, new_n24670, new_n24609);
nor_4  g22323(new_n24672, new_n24671, new_n24607);
nor_4  g22324(new_n24673, new_n24672, new_n24606);
nand_4 g22325(new_n24674, new_n24673, new_n24601);
not_3  g22326(new_n24675, new_n24607);
not_3  g22327(new_n24676, new_n24609);
xnor_3 g22328(new_n24677, new_n24608, new_n23705);
not_3  g22329(new_n24678, new_n24612);
not_3  g22330(new_n24679, new_n24613);
nand_4 g22331(new_n24680, new_n24666, new_n24679);
nand_4 g22332(new_n24681, new_n24680, new_n24678);
nand_4 g22333(new_n24682, new_n24681, new_n24677);
nand_4 g22334(new_n24683, new_n24682, new_n24676);
nand_4 g22335(new_n24684, new_n24683, new_n24675);
nand_4 g22336(new_n24685, new_n24684, new_n24605);
nand_4 g22337(new_n24686, new_n24685, new_n23695);
nand_4 g22338(new_n24687, new_n24686, new_n24674);
xnor_3 g22339(n6628, new_n24687, new_n24600);
not_3  g22340(new_n24689, new_n2969);
xor_3  g22341(n6630, new_n24689, new_n2946);
xor_3  g22342(new_n24691, n25331, n17911);
nand_4 g22343(new_n24692, new_n19389_1, new_n15190);
nand_4 g22344(new_n24693, new_n23801, new_n23793);
nand_4 g22345(new_n24694, new_n24693, new_n24692);
xnor_3 g22346(new_n24695, new_n24694, new_n24691);
xnor_3 g22347(new_n24696, new_n24695, new_n8861_1);
not_3  g22348(new_n24697, new_n24696);
not_3  g22349(new_n24698, new_n23804);
nand_4 g22350(new_n24699, new_n23821, new_n23807);
nand_4 g22351(new_n24700, new_n24699, new_n24698);
xnor_3 g22352(new_n24701, new_n24700, new_n24697);
not_3  g22353(new_n24702, new_n24701);
xor_3  g22354(new_n24703, n14130, new_n9834);
not_3  g22355(new_n24704, n16482);
nand_4 g22356(new_n24705, new_n24704, n5400);
xor_3  g22357(new_n24706, n16482, new_n9840);
nor_4  g22358(new_n24707, new_n8258, n9942);
not_3  g22359(new_n24708, new_n24707);
nor_4  g22360(new_n24709, n25643, new_n9849);
not_3  g22361(new_n24710, new_n24709);
xor_3  g22362(new_n24711, n25643, new_n9849);
nor_4  g22363(new_n24712, new_n9857, n9557);
xor_3  g22364(new_n24713, n24170, new_n2359);
nor_4  g22365(new_n24714, new_n2364, n2409);
xor_3  g22366(new_n24715_1, n3136, new_n9858);
not_3  g22367(new_n24716, new_n24715_1);
nor_4  g22368(new_n24717, n8869, new_n2366);
not_3  g22369(new_n24718, new_n23302);
not_3  g22370(new_n24719, new_n23305_1);
nor_4  g22371(new_n24720, new_n24719, new_n24718);
nor_4  g22372(new_n24721, new_n24720, new_n24717);
nor_4  g22373(new_n24722, new_n24721, new_n24716);
nor_4  g22374(new_n24723_1, new_n24722, new_n24714);
and_4  g22375(new_n24724, new_n24723_1, new_n24713);
nor_4  g22376(new_n24725, new_n24724, new_n24712);
not_3  g22377(new_n24726, new_n24725);
nand_4 g22378(new_n24727, new_n24726, new_n24711);
nand_4 g22379(new_n24728, new_n24727, new_n24710);
xor_3  g22380(new_n24729, n23923, new_n2349);
nand_4 g22381(new_n24730, new_n24729, new_n24728);
nand_4 g22382(new_n24731, new_n24730, new_n24708);
nand_4 g22383(new_n24732_1, new_n24731, new_n24706);
nand_4 g22384(new_n24733, new_n24732_1, new_n24705);
xnor_3 g22385(new_n24734, new_n24733, new_n24703);
xnor_3 g22386(new_n24735, new_n24734, new_n24702);
not_3  g22387(new_n24736, new_n24706);
xnor_3 g22388(new_n24737, new_n24731, new_n24736);
nor_4  g22389(new_n24738, new_n24737, new_n23824);
xnor_3 g22390(new_n24739, new_n24737, new_n23822);
not_3  g22391(new_n24740, new_n24739);
not_3  g22392(new_n24741, new_n24729);
xnor_3 g22393(new_n24742, new_n24741, new_n24728);
nor_4  g22394(new_n24743, new_n24742, new_n23828);
xnor_3 g22395(new_n24744, new_n24725, new_n24711);
nor_4  g22396(new_n24745, new_n24744, new_n23382);
not_3  g22397(new_n24746, new_n24744);
nor_4  g22398(new_n24747, new_n24746, new_n23356);
nor_4  g22399(new_n24748, new_n24747, new_n24745);
not_3  g22400(new_n24749_1, new_n24748);
not_3  g22401(new_n24750, new_n23389);
xor_3  g22402(new_n24751, new_n24723_1, new_n24713);
nor_4  g22403(new_n24752, new_n24751, new_n24750);
xnor_3 g22404(new_n24753, new_n24751, new_n23389);
not_3  g22405(new_n24754, new_n24753);
xnor_3 g22406(new_n24755, new_n24721, new_n24716);
nor_4  g22407(new_n24756, new_n24755, new_n23391);
xnor_3 g22408(new_n24757, new_n24755, new_n23391);
nor_4  g22409(new_n24758_1, new_n23306, new_n23301);
nor_4  g22410(new_n24759, new_n23310, new_n23307);
nor_4  g22411(new_n24760, new_n24759, new_n24758_1);
nor_4  g22412(new_n24761, new_n24760, new_n24757);
nor_4  g22413(new_n24762, new_n24761, new_n24756);
nor_4  g22414(new_n24763, new_n24762, new_n24754);
nor_4  g22415(new_n24764, new_n24763, new_n24752);
nor_4  g22416(new_n24765, new_n24764, new_n24749_1);
nor_4  g22417(new_n24766, new_n24765, new_n24745);
xnor_3 g22418(new_n24767, new_n24742, new_n23829);
not_3  g22419(new_n24768_1, new_n24767);
nor_4  g22420(new_n24769, new_n24768_1, new_n24766);
nor_4  g22421(new_n24770, new_n24769, new_n24743);
nor_4  g22422(new_n24771, new_n24770, new_n24740);
nor_4  g22423(new_n24772, new_n24771, new_n24738);
xor_3  g22424(n6634, new_n24772, new_n24735);
not_3  g22425(new_n24774, new_n7721_1);
xor_3  g22426(n6652, new_n24774, new_n7704);
not_3  g22427(new_n24776, new_n15121);
xor_3  g22428(n6655, new_n24776, new_n15106);
not_3  g22429(new_n24778, new_n14497);
xor_3  g22430(n6669, new_n14528, new_n24778);
not_3  g22431(new_n24780, new_n11287);
xor_3  g22432(n6671, new_n24780, new_n11265);
not_3  g22433(new_n24782, new_n16390);
xor_3  g22434(n6673, new_n16412, new_n24782);
nand_4 g22435(new_n24784_1, new_n24409, new_n24402);
nor_4  g22436(new_n24785, new_n13787, new_n13774);
nand_4 g22437(new_n24786_1, new_n24406_1, new_n24785);
nand_4 g22438(n6674, new_n24786_1, new_n24784_1);
not_3  g22439(new_n24788, new_n20223);
xor_3  g22440(n6684, new_n20235_1, new_n24788);
xnor_3 g22441(n6706, new_n14812, new_n14754);
xor_3  g22442(new_n24791, n12702, n8614);
nand_4 g22443(new_n24792, new_n6433, new_n6326);
xor_3  g22444(new_n24793, n26797, n15182);
nor_4  g22445(new_n24794, n27037, n23913);
not_3  g22446(new_n24795, new_n24794);
xor_3  g22447(new_n24796, n27037, n23913);
nor_4  g22448(new_n24797, n22554, n8964);
not_3  g22449(new_n24798, new_n24797);
xor_3  g22450(new_n24799, n22554, n8964);
nor_4  g22451(new_n24800, n20429, n20151);
not_3  g22452(new_n24801, new_n24800);
xor_3  g22453(new_n24802, n20429, n20151);
nor_4  g22454(new_n24803, n7693, n3909);
not_3  g22455(new_n24804, new_n24803);
xor_3  g22456(new_n24805, n7693, n3909);
nor_4  g22457(new_n24806, n23974, n10405);
not_3  g22458(new_n24807_1, new_n24806);
xor_3  g22459(new_n24808, n23974, n10405);
nand_4 g22460(new_n24809, n11302, n2146);
not_3  g22461(new_n24810, new_n24809);
nor_4  g22462(new_n24811, n11302, n2146);
not_3  g22463(new_n24812, new_n19069);
nand_4 g22464(new_n24813, new_n19072, new_n19068);
nand_4 g22465(new_n24814, new_n24813, new_n24812);
nor_4  g22466(new_n24815, new_n24814, new_n24811);
nor_4  g22467(new_n24816, new_n24815, new_n24810);
nand_4 g22468(new_n24817, new_n24816, new_n24808);
nand_4 g22469(new_n24818, new_n24817, new_n24807_1);
nand_4 g22470(new_n24819, new_n24818, new_n24805);
nand_4 g22471(new_n24820, new_n24819, new_n24804);
nand_4 g22472(new_n24821, new_n24820, new_n24802);
nand_4 g22473(new_n24822, new_n24821, new_n24801);
nand_4 g22474(new_n24823, new_n24822, new_n24799);
nand_4 g22475(new_n24824, new_n24823, new_n24798);
nand_4 g22476(new_n24825, new_n24824, new_n24796);
nand_4 g22477(new_n24826_1, new_n24825, new_n24795);
nand_4 g22478(new_n24827, new_n24826_1, new_n24793);
nand_4 g22479(new_n24828, new_n24827, new_n24792);
not_3  g22480(new_n24829, new_n24828);
xor_3  g22481(new_n24830, new_n24829, new_n24791);
not_3  g22482(new_n24831, new_n24830);
nand_4 g22483(new_n24832, new_n24831, n1831);
not_3  g22484(new_n24833, new_n24832);
xnor_3 g22485(new_n24834, new_n24830, new_n16881);
not_3  g22486(new_n24835, new_n24826_1);
xnor_3 g22487(new_n24836, new_n24835, new_n24793);
not_3  g22488(new_n24837, new_n24836);
nor_4  g22489(new_n24838, new_n24837, new_n16885_1);
nor_4  g22490(new_n24839, new_n24836, n13137);
nor_4  g22491(new_n24840_1, new_n24839, new_n24838);
xnor_3 g22492(new_n24841_1, new_n24824, new_n24796);
not_3  g22493(new_n24842, new_n24841_1);
nand_4 g22494(new_n24843, new_n24842, n18452);
xor_3  g22495(new_n24844, new_n24842, n18452);
xnor_3 g22496(new_n24845, new_n24822, new_n24799);
not_3  g22497(new_n24846, new_n24845);
nand_4 g22498(new_n24847, new_n24846, n21317);
xor_3  g22499(new_n24848, new_n24846, n21317);
not_3  g22500(new_n24849, new_n24821);
nor_4  g22501(new_n24850, new_n24820, new_n24802);
nor_4  g22502(new_n24851, new_n24850, new_n24849);
nand_4 g22503(new_n24852, new_n24851, n12398);
xnor_3 g22504(new_n24853_1, new_n24851, new_n4426_1);
not_3  g22505(new_n24854, new_n24805);
xnor_3 g22506(new_n24855, new_n24818, new_n24854);
nand_4 g22507(new_n24856, new_n24855, n19789);
xnor_3 g22508(new_n24857_1, new_n24855, new_n16899);
not_3  g22509(new_n24858, new_n24816);
xnor_3 g22510(new_n24859, new_n24858, new_n24808);
nand_4 g22511(new_n24860, new_n24859, n20169);
xnor_3 g22512(new_n24861, new_n24859, new_n4507);
not_3  g22513(new_n24862, new_n24814);
nor_4  g22514(new_n24863, new_n24811, new_n24810);
xnor_3 g22515(new_n24864, new_n24863, new_n24862);
nand_4 g22516(new_n24865, new_n24864, n8285);
xnor_3 g22517(new_n24866, new_n24864, new_n14688);
not_3  g22518(new_n24867, new_n19066);
nand_4 g22519(new_n24868, new_n19073, new_n19067);
nand_4 g22520(new_n24869, new_n24868, new_n24867);
nand_4 g22521(new_n24870, new_n24869, new_n24866);
nand_4 g22522(new_n24871, new_n24870, new_n24865);
nand_4 g22523(new_n24872, new_n24871, new_n24861);
nand_4 g22524(new_n24873, new_n24872, new_n24860);
nand_4 g22525(new_n24874, new_n24873, new_n24857_1);
nand_4 g22526(new_n24875, new_n24874, new_n24856);
nand_4 g22527(new_n24876, new_n24875, new_n24853_1);
nand_4 g22528(new_n24877, new_n24876, new_n24852);
nand_4 g22529(new_n24878, new_n24877, new_n24848);
nand_4 g22530(new_n24879_1, new_n24878, new_n24847);
nand_4 g22531(new_n24880, new_n24879_1, new_n24844);
nand_4 g22532(new_n24881, new_n24880, new_n24843);
nand_4 g22533(new_n24882, new_n24881, new_n24840_1);
not_3  g22534(new_n24883, new_n24882);
nor_4  g22535(new_n24884, new_n24883, new_n24838);
nor_4  g22536(new_n24885, new_n24884, new_n24834);
nor_4  g22537(new_n24886, new_n24885, new_n24833);
nor_4  g22538(new_n24887_1, n12702, n8614);
not_3  g22539(new_n24888, new_n24791);
nor_4  g22540(new_n24889, new_n24829, new_n24888);
nor_4  g22541(new_n24890, new_n24889, new_n24887_1);
xnor_3 g22542(new_n24891, new_n24890, new_n24886);
not_3  g22543(new_n24892, new_n24461);
nand_4 g22544(new_n24893, new_n24483_1, new_n24892);
not_3  g22545(new_n24894, new_n24458);
nor_4  g22546(new_n24895, new_n24894, n1536);
xnor_3 g22547(new_n24896, new_n24895, new_n5125);
xnor_3 g22548(new_n24897, new_n24896, new_n24893);
not_3  g22549(new_n24898, new_n24897);
xnor_3 g22550(new_n24899, new_n24898, new_n24891);
xnor_3 g22551(new_n24900, new_n24884, new_n24834);
nor_4  g22552(new_n24901, new_n24900, new_n24486);
xnor_3 g22553(new_n24902, new_n24900, new_n24486);
xnor_3 g22554(new_n24903, new_n24881, new_n24840_1);
nor_4  g22555(new_n24904, new_n24903, new_n24509);
xnor_3 g22556(new_n24905, new_n24903, new_n24509);
xnor_3 g22557(new_n24906, new_n24879_1, new_n24844);
nor_4  g22558(new_n24907, new_n24906, new_n24516);
xnor_3 g22559(new_n24908, new_n24906, new_n24515);
xnor_3 g22560(new_n24909, new_n24877, new_n24848);
not_3  g22561(new_n24910, new_n24909);
nand_4 g22562(new_n24911, new_n24910, new_n24521);
xnor_3 g22563(new_n24912, new_n24909, new_n24521);
xnor_3 g22564(new_n24913, new_n24875, new_n24853_1);
nor_4  g22565(new_n24914, new_n24913, new_n16585);
not_3  g22566(new_n24915, new_n24914);
not_3  g22567(new_n24916, new_n24913);
nor_4  g22568(new_n24917, new_n24916, new_n24526);
nor_4  g22569(new_n24918, new_n24917, new_n24914);
xnor_3 g22570(new_n24919, new_n24873, new_n24857_1);
not_3  g22571(new_n24920, new_n24919);
nand_4 g22572(new_n24921, new_n24920, new_n16614);
xnor_3 g22573(new_n24922, new_n24919, new_n16614);
not_3  g22574(new_n24923, new_n24861);
xnor_3 g22575(new_n24924, new_n24871, new_n24923);
nand_4 g22576(new_n24925, new_n24924, new_n16618);
xnor_3 g22577(new_n24926, new_n24924, new_n16617_1);
not_3  g22578(new_n24927, new_n24866);
xnor_3 g22579(new_n24928, new_n24869, new_n24927);
nor_4  g22580(new_n24929, new_n24928, new_n16623);
not_3  g22581(new_n24930, new_n19061);
nand_4 g22582(new_n24931, new_n19079, new_n24930);
nand_4 g22583(new_n24932, new_n24931, new_n19076);
xnor_3 g22584(new_n24933, new_n24928, new_n16623);
nor_4  g22585(new_n24934_1, new_n24933, new_n24932);
nor_4  g22586(new_n24935, new_n24934_1, new_n24929);
nand_4 g22587(new_n24936, new_n24935, new_n24926);
nand_4 g22588(new_n24937_1, new_n24936, new_n24925);
nand_4 g22589(new_n24938, new_n24937_1, new_n24922);
nand_4 g22590(new_n24939, new_n24938, new_n24921);
nand_4 g22591(new_n24940, new_n24939, new_n24918);
nand_4 g22592(new_n24941, new_n24940, new_n24915);
nand_4 g22593(new_n24942, new_n24941, new_n24912);
nand_4 g22594(new_n24943, new_n24942, new_n24911);
nand_4 g22595(new_n24944, new_n24943, new_n24908);
not_3  g22596(new_n24945, new_n24944);
nor_4  g22597(new_n24946, new_n24945, new_n24907);
nor_4  g22598(new_n24947, new_n24946, new_n24905);
nor_4  g22599(new_n24948, new_n24947, new_n24904);
nor_4  g22600(new_n24949, new_n24948, new_n24902);
nor_4  g22601(new_n24950, new_n24949, new_n24901);
xnor_3 g22602(n6707, new_n24950, new_n24899);
xor_3  g22603(n6736, new_n15837, new_n15496_1);
xor_3  g22604(new_n24953, n23895, new_n19418);
not_3  g22605(new_n24954, new_n24953);
nor_4  g22606(new_n24955, n17351, new_n19422);
xor_3  g22607(new_n24956, n17351, new_n19422);
nand_4 g22608(new_n24957, n22470, new_n6330_1);
xor_3  g22609(new_n24958, n22470, new_n6330_1);
nand_4 g22610(new_n24959, new_n8081, n19116);
nand_4 g22611(new_n24960, new_n6335, n6861);
nand_4 g22612(new_n24961, new_n21941, new_n21920);
nand_4 g22613(new_n24962, new_n24961, new_n24960);
xor_3  g22614(new_n24963, n23200, new_n3275);
nand_4 g22615(new_n24964, new_n24963, new_n24962);
nand_4 g22616(new_n24965, new_n24964, new_n24959);
nand_4 g22617(new_n24966, new_n24965, new_n24958);
nand_4 g22618(new_n24967, new_n24966, new_n24957);
nand_4 g22619(new_n24968, new_n24967, new_n24956);
not_3  g22620(new_n24969, new_n24968);
nor_4  g22621(new_n24970, new_n24969, new_n24955);
xor_3  g22622(new_n24971, new_n24970, new_n24954);
nor_4  g22623(new_n24972, new_n21946, n22660);
not_3  g22624(new_n24973, new_n24972);
nor_4  g22625(new_n24974, new_n24973, n13490);
not_3  g22626(new_n24975, new_n24974);
nor_4  g22627(new_n24976, new_n24975, n9655);
not_3  g22628(new_n24977, new_n24976);
nor_4  g22629(new_n24978, new_n24977, n25345);
not_3  g22630(new_n24979, new_n24978);
xor_3  g22631(new_n24980, new_n24979, n13494);
not_3  g22632(new_n24981, new_n24980);
xor_3  g22633(new_n24982, new_n24981, n12650);
xor_3  g22634(new_n24983, new_n24976, new_n6381_1);
nor_4  g22635(new_n24984, new_n24983, new_n22783);
not_3  g22636(new_n24985, new_n24984);
not_3  g22637(new_n24986, new_n24983);
xor_3  g22638(new_n24987, new_n24986, n10201);
xor_3  g22639(new_n24988, new_n24975, n9655);
nor_4  g22640(new_n24989, new_n24988, new_n10735);
not_3  g22641(new_n24990, new_n24989);
not_3  g22642(new_n24991, new_n24988);
xor_3  g22643(new_n24992, new_n24991, n10593);
xor_3  g22644(new_n24993, new_n24972, new_n7988);
nor_4  g22645(new_n24994, new_n24993, new_n10738);
not_3  g22646(new_n24995, new_n24994);
not_3  g22647(new_n24996, new_n24993);
xor_3  g22648(new_n24997, new_n24996, n18290);
nor_4  g22649(new_n24998_1, new_n21947, new_n10744);
not_3  g22650(new_n24999, new_n24998_1);
nand_4 g22651(new_n25000, new_n21989, new_n21988);
nand_4 g22652(new_n25001, new_n25000, new_n24999);
nand_4 g22653(new_n25002, new_n25001, new_n24997);
nand_4 g22654(new_n25003, new_n25002, new_n24995);
nand_4 g22655(new_n25004, new_n25003, new_n24992);
nand_4 g22656(new_n25005, new_n25004, new_n24990);
nand_4 g22657(new_n25006_1, new_n25005, new_n24987);
nand_4 g22658(new_n25007, new_n25006_1, new_n24985);
xnor_3 g22659(new_n25008, new_n25007, new_n24982);
nand_4 g22660(new_n25009, new_n25008, new_n19381);
not_3  g22661(new_n25010, new_n25009);
nor_4  g22662(new_n25011, new_n25008, new_n19381);
nor_4  g22663(new_n25012, new_n25011, new_n25010);
xnor_3 g22664(new_n25013, new_n25005, new_n24987);
nand_4 g22665(new_n25014, new_n25013, new_n19386);
not_3  g22666(new_n25015, new_n25014);
xnor_3 g22667(new_n25016, new_n25003, new_n24992);
nor_4  g22668(new_n25017, new_n25016, new_n19390);
not_3  g22669(new_n25018, new_n25017);
xnor_3 g22670(new_n25019, new_n25016, new_n19392);
xnor_3 g22671(new_n25020, new_n25001, new_n24997);
nand_4 g22672(new_n25021, new_n25020, new_n19396);
xnor_3 g22673(new_n25022, new_n25020, new_n19398);
not_3  g22674(new_n25023_1, new_n21991);
nand_4 g22675(new_n25024, new_n25023_1, new_n19402);
nand_4 g22676(new_n25025, new_n22014, new_n21992);
nand_4 g22677(new_n25026, new_n25025, new_n25024);
nand_4 g22678(new_n25027, new_n25026, new_n25022);
nand_4 g22679(new_n25028, new_n25027, new_n25021);
not_3  g22680(new_n25029, new_n25028);
nand_4 g22681(new_n25030, new_n25029, new_n25019);
nand_4 g22682(new_n25031, new_n25030, new_n25018);
nor_4  g22683(new_n25032_1, new_n25013, new_n19386);
nor_4  g22684(new_n25033, new_n25032_1, new_n25015);
not_3  g22685(new_n25034, new_n25033);
nor_4  g22686(new_n25035, new_n25034, new_n25031);
nor_4  g22687(new_n25036, new_n25035, new_n25015);
xnor_3 g22688(new_n25037, new_n25036, new_n25012);
xnor_3 g22689(new_n25038, new_n25037, new_n24971);
not_3  g22690(new_n25039, new_n24956);
xor_3  g22691(new_n25040, new_n24967, new_n25039);
xnor_3 g22692(new_n25041, new_n25033, new_n25031);
not_3  g22693(new_n25042, new_n25041);
nand_4 g22694(new_n25043, new_n25042, new_n25040);
xnor_3 g22695(new_n25044, new_n25042, new_n25040);
not_3  g22696(new_n25045, new_n25044);
xor_3  g22697(new_n25046, new_n24965, new_n24958);
xnor_3 g22698(new_n25047, new_n25029, new_n25019);
nor_4  g22699(new_n25048, new_n25047, new_n25046);
not_3  g22700(new_n25049, new_n25048);
not_3  g22701(new_n25050, new_n25046);
not_3  g22702(new_n25051, new_n25047);
nor_4  g22703(new_n25052, new_n25051, new_n25050);
nor_4  g22704(new_n25053, new_n25052, new_n25048);
xor_3  g22705(new_n25054, new_n24963, new_n24962);
not_3  g22706(new_n25055, new_n25054);
xnor_3 g22707(new_n25056, new_n25026, new_n25022);
nor_4  g22708(new_n25057, new_n25056, new_n25055);
not_3  g22709(new_n25058, new_n25056);
xnor_3 g22710(new_n25059, new_n25058, new_n25054);
not_3  g22711(new_n25060, new_n21942);
nor_4  g22712(new_n25061, new_n22015, new_n25060);
nor_4  g22713(new_n25062_1, new_n22056, new_n22017);
nor_4  g22714(new_n25063, new_n25062_1, new_n25061);
nor_4  g22715(new_n25064, new_n25063, new_n25059);
nor_4  g22716(new_n25065, new_n25064, new_n25057);
nand_4 g22717(new_n25066, new_n25065, new_n25053);
nand_4 g22718(new_n25067, new_n25066, new_n25049);
nand_4 g22719(new_n25068_1, new_n25067, new_n25045);
nand_4 g22720(new_n25069, new_n25068_1, new_n25043);
nor_4  g22721(new_n25070, new_n25069, new_n25038);
not_3  g22722(new_n25071, new_n25038);
not_3  g22723(new_n25072, new_n25069);
nor_4  g22724(new_n25073_1, new_n25072, new_n25071);
nor_4  g22725(n6791, new_n25073_1, new_n25070);
not_3  g22726(new_n25075, new_n4058);
xor_3  g22727(n6802, new_n25075, new_n4038);
not_3  g22728(new_n25077, new_n19818);
xor_3  g22729(n6826, new_n19846, new_n25077);
not_3  g22730(new_n25079, new_n12079);
xor_3  g22731(n6835, new_n25079, new_n12054);
nor_4  g22732(new_n25081, new_n22335_1, new_n22309_1);
and_4  g22733(new_n25082, new_n22335_1, new_n22309_1);
nor_4  g22734(new_n25083_1, new_n25082, new_n25081);
not_3  g22735(new_n25084, new_n3074);
nand_4 g22736(new_n25085, new_n25084, n22379);
xor_3  g22737(new_n25086, new_n3074, new_n22313);
nand_4 g22738(new_n25087, new_n3121, n1662);
xor_3  g22739(new_n25088, new_n3122, new_n2987);
nand_4 g22740(new_n25089, new_n3127, n12875);
xor_3  g22741(new_n25090, new_n3128, new_n2989);
nor_4  g22742(new_n25091, new_n3133, new_n2993);
not_3  g22743(new_n25092, new_n25091);
nor_4  g22744(new_n25093, new_n3137, n5213);
xor_3  g22745(new_n25094_1, new_n3138, n5213);
nor_4  g22746(new_n25095, new_n10145, n4665);
nor_4  g22747(new_n25096, new_n3143, new_n3002);
nor_4  g22748(new_n25097_1, new_n25096, new_n25095);
not_3  g22749(new_n25098, new_n25097_1);
nor_4  g22750(new_n25099, new_n3152, new_n3007);
not_3  g22751(new_n25100, new_n25099);
not_3  g22752(new_n25101, new_n3152);
nor_4  g22753(new_n25102, new_n25101, n19005);
nor_4  g22754(new_n25103, new_n25102, new_n25099);
nand_4 g22755(new_n25104, new_n3165, n5438);
not_3  g22756(new_n25105, new_n25104);
nor_4  g22757(new_n25106, new_n25105, n4326);
not_3  g22758(new_n25107, new_n25106);
xor_3  g22759(new_n25108, new_n25105, n4326);
nand_4 g22760(new_n25109, new_n25108, new_n3169);
nand_4 g22761(new_n25110, new_n25109, new_n25107);
not_3  g22762(new_n25111, new_n25110);
nand_4 g22763(new_n25112, new_n25111, new_n25103);
nand_4 g22764(new_n25113, new_n25112, new_n25100);
nor_4  g22765(new_n25114, new_n25113, new_n25098);
nor_4  g22766(new_n25115, new_n25114, new_n25095);
nor_4  g22767(new_n25116, new_n25115, new_n25094_1);
nor_4  g22768(new_n25117, new_n25116, new_n25093);
xor_3  g22769(new_n25118, new_n3133, new_n2993);
nand_4 g22770(new_n25119_1, new_n25118, new_n25117);
nand_4 g22771(new_n25120_1, new_n25119_1, new_n25092);
nand_4 g22772(new_n25121, new_n25120_1, new_n25090);
nand_4 g22773(new_n25122, new_n25121, new_n25089);
nand_4 g22774(new_n25123, new_n25122, new_n25088);
nand_4 g22775(new_n25124, new_n25123, new_n25087);
nand_4 g22776(new_n25125, new_n25124, new_n25086);
nand_4 g22777(new_n25126_1, new_n25125, new_n25085);
nand_4 g22778(new_n25127, new_n25126_1, new_n25083_1);
not_3  g22779(new_n25128, new_n25127);
nor_4  g22780(new_n25129, new_n25128, new_n25081);
nor_4  g22781(new_n25130, new_n25129, new_n22330);
nor_4  g22782(new_n25131, new_n25130, new_n21898_1);
not_3  g22783(new_n25132, new_n25130);
nor_4  g22784(new_n25133_1, new_n25132, new_n21896);
nor_4  g22785(new_n25134, new_n25133_1, new_n25131);
xnor_3 g22786(new_n25135, new_n25129, new_n22330);
nand_4 g22787(new_n25136, new_n25135, new_n21902);
xnor_3 g22788(new_n25137, new_n25135, new_n21901);
xnor_3 g22789(new_n25138, new_n25126_1, new_n25083_1);
nand_4 g22790(new_n25139, new_n25138, new_n7126);
xnor_3 g22791(new_n25140, new_n25138, new_n15524);
xnor_3 g22792(new_n25141, new_n25124, new_n25086);
nand_4 g22793(new_n25142, new_n25141, new_n7128);
xnor_3 g22794(new_n25143, new_n25141, new_n15565);
xnor_3 g22795(new_n25144, new_n25122, new_n25088);
nand_4 g22796(new_n25145, new_n25144, new_n15569);
xnor_3 g22797(new_n25146, new_n25144, new_n7136);
xnor_3 g22798(new_n25147, new_n25120_1, new_n25090);
nand_4 g22799(new_n25148, new_n25147, new_n15574);
xnor_3 g22800(new_n25149, new_n25147, new_n7141);
xnor_3 g22801(new_n25150, new_n25118, new_n25117);
nand_4 g22802(new_n25151, new_n25150, new_n7146);
xnor_3 g22803(new_n25152, new_n25150, new_n7150);
not_3  g22804(new_n25153, new_n25115);
xnor_3 g22805(new_n25154, new_n25153, new_n25094_1);
nand_4 g22806(new_n25155_1, new_n25154, new_n7157);
xnor_3 g22807(new_n25156, new_n25154, new_n7155);
not_3  g22808(new_n25157, new_n25113);
nor_4  g22809(new_n25158, new_n25157, new_n25097_1);
nor_4  g22810(new_n25159, new_n25158, new_n25114);
nand_4 g22811(new_n25160, new_n25159, new_n15586);
not_3  g22812(new_n25161, new_n25160);
nor_4  g22813(new_n25162, new_n25159, new_n15586);
nor_4  g22814(new_n25163, new_n25162, new_n25161);
not_3  g22815(new_n25164, new_n7169);
xnor_3 g22816(new_n25165, new_n25111, new_n25103);
nand_4 g22817(new_n25166, new_n25165, new_n25164);
not_3  g22818(new_n25167, new_n25166);
nor_4  g22819(new_n25168_1, new_n25165, new_n25164);
nor_4  g22820(new_n25169, new_n25168_1, new_n25167);
not_3  g22821(new_n25170, new_n25109);
nor_4  g22822(new_n25171, new_n25108, new_n3169);
nor_4  g22823(new_n25172, new_n25171, new_n25170);
nand_4 g22824(new_n25173, new_n25172, new_n15592);
not_3  g22825(new_n25174, new_n6771);
nor_4  g22826(new_n25175, new_n6773_1, new_n25174);
not_3  g22827(new_n25176, new_n25173);
nor_4  g22828(new_n25177, new_n25172, new_n15592);
nor_4  g22829(new_n25178, new_n25177, new_n25176);
nand_4 g22830(new_n25179, new_n25178, new_n25175);
nand_4 g22831(new_n25180, new_n25179, new_n25173);
nand_4 g22832(new_n25181_1, new_n25180, new_n25169);
nand_4 g22833(new_n25182, new_n25181_1, new_n25166);
nand_4 g22834(new_n25183, new_n25182, new_n25163);
nand_4 g22835(new_n25184, new_n25183, new_n25160);
nand_4 g22836(new_n25185, new_n25184, new_n25156);
nand_4 g22837(new_n25186, new_n25185, new_n25155_1);
nand_4 g22838(new_n25187, new_n25186, new_n25152);
nand_4 g22839(new_n25188, new_n25187, new_n25151);
nand_4 g22840(new_n25189, new_n25188, new_n25149);
nand_4 g22841(new_n25190, new_n25189, new_n25148);
nand_4 g22842(new_n25191, new_n25190, new_n25146);
nand_4 g22843(new_n25192, new_n25191, new_n25145);
nand_4 g22844(new_n25193, new_n25192, new_n25143);
nand_4 g22845(new_n25194, new_n25193, new_n25142);
nand_4 g22846(new_n25195, new_n25194, new_n25140);
nand_4 g22847(new_n25196, new_n25195, new_n25139);
nand_4 g22848(new_n25197, new_n25196, new_n25137);
nand_4 g22849(new_n25198, new_n25197, new_n25136);
xnor_3 g22850(n6853, new_n25198, new_n25134);
xnor_3 g22851(new_n25200_1, new_n18123, new_n13403);
nor_4  g22852(new_n25201, new_n18131, new_n13410);
not_3  g22853(new_n25202, new_n25201);
not_3  g22854(new_n25203, new_n15621);
nand_4 g22855(new_n25204, new_n15640, new_n15624);
nand_4 g22856(new_n25205, new_n25204, new_n25203);
not_3  g22857(new_n25206, new_n18131);
nor_4  g22858(new_n25207, new_n25206, new_n13406);
nor_4  g22859(new_n25208, new_n25207, new_n25201);
nand_4 g22860(new_n25209_1, new_n25208, new_n25205);
nand_4 g22861(new_n25210, new_n25209_1, new_n25202);
xor_3  g22862(n6862, new_n25210, new_n25200_1);
not_3  g22863(new_n25212, new_n19318);
nand_4 g22864(new_n25213, new_n19349, new_n25212);
not_3  g22865(new_n25214, new_n13604);
nand_4 g22866(new_n25215_1, new_n13637, new_n13605);
nand_4 g22867(new_n25216, new_n25215_1, new_n25214);
nor_4  g22868(new_n25217, new_n13584, n23717);
nor_4  g22869(new_n25218, new_n13600, new_n13586);
nor_4  g22870(new_n25219, new_n25218, new_n25217);
xor_3  g22871(new_n25220, new_n25219, new_n22535);
xnor_3 g22872(new_n25221, new_n25220, new_n25216);
not_3  g22873(new_n25222, n22253);
nor_4  g22874(new_n25223, new_n25222, n8305);
nor_4  g22875(new_n25224, new_n19315_1, new_n19297);
nor_4  g22876(new_n25225, new_n25224, new_n25223);
not_3  g22877(new_n25226, new_n25225);
nand_4 g22878(new_n25227, new_n25226, new_n25221);
nand_4 g22879(new_n25228, new_n25227, new_n25213);
not_3  g22880(new_n25229, new_n25219);
nand_4 g22881(new_n25230, new_n25229, new_n22656);
nand_4 g22882(new_n25231, new_n25220, new_n25216);
nand_4 g22883(new_n25232, new_n25231, new_n25230);
not_3  g22884(new_n25233, new_n25232);
nor_4  g22885(new_n25234, new_n25233, new_n25228);
nand_4 g22886(new_n25235, new_n25233, new_n25225);
nand_4 g22887(new_n25236, new_n25225, new_n25221);
nand_4 g22888(new_n25237, new_n25236, new_n25228);
nand_4 g22889(new_n25238, new_n25237, new_n25235);
nor_4  g22890(n6863, new_n25238, new_n25234);
xor_3  g22891(n6867, new_n7195, new_n7133);
not_3  g22892(new_n25241, new_n21833);
xor_3  g22893(n6965, new_n25241, new_n21826);
xnor_3 g22894(n6967, new_n8779, new_n8733);
xor_3  g22895(n6975, new_n17560, new_n17501);
xor_3  g22896(n6983, new_n24383, new_n24382);
xnor_3 g22897(new_n25246, new_n18090, new_n13381);
nor_4  g22898(new_n25247, new_n18095, new_n13383);
not_3  g22899(new_n25248, new_n25247);
nor_4  g22900(new_n25249, new_n18099, new_n13387);
nor_4  g22901(new_n25250, new_n25249, new_n25247);
nand_4 g22902(new_n25251, new_n18102, new_n13395);
xnor_3 g22903(new_n25252, new_n18102, new_n13391);
nand_4 g22904(new_n25253, new_n18108, new_n13398);
xnor_3 g22905(new_n25254_1, new_n18107, new_n13398);
nor_4  g22906(new_n25255, new_n18127, new_n13403);
not_3  g22907(new_n25256_1, new_n25255);
nand_4 g22908(new_n25257, new_n25210, new_n25200_1);
nand_4 g22909(new_n25258, new_n25257, new_n25256_1);
nand_4 g22910(new_n25259, new_n25258, new_n25254_1);
nand_4 g22911(new_n25260, new_n25259, new_n25253);
not_3  g22912(new_n25261, new_n25260);
nand_4 g22913(new_n25262, new_n25261, new_n25252);
nand_4 g22914(new_n25263, new_n25262, new_n25251);
nand_4 g22915(new_n25264, new_n25263, new_n25250);
nand_4 g22916(new_n25265, new_n25264, new_n25248);
xnor_3 g22917(n6985, new_n25265, new_n25246);
xnor_3 g22918(n6998, new_n17881, new_n17830);
xor_3  g22919(n7032, new_n14785, new_n10635);
xnor_3 g22920(n7038, new_n24210, new_n24170_1);
not_3  g22921(new_n25270, new_n21592);
xor_3  g22922(n7079, new_n21595, new_n25270);
not_3  g22923(new_n25272, new_n8765);
xor_3  g22924(n7190, new_n8768, new_n25272);
xnor_3 g22925(n7229, new_n19255, new_n19252);
not_3  g22926(new_n25275, new_n10216);
xor_3  g22927(n7230, new_n25275, new_n10202);
not_3  g22928(new_n25277, new_n23271);
xor_3  g22929(n7233, new_n25277, new_n23270_1);
not_3  g22930(new_n25279, new_n15976);
xor_3  g22931(n7236, new_n25279, new_n15966);
xor_3  g22932(n7253, new_n19704, new_n8177);
not_3  g22933(new_n25282, new_n23737);
nand_4 g22934(new_n25283, new_n23744, new_n25282);
nor_4  g22935(new_n25284, new_n23735, n17458);
nor_4  g22936(new_n25285, new_n23739, new_n25284);
nand_4 g22937(new_n25286, new_n25285, new_n25283);
not_3  g22938(new_n25287, new_n24301);
xnor_3 g22939(new_n25288, new_n25287, new_n17104_1);
nand_4 g22940(new_n25289, new_n25288, new_n12166);
xnor_3 g22941(new_n25290, new_n25288, new_n12228_1);
nor_4  g22942(new_n25291, new_n24303, new_n12172);
not_3  g22943(new_n25292, new_n25291);
not_3  g22944(new_n25293_1, new_n24304);
nand_4 g22945(new_n25294, new_n24346, new_n25293_1);
nand_4 g22946(new_n25295, new_n25294, new_n25292);
nand_4 g22947(new_n25296_1, new_n25295, new_n25290);
nand_4 g22948(new_n25297, new_n25296_1, new_n25289);
nor_4  g22949(new_n25298, new_n25287, new_n17104_1);
not_3  g22950(new_n25299, new_n25298);
nand_4 g22951(new_n25300, new_n25299, new_n17162);
nand_4 g22952(new_n25301, new_n25298, new_n17160);
nand_4 g22953(new_n25302, new_n25301, new_n25300);
not_3  g22954(new_n25303, new_n25302);
nor_4  g22955(new_n25304, new_n25303, new_n12161_1);
not_3  g22956(new_n25305, new_n12161_1);
nor_4  g22957(new_n25306, new_n25302, new_n25305);
nor_4  g22958(new_n25307, new_n25306, new_n25304);
not_3  g22959(new_n25308, new_n25307);
xnor_3 g22960(new_n25309, new_n25308, new_n25297);
nand_4 g22961(new_n25310, new_n25309, new_n25286);
not_3  g22962(new_n25311, new_n25286);
xnor_3 g22963(new_n25312, new_n25309, new_n25311);
not_3  g22964(new_n25313, new_n25290);
xnor_3 g22965(new_n25314, new_n25295, new_n25313);
nand_4 g22966(new_n25315, new_n25314, new_n23745);
nor_4  g22967(new_n25316_1, new_n24347_1, new_n20314);
nor_4  g22968(new_n25317, new_n24398, new_n24348);
nor_4  g22969(new_n25318, new_n25317, new_n25316_1);
xnor_3 g22970(new_n25319, new_n25314, new_n23746);
nand_4 g22971(new_n25320, new_n25319, new_n25318);
nand_4 g22972(new_n25321, new_n25320, new_n25315);
nand_4 g22973(new_n25322, new_n25321, new_n25312);
nand_4 g22974(new_n25323, new_n25322, new_n25310);
nor_4  g22975(new_n25324, new_n25304, new_n25297);
not_3  g22976(new_n25325, new_n25306);
nand_4 g22977(new_n25326, new_n25325, new_n25301);
nor_4  g22978(new_n25327, new_n25326, new_n25324);
xnor_3 g22979(n7256, new_n25327, new_n25323);
nor_4  g22980(new_n25329, new_n10424, n2416);
xor_3  g22981(new_n25330, n22764, new_n11802);
not_3  g22982(new_n25331_1, new_n25330);
not_3  g22983(new_n25332_1, n26264);
nor_4  g22984(new_n25333, new_n25332_1, n21905);
nand_4 g22985(new_n25334, new_n23857, new_n23846);
not_3  g22986(new_n25335, new_n25334);
nor_4  g22987(new_n25336_1, new_n25335, new_n25333);
nor_4  g22988(new_n25337_1, new_n25336_1, new_n25331_1);
nor_4  g22989(new_n25338, new_n25337_1, new_n25329);
not_3  g22990(new_n25339, new_n25338);
not_3  g22991(new_n25340, new_n25336_1);
nor_4  g22992(new_n25341, new_n25340, new_n25330);
nor_4  g22993(new_n25342, new_n25341, new_n25337_1);
nand_4 g22994(new_n25343, new_n25342, new_n18905);
xnor_3 g22995(new_n25344, new_n25342, new_n18902);
not_3  g22996(new_n25345_1, new_n23859);
nand_4 g22997(new_n25346, new_n23879, new_n25345_1);
nand_4 g22998(new_n25347, new_n25346, new_n25344);
nand_4 g22999(new_n25348, new_n25347, new_n25343);
xnor_3 g23000(new_n25349, new_n25348, new_n25339);
nand_4 g23001(new_n25350, new_n25349, new_n18964);
not_3  g23002(new_n25351, new_n18964);
xnor_3 g23003(new_n25352, new_n25348, new_n25338);
nand_4 g23004(new_n25353, new_n25352, new_n25351);
nand_4 g23005(new_n25354, new_n25353, new_n25350);
xnor_3 g23006(new_n25355, new_n25354, new_n23983);
not_3  g23007(new_n25356_1, new_n25347);
nor_4  g23008(new_n25357, new_n25346, new_n25344);
nor_4  g23009(new_n25358, new_n25357, new_n25356_1);
nor_4  g23010(new_n25359, new_n25358, new_n23997);
not_3  g23011(new_n25360, new_n25359);
not_3  g23012(new_n25361, new_n25358);
nor_4  g23013(new_n25362_1, new_n25361, new_n24000);
nor_4  g23014(new_n25363, new_n25362_1, new_n25359);
nor_4  g23015(new_n25364, new_n23882, new_n23845);
not_3  g23016(new_n25365_1, new_n25364);
not_3  g23017(new_n25366, new_n23883_1);
nand_4 g23018(new_n25367, new_n23901, new_n25366);
nand_4 g23019(new_n25368, new_n25367, new_n25365_1);
nand_4 g23020(new_n25369, new_n25368, new_n25363);
nand_4 g23021(new_n25370_1, new_n25369, new_n25360);
xnor_3 g23022(n7268, new_n25370_1, new_n25355);
not_3  g23023(new_n25372, new_n13083);
nor_4  g23024(new_n25373, new_n25372, n752);
not_3  g23025(new_n25374, new_n25373);
nor_4  g23026(new_n25375, new_n25374, n2175);
not_3  g23027(new_n25376, new_n25375);
nor_4  g23028(new_n25377, new_n25376, n13026);
not_3  g23029(new_n25378, new_n25377);
nor_4  g23030(new_n25379, new_n25378, n23912);
not_3  g23031(new_n25380, new_n25379);
not_3  g23032(new_n25381_1, n10514);
xor_3  g23033(new_n25382, new_n25378, n23912);
nor_4  g23034(new_n25383, new_n25382, new_n25381_1);
not_3  g23035(new_n25384, new_n25383);
not_3  g23036(new_n25385, new_n25382);
xor_3  g23037(new_n25386, new_n25385, n10514);
not_3  g23038(new_n25387, n18649);
xor_3  g23039(new_n25388, new_n25375, new_n13975);
nor_4  g23040(new_n25389, new_n25388, new_n25387);
not_3  g23041(new_n25390, new_n25389);
not_3  g23042(new_n25391, new_n25388);
xor_3  g23043(new_n25392, new_n25391, n18649);
not_3  g23044(new_n25393, n6218);
xor_3  g23045(new_n25394, new_n25374, n2175);
nor_4  g23046(new_n25395, new_n25394, new_n25393);
not_3  g23047(new_n25396, new_n25395);
not_3  g23048(new_n25397, new_n25394);
xor_3  g23049(new_n25398, new_n25397, n6218);
nor_4  g23050(new_n25399, new_n13084, new_n13724);
not_3  g23051(new_n25400, new_n25399);
not_3  g23052(new_n25401, new_n13084);
xor_3  g23053(new_n25402, new_n25401, n20470);
not_3  g23054(new_n25403, n21222);
nor_4  g23055(new_n25404, new_n13087, new_n25403);
not_3  g23056(new_n25405, new_n25404);
xor_3  g23057(new_n25406, new_n13088, n21222);
not_3  g23058(new_n25407, n9832);
nor_4  g23059(new_n25408, new_n13094, new_n25407);
not_3  g23060(new_n25409, new_n13094);
nor_4  g23061(new_n25410, new_n25409, n9832);
nor_4  g23062(new_n25411, new_n25410, new_n25408);
not_3  g23063(new_n25412_1, n1558);
nor_4  g23064(new_n25413, new_n13099, new_n25412_1);
not_3  g23065(new_n25414, new_n25413);
not_3  g23066(new_n25415, new_n13099);
nor_4  g23067(new_n25416, new_n25415, n1558);
nor_4  g23068(new_n25417, new_n25416, new_n25413);
not_3  g23069(new_n25418, n21749);
nor_4  g23070(new_n25419, new_n13103, new_n25418);
not_3  g23071(new_n25420, new_n25419);
not_3  g23072(new_n25421, new_n13103);
nor_4  g23073(new_n25422, new_n25421, n21749);
nor_4  g23074(new_n25423, new_n25422, new_n25419);
not_3  g23075(new_n25424, n7769);
nor_4  g23076(new_n25425, new_n13109, new_n25424);
not_3  g23077(new_n25426, new_n25425);
not_3  g23078(new_n25427, n21138);
nor_4  g23079(new_n25428, new_n25427, n15506);
nor_4  g23080(new_n25429, new_n13108, n7769);
nor_4  g23081(new_n25430, new_n25429, new_n25425);
nand_4 g23082(new_n25431, new_n25430, new_n25428);
nand_4 g23083(new_n25432, new_n25431, new_n25426);
nand_4 g23084(new_n25433, new_n25432, new_n25423);
nand_4 g23085(new_n25434, new_n25433, new_n25420);
nand_4 g23086(new_n25435_1, new_n25434, new_n25417);
nand_4 g23087(new_n25436, new_n25435_1, new_n25414);
nand_4 g23088(new_n25437, new_n25436, new_n25411);
not_3  g23089(new_n25438, new_n25437);
nor_4  g23090(new_n25439, new_n25438, new_n25408);
not_3  g23091(new_n25440, new_n25439);
nand_4 g23092(new_n25441, new_n25440, new_n25406);
nand_4 g23093(new_n25442, new_n25441, new_n25405);
nand_4 g23094(new_n25443, new_n25442, new_n25402);
nand_4 g23095(new_n25444, new_n25443, new_n25400);
nand_4 g23096(new_n25445, new_n25444, new_n25398);
nand_4 g23097(new_n25446, new_n25445, new_n25396);
nand_4 g23098(new_n25447, new_n25446, new_n25392);
nand_4 g23099(new_n25448, new_n25447, new_n25390);
nand_4 g23100(new_n25449, new_n25448, new_n25386);
nand_4 g23101(new_n25450, new_n25449, new_n25384);
nor_4  g23102(new_n25451, new_n25450, new_n25380);
not_3  g23103(new_n25452, new_n25449);
nor_4  g23104(new_n25453, new_n25448, new_n25386);
nor_4  g23105(new_n25454, new_n25453, new_n25452);
nor_4  g23106(new_n25455, new_n25454, n9872);
not_3  g23107(new_n25456, n9872);
xnor_3 g23108(new_n25457, new_n25454, new_n25456);
not_3  g23109(new_n25458, n5842);
xnor_3 g23110(new_n25459, new_n25446, new_n25392);
nand_4 g23111(new_n25460_1, new_n25459, new_n25458);
xnor_3 g23112(new_n25461, new_n25459, n5842);
not_3  g23113(new_n25462, n6379);
xnor_3 g23114(new_n25463, new_n25444, new_n25398);
nand_4 g23115(new_n25464_1, new_n25463, new_n25462);
xnor_3 g23116(new_n25465, new_n25463, n6379);
not_3  g23117(new_n25466, new_n25402);
xnor_3 g23118(new_n25467, new_n25442, new_n25466);
nor_4  g23119(new_n25468_1, new_n25467, n2102);
not_3  g23120(new_n25469, new_n25468_1);
not_3  g23121(new_n25470, n2102);
not_3  g23122(new_n25471_1, new_n25467);
nor_4  g23123(new_n25472, new_n25471_1, new_n25470);
nor_4  g23124(new_n25473, new_n25472, new_n25468_1);
xnor_3 g23125(new_n25474, new_n25439, new_n25406);
nor_4  g23126(new_n25475_1, new_n25474, n17954);
not_3  g23127(new_n25476, new_n25475_1);
not_3  g23128(new_n25477, n8256);
xnor_3 g23129(new_n25478, new_n25436, new_n25411);
nand_4 g23130(new_n25479, new_n25478, new_n25477);
xnor_3 g23131(new_n25480, new_n25478, n8256);
not_3  g23132(new_n25481, n24150);
xnor_3 g23133(new_n25482, new_n25434, new_n25417);
nand_4 g23134(new_n25483, new_n25482, new_n25481);
xnor_3 g23135(new_n25484, new_n25482, n24150);
xnor_3 g23136(new_n25485, new_n25432, new_n25423);
nand_4 g23137(new_n25486, new_n25485, new_n20082);
xnor_3 g23138(new_n25487, new_n25485, n19584);
xnor_3 g23139(new_n25488, new_n25430, new_n25428);
nor_4  g23140(new_n25489, new_n25488, new_n20097);
not_3  g23141(new_n25490, new_n25488);
nor_4  g23142(new_n25491, new_n25490, n5060);
xor_3  g23143(new_n25492, n21138, new_n13106);
nand_4 g23144(new_n25493, new_n25492, n15332);
nor_4  g23145(new_n25494_1, new_n25493, new_n25491);
nor_4  g23146(new_n25495, new_n25494_1, new_n25489);
nand_4 g23147(new_n25496, new_n25495, new_n25487);
nand_4 g23148(new_n25497, new_n25496, new_n25486);
nand_4 g23149(new_n25498, new_n25497, new_n25484);
nand_4 g23150(new_n25499_1, new_n25498, new_n25483);
nand_4 g23151(new_n25500, new_n25499_1, new_n25480);
nand_4 g23152(new_n25501, new_n25500, new_n25479);
not_3  g23153(new_n25502, n17954);
not_3  g23154(new_n25503, new_n25474);
nor_4  g23155(new_n25504, new_n25503, new_n25502);
nor_4  g23156(new_n25505, new_n25504, new_n25475_1);
nand_4 g23157(new_n25506, new_n25505, new_n25501);
nand_4 g23158(new_n25507, new_n25506, new_n25476);
nand_4 g23159(new_n25508, new_n25507, new_n25473);
nand_4 g23160(new_n25509, new_n25508, new_n25469);
nand_4 g23161(new_n25510, new_n25509, new_n25465);
nand_4 g23162(new_n25511, new_n25510, new_n25464_1);
nand_4 g23163(new_n25512, new_n25511, new_n25461);
nand_4 g23164(new_n25513_1, new_n25512, new_n25460_1);
nand_4 g23165(new_n25514, new_n25513_1, new_n25457);
not_3  g23166(new_n25515, new_n25514);
nor_4  g23167(new_n25516, new_n25515, new_n25455);
not_3  g23168(new_n25517, new_n25516);
nand_4 g23169(new_n25518_1, new_n25517, new_n25451);
not_3  g23170(new_n25519, new_n25450);
nor_4  g23171(new_n25520, new_n25519, new_n25379);
nand_4 g23172(new_n25521, new_n25520, new_n25516);
nand_4 g23173(new_n25522, new_n25521, new_n25518_1);
xnor_3 g23174(new_n25523_1, new_n25522, new_n17817);
nor_4  g23175(new_n25524, new_n25520, new_n25451);
xnor_3 g23176(new_n25525, new_n25524, new_n25516);
not_3  g23177(new_n25526, new_n25525);
nor_4  g23178(new_n25527, new_n25526, new_n17821);
xnor_3 g23179(new_n25528, new_n25525, new_n17820_1);
xnor_3 g23180(new_n25529, new_n25513_1, new_n25457);
nand_4 g23181(new_n25530, new_n25529, new_n17826);
xnor_3 g23182(new_n25531, new_n25529, new_n2756);
xnor_3 g23183(new_n25532_1, new_n25511, new_n25461);
nand_4 g23184(new_n25533, new_n25532_1, new_n2913);
xnor_3 g23185(new_n25534, new_n25509, new_n25465);
nand_4 g23186(new_n25535, new_n25534, new_n2917);
xnor_3 g23187(new_n25536, new_n25534, new_n2922);
xnor_3 g23188(new_n25537, new_n25507, new_n25473);
nand_4 g23189(new_n25538, new_n25537, new_n2924);
xnor_3 g23190(new_n25539_1, new_n25537, new_n2925);
xnor_3 g23191(new_n25540, new_n25505, new_n25501);
nand_4 g23192(new_n25541, new_n25540, new_n2931);
not_3  g23193(new_n25542, new_n25541);
nor_4  g23194(new_n25543, new_n25540, new_n2931);
nor_4  g23195(new_n25544, new_n25543, new_n25542);
xnor_3 g23196(new_n25545, new_n25499_1, new_n25480);
nand_4 g23197(new_n25546, new_n25545, new_n2937);
xnor_3 g23198(new_n25547, new_n25545, new_n2936);
xnor_3 g23199(new_n25548, new_n25497, new_n25484);
nand_4 g23200(new_n25549, new_n25548, new_n2944_1);
xnor_3 g23201(new_n25550_1, new_n25548, new_n17848);
not_3  g23202(new_n25551, new_n25487);
xnor_3 g23203(new_n25552, new_n25495, new_n25551);
nor_4  g23204(new_n25553, new_n25552, new_n2951);
not_3  g23205(new_n25554, new_n25553);
not_3  g23206(new_n25555, new_n25552);
nor_4  g23207(new_n25556, new_n25555, new_n2952);
nor_4  g23208(new_n25557, new_n25556, new_n25553);
not_3  g23209(new_n25558, new_n25493);
nor_4  g23210(new_n25559, new_n25491, new_n25489);
xnor_3 g23211(new_n25560, new_n25559, new_n25558);
nor_4  g23212(new_n25561, new_n25560, new_n2959);
not_3  g23213(new_n25562, new_n25561);
not_3  g23214(new_n25563, new_n25492);
xor_3  g23215(new_n25564, new_n25563, n15332);
nand_4 g23216(new_n25565_1, new_n25564, new_n2962);
not_3  g23217(new_n25566, new_n25560);
nor_4  g23218(new_n25567, new_n25566, new_n2960);
nor_4  g23219(new_n25568, new_n25567, new_n25561);
nand_4 g23220(new_n25569, new_n25568, new_n25565_1);
nand_4 g23221(new_n25570, new_n25569, new_n25562);
nand_4 g23222(new_n25571, new_n25570, new_n25557);
nand_4 g23223(new_n25572, new_n25571, new_n25554);
nand_4 g23224(new_n25573, new_n25572, new_n25550_1);
nand_4 g23225(new_n25574, new_n25573, new_n25549);
nand_4 g23226(new_n25575, new_n25574, new_n25547);
nand_4 g23227(new_n25576, new_n25575, new_n25546);
nand_4 g23228(new_n25577, new_n25576, new_n25544);
nand_4 g23229(new_n25578, new_n25577, new_n25541);
nand_4 g23230(new_n25579, new_n25578, new_n25539_1);
nand_4 g23231(new_n25580, new_n25579, new_n25538);
nand_4 g23232(new_n25581, new_n25580, new_n25536);
nand_4 g23233(new_n25582, new_n25581, new_n25535);
xnor_3 g23234(new_n25583, new_n25532_1, new_n2912);
nand_4 g23235(new_n25584, new_n25583, new_n25582);
nand_4 g23236(new_n25585, new_n25584, new_n25533);
nand_4 g23237(new_n25586_1, new_n25585, new_n25531);
nand_4 g23238(new_n25587, new_n25586_1, new_n25530);
not_3  g23239(new_n25588, new_n25587);
nor_4  g23240(new_n25589, new_n25588, new_n25528);
nor_4  g23241(new_n25590, new_n25589, new_n25527);
xnor_3 g23242(n7277, new_n25590, new_n25523_1);
xor_3  g23243(n7280, new_n16202, new_n16189);
not_3  g23244(new_n25593, new_n6669_1);
xor_3  g23245(n7298, new_n6705, new_n25593);
not_3  g23246(new_n25595, new_n23725);
xor_3  g23247(n7308, new_n25595, new_n23711);
not_3  g23248(new_n25597, new_n8546);
nor_4  g23249(new_n25598, new_n23992, new_n25597);
nand_4 g23250(new_n25599, new_n23992, new_n25597);
not_3  g23251(new_n25600, new_n25599);
nor_4  g23252(new_n25601, new_n25600, new_n25598);
nand_4 g23253(new_n25602, new_n23996, new_n8571);
xnor_3 g23254(new_n25603, new_n23995, new_n8571);
nand_4 g23255(new_n25604, new_n24004_1, new_n8578);
nand_4 g23256(new_n25605, new_n18226, new_n18189);
nand_4 g23257(new_n25606, new_n25605, new_n25604);
nand_4 g23258(new_n25607, new_n25606, new_n25603);
nand_4 g23259(new_n25608, new_n25607, new_n25602);
not_3  g23260(new_n25609, new_n25608);
nand_4 g23261(new_n25610, new_n25609, new_n25601);
not_3  g23262(new_n25611_1, new_n25610);
nor_4  g23263(new_n25612, new_n25609, new_n25601);
nor_4  g23264(new_n25613, new_n25612, new_n25611_1);
nor_4  g23265(new_n25614_1, new_n25613, new_n24031);
not_3  g23266(new_n25615, new_n25613);
nor_4  g23267(new_n25616, new_n25615, new_n24030);
nor_4  g23268(new_n25617, new_n25616, new_n25614_1);
not_3  g23269(new_n25618, new_n25603);
xnor_3 g23270(new_n25619_1, new_n25606, new_n25618);
nor_4  g23271(new_n25620, new_n25619_1, new_n24041);
not_3  g23272(new_n25621, new_n25620);
not_3  g23273(new_n25622, new_n18227_1);
nor_4  g23274(new_n25623, new_n24049, new_n25622);
nor_4  g23275(new_n25624, new_n23279, new_n23244);
nor_4  g23276(new_n25625, new_n25624, new_n25623);
xnor_3 g23277(new_n25626, new_n25606, new_n25603);
nor_4  g23278(new_n25627, new_n25626, new_n24042);
nor_4  g23279(new_n25628, new_n25627, new_n25620);
nand_4 g23280(new_n25629_1, new_n25628, new_n25625);
nand_4 g23281(new_n25630, new_n25629_1, new_n25621);
xnor_3 g23282(n7313, new_n25630, new_n25617);
not_3  g23283(new_n25632, new_n4024);
xor_3  g23284(n7346, new_n4062, new_n25632);
nor_4  g23285(new_n25634, new_n25229, new_n16983);
nor_4  g23286(new_n25635, new_n25219, new_n16986);
nor_4  g23287(new_n25636, new_n25635, new_n25634);
nor_4  g23288(new_n25637, new_n25219, new_n16993);
not_3  g23289(new_n25638, new_n25637);
nor_4  g23290(new_n25639, new_n25229, new_n16991);
nor_4  g23291(new_n25640, new_n25639, new_n25637);
nand_4 g23292(new_n25641, new_n16998, new_n13603);
xnor_3 g23293(new_n25642, new_n16998, new_n13601);
nor_4  g23294(new_n25643_1, new_n17003, new_n13608);
not_3  g23295(new_n25644, new_n25643_1);
nor_4  g23296(new_n25645, new_n17007, new_n13609);
nor_4  g23297(new_n25646, new_n25645, new_n25643_1);
nand_4 g23298(new_n25647, new_n17012, new_n13617);
nor_4  g23299(new_n25648, new_n7682, new_n7524_1);
nor_4  g23300(new_n25649, new_n7727, new_n7683);
nor_4  g23301(new_n25650, new_n25649, new_n25648);
xnor_3 g23302(new_n25651, new_n17012, new_n13618);
nand_4 g23303(new_n25652, new_n25651, new_n25650);
nand_4 g23304(new_n25653, new_n25652, new_n25647);
nand_4 g23305(new_n25654, new_n25653, new_n25646);
nand_4 g23306(new_n25655, new_n25654, new_n25644);
nand_4 g23307(new_n25656, new_n25655, new_n25642);
nand_4 g23308(new_n25657, new_n25656, new_n25641);
nand_4 g23309(new_n25658, new_n25657, new_n25640);
nand_4 g23310(new_n25659, new_n25658, new_n25638);
xnor_3 g23311(n7349, new_n25659, new_n25636);
xnor_3 g23312(n7363, new_n25585, new_n25531);
nor_4  g23313(new_n25662, n21839, new_n10728);
nor_4  g23314(new_n25663, new_n23968, new_n23964);
nor_4  g23315(new_n25664, new_n25663, new_n25662);
xnor_3 g23316(new_n25665_1, new_n25664, new_n12233);
nor_4  g23317(new_n25666, new_n23969, new_n12236);
nor_4  g23318(new_n25667, new_n23974_1, new_n23970);
nor_4  g23319(new_n25668, new_n25667, new_n25666);
xnor_3 g23320(n7390, new_n25668, new_n25665_1);
not_3  g23321(new_n25670, new_n10850);
xor_3  g23322(n7403, new_n10851_1, new_n25670);
xor_3  g23323(n7408, new_n11076, new_n11027);
not_3  g23324(new_n25673, new_n24392);
xor_3  g23325(n7432, new_n25673, new_n24363);
not_3  g23326(new_n25675, new_n21897);
nand_4 g23327(new_n25676, new_n21911, new_n21900);
nand_4 g23328(n7475, new_n25676, new_n25675);
xor_3  g23329(n7477, new_n5995, new_n5993);
not_3  g23330(new_n25679, new_n10616);
xor_3  g23331(n7507, new_n10652, new_n25679);
nor_4  g23332(new_n25681, new_n14412_1, new_n6319);
not_3  g23333(new_n25682, new_n25681);
nor_4  g23334(new_n25683, new_n14415, n23895);
nor_4  g23335(new_n25684, new_n25683, new_n25681);
nor_4  g23336(new_n25685, new_n8074, new_n6324);
not_3  g23337(new_n25686, new_n25685);
nand_4 g23338(new_n25687, new_n8133, new_n8075);
nand_4 g23339(new_n25688, new_n25687, new_n25686);
nand_4 g23340(new_n25689, new_n25688, new_n25684);
nand_4 g23341(new_n25690, new_n25689, new_n25682);
xnor_3 g23342(new_n25691, new_n25690, new_n14468);
xnor_3 g23343(new_n25692, new_n25691, new_n21048);
xnor_3 g23344(new_n25693, new_n25688, new_n25684);
nand_4 g23345(new_n25694_1, new_n25693, new_n21063);
xnor_3 g23346(new_n25695, new_n25693, new_n21064);
not_3  g23347(new_n25696, new_n8043);
nand_4 g23348(new_n25697, new_n8134, new_n25696);
nand_4 g23349(new_n25698, new_n8198, new_n8135_1);
nand_4 g23350(new_n25699, new_n25698, new_n25697);
nand_4 g23351(new_n25700, new_n25699, new_n25695);
nand_4 g23352(new_n25701, new_n25700, new_n25694_1);
xnor_3 g23353(n7514, new_n25701, new_n25692);
xnor_3 g23354(n7558, new_n13063, new_n13031);
not_3  g23355(new_n25704, new_n14519);
xor_3  g23356(n7572, new_n14522, new_n25704);
nor_4  g23357(new_n25706_1, new_n7335_1, new_n4447);
nor_4  g23358(new_n25707, new_n14941, n7693);
nor_4  g23359(new_n25708, new_n25707, new_n25706_1);
nand_4 g23360(new_n25709, new_n24428, new_n24418);
nand_4 g23361(new_n25710, new_n25709, new_n24415_1);
xnor_3 g23362(new_n25711, new_n25710, new_n25708);
nor_4  g23363(new_n25712, new_n25711, new_n11663);
not_3  g23364(new_n25713, new_n11581);
nor_4  g23365(new_n25714, new_n11580_1, new_n11560);
nor_4  g23366(new_n25715, new_n25714, new_n25713);
xnor_3 g23367(new_n25716, new_n14941, n7693);
xnor_3 g23368(new_n25717, new_n25710, new_n25716);
nor_4  g23369(new_n25718, new_n25717, new_n25715);
nor_4  g23370(new_n25719_1, new_n25718, new_n25712);
not_3  g23371(new_n25720, new_n25719_1);
nand_4 g23372(new_n25721, new_n24429, new_n11670);
nand_4 g23373(new_n25722, new_n24449, new_n24430);
nand_4 g23374(new_n25723, new_n25722, new_n25721);
xor_3  g23375(n7575, new_n25723, new_n25720);
xnor_3 g23376(new_n25725, new_n25388, new_n11592);
nor_4  g23377(new_n25726, new_n25397, new_n11647_1);
not_3  g23378(new_n25727, new_n25726);
nor_4  g23379(new_n25728, new_n25394, new_n11648);
nor_4  g23380(new_n25729, new_n25728, new_n25726);
not_3  g23381(new_n25730, new_n11653);
nor_4  g23382(new_n25731, new_n25401, new_n25730);
not_3  g23383(new_n25732, new_n25731);
nand_4 g23384(new_n25733, new_n13126, new_n13086);
nand_4 g23385(new_n25734, new_n25733, new_n25732);
nand_4 g23386(new_n25735, new_n25734, new_n25729);
nand_4 g23387(new_n25736, new_n25735, new_n25727);
xnor_3 g23388(new_n25737, new_n25736, new_n25725);
xnor_3 g23389(new_n25738_1, new_n25737, new_n13861);
xnor_3 g23390(new_n25739, new_n25734, new_n25729);
nor_4  g23391(new_n25740, new_n25739, new_n13869);
xnor_3 g23392(new_n25741, new_n25739, new_n13869);
not_3  g23393(new_n25742, new_n13127);
nor_4  g23394(new_n25743, new_n13138, new_n25742);
not_3  g23395(new_n25744, new_n25743);
nand_4 g23396(new_n25745, new_n13196, new_n13139);
nand_4 g23397(new_n25746, new_n25745, new_n25744);
nor_4  g23398(new_n25747, new_n25746, new_n25741);
nor_4  g23399(new_n25748, new_n25747, new_n25740);
xor_3  g23400(n7585, new_n25748, new_n25738_1);
xnor_3 g23401(new_n25750, new_n25037, new_n9129_1);
nor_4  g23402(new_n25751_1, new_n25041, new_n9139);
not_3  g23403(new_n25752, new_n25751_1);
nor_4  g23404(new_n25753, new_n25042, new_n9144);
nor_4  g23405(new_n25754, new_n25753, new_n25751_1);
nor_4  g23406(new_n25755, new_n25047, new_n9149);
not_3  g23407(new_n25756_1, new_n25755);
nor_4  g23408(new_n25757, new_n25051, new_n9154);
nor_4  g23409(new_n25758_1, new_n25757, new_n25755);
nor_4  g23410(new_n25759, new_n25058, new_n9159);
not_3  g23411(new_n25760, new_n25759);
nor_4  g23412(new_n25761, new_n25056, new_n9164_1);
nor_4  g23413(new_n25762, new_n25761, new_n25759);
nor_4  g23414(new_n25763, new_n22016_1, new_n9177);
not_3  g23415(new_n25764, new_n25763);
nor_4  g23416(new_n25765, new_n22015, new_n9176);
nor_4  g23417(new_n25766, new_n25765, new_n25763);
not_3  g23418(new_n25767, new_n22019);
nor_4  g23419(new_n25768, new_n25767, new_n9186);
not_3  g23420(new_n25769, new_n25768);
nor_4  g23421(new_n25770, new_n22019, new_n9185);
nor_4  g23422(new_n25771, new_n25770, new_n25768);
nor_4  g23423(new_n25772, new_n22023, new_n9195);
not_3  g23424(new_n25773_1, new_n25772);
not_3  g23425(new_n25774, new_n22023);
nor_4  g23426(new_n25775, new_n25774, new_n9194);
nor_4  g23427(new_n25776, new_n25775, new_n25772);
nand_4 g23428(new_n25777, new_n22035, new_n9204);
xnor_3 g23429(new_n25778, new_n22030, new_n9204);
nor_4  g23430(new_n25779, new_n22039, new_n9218);
nor_4  g23431(new_n25780, new_n25779, new_n9212);
not_3  g23432(new_n25781, new_n25780);
not_3  g23433(new_n25782, new_n22046);
not_3  g23434(new_n25783, new_n25779);
xor_3  g23435(new_n25784_1, new_n25783, new_n9213);
nand_4 g23436(new_n25785, new_n25784_1, new_n25782);
nand_4 g23437(new_n25786, new_n25785, new_n25781);
nand_4 g23438(new_n25787, new_n25786, new_n25778);
nand_4 g23439(new_n25788, new_n25787, new_n25777);
nand_4 g23440(new_n25789, new_n25788, new_n25776);
nand_4 g23441(new_n25790, new_n25789, new_n25773_1);
nand_4 g23442(new_n25791, new_n25790, new_n25771);
nand_4 g23443(new_n25792_1, new_n25791, new_n25769);
nand_4 g23444(new_n25793, new_n25792_1, new_n25766);
nand_4 g23445(new_n25794, new_n25793, new_n25764);
nand_4 g23446(new_n25795, new_n25794, new_n25762);
nand_4 g23447(new_n25796, new_n25795, new_n25760);
nand_4 g23448(new_n25797_1, new_n25796, new_n25758_1);
nand_4 g23449(new_n25798, new_n25797_1, new_n25756_1);
nand_4 g23450(new_n25799, new_n25798, new_n25754);
nand_4 g23451(new_n25800, new_n25799, new_n25752);
xnor_3 g23452(n7588, new_n25800, new_n25750);
nor_4  g23453(new_n25802, new_n17492, new_n17390);
nor_4  g23454(new_n25803, new_n25802, new_n17385);
nor_4  g23455(new_n25804, new_n24246, new_n25803);
not_3  g23456(new_n25805, new_n7853);
nor_4  g23457(new_n25806, new_n25805, n21832);
not_3  g23458(new_n25807, new_n25806);
nor_4  g23459(new_n25808, new_n25807, n21753);
not_3  g23460(new_n25809, new_n25808);
nor_4  g23461(new_n25810, new_n25809, n10739);
not_3  g23462(new_n25811, new_n25810);
nor_4  g23463(new_n25812, new_n25811, n13074);
xor_3  g23464(new_n25813, new_n25812, new_n13462);
not_3  g23465(new_n25814, new_n25813);
xor_3  g23466(new_n25815, new_n25814, new_n19420);
not_3  g23467(new_n25816_1, new_n25815);
xor_3  g23468(new_n25817, new_n25811, n13074);
nor_4  g23469(new_n25818, new_n25817, n11455);
not_3  g23470(new_n25819, new_n25817);
xor_3  g23471(new_n25820, new_n25819, new_n19425);
not_3  g23472(new_n25821, new_n25820);
xor_3  g23473(new_n25822, new_n25808, new_n13467);
nor_4  g23474(new_n25823, new_n25822, n3945);
not_3  g23475(new_n25824, new_n25822);
xor_3  g23476(new_n25825, new_n25824, new_n19429);
not_3  g23477(new_n25826_1, new_n25825);
xor_3  g23478(new_n25827, new_n25806, new_n2354);
nor_4  g23479(new_n25828, new_n25827, n5255);
xor_3  g23480(new_n25829, new_n25806, n21753);
nor_4  g23481(new_n25830, new_n25829, new_n19433);
nor_4  g23482(new_n25831, new_n25830, new_n25828);
not_3  g23483(new_n25832, new_n25831);
xor_3  g23484(new_n25833, new_n7853, new_n2356);
nor_4  g23485(new_n25834, new_n25833, n21649);
nor_4  g23486(new_n25835, new_n7854, new_n5941);
nor_4  g23487(new_n25836, new_n25835, new_n25834);
nand_4 g23488(new_n25837, new_n7877, new_n5945);
nand_4 g23489(new_n25838, new_n7895, new_n5818);
xor_3  g23490(new_n25839_1, new_n7896, n3828);
nand_4 g23491(new_n25840_1, new_n7889, new_n5795);
nand_4 g23492(new_n25841, n21654, n2387);
xor_3  g23493(new_n25842, new_n7889, new_n5795);
nand_4 g23494(new_n25843, new_n25842, new_n25841);
nand_4 g23495(new_n25844, new_n25843, new_n25840_1);
nand_4 g23496(new_n25845, new_n25844, new_n25839_1);
nand_4 g23497(new_n25846, new_n25845, new_n25838);
nor_4  g23498(new_n25847, new_n7872, n18274);
nor_4  g23499(new_n25848, new_n7877, new_n5945);
nor_4  g23500(new_n25849, new_n25848, new_n25847);
nand_4 g23501(new_n25850, new_n25849, new_n25846);
nand_4 g23502(new_n25851, new_n25850, new_n25837);
nand_4 g23503(new_n25852, new_n25851, new_n25836);
not_3  g23504(new_n25853, new_n25852);
nor_4  g23505(new_n25854, new_n25853, new_n25834);
nor_4  g23506(new_n25855, new_n25854, new_n25832);
nor_4  g23507(new_n25856, new_n25855, new_n25828);
nor_4  g23508(new_n25857, new_n25856, new_n25826_1);
nor_4  g23509(new_n25858, new_n25857, new_n25823);
nor_4  g23510(new_n25859, new_n25858, new_n25821);
nor_4  g23511(new_n25860, new_n25859, new_n25818);
xnor_3 g23512(new_n25861, new_n25860, new_n25816_1);
xnor_3 g23513(new_n25862, new_n25861, new_n25804);
xnor_3 g23514(new_n25863, new_n25858, new_n25821);
nor_4  g23515(new_n25864, new_n25863, new_n17494);
xnor_3 g23516(new_n25865, new_n25863, new_n17494);
not_3  g23517(new_n25866, new_n25856);
nor_4  g23518(new_n25867, new_n25866, new_n25825);
nor_4  g23519(new_n25868, new_n25867, new_n25857);
not_3  g23520(new_n25869, new_n25868);
nand_4 g23521(new_n25870, new_n25869, new_n17504);
xnor_3 g23522(new_n25871, new_n25868, new_n17504);
xnor_3 g23523(new_n25872_1, new_n25854, new_n25832);
nand_4 g23524(new_n25873_1, new_n25872_1, new_n17508);
xnor_3 g23525(new_n25874, new_n25851, new_n25836);
nand_4 g23526(new_n25875, new_n25874, new_n17515);
xnor_3 g23527(new_n25876, new_n25849, new_n25846);
nand_4 g23528(new_n25877_1, new_n25876, new_n17522);
xnor_3 g23529(new_n25878, new_n25876, new_n17519);
not_3  g23530(new_n25879, new_n25839_1);
xnor_3 g23531(new_n25880, new_n25844, new_n25879);
nor_4  g23532(new_n25881, new_n25880, new_n17532);
not_3  g23533(new_n25882, new_n25881);
not_3  g23534(new_n25883, new_n25880);
nor_4  g23535(new_n25884, new_n25883, new_n17531);
nor_4  g23536(new_n25885, new_n25884, new_n25881);
nor_4  g23537(new_n25886, new_n25842, new_n17538);
not_3  g23538(new_n25887, new_n25841);
xnor_3 g23539(new_n25888, new_n25842, new_n25887);
nor_4  g23540(new_n25889, new_n25888, new_n17537);
xor_3  g23541(new_n25890, n21654, new_n2571);
nor_4  g23542(new_n25891, new_n25890, new_n17546);
nor_4  g23543(new_n25892, new_n25891, new_n25889);
nor_4  g23544(new_n25893, new_n25892, new_n25886);
nand_4 g23545(new_n25894, new_n25893, new_n25885);
nand_4 g23546(new_n25895, new_n25894, new_n25882);
nand_4 g23547(new_n25896, new_n25895, new_n25878);
nand_4 g23548(new_n25897, new_n25896, new_n25877_1);
xnor_3 g23549(new_n25898, new_n25874, new_n17514);
nand_4 g23550(new_n25899, new_n25898, new_n25897);
nand_4 g23551(new_n25900, new_n25899, new_n25875);
not_3  g23552(new_n25901, new_n17508);
xnor_3 g23553(new_n25902, new_n25872_1, new_n25901);
nand_4 g23554(new_n25903, new_n25902, new_n25900);
nand_4 g23555(new_n25904, new_n25903, new_n25873_1);
nand_4 g23556(new_n25905, new_n25904, new_n25871);
nand_4 g23557(new_n25906, new_n25905, new_n25870);
nor_4  g23558(new_n25907, new_n25906, new_n25865);
nor_4  g23559(new_n25908, new_n25907, new_n25864);
xor_3  g23560(n7598, new_n25908, new_n25862);
xnor_3 g23561(n7607, new_n21909, new_n21906);
not_3  g23562(new_n25911, new_n5698);
xor_3  g23563(n7610, new_n5736, new_n25911);
not_3  g23564(new_n25913, new_n3626);
xor_3  g23565(n7616, new_n25913, new_n3611);
not_3  g23566(new_n25915, new_n19051);
xor_3  g23567(new_n25916, n10514, n6105);
not_3  g23568(new_n25917, new_n25916);
nand_4 g23569(new_n25918, new_n25387, new_n7393);
xor_3  g23570(new_n25919, n18649, n3795);
nand_4 g23571(new_n25920, new_n14823, new_n25393);
xor_3  g23572(new_n25921, n25464, n6218);
nand_4 g23573(new_n25922, new_n13724, new_n14827_1);
xor_3  g23574(new_n25923_1, n20470, n4590);
nand_4 g23575(new_n25924, new_n14831, new_n25403);
xor_3  g23576(new_n25925, n26752, n21222);
nor_4  g23577(new_n25926_1, n9832, n6513);
not_3  g23578(new_n25927, new_n25926_1);
xor_3  g23579(new_n25928, n9832, n6513);
nand_4 g23580(new_n25929, n3918, n1558);
not_3  g23581(new_n25930, new_n25929);
nor_4  g23582(new_n25931, n3918, n1558);
nor_4  g23583(new_n25932, n21749, n919);
not_3  g23584(new_n25933, new_n25932);
nand_4 g23585(new_n25934_1, new_n20093, new_n25933);
nor_4  g23586(new_n25935, new_n25934_1, new_n25931);
nor_4  g23587(new_n25936, new_n25935, new_n25930);
nand_4 g23588(new_n25937, new_n25936, new_n25928);
nand_4 g23589(new_n25938_1, new_n25937, new_n25927);
nand_4 g23590(new_n25939, new_n25938_1, new_n25925);
nand_4 g23591(new_n25940, new_n25939, new_n25924);
nand_4 g23592(new_n25941, new_n25940, new_n25923_1);
nand_4 g23593(new_n25942, new_n25941, new_n25922);
nand_4 g23594(new_n25943, new_n25942, new_n25921);
nand_4 g23595(new_n25944, new_n25943, new_n25920);
nand_4 g23596(new_n25945, new_n25944, new_n25919);
nand_4 g23597(new_n25946, new_n25945, new_n25918);
not_3  g23598(new_n25947, new_n25946);
xor_3  g23599(new_n25948, new_n25947, new_n25917);
nand_4 g23600(new_n25949, new_n25948, n9872);
not_3  g23601(new_n25950, new_n25949);
xnor_3 g23602(new_n25951, new_n25948, n9872);
xnor_3 g23603(new_n25952, new_n25944, new_n25919);
nor_4  g23604(new_n25953, new_n25952, new_n25458);
not_3  g23605(new_n25954, new_n25952);
xor_3  g23606(new_n25955, new_n25954, n5842);
xnor_3 g23607(new_n25956, new_n25942, new_n25921);
not_3  g23608(new_n25957, new_n25956);
nand_4 g23609(new_n25958, new_n25957, n6379);
xor_3  g23610(new_n25959, new_n25957, n6379);
xnor_3 g23611(new_n25960, new_n25940, new_n25923_1);
not_3  g23612(new_n25961, new_n25960);
nand_4 g23613(new_n25962, new_n25961, n2102);
xor_3  g23614(new_n25963, new_n25961, n2102);
not_3  g23615(new_n25964, new_n25925);
xnor_3 g23616(new_n25965, new_n25938_1, new_n25964);
nand_4 g23617(new_n25966, new_n25965, n17954);
xnor_3 g23618(new_n25967, new_n25965, new_n25502);
not_3  g23619(new_n25968, new_n25928);
xnor_3 g23620(new_n25969, new_n25936, new_n25968);
nand_4 g23621(new_n25970, new_n25969, n8256);
xnor_3 g23622(new_n25971, new_n25969, new_n25477);
not_3  g23623(new_n25972_1, new_n25934_1);
nor_4  g23624(new_n25973, new_n25931, new_n25930);
xnor_3 g23625(new_n25974_1, new_n25973, new_n25972_1);
nand_4 g23626(new_n25975, new_n25974_1, n24150);
xnor_3 g23627(new_n25976, new_n25974_1, new_n25481);
nand_4 g23628(new_n25977, new_n20095, n19584);
nand_4 g23629(new_n25978, new_n20105, new_n20096_1);
nand_4 g23630(new_n25979, new_n25978, new_n25977);
nand_4 g23631(new_n25980, new_n25979, new_n25976);
nand_4 g23632(new_n25981, new_n25980, new_n25975);
nand_4 g23633(new_n25982, new_n25981, new_n25971);
nand_4 g23634(new_n25983, new_n25982, new_n25970);
nand_4 g23635(new_n25984, new_n25983, new_n25967);
nand_4 g23636(new_n25985_1, new_n25984, new_n25966);
nand_4 g23637(new_n25986, new_n25985_1, new_n25963);
nand_4 g23638(new_n25987, new_n25986, new_n25962);
nand_4 g23639(new_n25988, new_n25987, new_n25959);
nand_4 g23640(new_n25989, new_n25988, new_n25958);
nand_4 g23641(new_n25990, new_n25989, new_n25955);
not_3  g23642(new_n25991, new_n25990);
nor_4  g23643(new_n25992, new_n25991, new_n25953);
nor_4  g23644(new_n25993, new_n25992, new_n25951);
nor_4  g23645(new_n25994_1, new_n25993, new_n25950);
nor_4  g23646(new_n25995, n10514, n6105);
nor_4  g23647(new_n25996, new_n25947, new_n25917);
nor_4  g23648(new_n25997, new_n25996, new_n25995);
nor_4  g23649(new_n25998, new_n25997, new_n25994_1);
xnor_3 g23650(new_n25999, new_n25998, new_n25915);
xnor_3 g23651(new_n26000, new_n25997, new_n25994_1);
nor_4  g23652(new_n26001, new_n26000, new_n18965);
not_3  g23653(new_n26002, new_n26001);
xnor_3 g23654(new_n26003, new_n26000, new_n18965);
not_3  g23655(new_n26004, new_n26003);
xnor_3 g23656(new_n26005, new_n25992, new_n25951);
nor_4  g23657(new_n26006, new_n26005, new_n18970_1);
not_3  g23658(new_n26007, new_n26006);
xnor_3 g23659(new_n26008, new_n26005, new_n18970_1);
not_3  g23660(new_n26009, new_n26008);
xnor_3 g23661(new_n26010, new_n25989, new_n25955);
nor_4  g23662(new_n26011, new_n26010, new_n18977_1);
not_3  g23663(new_n26012, new_n26011);
xnor_3 g23664(new_n26013, new_n26010, new_n18977_1);
not_3  g23665(new_n26014, new_n26013);
xnor_3 g23666(new_n26015, new_n25987, new_n25959);
nor_4  g23667(new_n26016, new_n26015, new_n18983);
not_3  g23668(new_n26017, new_n26016);
xnor_3 g23669(new_n26018, new_n26015, new_n18982_1);
xnor_3 g23670(new_n26019, new_n25985_1, new_n25963);
not_3  g23671(new_n26020, new_n26019);
nand_4 g23672(new_n26021, new_n26020, new_n18991);
xnor_3 g23673(new_n26022, new_n26019, new_n18991);
xnor_3 g23674(new_n26023, new_n25983, new_n25967);
not_3  g23675(new_n26024, new_n26023);
nand_4 g23676(new_n26025, new_n26024, new_n18996);
xnor_3 g23677(new_n26026, new_n26023, new_n18996);
xnor_3 g23678(new_n26027, new_n25981, new_n25971);
not_3  g23679(new_n26028, new_n26027);
nand_4 g23680(new_n26029, new_n26028, new_n19001);
xnor_3 g23681(new_n26030, new_n26027, new_n19001);
not_3  g23682(new_n26031, new_n25976);
xnor_3 g23683(new_n26032, new_n25979, new_n26031);
nand_4 g23684(new_n26033, new_n26032, new_n19007);
xnor_3 g23685(new_n26034, new_n26032, new_n19006);
not_3  g23686(new_n26035, new_n20106);
nand_4 g23687(new_n26036_1, new_n26035, new_n19012);
nand_4 g23688(new_n26037, new_n20116, new_n20107);
nand_4 g23689(new_n26038, new_n26037, new_n26036_1);
nand_4 g23690(new_n26039, new_n26038, new_n26034);
nand_4 g23691(new_n26040, new_n26039, new_n26033);
nand_4 g23692(new_n26041, new_n26040, new_n26030);
nand_4 g23693(new_n26042, new_n26041, new_n26029);
nand_4 g23694(new_n26043, new_n26042, new_n26026);
nand_4 g23695(new_n26044, new_n26043, new_n26025);
nand_4 g23696(new_n26045, new_n26044, new_n26022);
nand_4 g23697(new_n26046, new_n26045, new_n26021);
nand_4 g23698(new_n26047, new_n26046, new_n26018);
nand_4 g23699(new_n26048, new_n26047, new_n26017);
nand_4 g23700(new_n26049, new_n26048, new_n26014);
nand_4 g23701(new_n26050, new_n26049, new_n26012);
nand_4 g23702(new_n26051, new_n26050, new_n26009);
nand_4 g23703(new_n26052, new_n26051, new_n26007);
nand_4 g23704(new_n26053_1, new_n26052, new_n26004);
nand_4 g23705(new_n26054_1, new_n26053_1, new_n26002);
xnor_3 g23706(n7630, new_n26054_1, new_n25999);
nor_4  g23707(new_n26056, new_n22967, new_n22937);
nor_4  g23708(new_n26057, new_n22977, new_n22968);
nor_4  g23709(n7643, new_n26057, new_n26056);
not_3  g23710(new_n26059, new_n14641);
xor_3  g23711(n7647, new_n14679, new_n26059);
xnor_3 g23712(n7679, new_n12081, new_n12047);
not_3  g23713(new_n26062, new_n24625);
xor_3  g23714(n7686, new_n24660, new_n26062);
nor_4  g23715(new_n26064, new_n22367, new_n22346);
xnor_3 g23716(n7698, new_n26064, new_n22364);
xnor_3 g23717(n7708, new_n23727, new_n23706);
xor_3  g23718(new_n26067, new_n22335_1, new_n19353);
nor_4  g23719(new_n26068, new_n3074, new_n19385_1);
xor_3  g23720(new_n26069, new_n3074, n17911);
nor_4  g23721(new_n26070, new_n3121, n21997);
not_3  g23722(new_n26071, new_n26070);
xor_3  g23723(new_n26072, new_n3122, new_n19389_1);
nor_4  g23724(new_n26073, new_n3127, n25119);
not_3  g23725(new_n26074, new_n26073);
nand_4 g23726(new_n26075, new_n10168, new_n26074);
nand_4 g23727(new_n26076, new_n26075, new_n26072);
nand_4 g23728(new_n26077, new_n26076, new_n26071);
nor_4  g23729(new_n26078, new_n26077, new_n26069);
nor_4  g23730(new_n26079, new_n26078, new_n26068);
nand_4 g23731(new_n26080, new_n26079, new_n26067);
not_3  g23732(new_n26081, new_n26080);
nor_4  g23733(new_n26082, new_n26079, new_n26067);
nor_4  g23734(new_n26083, new_n26082, new_n26081);
xnor_3 g23735(new_n26084_1, new_n7068, new_n21148);
not_3  g23736(new_n26085, new_n26084_1);
nor_4  g23737(new_n26086, new_n7072, new_n17338);
not_3  g23738(new_n26087, new_n19791);
nor_4  g23739(new_n26088, new_n19799, new_n26087);
nor_4  g23740(new_n26089, new_n26088, new_n26086);
xnor_3 g23741(new_n26090, new_n26089, new_n26085);
not_3  g23742(new_n26091, new_n26090);
xnor_3 g23743(new_n26092, new_n26091, new_n26083);
xnor_3 g23744(new_n26093, new_n26077, new_n26069);
nand_4 g23745(new_n26094, new_n26093, new_n19800);
not_3  g23746(new_n26095, new_n19800);
xnor_3 g23747(new_n26096_1, new_n26093, new_n26095);
not_3  g23748(new_n26097, new_n19802);
not_3  g23749(new_n26098, new_n26076);
nor_4  g23750(new_n26099, new_n26075, new_n26072);
nor_4  g23751(new_n26100, new_n26099, new_n26098);
nand_4 g23752(new_n26101, new_n26100, new_n26097);
xnor_3 g23753(new_n26102, new_n26100, new_n19802);
nand_4 g23754(new_n26103, new_n10171, new_n10135);
nand_4 g23755(new_n26104, new_n10224, new_n10172);
nand_4 g23756(new_n26105, new_n26104, new_n26103);
nand_4 g23757(new_n26106, new_n26105, new_n26102);
nand_4 g23758(new_n26107_1, new_n26106, new_n26101);
nand_4 g23759(new_n26108, new_n26107_1, new_n26096_1);
nand_4 g23760(new_n26109, new_n26108, new_n26094);
xnor_3 g23761(n7780, new_n26109, new_n26092);
nor_4  g23762(new_n26111_1, new_n2666, new_n5035);
xnor_3 g23763(new_n26112, new_n2666, new_n5035);
nor_4  g23764(new_n26113_1, new_n2672, new_n5007);
nor_4  g23765(new_n26114, new_n11591_1, new_n11550);
nor_4  g23766(new_n26115, new_n26114, new_n26113_1);
nor_4  g23767(new_n26116, new_n26115, new_n26112);
nor_4  g23768(new_n26117, new_n26116, new_n26111_1);
xnor_3 g23769(new_n26118, new_n26117, new_n17814);
nor_4  g23770(new_n26119, new_n21163, new_n2819);
nor_4  g23771(new_n26120, new_n21162, new_n2821);
nor_4  g23772(new_n26121, new_n26120, new_n26119);
not_3  g23773(new_n26122, new_n26121);
nor_4  g23774(new_n26123, new_n11600, new_n12169);
not_3  g23775(new_n26124, new_n11601);
nor_4  g23776(new_n26125, new_n11644, new_n26124);
nor_4  g23777(new_n26126, new_n26125, new_n26123);
nor_4  g23778(new_n26127, new_n26126, new_n26122);
nor_4  g23779(new_n26128, new_n26127, new_n26119);
not_3  g23780(new_n26129, new_n21161);
nor_4  g23781(new_n26130, new_n26129, n21839);
nand_4 g23782(new_n26131, new_n26130, new_n19243);
not_3  g23783(new_n26132, new_n26130);
nand_4 g23784(new_n26133, new_n26132, new_n12164);
nand_4 g23785(new_n26134, new_n26133, new_n26131);
xnor_3 g23786(new_n26135, new_n26134, new_n26128);
xnor_3 g23787(new_n26136, new_n26135, new_n26118);
not_3  g23788(new_n26137, new_n26115);
xnor_3 g23789(new_n26138, new_n26137, new_n26112);
xnor_3 g23790(new_n26139, new_n26126, new_n26121);
nor_4  g23791(new_n26140, new_n26139, new_n26138);
xnor_3 g23792(new_n26141, new_n26139, new_n26138);
nor_4  g23793(new_n26142, new_n11645, new_n11593);
nor_4  g23794(new_n26143, new_n11710_1, new_n11646);
nor_4  g23795(new_n26144, new_n26143, new_n26142);
nor_4  g23796(new_n26145, new_n26144, new_n26141);
nor_4  g23797(new_n26146, new_n26145, new_n26140);
xnor_3 g23798(n7794, new_n26146, new_n26136);
not_3  g23799(new_n26148, new_n21375);
xor_3  g23800(n7811, new_n26148, new_n21367_1);
xor_3  g23801(n7830, new_n21311, new_n21304);
not_3  g23802(new_n26151, new_n25796);
xor_3  g23803(n7834, new_n26151, new_n25758_1);
not_3  g23804(new_n26153, new_n13190_1);
xor_3  g23805(n7884, new_n26153, new_n13171);
xor_3  g23806(n7937, new_n3248, new_n3244_1);
xnor_3 g23807(n7943, new_n3260_1, new_n3195);
xor_3  g23808(n7950, new_n11704, new_n11662);
xnor_3 g23809(new_n26158, new_n24038, new_n25351);
xnor_3 g23810(new_n26159_1, new_n24012, new_n24002_1);
nor_4  g23811(new_n26160, new_n26159_1, new_n18905);
not_3  g23812(new_n26161, new_n26160);
nor_4  g23813(new_n26162, new_n24046, new_n18911);
not_3  g23814(new_n26163, new_n26162);
nor_4  g23815(new_n26164, new_n24050, new_n18909);
nor_4  g23816(new_n26165, new_n26164, new_n26162);
not_3  g23817(new_n26166, new_n18553);
nand_4 g23818(new_n26167_1, new_n18607, new_n18554);
nand_4 g23819(new_n26168, new_n26167_1, new_n26166);
nand_4 g23820(new_n26169, new_n26168, new_n26165);
nand_4 g23821(new_n26170, new_n26169, new_n26163);
nor_4  g23822(new_n26171, new_n24044, new_n18902);
nor_4  g23823(new_n26172, new_n26171, new_n26160);
nand_4 g23824(new_n26173, new_n26172, new_n26170);
nand_4 g23825(new_n26174, new_n26173, new_n26161);
nor_4  g23826(new_n26175, new_n26174, new_n26158);
nor_4  g23827(new_n26176, new_n24038, new_n25351);
nor_4  g23828(new_n26177, new_n24035, new_n18964);
nor_4  g23829(new_n26178, new_n26177, new_n26176);
not_3  g23830(new_n26179_1, new_n26170);
xnor_3 g23831(new_n26180_1, new_n24044, new_n18902);
nor_4  g23832(new_n26181, new_n26180_1, new_n26179_1);
nor_4  g23833(new_n26182, new_n26181, new_n26160);
nor_4  g23834(new_n26183, new_n26182, new_n26178);
nor_4  g23835(n7959, new_n26183, new_n26175);
not_3  g23836(new_n26185, new_n21379);
xor_3  g23837(n7968, new_n26185, new_n21359);
xor_3  g23838(n7992, new_n22644, new_n22640);
xor_3  g23839(new_n26188, new_n15536, new_n9258);
nor_4  g23840(new_n26189, new_n15545, new_n21228);
not_3  g23841(new_n26190, new_n26189);
nor_4  g23842(new_n26191_1, new_n15544, n26408);
nor_4  g23843(new_n26192, new_n26191_1, new_n26189);
nand_4 g23844(new_n26193, new_n12688, n18227);
nand_4 g23845(new_n26194, new_n21343, new_n21331);
nand_4 g23846(new_n26195, new_n26194, new_n26193);
nand_4 g23847(new_n26196, new_n26195, new_n26192);
nand_4 g23848(new_n26197, new_n26196, new_n26190);
nand_4 g23849(new_n26198, new_n26197, new_n26188);
not_3  g23850(new_n26199, new_n26198);
nor_4  g23851(new_n26200, new_n26197, new_n26188);
nor_4  g23852(new_n26201, new_n26200, new_n26199);
xnor_3 g23853(new_n26202, new_n26201, new_n22847);
not_3  g23854(new_n26203, new_n26196);
nor_4  g23855(new_n26204, new_n26195, new_n26192);
nor_4  g23856(new_n26205, new_n26204, new_n26203);
nand_4 g23857(new_n26206, new_n26205, new_n22860);
xnor_3 g23858(new_n26207, new_n26205, new_n22855);
nand_4 g23859(new_n26208, new_n22867, new_n21344);
xnor_3 g23860(new_n26209, new_n22862, new_n21344);
nand_4 g23861(new_n26210, new_n22874, new_n21347);
xnor_3 g23862(new_n26211, new_n22869, new_n21347);
nand_4 g23863(new_n26212, new_n22881, new_n21351);
xnor_3 g23864(new_n26213, new_n22878, new_n21351);
nand_4 g23865(new_n26214, new_n22887, new_n15654);
nand_4 g23866(new_n26215, new_n15680, new_n15667);
nand_4 g23867(new_n26216, new_n26215, new_n26214);
nand_4 g23868(new_n26217, new_n26216, new_n26213);
nand_4 g23869(new_n26218, new_n26217, new_n26212);
nand_4 g23870(new_n26219, new_n26218, new_n26211);
nand_4 g23871(new_n26220_1, new_n26219, new_n26210);
nand_4 g23872(new_n26221, new_n26220_1, new_n26209);
nand_4 g23873(new_n26222, new_n26221, new_n26208);
nand_4 g23874(new_n26223, new_n26222, new_n26207);
nand_4 g23875(new_n26224_1, new_n26223, new_n26206);
xnor_3 g23876(n7999, new_n26224_1, new_n26202);
not_3  g23877(new_n26226, new_n22177);
xor_3  g23878(n8027, new_n22197, new_n26226);
nor_4  g23879(new_n26228, new_n26117, new_n17815);
nor_4  g23880(new_n26229_1, new_n7307, new_n6321);
not_3  g23881(new_n26230, new_n26229_1);
nor_4  g23882(new_n26231, new_n7308_1, n8614);
nor_4  g23883(new_n26232, new_n26231, new_n26229_1);
nor_4  g23884(new_n26233, new_n14927, new_n6326);
not_3  g23885(new_n26234, new_n26233);
nor_4  g23886(new_n26235, new_n7318, n27037);
xnor_3 g23887(new_n26236, new_n14932, new_n6328);
nor_4  g23888(new_n26237_1, new_n7374, n8964);
xnor_3 g23889(new_n26238, new_n7374, n8964);
nor_4  g23890(new_n26239, new_n7330_1, new_n7279);
not_3  g23891(new_n26240, new_n26239);
not_3  g23892(new_n26241, new_n25706_1);
nand_4 g23893(new_n26242, new_n25710, new_n25708);
nand_4 g23894(new_n26243, new_n26242, new_n26241);
nor_4  g23895(new_n26244, new_n7332, n20151);
nor_4  g23896(new_n26245, new_n26244, new_n26239);
nand_4 g23897(new_n26246, new_n26245, new_n26243);
nand_4 g23898(new_n26247, new_n26246, new_n26240);
nor_4  g23899(new_n26248, new_n26247, new_n26238);
nor_4  g23900(new_n26249, new_n26248, new_n26237_1);
nor_4  g23901(new_n26250_1, new_n26249, new_n26236);
nor_4  g23902(new_n26251, new_n26250_1, new_n26235);
nor_4  g23903(new_n26252, new_n7314, n15182);
nor_4  g23904(new_n26253, new_n26252, new_n26233);
nand_4 g23905(new_n26254, new_n26253, new_n26251);
nand_4 g23906(new_n26255, new_n26254, new_n26234);
nand_4 g23907(new_n26256, new_n26255, new_n26232);
nand_4 g23908(new_n26257, new_n26256, new_n26230);
nand_4 g23909(new_n26258, new_n26257, new_n7248);
nand_4 g23910(new_n26259, new_n26258, new_n26228);
xnor_3 g23911(new_n26260, new_n26257, new_n7248);
nand_4 g23912(new_n26261, new_n26260, new_n26118);
not_3  g23913(new_n26262, new_n26118);
xnor_3 g23914(new_n26263, new_n26260, new_n26262);
xnor_3 g23915(new_n26264_1, new_n26255, new_n26232);
nand_4 g23916(new_n26265, new_n26264_1, new_n26138);
not_3  g23917(new_n26266, new_n26138);
xnor_3 g23918(new_n26267, new_n26264_1, new_n26266);
xnor_3 g23919(new_n26268, new_n26253, new_n26251);
nand_4 g23920(new_n26269, new_n26268, new_n11593);
xnor_3 g23921(new_n26270, new_n26268, new_n11592);
not_3  g23922(new_n26271, new_n26236);
xnor_3 g23923(new_n26272, new_n26249, new_n26271);
nand_4 g23924(new_n26273, new_n26272, new_n11648);
xnor_3 g23925(new_n26274_1, new_n26272, new_n11647_1);
not_3  g23926(new_n26275, new_n26238);
xnor_3 g23927(new_n26276, new_n26247, new_n26275);
nand_4 g23928(new_n26277, new_n26276, new_n11653);
xnor_3 g23929(new_n26278, new_n26276, new_n25730);
xnor_3 g23930(new_n26279, new_n26245, new_n26243);
nand_4 g23931(new_n26280, new_n26279, new_n11659);
xnor_3 g23932(new_n26281, new_n26279, new_n11658);
not_3  g23933(new_n26282, new_n25718);
nand_4 g23934(new_n26283, new_n25723, new_n25719_1);
nand_4 g23935(new_n26284, new_n26283, new_n26282);
nand_4 g23936(new_n26285, new_n26284, new_n26281);
nand_4 g23937(new_n26286, new_n26285, new_n26280);
nand_4 g23938(new_n26287_1, new_n26286, new_n26278);
nand_4 g23939(new_n26288, new_n26287_1, new_n26277);
nand_4 g23940(new_n26289, new_n26288, new_n26274_1);
nand_4 g23941(new_n26290, new_n26289, new_n26273);
nand_4 g23942(new_n26291, new_n26290, new_n26270);
nand_4 g23943(new_n26292, new_n26291, new_n26269);
nand_4 g23944(new_n26293, new_n26292, new_n26267);
nand_4 g23945(new_n26294, new_n26293, new_n26265);
nand_4 g23946(new_n26295, new_n26294, new_n26263);
nand_4 g23947(new_n26296, new_n26295, new_n26261);
not_3  g23948(new_n26297, new_n26228);
xnor_3 g23949(new_n26298, new_n26258, new_n26297);
nand_4 g23950(new_n26299, new_n26298, new_n26296);
nand_4 g23951(n8031, new_n26299, new_n26259);
not_3  g23952(new_n26301, new_n21164);
nor_4  g23953(new_n26302, new_n21174, new_n21165);
nor_4  g23954(new_n26303, new_n26302, new_n26130);
nand_4 g23955(new_n26304, new_n26303, new_n26301);
nor_4  g23956(new_n26305, new_n26304, new_n24238);
not_3  g23957(new_n26306, new_n26305);
not_3  g23958(new_n26307, new_n26304);
nor_4  g23959(new_n26308, new_n26307, new_n24239);
nor_4  g23960(new_n26309, new_n26308, new_n26305);
nor_4  g23961(new_n26310, new_n21175, new_n21158);
not_3  g23962(new_n26311, new_n26310);
nand_4 g23963(new_n26312, new_n21209, new_n21176_1);
nand_4 g23964(new_n26313, new_n26312, new_n26311);
nand_4 g23965(new_n26314, new_n26313, new_n26309);
nand_4 g23966(new_n26315, new_n26314, new_n26306);
not_3  g23967(new_n26316, new_n21224);
nand_4 g23968(new_n26317_1, new_n21262, new_n26316);
nand_4 g23969(new_n26318_1, new_n26317_1, new_n24594);
nor_4  g23970(new_n26319, new_n26318_1, new_n21223);
nor_4  g23971(new_n26320, new_n26319, new_n26315);
xnor_3 g23972(new_n26321, new_n26319, new_n26315);
not_3  g23973(new_n26322, new_n26319);
xnor_3 g23974(new_n26323, new_n26313, new_n26309);
not_3  g23975(new_n26324, new_n26323);
nor_4  g23976(new_n26325, new_n26324, new_n26322);
xnor_3 g23977(new_n26326, new_n26323, new_n26319);
not_3  g23978(new_n26327, new_n21210);
nor_4  g23979(new_n26328, new_n21263, new_n26327);
nor_4  g23980(new_n26329, new_n21326, new_n26328);
nor_4  g23981(new_n26330, new_n26329, new_n26326);
nor_4  g23982(new_n26331, new_n26330, new_n26325);
nor_4  g23983(new_n26332, new_n26331, new_n26321);
nor_4  g23984(n8042, new_n26332, new_n26320);
nand_4 g23985(new_n26334, new_n12014, new_n11879);
nand_4 g23986(new_n26335, new_n12093, new_n12016);
nand_4 g23987(n8095, new_n26335, new_n26334);
nor_4  g23988(new_n26337, new_n21211, n4306);
xor_3  g23989(new_n26338, n23166, new_n10868);
not_3  g23990(new_n26339, new_n26338);
nor_4  g23991(new_n26340, new_n10886, n3279);
not_3  g23992(new_n26341, new_n26340);
xor_3  g23993(new_n26342, n10577, new_n10933);
nor_4  g23994(new_n26343, n13914, new_n10890);
not_3  g23995(new_n26344, new_n26343);
xor_3  g23996(new_n26345, n13914, new_n10890);
nor_4  g23997(new_n26346, n14702, new_n10893);
not_3  g23998(new_n26347, new_n26346);
nand_4 g23999(new_n26348, new_n23918, new_n23903_1);
nand_4 g24000(new_n26349, new_n26348, new_n26347);
nand_4 g24001(new_n26350, new_n26349, new_n26345);
nand_4 g24002(new_n26351, new_n26350, new_n26344);
nand_4 g24003(new_n26352, new_n26351, new_n26342);
nand_4 g24004(new_n26353_1, new_n26352, new_n26341);
not_3  g24005(new_n26354, new_n26353_1);
nor_4  g24006(new_n26355, new_n26354, new_n26339);
nor_4  g24007(new_n26356, new_n26355, new_n26337);
not_3  g24008(new_n26357, new_n26356);
xnor_3 g24009(new_n26358, new_n26357, new_n10727);
xor_3  g24010(new_n26359, new_n26354, new_n26339);
nor_4  g24011(new_n26360, new_n26359, new_n10788);
xnor_3 g24012(new_n26361, new_n26359, new_n10788);
not_3  g24013(new_n26362, new_n10792_1);
not_3  g24014(new_n26363, new_n26351);
xor_3  g24015(new_n26364, new_n26363, new_n26342);
nand_4 g24016(new_n26365, new_n26364, new_n26362);
xnor_3 g24017(new_n26366, new_n26364, new_n10792_1);
not_3  g24018(new_n26367, new_n26345);
xor_3  g24019(new_n26368, new_n26349, new_n26367);
nand_4 g24020(new_n26369, new_n26368, new_n10798);
xnor_3 g24021(new_n26370, new_n26368, new_n10799);
nor_4  g24022(new_n26371, new_n23919, new_n10804);
nor_4  g24023(new_n26372, new_n23935_1, new_n23920);
nor_4  g24024(new_n26373, new_n26372, new_n26371);
nand_4 g24025(new_n26374, new_n26373, new_n26370);
nand_4 g24026(new_n26375_1, new_n26374, new_n26369);
nand_4 g24027(new_n26376, new_n26375_1, new_n26366);
nand_4 g24028(new_n26377, new_n26376, new_n26365);
not_3  g24029(new_n26378, new_n26377);
nor_4  g24030(new_n26379, new_n26378, new_n26361);
nor_4  g24031(new_n26380, new_n26379, new_n26360);
xnor_3 g24032(n8103, new_n26380, new_n26358);
xnor_3 g24033(n8109, new_n23131, new_n23118);
nand_4 g24034(new_n26383, new_n24601, new_n23679);
nand_4 g24035(new_n26384, new_n23731, new_n23696);
nand_4 g24036(n8127, new_n26384, new_n26383);
not_3  g24037(new_n26386, new_n20566);
xor_3  g24038(n8130, new_n20572, new_n26386);
nor_4  g24039(new_n26388, n8856, new_n14181);
xor_3  g24040(new_n26389, n8856, new_n14181);
not_3  g24041(new_n26390, new_n26389);
nor_4  g24042(new_n26391, new_n13462, n14130);
xor_3  g24043(new_n26392, n23463, new_n9033);
nand_4 g24044(new_n26393, new_n24704, n13074);
xor_3  g24045(new_n26394, n16482, new_n3335);
nand_4 g24046(new_n26395, n10739, new_n2349);
nand_4 g24047(new_n26396_1, new_n2386, new_n2350);
nand_4 g24048(new_n26397, new_n26396_1, new_n26395);
nand_4 g24049(new_n26398, new_n26397, new_n26394);
nand_4 g24050(new_n26399, new_n26398, new_n26393);
nand_4 g24051(new_n26400, new_n26399, new_n26392);
not_3  g24052(new_n26401, new_n26400);
nor_4  g24053(new_n26402, new_n26401, new_n26391);
nor_4  g24054(new_n26403, new_n26402, new_n26390);
nor_4  g24055(new_n26404, new_n26403, new_n26388);
not_3  g24056(new_n26405, new_n26404);
xnor_3 g24057(new_n26406, new_n26405, new_n8936);
nand_4 g24058(new_n26407, new_n26405, new_n8943_1);
xnor_3 g24059(new_n26408_1, new_n26404, new_n8943_1);
xor_3  g24060(new_n26409, new_n26402, new_n26390);
not_3  g24061(new_n26410, new_n26409);
nand_4 g24062(new_n26411, new_n26410, new_n8952);
not_3  g24063(new_n26412, new_n26411);
nor_4  g24064(new_n26413, new_n26410, new_n8952);
nor_4  g24065(new_n26414, new_n26413, new_n26412);
xor_3  g24066(new_n26415, new_n26399, new_n26392);
nor_4  g24067(new_n26416, new_n26415, new_n8956);
not_3  g24068(new_n26417, new_n26416);
not_3  g24069(new_n26418, new_n26415);
nor_4  g24070(new_n26419, new_n26418, new_n8957);
nor_4  g24071(new_n26420, new_n26419, new_n26416);
not_3  g24072(new_n26421, new_n26394);
xor_3  g24073(new_n26422, new_n26397, new_n26421);
nor_4  g24074(new_n26423, new_n26422, new_n8963);
not_3  g24075(new_n26424, new_n26422);
xnor_3 g24076(new_n26425, new_n26424, new_n8965);
nor_4  g24077(new_n26426, new_n2539, new_n2387_1);
nor_4  g24078(new_n26427, new_n2591, new_n2540);
nor_4  g24079(new_n26428, new_n26427, new_n26426);
nor_4  g24080(new_n26429_1, new_n26428, new_n26425);
nor_4  g24081(new_n26430, new_n26429_1, new_n26423);
nand_4 g24082(new_n26431_1, new_n26430, new_n26420);
nand_4 g24083(new_n26432, new_n26431_1, new_n26417);
nand_4 g24084(new_n26433, new_n26432, new_n26414);
nand_4 g24085(new_n26434, new_n26433, new_n26411);
nand_4 g24086(new_n26435, new_n26434, new_n26408_1);
nand_4 g24087(new_n26436, new_n26435, new_n26407);
xnor_3 g24088(n8135, new_n26436, new_n26406);
xor_3  g24089(n8139, new_n9008, new_n2579);
nand_4 g24090(new_n26439_1, new_n22374, new_n9045);
nor_4  g24091(new_n26440, new_n26439_1, n26660);
xor_3  g24092(new_n26441, new_n26440, new_n8849_1);
xnor_3 g24093(new_n26442, new_n26441, new_n3129);
xor_3  g24094(new_n26443_1, new_n26439_1, n26660);
nand_4 g24095(new_n26444, new_n26443_1, new_n16140);
xnor_3 g24096(new_n26445, new_n26443_1, new_n3134);
nand_4 g24097(new_n26446, new_n22375, new_n16146);
nand_4 g24098(new_n26447, new_n22393, new_n22376);
nand_4 g24099(new_n26448, new_n26447, new_n26446);
nand_4 g24100(new_n26449, new_n26448, new_n26445);
nand_4 g24101(new_n26450, new_n26449, new_n26444);
xnor_3 g24102(new_n26451, new_n26450, new_n26442);
xnor_3 g24103(new_n26452_1, new_n26451, new_n8143);
xnor_3 g24104(new_n26453, new_n26448, new_n26445);
nand_4 g24105(new_n26454, new_n26453, new_n8150);
xnor_3 g24106(new_n26455, new_n26453, new_n8148_1);
nand_4 g24107(new_n26456, new_n22394, new_n8155);
nand_4 g24108(new_n26457, new_n22418, new_n22395);
nand_4 g24109(new_n26458, new_n26457, new_n26456);
nand_4 g24110(new_n26459, new_n26458, new_n26455);
nand_4 g24111(new_n26460, new_n26459, new_n26454);
xnor_3 g24112(n8148, new_n26460, new_n26452_1);
xor_3  g24113(n8149, new_n21602, new_n21601);
not_3  g24114(new_n26463, new_n4302);
xor_3  g24115(n8159, new_n4326_1, new_n26463);
xor_3  g24116(n8179, new_n14128, new_n2609);
not_3  g24117(new_n26466, new_n18137);
xor_3  g24118(n8215, new_n26466, new_n18135);
not_3  g24119(new_n26468, new_n23120_1);
xor_3  g24120(n8267, new_n23129, new_n26468);
not_3  g24121(new_n26470, new_n24442);
xor_3  g24122(n8276, new_n24445, new_n26470);
nand_4 g24123(new_n26472, new_n26440, new_n8849_1);
nor_4  g24124(new_n26473, new_n26472, n1654);
nand_4 g24125(new_n26474, new_n26473, new_n21167);
nor_4  g24126(new_n26475, new_n26474, n22626);
xor_3  g24127(new_n26476, new_n26474, n22626);
not_3  g24128(new_n26477, new_n26476);
nand_4 g24129(new_n26478, new_n26477, new_n18353);
xnor_3 g24130(new_n26479, new_n26477, new_n18350_1);
xor_3  g24131(new_n26480, new_n26473, n14440);
nand_4 g24132(new_n26481, new_n26480, new_n3119);
xnor_3 g24133(new_n26482, new_n26480, new_n18357);
xor_3  g24134(new_n26483_1, new_n26472, n1654);
nand_4 g24135(new_n26484, new_n26483_1, new_n3125_1);
nand_4 g24136(new_n26485, new_n26441, new_n18367);
nand_4 g24137(new_n26486, new_n26450, new_n26442);
nand_4 g24138(new_n26487, new_n26486, new_n26485);
xnor_3 g24139(new_n26488, new_n26483_1, new_n3123);
nand_4 g24140(new_n26489, new_n26488, new_n26487);
nand_4 g24141(new_n26490, new_n26489, new_n26484);
not_3  g24142(new_n26491, new_n26490);
nand_4 g24143(new_n26492_1, new_n26491, new_n26482);
nand_4 g24144(new_n26493, new_n26492_1, new_n26481);
nand_4 g24145(new_n26494, new_n26493, new_n26479);
nand_4 g24146(new_n26495, new_n26494, new_n26478);
nor_4  g24147(new_n26496, new_n26495, new_n18388);
and_4  g24148(new_n26497, new_n26496, new_n26475);
not_3  g24149(new_n26498, new_n26475);
xnor_3 g24150(new_n26499, new_n26495, new_n18388);
xnor_3 g24151(new_n26500, new_n26499, new_n26498);
nor_4  g24152(new_n26501, new_n26500, new_n21049);
not_3  g24153(new_n26502, new_n26501);
xnor_3 g24154(new_n26503, new_n26500, new_n21048);
xnor_3 g24155(new_n26504, new_n26493, new_n26479);
nor_4  g24156(new_n26505, new_n26504, new_n21063);
not_3  g24157(new_n26506, new_n26505);
xnor_3 g24158(new_n26507, new_n26504, new_n21063);
not_3  g24159(new_n26508, new_n26507);
xnor_3 g24160(new_n26509, new_n26490, new_n26482);
nand_4 g24161(new_n26510_1, new_n26509, new_n8043);
xnor_3 g24162(new_n26511, new_n26488, new_n26487);
nand_4 g24163(new_n26512_1, new_n26511, new_n8137);
xnor_3 g24164(new_n26513, new_n26511, new_n8138);
nand_4 g24165(new_n26514, new_n26451, new_n8142);
nand_4 g24166(new_n26515_1, new_n26460, new_n26452_1);
nand_4 g24167(new_n26516, new_n26515_1, new_n26514);
nand_4 g24168(new_n26517, new_n26516, new_n26513);
nand_4 g24169(new_n26518, new_n26517, new_n26512_1);
xnor_3 g24170(new_n26519, new_n26509, new_n25696);
nand_4 g24171(new_n26520, new_n26519, new_n26518);
nand_4 g24172(new_n26521, new_n26520, new_n26510_1);
nand_4 g24173(new_n26522, new_n26521, new_n26508);
nand_4 g24174(new_n26523, new_n26522, new_n26506);
nand_4 g24175(new_n26524, new_n26523, new_n26503);
nand_4 g24176(new_n26525, new_n26524, new_n26502);
not_3  g24177(new_n26526, new_n26525);
nand_4 g24178(new_n26527, new_n26526, new_n20979);
not_3  g24179(new_n26528, new_n20979);
nand_4 g24180(new_n26529, new_n26525, new_n26528);
not_3  g24181(new_n26530, new_n26495);
nor_4  g24182(new_n26531, new_n26530, new_n18389);
not_3  g24183(new_n26532, new_n26531);
nor_4  g24184(new_n26533, new_n26532, new_n26475);
not_3  g24185(new_n26534, new_n26533);
nand_4 g24186(new_n26535, new_n26534, new_n26529);
nand_4 g24187(new_n26536, new_n26535, new_n26527);
nor_4  g24188(n8288, new_n26536, new_n26497);
xor_3  g24189(n8306, new_n13533, new_n8758);
xor_3  g24190(n8320, new_n9388, new_n9333);
not_3  g24191(new_n26540, new_n15045);
xor_3  g24192(n8321, new_n15071, new_n26540);
xnor_3 g24193(n8339, new_n20043, new_n20026);
xnor_3 g24194(n8376, new_n10859, new_n10801);
xor_3  g24195(n8408, new_n23522, new_n12280);
xor_3  g24196(n8417, new_n17546, new_n17545);
not_3  g24197(new_n26546, new_n15584);
xor_3  g24198(n8432, new_n15604, new_n26546);
not_3  g24199(new_n26548, new_n12142);
nor_4  g24200(new_n26549, new_n12164, new_n25305);
not_3  g24201(new_n26550, new_n12232);
nor_4  g24202(new_n26551, new_n26550, new_n12165);
nor_4  g24203(new_n26552, new_n26551, new_n26549);
nor_4  g24204(new_n26553_1, new_n26552, new_n26548);
nor_4  g24205(new_n26554, new_n12233, new_n12142);
nor_4  g24206(new_n26555, new_n12314, new_n12234);
nor_4  g24207(new_n26556, new_n26555, new_n26554);
nor_4  g24208(new_n26557, new_n26556, new_n26553_1);
not_3  g24209(new_n26558, new_n26552);
nor_4  g24210(new_n26559, new_n26558, new_n12142);
nor_4  g24211(new_n26560, new_n26559, new_n26555);
nor_4  g24212(n8453, new_n26560, new_n26557);
xor_3  g24213(n8480, new_n19060, new_n16641);
xnor_3 g24214(n8489, new_n20239, new_n20214);
xnor_3 g24215(n8505, new_n26432, new_n26414);
xnor_3 g24216(n8510, new_n24060, new_n24040);
xor_3  g24217(n8519, new_n14669, new_n10309);
not_3  g24218(new_n26567, new_n11696);
xor_3  g24219(n8535, new_n26567, new_n11695);
xnor_3 g24220(n8550, new_n23723, new_n23719_1);
not_3  g24221(new_n26570, new_n25180);
xor_3  g24222(n8563, new_n26570, new_n25169);
xor_3  g24223(n8594, new_n16200, new_n16196_1);
not_3  g24224(new_n26573, new_n8164);
xor_3  g24225(n8608, new_n8188, new_n26573);
xor_3  g24226(n8620, new_n5198, new_n5195);
xnor_3 g24227(n8637, new_n8783, new_n8717);
xnor_3 g24228(n8662, new_n21081, new_n21080);
not_3  g24229(new_n26578, new_n23176);
xor_3  g24230(n8716, new_n23187, new_n26578);
nand_4 g24231(new_n26580, new_n9341, new_n9339);
xor_3  g24232(n8744, new_n26580, new_n9386);
nor_4  g24233(new_n26582, new_n15536, new_n9258);
not_3  g24234(new_n26583, new_n26582);
nand_4 g24235(new_n26584, new_n26198, new_n26583);
nand_4 g24236(new_n26585, new_n26584, new_n18755);
not_3  g24237(new_n26586, new_n26585);
nor_4  g24238(new_n26587, new_n26584, new_n18755);
nor_4  g24239(new_n26588, new_n26587, new_n26586);
nor_4  g24240(new_n26589, new_n7068, new_n21148);
nor_4  g24241(new_n26590_1, new_n26089, new_n26084_1);
nor_4  g24242(new_n26591, new_n26590_1, new_n26589);
xnor_3 g24243(new_n26592, new_n26591, new_n21894);
not_3  g24244(new_n26593, new_n26592);
nor_4  g24245(new_n26594, new_n26593, new_n26588);
xnor_3 g24246(new_n26595, new_n26584, new_n18755);
nor_4  g24247(new_n26596, new_n26592, new_n26595);
nor_4  g24248(new_n26597, new_n26596, new_n26594);
xnor_3 g24249(new_n26598_1, new_n26197, new_n26188);
nor_4  g24250(new_n26599, new_n26598_1, new_n26090);
not_3  g24251(new_n26600, new_n26599);
nor_4  g24252(new_n26601, new_n26201, new_n26091);
nor_4  g24253(new_n26602, new_n26601, new_n26599);
nor_4  g24254(new_n26603, new_n26205, new_n26095);
xnor_3 g24255(new_n26604, new_n26205, new_n26095);
nor_4  g24256(new_n26605_1, new_n21344, new_n19802);
nor_4  g24257(new_n26606, new_n21385, new_n21345);
nor_4  g24258(new_n26607, new_n26606, new_n26605_1);
nor_4  g24259(new_n26608, new_n26607, new_n26604);
nor_4  g24260(new_n26609, new_n26608, new_n26603);
nand_4 g24261(new_n26610, new_n26609, new_n26602);
nand_4 g24262(new_n26611, new_n26610, new_n26600);
xnor_3 g24263(n8803, new_n26611, new_n26597);
nor_4  g24264(new_n26613, new_n24979, n13494);
nor_4  g24265(new_n26614, new_n24980, new_n6510);
not_3  g24266(new_n26615, new_n26614);
nand_4 g24267(new_n26616, new_n25007, new_n24982);
nand_4 g24268(new_n26617, new_n26616, new_n26615);
xnor_3 g24269(new_n26618, new_n26617, new_n26613);
not_3  g24270(new_n26619, new_n26618);
nor_4  g24271(new_n26620, n16544, n4319);
not_3  g24272(new_n26621, new_n26620);
nand_4 g24273(new_n26622, new_n19378, new_n26621);
nor_4  g24274(new_n26623, new_n26622, new_n26619);
not_3  g24275(new_n26624, new_n26623);
not_3  g24276(new_n26625_1, new_n26622);
nor_4  g24277(new_n26626, new_n26625_1, new_n26618);
not_3  g24278(new_n26627, new_n26626);
nand_4 g24279(new_n26628, new_n26627, new_n26624);
not_3  g24280(new_n26629, new_n25012);
nor_4  g24281(new_n26630, new_n25036, new_n26629);
nor_4  g24282(new_n26631, new_n26630, new_n25010);
not_3  g24283(new_n26632, new_n26631);
xnor_3 g24284(new_n26633, new_n26632, new_n26628);
nor_4  g24285(new_n26634, new_n26633, new_n9127);
not_3  g24286(new_n26635, new_n9127);
xnor_3 g24287(new_n26636, new_n26631, new_n26628);
nor_4  g24288(new_n26637, new_n26636, new_n26635);
nor_4  g24289(new_n26638, new_n26637, new_n26634);
nor_4  g24290(new_n26639, new_n25037, new_n9130);
not_3  g24291(new_n26640, new_n26639);
nand_4 g24292(new_n26641, new_n25800, new_n25750);
nand_4 g24293(new_n26642, new_n26641, new_n26640);
xnor_3 g24294(n8809, new_n26642, new_n26638);
nor_4  g24295(new_n26644, new_n26591, new_n21895);
not_3  g24296(new_n26645, new_n26644);
nand_4 g24297(new_n26646, new_n22335_1, new_n19353);
nand_4 g24298(new_n26647, new_n26080, new_n26646);
nor_4  g24299(new_n26648, new_n26647, new_n22330);
nor_4  g24300(new_n26649, new_n26648, new_n26645);
not_3  g24301(new_n26650, new_n26648);
nor_4  g24302(new_n26651, new_n26650, new_n26644);
nor_4  g24303(new_n26652, new_n26651, new_n26649);
xnor_3 g24304(new_n26653, new_n26647, new_n22330);
nand_4 g24305(new_n26654, new_n26653, new_n26592);
xnor_3 g24306(new_n26655, new_n26653, new_n26593);
nand_4 g24307(new_n26656_1, new_n26090, new_n26083);
nand_4 g24308(new_n26657, new_n26109, new_n26092);
nand_4 g24309(new_n26658, new_n26657, new_n26656_1);
nand_4 g24310(new_n26659, new_n26658, new_n26655);
nand_4 g24311(new_n26660_1, new_n26659, new_n26654);
xnor_3 g24312(n8821, new_n26660_1, new_n26652);
not_3  g24313(new_n26662, new_n19030);
xor_3  g24314(n8824, new_n26662, new_n19027);
xor_3  g24315(n8849, new_n21831, new_n21830);
xnor_3 g24316(n8861, new_n16804, new_n16795);
xor_3  g24317(new_n26666, n22442, new_n3662);
not_3  g24318(new_n26667, new_n26666);
nand_4 g24319(new_n26668, new_n9033, n468);
nand_4 g24320(new_n26669, new_n24733, new_n24703);
nand_4 g24321(new_n26670, new_n26669, new_n26668);
xnor_3 g24322(new_n26671, new_n26670, new_n26667);
not_3  g24323(new_n26672, new_n8869_1);
xor_3  g24324(new_n26673, n3324, n2272);
nand_4 g24325(new_n26674_1, new_n8203, new_n19385_1);
nand_4 g24326(new_n26675_1, new_n24694, new_n24691);
nand_4 g24327(new_n26676, new_n26675_1, new_n26674_1);
not_3  g24328(new_n26677, new_n26676);
xor_3  g24329(new_n26678, new_n26677, new_n26673);
nand_4 g24330(new_n26679, new_n26678, new_n26672);
not_3  g24331(new_n26680, new_n26679);
nor_4  g24332(new_n26681_1, new_n26678, new_n26672);
nor_4  g24333(new_n26682, new_n26681_1, new_n26680);
not_3  g24334(new_n26683, new_n8861_1);
not_3  g24335(new_n26684, new_n24695);
nor_4  g24336(new_n26685, new_n26684, new_n26683);
not_3  g24337(new_n26686, new_n26685);
nand_4 g24338(new_n26687, new_n24700, new_n24697);
nand_4 g24339(new_n26688, new_n26687, new_n26686);
xnor_3 g24340(new_n26689, new_n26688, new_n26682);
xnor_3 g24341(new_n26690, new_n26689, new_n26671);
nor_4  g24342(new_n26691, new_n24734, new_n24701);
not_3  g24343(new_n26692, new_n26691);
nand_4 g24344(new_n26693, new_n24772, new_n24735);
nand_4 g24345(new_n26694, new_n26693, new_n26692);
nand_4 g24346(new_n26695, new_n26694, new_n26690);
not_3  g24347(new_n26696_1, new_n26695);
nor_4  g24348(new_n26697, new_n26694, new_n26690);
nor_4  g24349(n8862, new_n26697, new_n26696_1);
xor_3  g24350(n8884, new_n16649, new_n16648);
xor_3  g24351(n8909, new_n23402, new_n22428);
not_3  g24352(new_n26701, new_n14150);
xor_3  g24353(n8911, new_n26701, new_n14090_1);
xnor_3 g24354(n8971, new_n13457_1, new_n13456_1);
xnor_3 g24355(n8982, new_n26292, new_n26267);
not_3  g24356(new_n26705, new_n6304);
xor_3  g24357(n8993, new_n26705, new_n6274);
xor_3  g24358(n9012, new_n17554, new_n17553);
nor_4  g24359(new_n26708, new_n24890, new_n24886);
nor_4  g24360(new_n26709, new_n24895, new_n5125);
not_3  g24361(new_n26710, new_n26709);
nor_4  g24362(new_n26711, new_n26710, new_n24893);
xnor_3 g24363(new_n26712, new_n26711, new_n26708);
nor_4  g24364(new_n26713, new_n24898, new_n24891);
nor_4  g24365(new_n26714, new_n24950, new_n24899);
nor_4  g24366(new_n26715, new_n26714, new_n26713);
xnor_3 g24367(n9032, new_n26715, new_n26712);
not_3  g24368(new_n26717, new_n19709);
xor_3  g24369(n9042, new_n26717, new_n19705);
xnor_3 g24370(n9046, new_n21319, new_n21282);
xnor_3 g24371(n9047, new_n9741, new_n9665);
not_3  g24372(new_n26721, new_n18685);
xor_3  g24373(n9104, new_n26721, new_n18684);
not_3  g24374(new_n26723, new_n25348);
nor_4  g24375(new_n26724, new_n26723, new_n25338);
nand_4 g24376(new_n26725_1, new_n26724, new_n18964);
nor_4  g24377(new_n26726, new_n25348, new_n25339);
nand_4 g24378(new_n26727_1, new_n26726, new_n25351);
nand_4 g24379(new_n26728, new_n26727_1, new_n26725_1);
nor_4  g24380(new_n26729_1, new_n26728, new_n23983);
not_3  g24381(new_n26730, new_n26728);
nor_4  g24382(new_n26731, new_n26730, new_n24015);
nor_4  g24383(new_n26732, new_n26731, new_n26729_1);
nand_4 g24384(new_n26733, new_n25354, new_n24015);
nand_4 g24385(new_n26734, new_n25370_1, new_n25355);
nand_4 g24386(new_n26735, new_n26734, new_n26733);
xnor_3 g24387(n9129, new_n26735, new_n26732);
xor_3  g24388(n9146, new_n23652, new_n23614);
xor_3  g24389(n9164, new_n10309, new_n7886);
xor_3  g24390(n9166, new_n15498, new_n15497);
xnor_3 g24391(new_n26740, new_n22347, new_n22320);
xnor_3 g24392(n9182, new_n26740, new_n22362);
xnor_3 g24393(n9191, new_n8453_1, new_n8416);
xnor_3 g24394(n9217, new_n14154, new_n14076);
xor_3  g24395(n9220, new_n19915, new_n19914);
not_3  g24396(new_n26745_1, new_n23634);
xor_3  g24397(n9261, new_n23642, new_n26745_1);
xor_3  g24398(new_n26747, n22626, new_n19353);
not_3  g24399(new_n26748_1, new_n26747);
nor_4  g24400(new_n26749, new_n19385_1, n14440);
not_3  g24401(new_n26750, new_n26749);
nand_4 g24402(new_n26751, new_n23159, new_n23135);
nand_4 g24403(new_n26752_1, new_n26751, new_n26750);
not_3  g24404(new_n26753, new_n26752_1);
xor_3  g24405(new_n26754, new_n26753, new_n26748_1);
not_3  g24406(new_n26755, new_n26754);
nor_4  g24407(new_n26756, new_n26755, new_n22352);
not_3  g24408(new_n26757, new_n26756);
nor_4  g24409(new_n26758, new_n26754, new_n22353_1);
nor_4  g24410(new_n26759, new_n26758, new_n26756);
not_3  g24411(new_n26760, new_n23162);
nand_4 g24412(new_n26761, new_n23193, new_n23165);
nand_4 g24413(new_n26762, new_n26761, new_n26760);
nand_4 g24414(new_n26763, new_n26762, new_n26759);
nand_4 g24415(new_n26764, new_n26763, new_n26757);
nor_4  g24416(new_n26765, n22626, new_n19353);
nor_4  g24417(new_n26766, new_n26753, new_n26748_1);
nor_4  g24418(new_n26767, new_n26766, new_n26765);
not_3  g24419(new_n26768, new_n26767);
nor_4  g24420(new_n26769, new_n26768, new_n22348);
nor_4  g24421(new_n26770, new_n26767, new_n22347);
nor_4  g24422(new_n26771, new_n26770, new_n26769);
xnor_3 g24423(n9287, new_n26771, new_n26764);
xor_3  g24424(n9308, new_n17315, new_n17302_1);
xnor_3 g24425(n9344, new_n5740, new_n5684);
not_3  g24426(new_n26775_1, new_n4032);
xor_3  g24427(n9364, new_n4060, new_n26775_1);
not_3  g24428(new_n26777, new_n26764);
not_3  g24429(new_n26778, new_n26770);
nor_4  g24430(new_n26779, new_n26778, new_n26777);
nand_4 g24431(new_n26780_1, new_n26779, new_n22345);
not_3  g24432(new_n26781, new_n26769);
nor_4  g24433(new_n26782, new_n26781, new_n26764);
nand_4 g24434(new_n26783, new_n26782, new_n22366);
nand_4 g24435(n9371, new_n26783, new_n26780_1);
xor_3  g24436(n9382, new_n12282, new_n12280);
not_3  g24437(new_n26786, new_n26325);
not_3  g24438(new_n26787, new_n26326);
not_3  g24439(new_n26788, new_n26328);
not_3  g24440(new_n26789, new_n21326);
nand_4 g24441(new_n26790, new_n26789, new_n26788);
nand_4 g24442(new_n26791, new_n26790, new_n26787);
nand_4 g24443(new_n26792, new_n26791, new_n26786);
xnor_3 g24444(n9403, new_n26792, new_n26321);
not_3  g24445(new_n26794_1, new_n15477_1);
xor_3  g24446(n9419, new_n15504, new_n26794_1);
xnor_3 g24447(new_n26796, new_n26015, new_n18983);
xor_3  g24448(n9423, new_n26046, new_n26796);
not_3  g24449(new_n26798, new_n23173);
xor_3  g24450(n9430, new_n23189, new_n26798);
xor_3  g24451(new_n26800, n25120, new_n4907);
nand_4 g24452(new_n26801_1, new_n22700, n8363);
xor_3  g24453(new_n26802, n11481, new_n22667);
nand_4 g24454(new_n26803, new_n22702, n14680);
nand_4 g24455(new_n26804, new_n19266, new_n19262);
nand_4 g24456(new_n26805, new_n26804, new_n26803);
nand_4 g24457(new_n26806, new_n26805, new_n26802);
nand_4 g24458(new_n26807, new_n26806, new_n26801_1);
xnor_3 g24459(new_n26808_1, new_n26807, new_n26800);
xnor_3 g24460(new_n26809, new_n26808_1, new_n21175);
xnor_3 g24461(new_n26810, new_n26805, new_n26802);
nor_4  g24462(new_n26811, new_n26810, new_n21178);
not_3  g24463(new_n26812, new_n26811);
not_3  g24464(new_n26813, new_n26810);
nor_4  g24465(new_n26814, new_n26813, new_n21204);
nor_4  g24466(new_n26815_1, new_n26814, new_n26811);
nand_4 g24467(new_n26816, new_n19275, new_n19268);
not_3  g24468(new_n26817, new_n19276);
nand_4 g24469(new_n26818, new_n19287, new_n26817);
nand_4 g24470(new_n26819, new_n26818, new_n26816);
nand_4 g24471(new_n26820, new_n26819, new_n26815_1);
nand_4 g24472(new_n26821, new_n26820, new_n26812);
xnor_3 g24473(new_n26822, new_n26821, new_n26809);
xnor_3 g24474(new_n26823_1, new_n26822, new_n21263);
not_3  g24475(new_n26824, new_n26823_1);
not_3  g24476(new_n26825, new_n26815_1);
xnor_3 g24477(new_n26826, new_n26819, new_n26825);
nor_4  g24478(new_n26827, new_n26826, new_n21266);
not_3  g24479(new_n26828, new_n26827);
xnor_3 g24480(new_n26829, new_n26819, new_n26815_1);
nor_4  g24481(new_n26830, new_n26829, new_n21267);
nor_4  g24482(new_n26831, new_n26830, new_n26827);
nor_4  g24483(new_n26832, new_n21272, new_n19288);
not_3  g24484(new_n26833, new_n26832);
xnor_3 g24485(new_n26834, new_n19287, new_n26817);
nor_4  g24486(new_n26835, new_n21273, new_n26834);
nor_4  g24487(new_n26836, new_n26835, new_n26832);
nand_4 g24488(new_n26837, new_n21278, new_n19290);
xnor_3 g24489(new_n26838, new_n21278, new_n12835);
nand_4 g24490(new_n26839, new_n21288, new_n12837);
not_3  g24491(new_n26840, new_n26839);
nor_4  g24492(new_n26841, new_n21288, new_n12837);
nor_4  g24493(new_n26842, new_n26841, new_n26840);
nor_4  g24494(new_n26843, new_n21292, new_n12844);
not_3  g24495(new_n26844, new_n12849);
nor_4  g24496(new_n26845, new_n21300, new_n26844);
nor_4  g24497(new_n26846, new_n18343_1, new_n18327);
nor_4  g24498(new_n26847_1, new_n26846, new_n26845);
xnor_3 g24499(new_n26848, new_n21292, new_n12844);
nor_4  g24500(new_n26849, new_n26848, new_n26847_1);
nor_4  g24501(new_n26850, new_n26849, new_n26843);
nand_4 g24502(new_n26851, new_n26850, new_n26842);
nand_4 g24503(new_n26852, new_n26851, new_n26839);
nand_4 g24504(new_n26853, new_n26852, new_n26838);
nand_4 g24505(new_n26854, new_n26853, new_n26837);
nand_4 g24506(new_n26855, new_n26854, new_n26836);
nand_4 g24507(new_n26856, new_n26855, new_n26833);
nand_4 g24508(new_n26857, new_n26856, new_n26831);
nand_4 g24509(new_n26858, new_n26857, new_n26828);
xnor_3 g24510(n9435, new_n26858, new_n26824);
xnor_3 g24511(n9451, new_n19848, new_n19813);
xor_3  g24512(new_n26861, n12657, new_n20487);
not_3  g24513(new_n26862, new_n26861);
nand_4 g24514(new_n26863, new_n8555, n7437);
nand_4 g24515(new_n26864, new_n23790, new_n23782);
nand_4 g24516(new_n26865, new_n26864, new_n26863);
xor_3  g24517(new_n26866, new_n26865, new_n26862);
xnor_3 g24518(new_n26867, new_n26866, new_n24702);
not_3  g24519(new_n26868, new_n23825);
nand_4 g24520(new_n26869, new_n23836, new_n23826);
nand_4 g24521(new_n26870, new_n26869, new_n26868);
xnor_3 g24522(n9458, new_n26870, new_n26867);
nor_4  g24523(new_n26872, n12507, new_n22309_1);
xor_3  g24524(new_n26873, n12507, new_n22309_1);
not_3  g24525(new_n26874, new_n26873);
nor_4  g24526(new_n26875, new_n22313, n15077);
not_3  g24527(new_n26876, new_n26875);
nand_4 g24528(new_n26877, new_n18253, new_n18228);
nand_4 g24529(new_n26878, new_n26877, new_n26876);
not_3  g24530(new_n26879, new_n26878);
nor_4  g24531(new_n26880, new_n26879, new_n26874);
nor_4  g24532(new_n26881, new_n26880, new_n26872);
nor_4  g24533(new_n26882_1, new_n26881, new_n25615);
nand_4 g24534(new_n26883, new_n26881, new_n25615);
not_3  g24535(new_n26884, new_n26883);
nor_4  g24536(new_n26885, new_n26884, new_n26882_1);
xor_3  g24537(new_n26886, new_n26879, new_n26874);
nor_4  g24538(new_n26887, new_n26886, new_n25619_1);
not_3  g24539(new_n26888, new_n26886);
nor_4  g24540(new_n26889, new_n26888, new_n25626);
nor_4  g24541(new_n26890, new_n26889, new_n26887);
not_3  g24542(new_n26891, new_n26890);
nand_4 g24543(new_n26892, new_n18255, new_n25622);
nand_4 g24544(new_n26893, new_n18292, new_n18256);
nand_4 g24545(new_n26894, new_n26893, new_n26892);
not_3  g24546(new_n26895, new_n26894);
nor_4  g24547(new_n26896, new_n26895, new_n26891);
nor_4  g24548(new_n26897, new_n26896, new_n26887);
not_3  g24549(new_n26898, new_n26897);
xnor_3 g24550(n9459, new_n26898, new_n26885);
xnor_3 g24551(n9508, new_n18605, new_n18600);
not_3  g24552(new_n26901, new_n15466);
xor_3  g24553(n9552, new_n15509, new_n26901);
xor_3  g24554(n9556, new_n5205, new_n5200);
xor_3  g24555(n9558, new_n13426, new_n10560);
xor_3  g24556(n9616, new_n25890, new_n17546);
not_3  g24557(new_n26906, new_n10220);
xor_3  g24558(n9622, new_n26906, new_n10184);
not_3  g24559(new_n26908, new_n20463);
xor_3  g24560(n9626, new_n20481, new_n26908);
not_3  g24561(new_n26910, new_n5184_1);
xor_3  g24562(n9633, new_n5210, new_n26910);
nand_4 g24563(new_n26912, n25120, new_n4907);
nand_4 g24564(new_n26913_1, new_n26807, new_n26800);
nand_4 g24565(new_n26914, new_n26913_1, new_n26912);
nor_4  g24566(new_n26915, new_n26914, new_n26304);
not_3  g24567(new_n26916, new_n26915);
not_3  g24568(new_n26917, new_n26914);
nor_4  g24569(new_n26918, new_n26917, new_n26307);
nor_4  g24570(new_n26919, new_n26918, new_n26915);
not_3  g24571(new_n26920, new_n26808_1);
nand_4 g24572(new_n26921_1, new_n26920, new_n21175);
nand_4 g24573(new_n26922, new_n26821, new_n26809);
nand_4 g24574(new_n26923_1, new_n26922, new_n26921_1);
not_3  g24575(new_n26924, new_n26923_1);
nand_4 g24576(new_n26925, new_n26924, new_n26919);
nand_4 g24577(new_n26926, new_n26925, new_n26916);
nor_4  g24578(new_n26927, new_n26926, new_n6430);
xnor_3 g24579(new_n26928, new_n26926, new_n6430);
xnor_3 g24580(new_n26929_1, new_n26923_1, new_n26919);
nor_4  g24581(new_n26930_1, new_n26929_1, new_n6431_1);
xnor_3 g24582(new_n26931, new_n26929_1, new_n6431_1);
not_3  g24583(new_n26932, new_n26809);
xnor_3 g24584(new_n26933, new_n26821, new_n26932);
nor_4  g24585(new_n26934, new_n26933, new_n6432);
not_3  g24586(new_n26935, new_n26934);
nor_4  g24587(new_n26936, new_n26829, new_n6519);
xnor_3 g24588(new_n26937, new_n26829, new_n6519);
nor_4  g24589(new_n26938, new_n26834, new_n6524);
nor_4  g24590(new_n26939, new_n19293, new_n19289);
nor_4  g24591(new_n26940, new_n26939, new_n26938);
nor_4  g24592(new_n26941, new_n26940, new_n26937);
nor_4  g24593(new_n26942, new_n26941, new_n26936);
nor_4  g24594(new_n26943_1, new_n26822, new_n6517);
nor_4  g24595(new_n26944, new_n26943_1, new_n26934);
nand_4 g24596(new_n26945, new_n26944, new_n26942);
nand_4 g24597(new_n26946, new_n26945, new_n26935);
nor_4  g24598(new_n26947, new_n26946, new_n26931);
nor_4  g24599(new_n26948, new_n26947, new_n26930_1);
nor_4  g24600(new_n26949, new_n26948, new_n26928);
nor_4  g24601(n9635, new_n26949, new_n26927);
xnor_3 g24602(n9648, new_n24089, new_n24086);
xor_3  g24603(n9689, new_n5720, new_n5718);
not_3  g24604(new_n26953, new_n13061);
xor_3  g24605(n9695, new_n26953, new_n13035);
xnor_3 g24606(n9699, new_n9022, new_n8959);
nor_4  g24607(new_n26956, new_n20600, new_n19854);
nor_4  g24608(new_n26957, new_n20589, new_n18003);
nor_4  g24609(new_n26958, new_n26957, new_n26956);
not_3  g24610(new_n26959, new_n19876);
nand_4 g24611(new_n26960, new_n19921, new_n19877);
nand_4 g24612(new_n26961, new_n26960, new_n26959);
xnor_3 g24613(n9726, new_n26961, new_n26958);
xor_3  g24614(n9753, new_n16213, new_n12071);
not_3  g24615(new_n26964, new_n3628);
xor_3  g24616(n9761, new_n26964, new_n3604);
xnor_3 g24617(n9763, new_n12085, new_n12037);
xor_3  g24618(n9767, new_n16646, new_n16642);
xor_3  g24619(n9771, new_n16863, new_n16513);
xor_3  g24620(n9778, new_n26428, new_n26425);
not_3  g24621(new_n26970_1, new_n19560);
xor_3  g24622(n9783, new_n19568, new_n26970_1);
not_3  g24623(new_n26972, new_n7923);
xor_3  g24624(n9803, new_n26972, new_n7919);
not_3  g24625(new_n26974, new_n25812);
nor_4  g24626(new_n26975, new_n26974, n23463);
not_3  g24627(new_n26976, new_n26975);
nor_4  g24628(new_n26977, new_n26976, n4319);
not_3  g24629(new_n26978, new_n26977);
xor_3  g24630(new_n26979_1, new_n26975, new_n14181);
not_3  g24631(new_n26980, new_n26979_1);
nand_4 g24632(new_n26981, new_n26980, new_n22279);
xnor_3 g24633(new_n26982, new_n26979_1, new_n22279);
nand_4 g24634(new_n26983, new_n25814, new_n22287);
nand_4 g24635(new_n26984, new_n25819, new_n20676);
xnor_3 g24636(new_n26985, new_n25819, new_n20675);
nand_4 g24637(new_n26986_1, new_n25824, new_n20683);
nor_4  g24638(new_n26987, new_n25829, new_n20687);
xnor_3 g24639(new_n26988, new_n25829, new_n20687);
nor_4  g24640(new_n26989, new_n7870, new_n7854);
nor_4  g24641(new_n26990, new_n7904, new_n7871);
nor_4  g24642(new_n26991, new_n26990, new_n26989);
nor_4  g24643(new_n26992, new_n26991, new_n26988);
nor_4  g24644(new_n26993, new_n26992, new_n26987);
xnor_3 g24645(new_n26994, new_n25824, new_n20682);
nand_4 g24646(new_n26995, new_n26994, new_n26993);
nand_4 g24647(new_n26996, new_n26995, new_n26986_1);
nand_4 g24648(new_n26997, new_n26996, new_n26985);
nand_4 g24649(new_n26998, new_n26997, new_n26984);
xnor_3 g24650(new_n26999, new_n25813, new_n22287);
nand_4 g24651(new_n27000, new_n26999, new_n26998);
nand_4 g24652(new_n27001, new_n27000, new_n26983);
nand_4 g24653(new_n27002, new_n27001, new_n26982);
nand_4 g24654(new_n27003, new_n27002, new_n26981);
xnor_3 g24655(new_n27004_1, new_n27003, new_n22273);
nand_4 g24656(new_n27005, new_n27004_1, new_n26978);
xnor_3 g24657(new_n27006, new_n27003, new_n22272);
nand_4 g24658(new_n27007, new_n27006, new_n26977);
nand_4 g24659(new_n27008, new_n27007, new_n27005);
not_3  g24660(new_n27009, new_n27008);
nand_4 g24661(new_n27010, new_n27009, new_n3644);
xnor_3 g24662(new_n27011_1, new_n27008, new_n3644);
xnor_3 g24663(new_n27012, new_n27001, new_n26982);
nor_4  g24664(new_n27013, new_n27012, new_n3559);
not_3  g24665(new_n27014, new_n27013);
not_3  g24666(new_n27015, new_n27012);
xnor_3 g24667(new_n27016, new_n27015, new_n3559);
not_3  g24668(new_n27017, new_n3565);
not_3  g24669(new_n27018, new_n27000);
nor_4  g24670(new_n27019_1, new_n26999, new_n26998);
nor_4  g24671(new_n27020, new_n27019_1, new_n27018);
nand_4 g24672(new_n27021, new_n27020, new_n27017);
xnor_3 g24673(new_n27022, new_n27020, new_n3565);
not_3  g24674(new_n27023, new_n3571);
not_3  g24675(new_n27024, new_n26985);
xnor_3 g24676(new_n27025, new_n26996, new_n27024);
nand_4 g24677(new_n27026, new_n27025, new_n27023);
xnor_3 g24678(new_n27027, new_n27025, new_n3571);
not_3  g24679(new_n27028, new_n26993);
xnor_3 g24680(new_n27029, new_n26994, new_n27028);
nand_4 g24681(new_n27030, new_n27029, new_n3577);
xnor_3 g24682(new_n27031_1, new_n27029, new_n3576);
xnor_3 g24683(new_n27032, new_n26991, new_n26988);
nand_4 g24684(new_n27033, new_n27032, new_n3585);
xnor_3 g24685(new_n27034, new_n27032, new_n3584);
nand_4 g24686(new_n27035, new_n7905, new_n3591);
nand_4 g24687(new_n27036, new_n7930, new_n7906);
nand_4 g24688(new_n27037_1, new_n27036, new_n27035);
nand_4 g24689(new_n27038, new_n27037_1, new_n27034);
nand_4 g24690(new_n27039, new_n27038, new_n27033);
nand_4 g24691(new_n27040, new_n27039, new_n27031_1);
nand_4 g24692(new_n27041, new_n27040, new_n27030);
nand_4 g24693(new_n27042, new_n27041, new_n27027);
nand_4 g24694(new_n27043, new_n27042, new_n27026);
nand_4 g24695(new_n27044, new_n27043, new_n27022);
nand_4 g24696(new_n27045, new_n27044, new_n27021);
nand_4 g24697(new_n27046, new_n27045, new_n27016);
nand_4 g24698(new_n27047, new_n27046, new_n27014);
nand_4 g24699(new_n27048, new_n27047, new_n27011_1);
nand_4 g24700(new_n27049, new_n27048, new_n27010);
not_3  g24701(new_n27050, new_n27003);
nor_4  g24702(new_n27051_1, new_n27050, new_n22272);
xor_3  g24703(new_n27052, new_n26978, new_n22270_1);
nand_4 g24704(new_n27053, new_n27052, new_n27051_1);
nor_4  g24705(new_n27054, new_n27052, new_n27003);
not_3  g24706(new_n27055, new_n27054);
nand_4 g24707(new_n27056, new_n27055, new_n27053);
nor_4  g24708(new_n27057, new_n27056, new_n27049);
nor_4  g24709(new_n27058, new_n26977, new_n22222);
nand_4 g24710(new_n27059, new_n27058, new_n27003);
xnor_3 g24711(n9833, new_n27059, new_n27057);
nand_4 g24712(new_n27061, new_n21547, new_n10445);
nor_4  g24713(new_n27062, new_n27061, n15077);
xor_3  g24714(new_n27063, new_n27062, new_n10423);
nor_4  g24715(new_n27064, new_n27063, new_n15734);
not_3  g24716(new_n27065, new_n27064);
xor_3  g24717(new_n27066, new_n27061, n15077);
nor_4  g24718(new_n27067, new_n27066, new_n6112);
not_3  g24719(new_n27068, new_n27067);
not_3  g24720(new_n27069, new_n27066);
nor_4  g24721(new_n27070, new_n27069, new_n6111);
nor_4  g24722(new_n27071, new_n27070, new_n27067);
nor_4  g24723(new_n27072_1, new_n21548, new_n6159);
nor_4  g24724(new_n27073, new_n21554, new_n27072_1);
nand_4 g24725(new_n27074, new_n27073, new_n27071);
nand_4 g24726(new_n27075, new_n27074, new_n27068);
not_3  g24727(new_n27076, new_n15734);
not_3  g24728(new_n27077, new_n27063);
nor_4  g24729(new_n27078, new_n27077, new_n27076);
nor_4  g24730(new_n27079_1, new_n27078, new_n27064);
nand_4 g24731(new_n27080, new_n27079_1, new_n27075);
nand_4 g24732(new_n27081, new_n27080, new_n27065);
not_3  g24733(new_n27082, new_n27062);
nor_4  g24734(new_n27083, new_n27082, n12507);
xor_3  g24735(new_n27084, new_n27083, new_n19857);
xnor_3 g24736(new_n27085, new_n27084, new_n27081);
nand_4 g24737(new_n27086, new_n21501, new_n8045);
nor_4  g24738(new_n27087, new_n27086, n21915);
xor_3  g24739(new_n27088, new_n27087, new_n20945);
nand_4 g24740(new_n27089_1, new_n27088, new_n22244);
not_3  g24741(new_n27090, new_n27089_1);
nor_4  g24742(new_n27091, new_n27088, new_n22244);
nor_4  g24743(new_n27092, new_n27091, new_n27090);
xor_3  g24744(new_n27093, new_n27086, n21915);
not_3  g24745(new_n27094, new_n27093);
nor_4  g24746(new_n27095, new_n27094, new_n22250);
not_3  g24747(new_n27096_1, new_n27095);
not_3  g24748(new_n27097, new_n22250);
nor_4  g24749(new_n27098, new_n27093, new_n27097);
nor_4  g24750(new_n27099, new_n27098, new_n27095);
not_3  g24751(new_n27100, new_n21504);
nand_4 g24752(new_n27101, new_n21545, new_n21507);
nand_4 g24753(new_n27102, new_n27101, new_n27100);
nand_4 g24754(new_n27103, new_n27102, new_n27099);
nand_4 g24755(new_n27104_1, new_n27103, new_n27096_1);
nand_4 g24756(new_n27105, new_n27104_1, new_n27092);
nand_4 g24757(new_n27106, new_n27105, new_n27089_1);
not_3  g24758(new_n27107, new_n27087);
nor_4  g24759(new_n27108, new_n27107, n25972);
xnor_3 g24760(new_n27109, new_n27108, new_n22267);
xnor_3 g24761(new_n27110_1, new_n27109, new_n27106);
nand_4 g24762(new_n27111, new_n27110_1, new_n27085);
not_3  g24763(new_n27112_1, new_n27080);
nor_4  g24764(new_n27113, new_n27112_1, new_n27064);
xnor_3 g24765(new_n27114, new_n27084, new_n27113);
xnor_3 g24766(new_n27115, new_n27110_1, new_n27114);
xnor_3 g24767(new_n27116, new_n27104_1, new_n27092);
xnor_3 g24768(new_n27117, new_n27079_1, new_n27075);
not_3  g24769(new_n27118, new_n27117);
nand_4 g24770(new_n27119, new_n27118, new_n27116);
xnor_3 g24771(new_n27120_1, new_n27117, new_n27116);
not_3  g24772(new_n27121, new_n27071);
xnor_3 g24773(new_n27122, new_n27073, new_n27121);
xnor_3 g24774(new_n27123, new_n27102, new_n27099);
nand_4 g24775(new_n27124, new_n27123, new_n27122);
xnor_3 g24776(new_n27125, new_n27073, new_n27071);
xnor_3 g24777(new_n27126, new_n27123, new_n27125);
not_3  g24778(new_n27127, new_n21557);
nand_4 g24779(new_n27128, new_n27127, new_n21546);
nand_4 g24780(new_n27129, new_n21608, new_n21558);
nand_4 g24781(new_n27130_1, new_n27129, new_n27128);
nand_4 g24782(new_n27131, new_n27130_1, new_n27126);
nand_4 g24783(new_n27132, new_n27131, new_n27124);
nand_4 g24784(new_n27133, new_n27132, new_n27120_1);
nand_4 g24785(new_n27134_1, new_n27133, new_n27119);
nand_4 g24786(new_n27135, new_n27134_1, new_n27115);
nand_4 g24787(new_n27136, new_n27135, new_n27111);
nor_4  g24788(new_n27137, new_n27108, new_n22267);
not_3  g24789(new_n27138, new_n27137);
nor_4  g24790(new_n27139, new_n27138, new_n27106);
nand_4 g24791(new_n27140, new_n27139, new_n27136);
xnor_3 g24792(new_n27141, new_n27139, new_n27136);
nor_4  g24793(new_n27142, new_n27083, new_n19857);
and_4  g24794(new_n27143, new_n27142, new_n27081);
nand_4 g24795(new_n27144, new_n27143, new_n27141);
nand_4 g24796(n9838, new_n27144, new_n27140);
xnor_3 g24797(n9867, new_n24280, new_n24277);
not_3  g24798(new_n27147, new_n23749);
nor_4  g24799(new_n27148, new_n23752, new_n27147);
nor_4  g24800(new_n27149, new_n27148, new_n23748_1);
nor_4  g24801(new_n27150, new_n27149, new_n25286);
xnor_3 g24802(new_n27151, new_n27149, new_n25286);
nand_4 g24803(new_n27152, new_n27151, new_n9652);
not_3  g24804(new_n27153, new_n23753);
nand_4 g24805(new_n27154, new_n27153, new_n9660);
nand_4 g24806(new_n27155, new_n23758, new_n23754);
nand_4 g24807(new_n27156, new_n27155, new_n27154);
nor_4  g24808(new_n27157, new_n9651, new_n9521);
nor_4  g24809(new_n27158_1, new_n27157, new_n9525);
xnor_3 g24810(new_n27159, new_n27151, new_n27158_1);
nand_4 g24811(new_n27160, new_n27159, new_n27156);
nand_4 g24812(new_n27161, new_n27160, new_n27152);
not_3  g24813(new_n27162, new_n27161);
nor_4  g24814(new_n27163_1, new_n27162, new_n27150);
nor_4  g24815(n9890, new_n27163_1, new_n9525);
and_4  g24816(new_n27165, new_n22302, new_n22286);
nor_4  g24817(new_n27166, new_n22302, new_n22286);
nor_4  g24818(n9917, new_n27166, new_n27165);
xnor_3 g24819(n9919, new_n25653, new_n25646);
not_3  g24820(new_n27169, new_n22509);
xor_3  g24821(n9938, new_n27169, new_n22490);
xor_3  g24822(n9946, new_n22047, new_n25782);
xor_3  g24823(new_n27172, n21784, n3740);
not_3  g24824(new_n27173, new_n27172);
nand_4 g24825(new_n27174, new_n14323_1, new_n17338);
xor_3  g24826(new_n27175, n5521, n2858);
nand_4 g24827(new_n27176, new_n14330, new_n5602);
xor_3  g24828(new_n27177, n11926, n2659);
nand_4 g24829(new_n27178, new_n5606, new_n4219);
xor_3  g24830(new_n27179, n24327, n4325);
nand_4 g24831(new_n27180, n22198, n5337);
not_3  g24832(new_n27181, new_n27180);
nor_4  g24833(new_n27182, n22198, n5337);
nor_4  g24834(new_n27183, n20826, n626);
not_3  g24835(new_n27184, new_n27183);
nand_4 g24836(new_n27185, new_n15705, new_n15702);
nand_4 g24837(new_n27186, new_n27185, new_n27184);
nor_4  g24838(new_n27187, new_n27186, new_n27182);
nor_4  g24839(new_n27188_1, new_n27187, new_n27181);
nand_4 g24840(new_n27189, new_n27188_1, new_n27179);
nand_4 g24841(new_n27190, new_n27189, new_n27178);
nand_4 g24842(new_n27191, new_n27190, new_n27177);
nand_4 g24843(new_n27192, new_n27191, new_n27176);
nand_4 g24844(new_n27193, new_n27192, new_n27175);
nand_4 g24845(new_n27194_1, new_n27193, new_n27174);
not_3  g24846(new_n27195, new_n27194_1);
xor_3  g24847(new_n27196, new_n27195, new_n27173);
xnor_3 g24848(new_n27197, new_n27196, new_n5519);
xnor_3 g24849(new_n27198, new_n27192, new_n27175);
nor_4  g24850(new_n27199, new_n27198, new_n17175);
not_3  g24851(new_n27200, new_n27199);
not_3  g24852(new_n27201, new_n27198);
xor_3  g24853(new_n27202, new_n27201, new_n5522);
xnor_3 g24854(new_n27203, new_n27190, new_n27177);
nor_4  g24855(new_n27204, new_n27203, new_n17182);
not_3  g24856(new_n27205, new_n27204);
xnor_3 g24857(new_n27206, new_n27188_1, new_n27179);
nor_4  g24858(new_n27207, new_n27206, new_n5532_1);
not_3  g24859(new_n27208, new_n27207);
xnor_3 g24860(new_n27209, new_n27206, new_n5532_1);
not_3  g24861(new_n27210, new_n27209);
nor_4  g24862(new_n27211, new_n27182, new_n27181);
xnor_3 g24863(new_n27212, new_n27211, new_n27186);
nor_4  g24864(new_n27213, new_n27212, new_n5537);
not_3  g24865(new_n27214, new_n27213);
nor_4  g24866(new_n27215, new_n15707, new_n15701);
nor_4  g24867(new_n27216, new_n15708, new_n5541);
nor_4  g24868(new_n27217, new_n27216, new_n27215);
xnor_3 g24869(new_n27218, new_n27212, new_n5537);
not_3  g24870(new_n27219, new_n27218);
nand_4 g24871(new_n27220, new_n27219, new_n27217);
nand_4 g24872(new_n27221, new_n27220, new_n27214);
nand_4 g24873(new_n27222, new_n27221, new_n27210);
nand_4 g24874(new_n27223, new_n27222, new_n27208);
not_3  g24875(new_n27224, new_n27203);
nor_4  g24876(new_n27225, new_n27224, new_n5527);
nor_4  g24877(new_n27226, new_n27225, new_n27204);
nand_4 g24878(new_n27227, new_n27226, new_n27223);
nand_4 g24879(new_n27228, new_n27227, new_n27205);
nand_4 g24880(new_n27229, new_n27228, new_n27202);
nand_4 g24881(new_n27230, new_n27229, new_n27200);
xnor_3 g24882(new_n27231, new_n27230, new_n27197);
xnor_3 g24883(new_n27232, new_n27231, new_n21395);
xnor_3 g24884(new_n27233, new_n27228, new_n27202);
nor_4  g24885(new_n27234, new_n27233, new_n20541);
not_3  g24886(new_n27235, new_n27234);
xnor_3 g24887(new_n27236, new_n27233, new_n20543);
xnor_3 g24888(new_n27237, new_n27226, new_n27223);
nor_4  g24889(new_n27238, new_n27237, new_n20546);
not_3  g24890(new_n27239, new_n27238);
xnor_3 g24891(new_n27240, new_n27237, new_n20547);
xnor_3 g24892(new_n27241, new_n27221, new_n27210);
nor_4  g24893(new_n27242, new_n27241, new_n4134_1);
not_3  g24894(new_n27243, new_n27242);
xnor_3 g24895(new_n27244, new_n27241, new_n20550);
not_3  g24896(new_n27245, new_n27215);
xnor_3 g24897(new_n27246, new_n15706, new_n15701);
nand_4 g24898(new_n27247, new_n27246, new_n5542);
nand_4 g24899(new_n27248, new_n27247, new_n27245);
xnor_3 g24900(new_n27249, new_n27219, new_n27248);
nor_4  g24901(new_n27250, new_n27249, new_n4138);
nor_4  g24902(new_n27251, new_n15709, new_n4143);
nor_4  g24903(new_n27252, new_n15722, new_n15710);
nor_4  g24904(new_n27253, new_n27252, new_n27251);
xnor_3 g24905(new_n27254, new_n27249, new_n4138);
nor_4  g24906(new_n27255, new_n27254, new_n27253);
nor_4  g24907(new_n27256, new_n27255, new_n27250);
nand_4 g24908(new_n27257, new_n27256, new_n27244);
nand_4 g24909(new_n27258, new_n27257, new_n27243);
nand_4 g24910(new_n27259, new_n27258, new_n27240);
nand_4 g24911(new_n27260, new_n27259, new_n27239);
nand_4 g24912(new_n27261, new_n27260, new_n27236);
nand_4 g24913(new_n27262, new_n27261, new_n27235);
nor_4  g24914(new_n27263, new_n27262, new_n27232);
not_3  g24915(new_n27264, new_n27232);
not_3  g24916(new_n27265, new_n27262);
nor_4  g24917(new_n27266, new_n27265, new_n27264);
nor_4  g24918(n9968, new_n27266, new_n27263);
nor_4  g24919(new_n27268, new_n25233, new_n16922);
xnor_3 g24920(new_n27269, new_n25232, new_n16923);
not_3  g24921(new_n27270, new_n25221);
nor_4  g24922(new_n27271, new_n27270, new_n16922);
not_3  g24923(new_n27272, new_n27271);
nor_4  g24924(new_n27273, new_n25221, new_n16923);
nor_4  g24925(new_n27274, new_n27273, new_n27271);
nor_4  g24926(new_n27275, new_n13638, new_n13562);
nor_4  g24927(new_n27276, new_n13707, new_n27275);
nand_4 g24928(new_n27277, new_n27276, new_n27274);
nand_4 g24929(new_n27278, new_n27277, new_n27272);
nor_4  g24930(new_n27279, new_n27278, new_n27269);
nor_4  g24931(n10009, new_n27279, new_n27268);
xnor_3 g24932(n10010, new_n26144, new_n26141);
not_3  g24933(new_n27282, new_n13288);
nand_4 g24934(new_n27283, new_n18003, new_n27282);
nand_4 g24935(new_n27284, new_n18149, new_n27283);
nor_4  g24936(new_n27285, new_n27284, new_n18090);
xnor_3 g24937(new_n27286, new_n27284, new_n18090);
nor_4  g24938(new_n27287, new_n18148, new_n18154);
nor_4  g24939(new_n27288, new_n27287, new_n27286);
nor_4  g24940(n10019, new_n27288, new_n27285);
xnor_3 g24941(n10021, new_n17885, new_n17823);
xor_3  g24942(n10055, new_n11544, new_n11531);
not_3  g24943(new_n27292, new_n12866);
xor_3  g24944(n10101, new_n27292, new_n12842);
xnor_3 g24945(n10111, new_n5218, new_n5157);
nor_4  g24946(new_n27295, n16544, new_n19353);
xor_3  g24947(new_n27296, n16544, new_n19353);
not_3  g24948(new_n27297, new_n27296);
nor_4  g24949(new_n27298, new_n19385_1, n6814);
xor_3  g24950(new_n27299, n17911, new_n10732);
not_3  g24951(new_n27300, new_n27299);
nor_4  g24952(new_n27301, new_n19389_1, n19701);
xor_3  g24953(new_n27302, n21997, new_n23667);
not_3  g24954(new_n27303, new_n27302);
nor_4  g24955(new_n27304, new_n10137, n23529);
xor_3  g24956(new_n27305, n25119, new_n3038);
not_3  g24957(new_n27306, new_n27305);
nor_4  g24958(new_n27307, n24620, new_n10139);
xor_3  g24959(new_n27308, n24620, new_n10139);
not_3  g24960(new_n27309, new_n27308);
nor_4  g24961(new_n27310, new_n10143, n5211);
nor_4  g24962(new_n27311, n18537, new_n10746);
nor_4  g24963(new_n27312, new_n10750, n7057);
not_3  g24964(new_n27313, new_n27312);
nand_4 g24965(new_n27314, new_n11387, new_n11374);
nand_4 g24966(new_n27315, new_n27314, new_n27313);
nor_4  g24967(new_n27316, new_n27315, new_n27311);
nor_4  g24968(new_n27317, new_n27316, new_n27310);
nor_4  g24969(new_n27318, new_n27317, new_n27309);
nor_4  g24970(new_n27319, new_n27318, new_n27307);
nor_4  g24971(new_n27320, new_n27319, new_n27306);
nor_4  g24972(new_n27321, new_n27320, new_n27304);
nor_4  g24973(new_n27322, new_n27321, new_n27303);
nor_4  g24974(new_n27323, new_n27322, new_n27301);
nor_4  g24975(new_n27324, new_n27323, new_n27300);
nor_4  g24976(new_n27325, new_n27324, new_n27298);
nor_4  g24977(new_n27326, new_n27325, new_n27297);
nor_4  g24978(new_n27327, new_n27326, new_n27295);
xnor_3 g24979(new_n27328, new_n27327, new_n26315);
not_3  g24980(new_n27329, new_n27327);
nor_4  g24981(new_n27330, new_n27329, new_n26324);
not_3  g24982(new_n27331, new_n27330);
nand_4 g24983(new_n27332, new_n27329, new_n26324);
xor_3  g24984(new_n27333, new_n27325, new_n27296);
nand_4 g24985(new_n27334, new_n27333, new_n26327);
xnor_3 g24986(new_n27335, new_n27333, new_n21210);
xor_3  g24987(new_n27336, new_n27323, new_n27299);
nand_4 g24988(new_n27337, new_n27336, new_n21268);
not_3  g24989(new_n27338, new_n21268);
xnor_3 g24990(new_n27339, new_n27336, new_n27338);
xor_3  g24991(new_n27340, new_n27321, new_n27303);
not_3  g24992(new_n27341, new_n27340);
nand_4 g24993(new_n27342, new_n27341, new_n21274);
xnor_3 g24994(new_n27343, new_n27340, new_n21274);
xor_3  g24995(new_n27344, new_n27319, new_n27305);
nand_4 g24996(new_n27345, new_n27344, new_n21279);
xnor_3 g24997(new_n27346, new_n27344, new_n21281);
xor_3  g24998(new_n27347, new_n27317, new_n27308);
nand_4 g24999(new_n27348, new_n27347, new_n21287_1);
nor_4  g25000(new_n27349, new_n27311, new_n27310);
xor_3  g25001(new_n27350, new_n27349, new_n27315);
nor_4  g25002(new_n27351, new_n27350, new_n21293);
xnor_3 g25003(new_n27352, new_n27350, new_n21293);
nor_4  g25004(new_n27353, new_n11388, new_n11373);
nor_4  g25005(new_n27354, new_n11415, new_n11389);
nor_4  g25006(new_n27355, new_n27354, new_n27353);
nor_4  g25007(new_n27356, new_n27355, new_n27352);
nor_4  g25008(new_n27357, new_n27356, new_n27351);
not_3  g25009(new_n27358, new_n27348);
nor_4  g25010(new_n27359, new_n27347, new_n21287_1);
nor_4  g25011(new_n27360, new_n27359, new_n27358);
nand_4 g25012(new_n27361, new_n27360, new_n27357);
nand_4 g25013(new_n27362, new_n27361, new_n27348);
nand_4 g25014(new_n27363, new_n27362, new_n27346);
nand_4 g25015(new_n27364, new_n27363, new_n27345);
nand_4 g25016(new_n27365, new_n27364, new_n27343);
nand_4 g25017(new_n27366, new_n27365, new_n27342);
nand_4 g25018(new_n27367, new_n27366, new_n27339);
nand_4 g25019(new_n27368, new_n27367, new_n27337);
nand_4 g25020(new_n27369, new_n27368, new_n27335);
nand_4 g25021(new_n27370, new_n27369, new_n27334);
not_3  g25022(new_n27371, new_n27370);
nand_4 g25023(new_n27372, new_n27371, new_n27332);
nand_4 g25024(new_n27373, new_n27372, new_n27331);
xnor_3 g25025(n10165, new_n27373, new_n27328);
xor_3  g25026(n10236, new_n15843, new_n15839);
not_3  g25027(new_n27376, new_n17703);
xor_3  g25028(n10239, new_n17729, new_n27376);
xnor_3 g25029(n10244, new_n7508, new_n7448);
not_3  g25030(new_n27379, new_n22400);
xor_3  g25031(n10261, new_n22416, new_n27379);
xor_3  g25032(n10262, new_n19346, new_n19326);
xor_3  g25033(n10287, new_n20872, new_n20871);
nor_4  g25034(new_n27383, new_n26644, new_n26585);
nor_4  g25035(new_n27384, new_n26645, new_n26586);
nor_4  g25036(new_n27385, new_n27384, new_n27383);
not_3  g25037(new_n27386, new_n26596);
nand_4 g25038(new_n27387, new_n26611, new_n26597);
nand_4 g25039(new_n27388, new_n27387, new_n27386);
xnor_3 g25040(n10295, new_n27388, new_n27385);
not_3  g25041(new_n27390, new_n18279);
xor_3  g25042(n10321, new_n18283, new_n27390);
not_3  g25043(new_n27392, new_n17731);
xor_3  g25044(n10326, new_n27392, new_n17697);
xor_3  g25045(n10327, new_n2967, new_n2954);
nor_4  g25046(new_n27395, new_n25226, new_n25221);
not_3  g25047(new_n27396, new_n27395);
nand_4 g25048(new_n27397, new_n27396, new_n25227);
xnor_3 g25049(n10330, new_n27397, new_n25213);
xnor_3 g25050(n10340, new_n26050, new_n26009);
xor_3  g25051(new_n27400, new_n20869_1, new_n24538);
xor_3  g25052(n10345, new_n27400, new_n20873);
nor_4  g25053(new_n27402, new_n23695, new_n5593_1);
nor_4  g25054(new_n27403, new_n23699, new_n5595);
not_3  g25055(new_n27404, new_n27403);
xnor_3 g25056(new_n27405, new_n23698, new_n5594);
not_3  g25057(new_n27406, new_n27405);
nor_4  g25058(new_n27407, new_n23703, new_n5596);
not_3  g25059(new_n27408, new_n27407);
xnor_3 g25060(new_n27409, new_n23705, new_n5596);
nor_4  g25061(new_n27410, new_n23708, new_n5599);
not_3  g25062(new_n27411, new_n27410);
xnor_3 g25063(new_n27412, new_n23708, new_n5599);
not_3  g25064(new_n27413, new_n27412);
nand_4 g25065(new_n27414, new_n23716, new_n5603_1);
xnor_3 g25066(new_n27415, new_n23717_1, new_n5603_1);
nand_4 g25067(new_n27416, new_n11242, new_n5607);
xnor_3 g25068(new_n27417, new_n11243, new_n5607);
nand_4 g25069(new_n27418, new_n11247, new_n5611);
xnor_3 g25070(new_n27419, new_n11248, new_n5611);
nor_4  g25071(new_n27420, new_n11254, new_n5615);
not_3  g25072(new_n27421, new_n27420);
nor_4  g25073(new_n27422, new_n11253, new_n5614);
nor_4  g25074(new_n27423, new_n27422, new_n27420);
nand_4 g25075(new_n27424, new_n24630, new_n5619);
xnor_3 g25076(new_n27425, new_n11261_1, new_n5619);
nor_4  g25077(new_n27426, new_n11269, new_n5622);
not_3  g25078(new_n27427, new_n27426);
xor_3  g25079(new_n27428, new_n11268, new_n5621);
nor_4  g25080(new_n27429, new_n11277, new_n5631);
nand_4 g25081(new_n27430, new_n27429, new_n24650);
not_3  g25082(new_n27431, new_n27430);
nor_4  g25083(new_n27432, new_n27429, new_n24650);
nor_4  g25084(new_n27433, new_n27432, new_n27431);
nand_4 g25085(new_n27434, new_n27433, new_n5629);
nand_4 g25086(new_n27435, new_n27434, new_n27430);
nand_4 g25087(new_n27436, new_n27435, new_n27428);
nand_4 g25088(new_n27437, new_n27436, new_n27427);
nand_4 g25089(new_n27438, new_n27437, new_n27425);
nand_4 g25090(new_n27439, new_n27438, new_n27424);
nand_4 g25091(new_n27440, new_n27439, new_n27423);
nand_4 g25092(new_n27441, new_n27440, new_n27421);
nand_4 g25093(new_n27442, new_n27441, new_n27419);
nand_4 g25094(new_n27443, new_n27442, new_n27418);
nand_4 g25095(new_n27444, new_n27443, new_n27417);
nand_4 g25096(new_n27445, new_n27444, new_n27416);
nand_4 g25097(new_n27446, new_n27445, new_n27415);
nand_4 g25098(new_n27447, new_n27446, new_n27414);
nand_4 g25099(new_n27448, new_n27447, new_n27413);
nand_4 g25100(new_n27449, new_n27448, new_n27411);
nand_4 g25101(new_n27450, new_n27449, new_n27409);
nand_4 g25102(new_n27451, new_n27450, new_n27408);
nand_4 g25103(new_n27452, new_n27451, new_n27406);
nand_4 g25104(new_n27453, new_n27452, new_n27404);
xor_3  g25105(new_n27454, new_n24601, new_n5592);
not_3  g25106(new_n27455, new_n27454);
nor_4  g25107(new_n27456, new_n27455, new_n27453);
nor_4  g25108(n10356, new_n27456, new_n27402);
xor_3  g25109(n10385, new_n24390, new_n24389);
not_3  g25110(new_n27459, new_n24599);
nand_4 g25111(new_n27460, new_n24686, new_n27459);
nand_4 g25112(new_n27461, new_n27460, new_n24674);
nor_4  g25113(n10387, new_n27461, new_n24596);
not_3  g25114(new_n27463, new_n24922);
xor_3  g25115(n10388, new_n24937_1, new_n27463);
xnor_3 g25116(n10390, new_n19040, new_n18988);
xor_3  g25117(n10404, new_n11401, new_n11400);
not_3  g25118(new_n27467, new_n19563);
xor_3  g25119(n10409, new_n19566, new_n27467);
xor_3  g25120(n10420, new_n19836, new_n10207);
xor_3  g25121(n10432, new_n22409, new_n8177);
xnor_3 g25122(new_n27471, new_n26138, new_n25385);
nand_4 g25123(new_n27472, new_n25388, new_n11593);
nand_4 g25124(new_n27473, new_n25736, new_n25725);
nand_4 g25125(new_n27474, new_n27473, new_n27472);
nand_4 g25126(new_n27475, new_n27474, new_n27471);
not_3  g25127(new_n27476, new_n27475);
nor_4  g25128(new_n27477, new_n27474, new_n27471);
nor_4  g25129(new_n27478, new_n27477, new_n27476);
xnor_3 g25130(new_n27479, new_n27478, new_n13854);
nor_4  g25131(new_n27480, new_n25737, new_n13861);
nor_4  g25132(new_n27481, new_n25748, new_n25738_1);
nor_4  g25133(new_n27482, new_n27481, new_n27480);
nor_4  g25134(new_n27483, new_n27482, new_n27479);
not_3  g25135(new_n27484, new_n27479);
not_3  g25136(new_n27485, new_n27482);
nor_4  g25137(new_n27486, new_n27485, new_n27484);
nor_4  g25138(n10484, new_n27486, new_n27483);
not_3  g25139(new_n27488, new_n13671);
xor_3  g25140(n10489, new_n13694, new_n27488);
xor_3  g25141(n10525, new_n16402, new_n3959_1);
not_3  g25142(new_n27491, new_n21597);
nor_4  g25143(new_n27492, new_n21589, new_n21587);
xor_3  g25144(n10540, new_n27492, new_n27491);
not_3  g25145(new_n27494, new_n19682);
xor_3  g25146(n10561, new_n19717, new_n27494);
xnor_3 g25147(n10564, new_n19044_1, new_n18973);
not_3  g25148(new_n27497, new_n12071);
xor_3  g25149(n10588, new_n27497, new_n12070);
not_3  g25150(new_n27499, new_n12072_1);
xor_3  g25151(n10595, new_n12073, new_n27499);
xor_3  g25152(n10617, new_n25895, new_n25878);
xnor_3 g25153(n10628, new_n15083, new_n15005);
xnor_3 g25154(new_n27503, new_n12802, new_n6667);
not_3  g25155(new_n27504, new_n27503);
not_3  g25156(new_n27505, new_n12812_1);
nand_4 g25157(new_n27506, new_n27505, new_n6672);
xnor_3 g25158(new_n27507, new_n12812_1, new_n6672);
nor_4  g25159(new_n27508, new_n12817, new_n6680);
not_3  g25160(new_n27509, new_n27508);
nor_4  g25161(new_n27510, new_n12818, new_n6681);
nor_4  g25162(new_n27511, new_n27510, new_n27508);
nor_4  g25163(new_n27512, new_n6725, new_n6687);
nor_4  g25164(new_n27513, new_n27512, new_n6741);
not_3  g25165(new_n27514, new_n27513);
not_3  g25166(new_n27515, new_n27512);
xor_3  g25167(new_n27516, new_n27515, new_n6742);
nand_4 g25168(new_n27517, new_n27516, new_n6696);
nand_4 g25169(new_n27518, new_n27517, new_n27514);
nand_4 g25170(new_n27519, new_n27518, new_n27511);
nand_4 g25171(new_n27520, new_n27519, new_n27509);
nand_4 g25172(new_n27521, new_n27520, new_n27507);
nand_4 g25173(new_n27522, new_n27521, new_n27506);
xor_3  g25174(n10647, new_n27522, new_n27504);
nand_4 g25175(new_n27524, new_n9924, new_n9917_1);
nor_4  g25176(new_n27525, new_n24253, new_n16353);
nor_4  g25177(new_n27526, new_n3983_1, new_n3895);
nor_4  g25178(new_n27527, new_n27526, new_n27525);
nor_4  g25179(new_n27528, new_n16348, new_n24255);
nand_4 g25180(new_n27529, new_n27528, new_n27527);
not_3  g25181(new_n27530, new_n27529);
nor_4  g25182(new_n27531, new_n27530, new_n27524);
not_3  g25183(new_n27532, new_n27524);
nor_4  g25184(new_n27533, new_n27529, new_n27532);
nor_4  g25185(new_n27534, new_n27533, new_n27531);
xor_3  g25186(new_n27535, new_n16348, new_n24256);
not_3  g25187(new_n27536, new_n27535);
xnor_3 g25188(new_n27537, new_n27536, new_n27527);
nand_4 g25189(new_n27538, new_n27537, new_n9925);
nand_4 g25190(new_n27539, new_n3984_1, new_n3823);
nand_4 g25191(new_n27540, new_n4072, new_n3985);
nand_4 g25192(new_n27541, new_n27540, new_n27539);
not_3  g25193(new_n27542, new_n9925);
xnor_3 g25194(new_n27543, new_n27537, new_n27542);
nand_4 g25195(new_n27544, new_n27543, new_n27541);
nand_4 g25196(new_n27545, new_n27544, new_n27538);
not_3  g25197(new_n27546, new_n27545);
xnor_3 g25198(n10653, new_n27546, new_n27534);
xor_3  g25199(n10692, new_n10834_1, new_n10833);
xor_3  g25200(n10694, new_n17945, new_n4842);
xor_3  g25201(n10701, new_n24770, new_n24739);
not_3  g25202(new_n27551, new_n7185);
xor_3  g25203(n10756, new_n27551, new_n7165);
not_3  g25204(new_n27553, new_n3650);
nor_4  g25205(new_n27554, new_n21610, n5101);
nor_4  g25206(new_n27555, new_n19461, new_n27554);
not_3  g25207(new_n27556, new_n19474);
not_3  g25208(new_n27557, new_n19472_1);
nand_4 g25209(new_n27558, new_n23605, new_n27557);
nand_4 g25210(new_n27559, new_n27558, new_n27556);
nor_4  g25211(new_n27560, new_n27559, new_n19466);
not_3  g25212(new_n27561, new_n27560);
nand_4 g25213(new_n27562, new_n27559, new_n19417);
nand_4 g25214(new_n27563, new_n27562, new_n19463);
nand_4 g25215(new_n27564, new_n27563, new_n27561);
not_3  g25216(new_n27565, new_n27564);
nor_4  g25217(new_n27566, new_n27565, new_n27555);
xnor_3 g25218(new_n27567, new_n27566, new_n27553);
xnor_3 g25219(new_n27568, new_n27564, new_n27555);
not_3  g25220(new_n27569, new_n27568);
nor_4  g25221(new_n27570, new_n27569, new_n3548);
not_3  g25222(new_n27571, new_n27570);
nor_4  g25223(new_n27572, new_n27568, new_n3549);
not_3  g25224(new_n27573, new_n27572);
xnor_3 g25225(new_n27574, new_n27559, new_n19466);
nor_4  g25226(new_n27575, new_n27574, new_n3460_1);
not_3  g25227(new_n27576, new_n27575);
xnor_3 g25228(new_n27577, new_n27574, new_n3460_1);
not_3  g25229(new_n27578, new_n27577);
not_3  g25230(new_n27579, new_n23598);
nand_4 g25231(new_n27580, new_n23597, new_n19518);
nand_4 g25232(new_n27581, new_n27580, n15602);
nand_4 g25233(new_n27582, new_n27581, new_n27579);
nor_4  g25234(new_n27583, new_n27582, new_n19475);
nor_4  g25235(new_n27584, new_n23605, new_n19476);
nor_4  g25236(new_n27585, new_n27584, new_n27583);
nor_4  g25237(new_n27586, new_n27585, new_n3466);
not_3  g25238(new_n27587, new_n23614);
nor_4  g25239(new_n27588, new_n23652, new_n27587);
nor_4  g25240(new_n27589, new_n27588, new_n23609);
nor_4  g25241(new_n27590, new_n27589, new_n23607);
nor_4  g25242(new_n27591, new_n27590, new_n27586);
nand_4 g25243(new_n27592, new_n27591, new_n27578);
nand_4 g25244(new_n27593, new_n27592, new_n27576);
nand_4 g25245(new_n27594, new_n27593, new_n27573);
nand_4 g25246(new_n27595, new_n27594, new_n27571);
xnor_3 g25247(n10775, new_n27595, new_n27567);
not_3  g25248(new_n27597, new_n25786);
xor_3  g25249(n10780, new_n27597, new_n25778);
xor_3  g25250(new_n27599, n17095, n1689);
nor_4  g25251(new_n27600, n22591, n22274);
not_3  g25252(new_n27601, new_n27600);
nand_4 g25253(new_n27602, n26167, n24129);
nand_4 g25254(new_n27603, n22591, n22274);
not_3  g25255(new_n27604, new_n27603);
nor_4  g25256(new_n27605, new_n27604, new_n27600);
nand_4 g25257(new_n27606, new_n27605, new_n27602);
nand_4 g25258(new_n27607, new_n27606, new_n27601);
nor_4  g25259(new_n27608, new_n27607, new_n27599);
nand_4 g25260(new_n27609, new_n27607, new_n27599);
not_3  g25261(new_n27610, new_n27609);
nor_4  g25262(new_n27611, new_n27610, new_n27608);
xnor_3 g25263(new_n27612, new_n27611, n21749);
nand_4 g25264(new_n27613, new_n10673, n21138);
nand_4 g25265(new_n27614, new_n27613, new_n25424);
not_3  g25266(new_n27615, new_n27614);
xor_3  g25267(new_n27616, new_n27605, new_n27602);
xor_3  g25268(new_n27617, new_n27613, n7769);
nor_4  g25269(new_n27618, new_n27617, new_n27616);
nor_4  g25270(new_n27619, new_n27618, new_n27615);
xnor_3 g25271(new_n27620, new_n27619, new_n27612);
xnor_3 g25272(new_n27621, new_n27620, new_n22628);
not_3  g25273(new_n27622, new_n27616);
not_3  g25274(new_n27623, new_n27617);
xor_3  g25275(new_n27624, new_n27623, new_n27622);
not_3  g25276(new_n27625, new_n27624);
nor_4  g25277(new_n27626, new_n27625, new_n22642);
nor_4  g25278(new_n27627, new_n10674, new_n10672);
not_3  g25279(new_n27628, new_n27627);
xnor_3 g25280(new_n27629, new_n27624, new_n22633);
nor_4  g25281(new_n27630, new_n27629, new_n27628);
nor_4  g25282(new_n27631, new_n27630, new_n27626);
xor_3  g25283(n10817, new_n27631, new_n27621);
not_3  g25284(new_n27633, new_n26613);
nor_4  g25285(new_n27634, new_n26617, new_n27633);
nor_4  g25286(new_n27635, new_n26631, new_n26626);
nor_4  g25287(new_n27636, new_n27635, new_n27634);
nand_4 g25288(new_n27637, new_n27636, new_n26624);
not_3  g25289(new_n27638, new_n27637);
nor_4  g25290(new_n27639, new_n27638, new_n9127);
not_3  g25291(new_n27640, new_n26634);
nand_4 g25292(new_n27641, new_n26642, new_n26638);
nand_4 g25293(new_n27642, new_n27641, new_n27640);
xnor_3 g25294(new_n27643, new_n27637, new_n26635);
nor_4  g25295(new_n27644, new_n27643, new_n27642);
nor_4  g25296(n10834, new_n27644, new_n27639);
not_3  g25297(new_n27646, new_n26930_1);
not_3  g25298(new_n27647, new_n26931);
not_3  g25299(new_n27648, new_n26936);
nor_4  g25300(new_n27649, new_n26826, new_n6520);
nor_4  g25301(new_n27650, new_n27649, new_n26936);
not_3  g25302(new_n27651, new_n26938);
not_3  g25303(new_n27652, new_n26939);
nand_4 g25304(new_n27653, new_n27652, new_n27651);
nand_4 g25305(new_n27654, new_n27653, new_n27650);
nand_4 g25306(new_n27655, new_n27654, new_n27648);
xnor_3 g25307(new_n27656, new_n26822, new_n6517);
nor_4  g25308(new_n27657, new_n27656, new_n27655);
nor_4  g25309(new_n27658, new_n27657, new_n26934);
nand_4 g25310(new_n27659, new_n27658, new_n27647);
nand_4 g25311(new_n27660, new_n27659, new_n27646);
xnor_3 g25312(n10851, new_n27660, new_n26928);
xnor_3 g25313(n10874, new_n26375_1, new_n26366);
xnor_3 g25314(new_n27663, new_n27161, new_n27150);
xnor_3 g25315(n10924, new_n27663, new_n9525);
not_3  g25316(new_n27665, new_n13375);
nor_4  g25317(new_n27666, new_n13378, new_n27665);
nor_4  g25318(new_n27667, new_n13459, new_n13380);
nor_4  g25319(n10943, new_n27667, new_n27666);
xnor_3 g25320(n10961, new_n14394, new_n14357);
not_3  g25321(new_n27670, new_n12724);
xor_3  g25322(n11005, new_n12737, new_n27670);
xnor_3 g25323(n11023, new_n26107_1, new_n26096_1);
nor_4  g25324(new_n27673, new_n22226, new_n8571);
xnor_3 g25325(new_n27674, new_n22226, new_n8571);
nor_4  g25326(new_n27675, new_n22232, new_n8578);
xnor_3 g25327(new_n27676, new_n22232, new_n8578);
nand_4 g25328(new_n27677, new_n20606, new_n8588);
not_3  g25329(new_n27678, new_n27677);
nor_4  g25330(new_n27679, new_n20606, new_n8588);
nor_4  g25331(new_n27680, new_n27679, new_n27678);
nand_4 g25332(new_n27681, new_n14621, new_n14589);
nand_4 g25333(new_n27682, new_n27681, new_n27680);
nand_4 g25334(new_n27683, new_n27682, new_n27677);
nor_4  g25335(new_n27684, new_n27683, new_n27676);
nor_4  g25336(new_n27685, new_n27684, new_n27675);
nor_4  g25337(new_n27686, new_n27685, new_n27674);
nor_4  g25338(new_n27687, new_n27686, new_n27673);
nor_4  g25339(new_n27688, new_n27687, new_n8546);
not_3  g25340(new_n27689, new_n27688);
nor_4  g25341(new_n27690, new_n27689, new_n22264);
not_3  g25342(new_n27691, new_n27687);
nor_4  g25343(new_n27692, new_n27691, new_n25597);
nor_4  g25344(new_n27693, new_n27692, new_n27688);
xnor_3 g25345(new_n27694, new_n27693, new_n22264);
not_3  g25346(new_n27695, new_n27694);
nand_4 g25347(new_n27696, new_n27695, new_n27085);
xnor_3 g25348(new_n27697, new_n27694, new_n27085);
not_3  g25349(new_n27698, new_n27674);
not_3  g25350(new_n27699, new_n27685);
nor_4  g25351(new_n27700, new_n27699, new_n27698);
nor_4  g25352(new_n27701, new_n27700, new_n27686);
nand_4 g25353(new_n27702, new_n27701, new_n27118);
xnor_3 g25354(new_n27703, new_n27701, new_n27117);
not_3  g25355(new_n27704, new_n27676);
not_3  g25356(new_n27705, new_n27683);
nor_4  g25357(new_n27706, new_n27705, new_n27704);
nor_4  g25358(new_n27707, new_n27706, new_n27684);
nand_4 g25359(new_n27708, new_n27707, new_n27122);
not_3  g25360(new_n27709, new_n27708);
nor_4  g25361(new_n27710, new_n27707, new_n27122);
nor_4  g25362(new_n27711, new_n27710, new_n27709);
xnor_3 g25363(new_n27712, new_n27681, new_n27680);
nand_4 g25364(new_n27713, new_n27712, new_n27127);
xnor_3 g25365(new_n27714, new_n27712, new_n21557);
not_3  g25366(new_n27715, new_n14625);
nand_4 g25367(new_n27716, new_n14683, new_n14630);
nand_4 g25368(new_n27717, new_n27716, new_n27715);
nand_4 g25369(new_n27718, new_n27717, new_n27714);
nand_4 g25370(new_n27719, new_n27718, new_n27713);
nand_4 g25371(new_n27720, new_n27719, new_n27711);
nand_4 g25372(new_n27721, new_n27720, new_n27708);
nand_4 g25373(new_n27722, new_n27721, new_n27703);
nand_4 g25374(new_n27723, new_n27722, new_n27702);
nand_4 g25375(new_n27724, new_n27723, new_n27697);
nand_4 g25376(new_n27725, new_n27724, new_n27696);
nand_4 g25377(new_n27726, new_n27725, new_n27690);
xnor_3 g25378(new_n27727, new_n27725, new_n27690);
nand_4 g25379(new_n27728, new_n27727, new_n27143);
nand_4 g25380(n11025, new_n27728, new_n27726);
xor_3  g25381(new_n27730, new_n20158, new_n10327_1);
nand_4 g25382(new_n27731, new_n20163, n13775);
xnor_3 g25383(new_n27732, new_n20163, new_n8045);
nand_4 g25384(new_n27733, new_n20166, n1293);
xnor_3 g25385(new_n27734, new_n20166, new_n10335);
nand_4 g25386(new_n27735, new_n20169_1, n19042);
nand_4 g25387(new_n27736, new_n23434_1, new_n23430_1);
nand_4 g25388(new_n27737, new_n27736, new_n27735);
nand_4 g25389(new_n27738, new_n27737, new_n27734);
nand_4 g25390(new_n27739, new_n27738, new_n27733);
nand_4 g25391(new_n27740, new_n27739, new_n27732);
nand_4 g25392(new_n27741, new_n27740, new_n27731);
xnor_3 g25393(new_n27742, new_n27741, new_n27730);
not_3  g25394(new_n27743, new_n23437);
nor_4  g25395(new_n27744, new_n27743, n26752);
not_3  g25396(new_n27745, new_n27744);
nor_4  g25397(new_n27746, new_n27745, n4590);
not_3  g25398(new_n27747, new_n27746);
nor_4  g25399(new_n27748, new_n27747, n25464);
xor_3  g25400(new_n27749, new_n27748, new_n7393);
not_3  g25401(new_n27750, new_n27749);
nor_4  g25402(new_n27751, new_n27750, new_n10510);
nor_4  g25403(new_n27752, new_n27749, new_n13390);
nor_4  g25404(new_n27753, new_n27752, new_n27751);
xor_3  g25405(new_n27754, new_n27746, new_n14823);
nor_4  g25406(new_n27755, new_n27754, new_n10522);
not_3  g25407(new_n27756, new_n27755);
not_3  g25408(new_n27757, new_n27754);
nor_4  g25409(new_n27758, new_n27757, new_n10517);
nor_4  g25410(new_n27759, new_n27758, new_n27755);
xor_3  g25411(new_n27760, new_n27744, new_n14827_1);
nor_4  g25412(new_n27761, new_n27760, new_n10527);
not_3  g25413(new_n27762, new_n27761);
not_3  g25414(new_n27763, new_n27760);
xor_3  g25415(new_n27764, new_n27763, new_n10527);
not_3  g25416(new_n27765, new_n27764);
nor_4  g25417(new_n27766, new_n23438, new_n10533);
not_3  g25418(new_n27767, new_n27766);
not_3  g25419(new_n27768, new_n23440);
nand_4 g25420(new_n27769, new_n23443, new_n27768);
nand_4 g25421(new_n27770, new_n27769, new_n27767);
nand_4 g25422(new_n27771, new_n27770, new_n27765);
nand_4 g25423(new_n27772, new_n27771, new_n27762);
nand_4 g25424(new_n27773, new_n27772, new_n27759);
nand_4 g25425(new_n27774, new_n27773, new_n27756);
xnor_3 g25426(new_n27775, new_n27774, new_n27753);
xnor_3 g25427(new_n27776, new_n27775, new_n27742);
not_3  g25428(new_n27777, new_n27732);
xnor_3 g25429(new_n27778, new_n27739, new_n27777);
not_3  g25430(new_n27779, new_n27778);
not_3  g25431(new_n27780, new_n27772);
xnor_3 g25432(new_n27781, new_n27780, new_n27759);
nand_4 g25433(new_n27782, new_n27781, new_n27779);
xnor_3 g25434(new_n27783, new_n27781, new_n27778);
xnor_3 g25435(new_n27784, new_n27737, new_n27734);
xnor_3 g25436(new_n27785, new_n27770, new_n27764);
nand_4 g25437(new_n27786, new_n27785, new_n27784);
not_3  g25438(new_n27787, new_n27786);
nor_4  g25439(new_n27788, new_n27785, new_n27784);
nor_4  g25440(new_n27789, new_n27788, new_n27787);
not_3  g25441(new_n27790, new_n23449);
nand_4 g25442(new_n27791, new_n23455, new_n23450_1);
nand_4 g25443(new_n27792, new_n27791, new_n27790);
nand_4 g25444(new_n27793, new_n27792, new_n27789);
nand_4 g25445(new_n27794, new_n27793, new_n27786);
nand_4 g25446(new_n27795, new_n27794, new_n27783);
nand_4 g25447(new_n27796, new_n27795, new_n27782);
xnor_3 g25448(n11063, new_n27796, new_n27776);
not_3  g25449(new_n27798, new_n24926);
xor_3  g25450(n11078, new_n24935, new_n27798);
not_3  g25451(new_n27800, new_n25776);
xor_3  g25452(n11080, new_n25788, new_n27800);
not_3  g25453(new_n27802, new_n16806);
xor_3  g25454(n11094, new_n27802, new_n16791);
not_3  g25455(new_n27804, new_n27357);
xor_3  g25456(n11101, new_n27360, new_n27804);
xor_3  g25457(new_n27806, new_n25888, new_n17537);
xor_3  g25458(n11103, new_n27806, new_n25891);
not_3  g25459(new_n27808, new_n7691);
xor_3  g25460(n11120, new_n7725, new_n27808);
xor_3  g25461(n11127, new_n5730, new_n5724);
not_3  g25462(new_n27811, new_n18286);
xor_3  g25463(n11132, new_n27811, new_n18285);
xnor_3 g25464(n11134, new_n13452, new_n13397);
xor_3  g25465(n11138, new_n4056, new_n4052);
xor_3  g25466(n11182, new_n12621_1, new_n12607_1);
xnor_3 g25467(n11234, new_n16816, new_n16755);
nor_4  g25468(new_n27817, new_n26588, new_n22842);
nor_4  g25469(new_n27818, new_n26595, new_n22843_1);
nor_4  g25470(new_n27819, new_n27818, new_n27817);
nand_4 g25471(new_n27820, new_n26201, new_n22853);
nand_4 g25472(new_n27821, new_n26224_1, new_n26202);
nand_4 g25473(new_n27822, new_n27821, new_n27820);
xnor_3 g25474(n11245, new_n27822, new_n27819);
not_3  g25475(new_n27824, new_n10302);
xor_3  g25476(n11261, new_n10320, new_n27824);
xnor_3 g25477(n11275, new_n27794, new_n27783);
not_3  g25478(new_n27827, new_n16426);
nand_4 g25479(n11290, new_n27827, new_n16344);
not_3  g25480(new_n27829, new_n11280);
xor_3  g25481(n11313, new_n11283, new_n27829);
not_3  g25482(new_n27831, new_n20596);
nor_4  g25483(new_n27832, new_n20593, new_n20592);
xnor_3 g25484(n11325, new_n27832, new_n27831);
not_3  g25485(new_n27834, new_n16870);
xor_3  g25486(n11326, new_n16873, new_n27834);
not_3  g25487(new_n27836, new_n20845);
xor_3  g25488(n11330, new_n20881, new_n27836);
xnor_3 g25489(n11347, new_n13446, new_n13412);
not_3  g25490(new_n27839, new_n27428);
xor_3  g25491(n11348, new_n27435, new_n27839);
xnor_3 g25492(n11352, new_n18422, new_n18414_1);
nor_4  g25493(new_n27842, new_n9752, n3324);
xor_3  g25494(new_n27843, n22442, new_n19353);
not_3  g25495(new_n27844, new_n27843);
nor_4  g25496(new_n27845, n17911, new_n9834);
nand_4 g25497(new_n27846, new_n19389_1, n5400);
nand_4 g25498(new_n27847, new_n21129, new_n21122);
nand_4 g25499(new_n27848, new_n27847, new_n27846);
xor_3  g25500(new_n27849, n17911, new_n9834);
nand_4 g25501(new_n27850, new_n27849, new_n27848);
not_3  g25502(new_n27851, new_n27850);
nor_4  g25503(new_n27852, new_n27851, new_n27845);
nor_4  g25504(new_n27853, new_n27852, new_n27844);
nor_4  g25505(new_n27854, new_n27853, new_n27842);
nor_4  g25506(new_n27855, new_n21800_1, new_n21794);
nor_4  g25507(new_n27856, new_n27855, new_n9075);
nand_4 g25508(new_n27857, new_n21800_1, new_n21794);
nand_4 g25509(new_n27858, new_n27857, new_n9075);
not_3  g25510(new_n27859, new_n27858);
nor_4  g25511(new_n27860, new_n27859, new_n27856);
xnor_3 g25512(new_n27861, new_n27860, new_n27854);
nand_4 g25513(new_n27862, new_n27854, new_n21807);
not_3  g25514(new_n27863, new_n27854);
nand_4 g25515(new_n27864, new_n27863, new_n21847);
xor_3  g25516(new_n27865, new_n27852, new_n27844);
nor_4  g25517(new_n27866, new_n27865, new_n21811);
xnor_3 g25518(new_n27867, new_n27865, new_n21811);
xor_3  g25519(new_n27868, new_n27849, new_n27848);
nand_4 g25520(new_n27869, new_n27868, new_n21815);
xnor_3 g25521(new_n27870, new_n27868, new_n21815);
not_3  g25522(new_n27871, new_n27870);
nand_4 g25523(new_n27872, new_n21130, new_n21121);
not_3  g25524(new_n27873, new_n21131);
not_3  g25525(new_n27874, new_n21145);
nand_4 g25526(new_n27875, new_n27874, new_n21135);
nand_4 g25527(new_n27876, new_n27875, new_n27873);
nand_4 g25528(new_n27877, new_n27876, new_n27872);
nand_4 g25529(new_n27878, new_n27877, new_n27871);
nand_4 g25530(new_n27879, new_n27878, new_n27869);
nor_4  g25531(new_n27880, new_n27879, new_n27867);
nor_4  g25532(new_n27881, new_n27880, new_n27866);
nand_4 g25533(new_n27882, new_n27881, new_n27864);
nand_4 g25534(new_n27883, new_n27882, new_n27862);
xnor_3 g25535(n11375, new_n27883, new_n27861);
xor_3  g25536(n11379, new_n15114, new_n8443);
nor_4  g25537(new_n27886, new_n10324, n2570);
nor_4  g25538(new_n27887, new_n20152, new_n20121);
nor_4  g25539(new_n27888, new_n27887, new_n27886);
xor_3  g25540(new_n27889, new_n27888, new_n14468);
nand_4 g25541(new_n27890, new_n20154, new_n14412_1);
not_3  g25542(new_n27891, new_n27890);
nor_4  g25543(new_n27892, new_n20202, new_n20159);
nor_4  g25544(new_n27893, new_n27892, new_n20155);
nor_4  g25545(new_n27894, new_n27893, new_n27891);
xnor_3 g25546(new_n27895, new_n27894, new_n27889);
xnor_3 g25547(new_n27896, new_n27895, new_n7429);
not_3  g25548(new_n27897, new_n27896);
nor_4  g25549(new_n27898, new_n20200, new_n7433);
not_3  g25550(new_n27899, new_n27898);
nand_4 g25551(new_n27900, new_n20245, new_n20201);
nand_4 g25552(new_n27901, new_n27900, new_n27899);
xnor_3 g25553(n11386, new_n27901, new_n27897);
not_3  g25554(new_n27903, new_n23631);
xor_3  g25555(n11391, new_n23644, new_n27903);
xnor_3 g25556(n11398, new_n26180_1, new_n26179_1);
xor_3  g25557(n11403, new_n15496_1, new_n15494);
not_3  g25558(new_n27907, new_n14792);
xor_3  g25559(n11419, new_n27907, new_n14783);
not_3  g25560(new_n27909, new_n23395);
xor_3  g25561(n11439, new_n23416, new_n27909);
xor_3  g25562(new_n27911, n7569, n2570);
nand_4 g25563(new_n27912, new_n19973, new_n13804);
xor_3  g25564(new_n27913, n19033, n17037);
nor_4  g25565(new_n27914, n5386, n655);
not_3  g25566(new_n27915, new_n27914);
xor_3  g25567(new_n27916, n5386, n655);
nor_4  g25568(new_n27917, n26191, n18145);
not_3  g25569(new_n27918, new_n27917);
xor_3  g25570(new_n27919, n26191, n18145);
nor_4  g25571(new_n27920, n26512, n10712);
not_3  g25572(new_n27921, new_n27920);
xor_3  g25573(new_n27922, n26512, n10712);
nor_4  g25574(new_n27923, n25126, n19575);
not_3  g25575(new_n27924, new_n27923);
xor_3  g25576(new_n27925, n25126, n19575);
nand_4 g25577(new_n27926, n19608, n15378);
not_3  g25578(new_n27927, new_n27926);
nor_4  g25579(new_n27928, n19608, n15378);
nor_4  g25580(new_n27929, n17095, n1689);
not_3  g25581(new_n27930, new_n27929);
nand_4 g25582(new_n27931, new_n27609, new_n27930);
nor_4  g25583(new_n27932, new_n27931, new_n27928);
nor_4  g25584(new_n27933, new_n27932, new_n27927);
nand_4 g25585(new_n27934, new_n27933, new_n27925);
nand_4 g25586(new_n27935, new_n27934, new_n27924);
nand_4 g25587(new_n27936, new_n27935, new_n27922);
nand_4 g25588(new_n27937, new_n27936, new_n27921);
nand_4 g25589(new_n27938, new_n27937, new_n27919);
nand_4 g25590(new_n27939, new_n27938, new_n27918);
nand_4 g25591(new_n27940, new_n27939, new_n27916);
nand_4 g25592(new_n27941, new_n27940, new_n27915);
nand_4 g25593(new_n27942, new_n27941, new_n27913);
nand_4 g25594(new_n27943, new_n27942, new_n27912);
not_3  g25595(new_n27944, new_n27943);
xor_3  g25596(new_n27945, new_n27944, new_n27911);
nand_4 g25597(new_n27946, new_n27945, new_n25381_1);
xnor_3 g25598(new_n27947, new_n27945, n10514);
not_3  g25599(new_n27948, new_n27941);
xnor_3 g25600(new_n27949, new_n27948, new_n27913);
nand_4 g25601(new_n27950, new_n27949, n18649);
xor_3  g25602(new_n27951, new_n27949, n18649);
not_3  g25603(new_n27952, new_n27939);
xor_3  g25604(new_n27953, new_n27952, new_n27916);
nor_4  g25605(new_n27954, new_n27953, new_n25393);
not_3  g25606(new_n27955, new_n27954);
not_3  g25607(new_n27956, new_n27916);
xor_3  g25608(new_n27957, new_n27952, new_n27956);
nor_4  g25609(new_n27958, new_n27957, n6218);
nor_4  g25610(new_n27959, new_n27958, new_n27954);
xnor_3 g25611(new_n27960, new_n27937, new_n27919);
not_3  g25612(new_n27961, new_n27960);
nand_4 g25613(new_n27962, new_n27961, n20470);
xor_3  g25614(new_n27963, new_n27961, n20470);
not_3  g25615(new_n27964, new_n27922);
xnor_3 g25616(new_n27965, new_n27935, new_n27964);
nand_4 g25617(new_n27966, new_n27965, n21222);
xnor_3 g25618(new_n27967, new_n27965, new_n25403);
not_3  g25619(new_n27968, new_n27925);
xnor_3 g25620(new_n27969, new_n27933, new_n27968);
nand_4 g25621(new_n27970, new_n27969, n9832);
xnor_3 g25622(new_n27971, new_n27969, new_n25407);
nor_4  g25623(new_n27972, new_n27928, new_n27927);
not_3  g25624(new_n27973, new_n27972);
xnor_3 g25625(new_n27974, new_n27973, new_n27931);
nor_4  g25626(new_n27975, new_n27974, n1558);
xnor_3 g25627(new_n27976, new_n27974, n1558);
nor_4  g25628(new_n27977, new_n27611, n21749);
nor_4  g25629(new_n27978, new_n27619, new_n27612);
nor_4  g25630(new_n27979, new_n27978, new_n27977);
nor_4  g25631(new_n27980, new_n27979, new_n27976);
nor_4  g25632(new_n27981, new_n27980, new_n27975);
nand_4 g25633(new_n27982, new_n27981, new_n27971);
nand_4 g25634(new_n27983, new_n27982, new_n27970);
nand_4 g25635(new_n27984, new_n27983, new_n27967);
nand_4 g25636(new_n27985, new_n27984, new_n27966);
nand_4 g25637(new_n27986, new_n27985, new_n27963);
nand_4 g25638(new_n27987, new_n27986, new_n27962);
nand_4 g25639(new_n27988, new_n27987, new_n27959);
nand_4 g25640(new_n27989, new_n27988, new_n27955);
nand_4 g25641(new_n27990, new_n27989, new_n27951);
nand_4 g25642(new_n27991, new_n27990, new_n27950);
not_3  g25643(new_n27992, new_n27991);
nand_4 g25644(new_n27993, new_n27992, new_n27947);
nand_4 g25645(new_n27994, new_n27993, new_n27946);
nor_4  g25646(new_n27995, n7569, n2570);
not_3  g25647(new_n27996, new_n27911);
nor_4  g25648(new_n27997, new_n27944, new_n27996);
nor_4  g25649(new_n27998, new_n27997, new_n27995);
xnor_3 g25650(new_n27999, new_n27998, new_n27994);
not_3  g25651(new_n28000, new_n27748);
nor_4  g25652(new_n28001, new_n28000, n3795);
not_3  g25653(new_n28002, new_n28001);
nor_4  g25654(new_n28003, new_n28002, n6105);
xor_3  g25655(new_n28004, new_n28003, new_n13378);
xor_3  g25656(new_n28005, new_n28001, n6105);
nand_4 g25657(new_n28006, new_n28005, new_n10422);
xnor_3 g25658(new_n28007, new_n28005, new_n10421);
not_3  g25659(new_n28008, new_n27752);
nand_4 g25660(new_n28009, new_n27774, new_n27753);
nand_4 g25661(new_n28010, new_n28009, new_n28008);
nand_4 g25662(new_n28011, new_n28010, new_n28007);
nand_4 g25663(new_n28012, new_n28011, new_n28006);
xnor_3 g25664(new_n28013, new_n28012, new_n28004);
xnor_3 g25665(new_n28014, new_n28013, new_n27999);
not_3  g25666(new_n28015, new_n28014);
xnor_3 g25667(new_n28016, new_n27991, new_n27947);
xnor_3 g25668(new_n28017, new_n28010, new_n28007);
nor_4  g25669(new_n28018, new_n28017, new_n28016);
xnor_3 g25670(new_n28019, new_n27992, new_n27947);
not_3  g25671(new_n28020, new_n28017);
xnor_3 g25672(new_n28021, new_n28020, new_n28019);
not_3  g25673(new_n28022, new_n27775);
not_3  g25674(new_n28023, new_n27951);
xnor_3 g25675(new_n28024, new_n27989, new_n28023);
nand_4 g25676(new_n28025, new_n28024, new_n28022);
xnor_3 g25677(new_n28026, new_n28024, new_n27775);
xnor_3 g25678(new_n28027, new_n27987, new_n27959);
not_3  g25679(new_n28028, new_n28027);
nand_4 g25680(new_n28029, new_n28028, new_n27781);
xnor_3 g25681(new_n28030, new_n28027, new_n27781);
not_3  g25682(new_n28031, new_n27963);
xnor_3 g25683(new_n28032, new_n27985, new_n28031);
nand_4 g25684(new_n28033, new_n28032, new_n27785);
not_3  g25685(new_n28034, new_n27785);
xnor_3 g25686(new_n28035, new_n28032, new_n28034);
not_3  g25687(new_n28036, new_n27967);
xnor_3 g25688(new_n28037, new_n27983, new_n28036);
nand_4 g25689(new_n28038, new_n28037, new_n23444);
xnor_3 g25690(new_n28039, new_n28037, new_n23448);
not_3  g25691(new_n28040, new_n27981);
xnor_3 g25692(new_n28041, new_n28040, new_n27971);
nand_4 g25693(new_n28042, new_n28041, new_n23452);
xnor_3 g25694(new_n28043, new_n28041, new_n22598);
xnor_3 g25695(new_n28044, new_n27979, new_n27976);
nand_4 g25696(new_n28045, new_n28044, new_n22623_1);
nor_4  g25697(new_n28046, new_n27620, new_n22628);
nor_4  g25698(new_n28047, new_n27631, new_n27621);
nor_4  g25699(new_n28048, new_n28047, new_n28046);
not_3  g25700(new_n28049, new_n28045);
nor_4  g25701(new_n28050, new_n28044, new_n22623_1);
nor_4  g25702(new_n28051, new_n28050, new_n28049);
nand_4 g25703(new_n28052, new_n28051, new_n28048);
nand_4 g25704(new_n28053, new_n28052, new_n28045);
nand_4 g25705(new_n28054, new_n28053, new_n28043);
nand_4 g25706(new_n28055, new_n28054, new_n28042);
nand_4 g25707(new_n28056, new_n28055, new_n28039);
nand_4 g25708(new_n28057, new_n28056, new_n28038);
nand_4 g25709(new_n28058, new_n28057, new_n28035);
nand_4 g25710(new_n28059, new_n28058, new_n28033);
nand_4 g25711(new_n28060, new_n28059, new_n28030);
nand_4 g25712(new_n28061, new_n28060, new_n28029);
nand_4 g25713(new_n28062, new_n28061, new_n28026);
nand_4 g25714(new_n28063, new_n28062, new_n28025);
not_3  g25715(new_n28064, new_n28063);
nor_4  g25716(new_n28065, new_n28064, new_n28021);
nor_4  g25717(new_n28066, new_n28065, new_n28018);
xnor_3 g25718(n11462, new_n28066, new_n28015);
xnor_3 g25719(n11470, new_n24941, new_n24912);
xnor_3 g25720(n11472, new_n18831_1, new_n18815);
xnor_3 g25721(n11496, new_n23224, new_n23223);
xnor_3 g25722(n11506, new_n24664, new_n24617);
nor_4  g25723(new_n28072, new_n26810, new_n6641);
nor_4  g25724(new_n28073, new_n26813, new_n6638);
nor_4  g25725(new_n28074, new_n28073, new_n28072);
not_3  g25726(new_n28075, new_n28074);
nor_4  g25727(new_n28076, new_n19268, new_n6646);
not_3  g25728(new_n28077, new_n28076);
not_3  g25729(new_n28078, new_n19268);
nor_4  g25730(new_n28079, new_n28078, new_n6649);
nor_4  g25731(new_n28080, new_n28079, new_n28076);
nand_4 g25732(new_n28081, new_n12769, new_n6655_1);
xnor_3 g25733(new_n28082, new_n19277, new_n6655_1);
nand_4 g25734(new_n28083, new_n12798, new_n6661);
not_3  g25735(new_n28084, new_n12798);
xnor_3 g25736(new_n28085, new_n28084, new_n6661);
nand_4 g25737(new_n28086, new_n12801_1, new_n6667);
nand_4 g25738(new_n28087, new_n27522, new_n27503);
nand_4 g25739(new_n28088, new_n28087, new_n28086);
nand_4 g25740(new_n28089, new_n28088, new_n28085);
nand_4 g25741(new_n28090, new_n28089, new_n28083);
nand_4 g25742(new_n28091, new_n28090, new_n28082);
nand_4 g25743(new_n28092, new_n28091, new_n28081);
nand_4 g25744(new_n28093, new_n28092, new_n28080);
nand_4 g25745(new_n28094, new_n28093, new_n28077);
xor_3  g25746(n11515, new_n28094, new_n28075);
xnor_3 g25747(n11538, new_n25798, new_n25754);
xnor_3 g25748(n11548, new_n22975, new_n22974);
not_3  g25749(new_n28098, new_n23266);
xor_3  g25750(n11564, new_n28098, new_n23257);
nand_4 g25751(new_n28100, n22442, new_n3662);
nand_4 g25752(new_n28101, new_n26670, new_n26666);
nand_4 g25753(new_n28102, new_n28101, new_n28100);
nor_4  g25754(new_n28103, n3324, n2272);
not_3  g25755(new_n28104, new_n26673);
nor_4  g25756(new_n28105, new_n26677, new_n28104);
nor_4  g25757(new_n28106, new_n28105, new_n28103);
nor_4  g25758(new_n28107, new_n28106, new_n8875);
nand_4 g25759(new_n28108, new_n26688, new_n26682);
nand_4 g25760(new_n28109, new_n28108, new_n26679);
xor_3  g25761(new_n28110, new_n28106, new_n8874);
nor_4  g25762(new_n28111, new_n28110, new_n28109);
nor_4  g25763(new_n28112, new_n28111, new_n28107);
not_3  g25764(new_n28113, new_n28112);
nor_4  g25765(new_n28114, new_n28113, new_n28102);
not_3  g25766(new_n28115, new_n28102);
nor_4  g25767(new_n28116, new_n28112, new_n28115);
nor_4  g25768(new_n28117, new_n28116, new_n28114);
xnor_3 g25769(new_n28118, new_n28110, new_n28109);
nor_4  g25770(new_n28119, new_n28118, new_n28115);
xnor_3 g25771(new_n28120, new_n28118, new_n28115);
not_3  g25772(new_n28121, new_n26689);
nand_4 g25773(new_n28122, new_n28121, new_n26671);
nand_4 g25774(new_n28123, new_n26695, new_n28122);
nor_4  g25775(new_n28124, new_n28123, new_n28120);
nor_4  g25776(new_n28125, new_n28124, new_n28119);
xnor_3 g25777(n11591, new_n28125, new_n28117);
not_3  g25778(new_n28127, new_n9905);
nor_4  g25779(new_n28128, new_n9912, new_n28127);
nand_4 g25780(new_n28129, new_n9997, new_n9927);
nand_4 g25781(new_n28130, new_n28129, new_n27524);
nor_4  g25782(new_n28131, new_n28130, new_n9926_1);
not_3  g25783(new_n28132, new_n28131);
nor_4  g25784(n11607, new_n28132, new_n28128);
xnor_3 g25785(n11647, new_n22908, new_n22875);
xor_3  g25786(n11674, new_n27877, new_n27871);
xnor_3 g25787(new_n28136, new_n24019, new_n18964);
not_3  g25788(new_n28137, new_n26176);
nand_4 g25789(new_n28138, new_n26182, new_n26178);
nand_4 g25790(new_n28139, new_n28138, new_n28137);
xnor_3 g25791(n11682, new_n28139, new_n28136);
nor_4  g25792(new_n28141, new_n27658, new_n27647);
nor_4  g25793(n11710, new_n28141, new_n26947);
xnor_3 g25794(n11712, new_n16810, new_n16768);
xor_3  g25795(n11724, new_n26521, new_n26507);
not_3  g25796(new_n28145, new_n22193);
xor_3  g25797(n11741, new_n28145, new_n22191);
xor_3  g25798(n11770, new_n21872, new_n3237);
not_3  g25799(new_n28148, new_n9983);
nor_4  g25800(new_n28149, new_n9955, new_n9954);
xor_3  g25801(n11771, new_n28149, new_n28148);
xnor_3 g25802(n11818, new_n23101, new_n23068_1);
not_3  g25803(new_n28152, new_n27518);
xor_3  g25804(n11837, new_n28152, new_n27511);
not_3  g25805(new_n28154, new_n19732);
nor_4  g25806(new_n28155, new_n28154, n7026);
xor_3  g25807(new_n28156, new_n28155, new_n3825);
not_3  g25808(new_n28157, new_n28156);
nor_4  g25809(new_n28158, new_n28157, new_n6925);
xnor_3 g25810(new_n28159, new_n28157, new_n6925);
nor_4  g25811(new_n28160, new_n19734, new_n6930);
nor_4  g25812(new_n28161, new_n19788, new_n19735);
nor_4  g25813(new_n28162, new_n28161, new_n28160);
nor_4  g25814(new_n28163, new_n28162, new_n28159);
nor_4  g25815(new_n28164, new_n28163, new_n28158);
not_3  g25816(new_n28165, new_n28164);
not_3  g25817(new_n28166, new_n28155);
nor_4  g25818(new_n28167, new_n28166, n2743);
not_3  g25819(new_n28168, new_n28167);
nor_4  g25820(new_n28169, new_n28168, new_n16277);
nor_4  g25821(new_n28170, new_n28167, new_n16278);
nor_4  g25822(new_n28171, new_n28170, new_n28169);
xnor_3 g25823(new_n28172, new_n28171, new_n28165);
xnor_3 g25824(new_n28173, new_n28172, new_n26592);
not_3  g25825(new_n28174, new_n28159);
not_3  g25826(new_n28175, new_n28162);
nor_4  g25827(new_n28176, new_n28175, new_n28174);
nor_4  g25828(new_n28177, new_n28176, new_n28163);
nor_4  g25829(new_n28178, new_n28177, new_n26090);
xnor_3 g25830(new_n28179, new_n28177, new_n26090);
nor_4  g25831(new_n28180, new_n19800, new_n19790);
not_3  g25832(new_n28181, new_n19852);
nor_4  g25833(new_n28182, new_n28181, new_n19801);
nor_4  g25834(new_n28183, new_n28182, new_n28180);
nor_4  g25835(new_n28184, new_n28183, new_n28179);
nor_4  g25836(new_n28185, new_n28184, new_n28178);
xnor_3 g25837(n11842, new_n28185, new_n28173);
not_3  g25838(new_n28187, new_n19204);
xor_3  g25839(n11843, new_n19227, new_n28187);
not_3  g25840(new_n28189, new_n22625);
xor_3  g25841(n11905, new_n22648, new_n28189);
not_3  g25842(new_n28191, new_n13687);
xor_3  g25843(n11965, new_n28191, new_n13678);
not_3  g25844(new_n28193, new_n22502);
xor_3  g25845(n12000, new_n22505, new_n28193);
xor_3  g25846(n12003, new_n19957, new_n19944);
not_3  g25847(new_n28196, new_n20694);
xor_3  g25848(n12011, new_n20695, new_n28196);
not_3  g25849(new_n28198, new_n21296);
xor_3  g25850(n12072, new_n21315, new_n28198);
xor_3  g25851(n12131, new_n12864_1, new_n12863);
xor_3  g25852(n12146, new_n19917, new_n19882);
not_3  g25853(new_n28202, new_n20230);
xor_3  g25854(n12157, new_n20233, new_n28202);
xnor_3 g25855(n12158, new_n12309, new_n12243);
xnor_3 g25856(n12179, new_n27043, new_n27022);
xor_3  g25857(n12192, new_n7510, new_n7442);
not_3  g25858(new_n28207, new_n27437);
xor_3  g25859(n12223, new_n28207, new_n27425);
xnor_3 g25860(n12225, new_n12307, new_n12248);
not_3  g25861(new_n28210, new_n27507);
xor_3  g25862(n12228, new_n27520, new_n28210);
xor_3  g25863(n12235, new_n16194, new_n8493);
not_3  g25864(new_n28213, new_n10818);
xor_3  g25865(n12302, new_n10853, new_n28213);
not_3  g25866(new_n28215, new_n20381);
xor_3  g25867(n12304, new_n20413, new_n28215);
xor_3  g25868(new_n28217, n19196, new_n14829);
nand_4 g25869(new_n28218, n23586, new_n7579);
xor_3  g25870(new_n28219, n23586, new_n7579);
nor_4  g25871(new_n28220, new_n14431, n8244);
not_3  g25872(new_n28221, new_n28220);
xor_3  g25873(new_n28222, n21226, new_n7583);
nor_4  g25874(new_n28223, n9493, new_n14435);
not_3  g25875(new_n28224, new_n28223);
nor_4  g25876(new_n28225, n20036, new_n7599);
nor_4  g25877(new_n28226, new_n23942_1, new_n23937);
nor_4  g25878(new_n28227, new_n28226, new_n28225);
xor_3  g25879(new_n28228, n9493, new_n14435);
nand_4 g25880(new_n28229, new_n28228, new_n28227);
nand_4 g25881(new_n28230, new_n28229, new_n28224);
nand_4 g25882(new_n28231, new_n28230, new_n28222);
nand_4 g25883(new_n28232, new_n28231, new_n28221);
nand_4 g25884(new_n28233, new_n28232, new_n28219);
nand_4 g25885(new_n28234, new_n28233, new_n28218);
xnor_3 g25886(new_n28235, new_n28234, new_n28217);
xnor_3 g25887(new_n28236, new_n28235, new_n23891);
not_3  g25888(new_n28237, new_n28232);
xor_3  g25889(new_n28238, new_n28237, new_n28219);
nand_4 g25890(new_n28239, new_n28238, new_n22163);
not_3  g25891(new_n28240, new_n28238);
xnor_3 g25892(new_n28241, new_n28240, new_n22163);
xor_3  g25893(new_n28242, new_n28230, new_n28222);
not_3  g25894(new_n28243, new_n28242);
nand_4 g25895(new_n28244, new_n28243, new_n22169);
xnor_3 g25896(new_n28245, new_n28242, new_n22169);
xor_3  g25897(new_n28246, new_n28228, new_n28227);
not_3  g25898(new_n28247, new_n28246);
nand_4 g25899(new_n28248, new_n28247, new_n22175);
xnor_3 g25900(new_n28249, new_n28246, new_n22175);
nand_4 g25901(new_n28250, new_n23943, new_n22183);
nand_4 g25902(new_n28251, new_n23955, new_n23944);
nand_4 g25903(new_n28252, new_n28251, new_n28250);
nand_4 g25904(new_n28253, new_n28252, new_n28249);
nand_4 g25905(new_n28254, new_n28253, new_n28248);
nand_4 g25906(new_n28255, new_n28254, new_n28245);
nand_4 g25907(new_n28256, new_n28255, new_n28244);
nand_4 g25908(new_n28257, new_n28256, new_n28241);
nand_4 g25909(new_n28258, new_n28257, new_n28239);
xnor_3 g25910(n12324, new_n28258, new_n28236);
xnor_3 g25911(n12325, new_n26168, new_n26165);
xor_3  g25912(n12329, new_n12624, new_n12599);
not_3  g25913(new_n28262, new_n10315);
nor_4  g25914(new_n28263, new_n28262, new_n10313);
xor_3  g25915(n12330, new_n28263, new_n10318);
xnor_3 g25916(n12346, new_n6711, new_n6651);
not_3  g25917(new_n28266, new_n9014);
xor_3  g25918(n12349, new_n28266, new_n8983);
not_3  g25919(new_n28268, new_n23640);
xor_3  g25920(n12364, new_n28268, new_n23639);
nor_4  g25921(new_n28270, new_n26917, new_n6623);
xnor_3 g25922(new_n28271, new_n26914, new_n6620);
nor_4  g25923(new_n28272, new_n26917, new_n6630_1);
not_3  g25924(new_n28273, new_n28272);
nor_4  g25925(new_n28274, new_n26914, new_n6627);
nor_4  g25926(new_n28275, new_n28274, new_n28272);
nor_4  g25927(new_n28276, new_n26920, new_n6634_1);
not_3  g25928(new_n28277, new_n28276);
nor_4  g25929(new_n28278, new_n26808_1, new_n11745);
nor_4  g25930(new_n28279, new_n28278, new_n28276);
not_3  g25931(new_n28280, new_n28073);
nand_4 g25932(new_n28281, new_n28094, new_n28074);
nand_4 g25933(new_n28282, new_n28281, new_n28280);
nand_4 g25934(new_n28283, new_n28282, new_n28279);
nand_4 g25935(new_n28284, new_n28283, new_n28277);
nand_4 g25936(new_n28285, new_n28284, new_n28275);
nand_4 g25937(new_n28286, new_n28285, new_n28273);
nor_4  g25938(new_n28287, new_n28286, new_n28271);
nor_4  g25939(n12383, new_n28287, new_n28270);
xor_3  g25940(n12397, new_n10210, new_n10207);
xor_3  g25941(n12408, new_n20875, new_n20864);
nor_4  g25942(new_n28291, new_n24019, new_n18964);
nor_4  g25943(new_n28292, new_n26175, new_n26176);
nor_4  g25944(new_n28293, new_n28292, new_n28136);
nor_4  g25945(n12449, new_n28293, new_n28291);
xnor_3 g25946(n12461, new_n25906, new_n25865);
nand_4 g25947(new_n28296, new_n25690, new_n14468);
nand_4 g25948(new_n28297, new_n28296, new_n20979);
nand_4 g25949(new_n28298, new_n25691, new_n21049);
nand_4 g25950(new_n28299, new_n25701, new_n25692);
nand_4 g25951(new_n28300, new_n28299, new_n28298);
xnor_3 g25952(new_n28301, new_n28296, new_n26528);
nand_4 g25953(new_n28302, new_n28301, new_n28300);
nand_4 g25954(n12462, new_n28302, new_n28297);
not_3  g25955(new_n28304, new_n27056);
xnor_3 g25956(n12467, new_n28304, new_n27049);
nand_4 g25957(new_n28306, new_n19415, new_n19384);
not_3  g25958(new_n28307, new_n28306);
nor_4  g25959(new_n28308, new_n28307, new_n19383);
not_3  g25960(new_n28309, new_n28308);
nor_4  g25961(new_n28310, new_n28309, new_n26625_1);
not_3  g25962(new_n28311, new_n27555);
not_3  g25963(new_n28312, new_n19465);
nand_4 g25964(new_n28313, new_n19524, new_n28312);
nor_4  g25965(new_n28314, new_n28313, new_n28311);
not_3  g25966(new_n28315, new_n28314);
xnor_3 g25967(new_n28316, new_n28308, new_n26622);
xnor_3 g25968(new_n28317, new_n28313, new_n28311);
nand_4 g25969(new_n28318, new_n28317, new_n28316);
not_3  g25970(new_n28319, new_n28318);
xnor_3 g25971(new_n28320, new_n28317, new_n28316);
nor_4  g25972(new_n28321, new_n19527, new_n22449);
not_3  g25973(new_n28322, new_n28321);
nand_4 g25974(new_n28323, new_n19579, new_n19528);
nand_4 g25975(new_n28324, new_n28323, new_n28322);
nor_4  g25976(new_n28325, new_n28324, new_n28320);
nor_4  g25977(new_n28326, new_n28325, new_n28319);
xnor_3 g25978(new_n28327, new_n28326, new_n28315);
xnor_3 g25979(n12469, new_n28327, new_n28310);
not_3  g25980(new_n28329, new_n13194);
xor_3  g25981(n12515, new_n28329, new_n13159);
nor_4  g25982(new_n28331, new_n10324, n5140);
xor_3  g25983(new_n28332, n10250, new_n14816);
not_3  g25984(new_n28333, new_n28332);
nor_4  g25985(new_n28334, new_n10329, n6204);
xor_3  g25986(new_n28335, n7674, new_n14820);
nand_4 g25987(new_n28336, n6397, new_n14825);
xor_3  g25988(new_n28337, n6397, new_n14825);
nand_4 g25989(new_n28338, n19196, new_n14829);
nand_4 g25990(new_n28339, new_n28234, new_n28217);
nand_4 g25991(new_n28340, new_n28339, new_n28338);
nand_4 g25992(new_n28341, new_n28340, new_n28337);
nand_4 g25993(new_n28342, new_n28341, new_n28336);
nand_4 g25994(new_n28343, new_n28342, new_n28335);
not_3  g25995(new_n28344, new_n28343);
nor_4  g25996(new_n28345, new_n28344, new_n28334);
nor_4  g25997(new_n28346, new_n28345, new_n28333);
nor_4  g25998(new_n28347, new_n28346, new_n28331);
nor_4  g25999(new_n28348, new_n28347, new_n26730);
not_3  g26000(new_n28349, new_n28347);
nor_4  g26001(new_n28350, new_n28349, new_n26728);
nor_4  g26002(new_n28351, new_n28350, new_n28348);
not_3  g26003(new_n28352, new_n25354);
nor_4  g26004(new_n28353, new_n28347, new_n28352);
nor_4  g26005(new_n28354, new_n28349, new_n25354);
xor_3  g26006(new_n28355, new_n28345, new_n28333);
nor_4  g26007(new_n28356, new_n28355, new_n25358);
xnor_3 g26008(new_n28357, new_n28355, new_n25358);
nor_4  g26009(new_n28358, new_n28342, new_n28335);
nor_4  g26010(new_n28359, new_n28358, new_n28344);
nor_4  g26011(new_n28360, new_n28359, new_n23882);
xnor_3 g26012(new_n28361, new_n28359, new_n23882);
not_3  g26013(new_n28362, new_n28337);
xnor_3 g26014(new_n28363, new_n28340, new_n28362);
not_3  g26015(new_n28364, new_n28363);
nand_4 g26016(new_n28365, new_n28364, new_n23886);
xnor_3 g26017(new_n28366, new_n28363, new_n23886);
nand_4 g26018(new_n28367, new_n28235, new_n23892);
nand_4 g26019(new_n28368, new_n28258, new_n28236);
nand_4 g26020(new_n28369, new_n28368, new_n28367);
nand_4 g26021(new_n28370, new_n28369, new_n28366);
nand_4 g26022(new_n28371, new_n28370, new_n28365);
not_3  g26023(new_n28372, new_n28371);
nor_4  g26024(new_n28373, new_n28372, new_n28361);
nor_4  g26025(new_n28374, new_n28373, new_n28360);
nor_4  g26026(new_n28375, new_n28374, new_n28357);
nor_4  g26027(new_n28376, new_n28375, new_n28356);
nor_4  g26028(new_n28377, new_n28376, new_n28354);
nor_4  g26029(new_n28378, new_n28377, new_n28353);
xnor_3 g26030(n12516, new_n28378, new_n28351);
not_3  g26031(new_n28380, new_n8770);
xor_3  g26032(n12540, new_n28380, new_n8756);
not_3  g26033(new_n28382, new_n14137);
xor_3  g26034(n12545, new_n28382, new_n14134);
not_3  g26035(new_n28384, new_n24918);
xor_3  g26036(n12552, new_n24939, new_n28384);
not_3  g26037(new_n28386, new_n9731);
xor_3  g26038(n12566, new_n28386, new_n9701);
xnor_3 g26039(n12569, new_n16132, new_n16110_1);
xnor_3 g26040(n12607, new_n7515, new_n7432_1);
xnor_3 g26041(n12620, new_n12091, new_n12021);
not_3  g26042(new_n28391, new_n4008);
xor_3  g26043(n12621, new_n4066, new_n28391);
not_3  g26044(new_n28393, new_n22410);
xor_3  g26045(n12654, new_n22411, new_n28393);
xor_3  g26046(n12665, new_n23945, new_n18304_1);
not_3  g26047(new_n28396, new_n20905);
xor_3  g26048(n12670, new_n20919, new_n28396);
xor_3  g26049(n12707, new_n8998, new_n2574);
not_3  g26050(new_n28399, new_n8434);
xor_3  g26051(n12725, new_n8446, new_n28399);
xnor_3 g26052(n12727, new_n19576, new_n19533);
xor_3  g26053(n12740, new_n11702, new_n11668);
xnor_3 g26054(n12742, new_n25319, new_n25318);
xor_3  g26055(n12746, new_n25564, new_n2962);
xor_3  g26056(n12756, new_n11062, new_n11061);
xor_3  g26057(n12783, new_n8459, new_n8399_1);
not_3  g26058(new_n28407, new_n28376);
nor_4  g26059(new_n28408, new_n28354, new_n28353);
xnor_3 g26060(n12801, new_n28408, new_n28407);
xnor_3 g26061(n12812, new_n21746, new_n21743);
xnor_3 g26062(n12816, new_n19850, new_n19808);
nor_4  g26063(new_n28412, new_n21158, n6659);
nor_4  g26064(new_n28413, new_n22472, new_n22450);
nor_4  g26065(new_n28414, new_n28413, new_n28412);
not_3  g26066(new_n28415, new_n28414);
nor_4  g26067(new_n28416, new_n28415, new_n24238);
nor_4  g26068(new_n28417, new_n28414, new_n24239);
nor_4  g26069(new_n28418, new_n28417, new_n28416);
not_3  g26070(new_n28419, new_n28418);
nand_4 g26071(new_n28420, new_n28419, new_n28316);
xnor_3 g26072(new_n28421, new_n28418, new_n28316);
nand_4 g26073(new_n28422, new_n22513, new_n22478);
nand_4 g26074(new_n28423, new_n28422, new_n22475);
nand_4 g26075(new_n28424, new_n28423, new_n28421);
nand_4 g26076(new_n28425, new_n28424, new_n28420);
not_3  g26077(new_n28426, new_n28425);
nor_4  g26078(new_n28427, new_n28426, new_n28416);
nor_4  g26079(n12843, new_n28427, new_n28310);
xnor_3 g26080(n12864, new_n25628, new_n25625);
nor_4  g26081(new_n28430, new_n27196, new_n5519);
nor_4  g26082(new_n28431, new_n27230, new_n27197);
nor_4  g26083(new_n28432, new_n28431, new_n28430);
nor_4  g26084(new_n28433, n21784, n3740);
nor_4  g26085(new_n28434, new_n27195, new_n27173);
nor_4  g26086(new_n28435, new_n28434, new_n28433);
nor_4  g26087(new_n28436, new_n28435, new_n17239);
not_3  g26088(new_n28437, new_n28435);
nor_4  g26089(new_n28438, new_n28437, new_n5590);
nor_4  g26090(new_n28439, new_n28438, new_n28436);
not_3  g26091(new_n28440, new_n28439);
xnor_3 g26092(new_n28441, new_n28440, new_n28432);
nor_4  g26093(new_n28442, new_n28441, new_n22966);
nor_4  g26094(new_n28443, new_n27231, new_n21395);
nor_4  g26095(new_n28444, new_n27263, new_n28443);
xnor_3 g26096(new_n28445, new_n28441, new_n22966);
nor_4  g26097(new_n28446, new_n28445, new_n28444);
nor_4  g26098(new_n28447, new_n28446, new_n28442);
not_3  g26099(new_n28448, new_n28447);
nor_4  g26100(new_n28449, new_n28436, new_n28432);
nor_4  g26101(new_n28450, new_n28449, new_n28438);
not_3  g26102(new_n28451, new_n28450);
nor_4  g26103(n12865, new_n28451, new_n28448);
xnor_3 g26104(n12870, new_n15606, new_n15580);
not_3  g26105(new_n28454, new_n25547);
xor_3  g26106(n12873, new_n25574, new_n28454);
nor_4  g26107(new_n28456, new_n26585, new_n22734);
not_3  g26108(new_n28457, new_n28456);
nor_4  g26109(new_n28458, new_n26586, new_n22735);
nor_4  g26110(new_n28459, new_n28458, new_n28456);
nand_4 g26111(new_n28460, new_n26588, new_n22842);
nand_4 g26112(new_n28461, new_n27822, new_n27819);
nand_4 g26113(new_n28462, new_n28461, new_n28460);
nand_4 g26114(new_n28463, new_n28462, new_n28459);
nand_4 g26115(n12904, new_n28463, new_n28457);
xor_3  g26116(n12941, new_n12629, new_n12628);
not_3  g26117(new_n28466, new_n13522);
xor_3  g26118(n12942, new_n28466, new_n13512);
xor_3  g26119(new_n28468, new_n6849, new_n4164);
xor_3  g26120(n12978, new_n28468, new_n6857);
xor_3  g26121(n12980, new_n20913, new_n9367);
xor_3  g26122(n12985, new_n7711, new_n5358);
xnor_3 g26123(n12987, new_n17733, new_n17690);
nor_4  g26124(new_n28473, n11220, new_n14210);
nor_4  g26125(new_n28474, new_n20507, new_n20486);
nor_4  g26126(new_n28475, new_n28474, new_n28473);
not_3  g26127(new_n28476, new_n28475);
nor_4  g26128(new_n28477, new_n28476, new_n18152_1);
nor_4  g26129(new_n28478, new_n28475, new_n18044);
nor_4  g26130(new_n28479, new_n28478, new_n28477);
not_3  g26131(new_n28480, new_n20508);
nor_4  g26132(new_n28481, new_n28480, new_n18098);
nor_4  g26133(new_n28482, new_n20530, new_n20509);
nor_4  g26134(new_n28483, new_n28482, new_n28481);
xnor_3 g26135(n12992, new_n28483, new_n28479);
nor_4  g26136(new_n28485, new_n26979_1, n6659);
nor_4  g26137(new_n28486, new_n25813, n23250);
nor_4  g26138(new_n28487, new_n25860, new_n25816_1);
nor_4  g26139(new_n28488, new_n28487, new_n28486);
nor_4  g26140(new_n28489, new_n26980, new_n21610);
nor_4  g26141(new_n28490, new_n28489, new_n28488);
nor_4  g26142(new_n28491, new_n28490, new_n28485);
nor_4  g26143(new_n28492, new_n28491, new_n26977);
not_3  g26144(new_n28493, new_n28492);
xnor_3 g26145(new_n28494, new_n28493, new_n24252);
nor_4  g26146(new_n28495, new_n28489, new_n28485);
xnor_3 g26147(new_n28496, new_n28495, new_n28488);
nor_4  g26148(new_n28497, new_n28496, new_n24275);
not_3  g26149(new_n28498, new_n28497);
not_3  g26150(new_n28499, new_n28496);
nor_4  g26151(new_n28500, new_n28499, new_n24270);
nor_4  g26152(new_n28501, new_n28500, new_n28497);
nand_4 g26153(new_n28502, new_n25861, new_n17444);
nand_4 g26154(new_n28503, new_n25908, new_n25862);
nand_4 g26155(new_n28504, new_n28503, new_n28502);
nand_4 g26156(new_n28505, new_n28504, new_n28501);
nand_4 g26157(new_n28506, new_n28505, new_n28498);
xnor_3 g26158(n13005, new_n28506, new_n28494);
xor_3  g26159(n13043, new_n24380, new_n20351);
xnor_3 g26160(n13048, new_n21840, new_n21839_1);
xnor_3 g26161(n13054, new_n18778, new_n18775);
xor_3  g26162(n13082, new_n22049, new_n22038);
not_3  g26163(new_n28512, new_n8451);
xor_3  g26164(n13096, new_n28512, new_n8422);
xor_3  g26165(n13116, new_n22052, new_n22027_1);
xnor_3 g26166(n13122, new_n24396, new_n24353);
not_3  g26167(new_n28516, new_n7496);
xor_3  g26168(n13141, new_n28516, new_n7494);
xor_3  g26169(n13144, new_n24200, new_n24191);
xnor_3 g26170(n13168, new_n24946, new_n24905);
not_3  g26171(new_n28520, new_n25766);
xor_3  g26172(n13198, new_n25792_1, new_n28520);
not_3  g26173(new_n28522, new_n17706);
xor_3  g26174(n13199, new_n17727, new_n28522);
not_3  g26175(new_n28524, new_n17871);
xor_3  g26176(n13204, new_n28524, new_n17853);
not_3  g26177(new_n28526, new_n12300);
xor_3  g26178(n13209, new_n28526, new_n12264);
not_3  g26179(new_n28528, new_n23924_1);
xor_3  g26180(n13270, new_n23933, new_n28528);
xnor_3 g26181(n13273, new_n15980, new_n15952);
not_3  g26182(new_n28531, new_n27045);
xor_3  g26183(n13285, new_n28531, new_n27016);
xnor_3 g26184(n13338, new_n26290, new_n26270);
not_3  g26185(new_n28534, new_n9353);
xor_3  g26186(n13407, new_n9382_1, new_n28534);
xor_3  g26187(new_n28536, new_n6288, new_n4798);
xor_3  g26188(n13409, new_n28536, new_n19902);
not_3  g26189(new_n28538, new_n6307);
nand_4 g26190(new_n28539, new_n28538, new_n6266);
xor_3  g26191(n13456, new_n28539, new_n6261);
nor_4  g26192(new_n28541, new_n26228, new_n25379);
nand_4 g26193(new_n28542, new_n26138, new_n25382);
nand_4 g26194(new_n28543, new_n27475, new_n28542);
nor_4  g26195(new_n28544, new_n26262, new_n25379);
nor_4  g26196(new_n28545, new_n28544, new_n28543);
nand_4 g26197(new_n28546, new_n28545, new_n28541);
not_3  g26198(new_n28547, new_n28543);
xnor_3 g26199(new_n28548, new_n26118, new_n25379);
xnor_3 g26200(new_n28549, new_n28548, new_n28547);
nor_4  g26201(new_n28550, new_n28549, new_n13735);
not_3  g26202(new_n28551, new_n28550);
xnor_3 g26203(new_n28552, new_n28548, new_n28543);
nor_4  g26204(new_n28553, new_n28552, new_n13734);
nor_4  g26205(new_n28554, new_n28553, new_n28550);
not_3  g26206(new_n28555, new_n27478);
nor_4  g26207(new_n28556, new_n28555, new_n13855);
nor_4  g26208(new_n28557, new_n27483, new_n28556);
nand_4 g26209(new_n28558, new_n28557, new_n28554);
nand_4 g26210(new_n28559, new_n28558, new_n28551);
xor_3  g26211(new_n28560, new_n26297, new_n25380);
nand_4 g26212(new_n28561, new_n28560, new_n28547);
not_3  g26213(new_n28562, new_n28545);
xor_3  g26214(new_n28563, new_n26297, new_n25379);
nand_4 g26215(new_n28564, new_n28563, new_n28562);
nand_4 g26216(new_n28565, new_n28564, new_n28561);
nand_4 g26217(new_n28566, new_n28565, new_n28559);
nand_4 g26218(n13457, new_n28566, new_n28546);
not_3  g26219(new_n28568, new_n14710);
xor_3  g26220(n13477, new_n14722, new_n28568);
xnor_3 g26221(n13484, new_n15126, new_n15125);
xnor_3 g26222(n13486, new_n25188, new_n25149);
xnor_3 g26223(new_n28572, new_n26929_1, new_n26322);
not_3  g26224(new_n28573, new_n28572);
nor_4  g26225(new_n28574, new_n26822, new_n21263);
nor_4  g26226(new_n28575, new_n26858, new_n26823_1);
nor_4  g26227(new_n28576, new_n28575, new_n28574);
xnor_3 g26228(n13487, new_n28576, new_n28573);
not_3  g26229(new_n28578, new_n5976);
xor_3  g26230(n13500, new_n5999, new_n28578);
xor_3  g26231(n13501, new_n5208, new_n5207);
not_3  g26232(new_n28581, new_n7468);
xor_3  g26233(n13506, new_n7502, new_n28581);
not_3  g26234(new_n28583, new_n7171);
xor_3  g26235(n13548, new_n7183, new_n28583);
xnor_3 g26236(n13551, new_n28057, new_n28035);
not_3  g26237(new_n28586, new_n5734);
xor_3  g26238(n13602, new_n28586, new_n5707);
not_3  g26239(new_n28588, new_n21377);
xor_3  g26240(n13626, new_n28588, new_n21363);
not_3  g26241(new_n28590, new_n9727);
xor_3  g26242(n13683, new_n28590, new_n9718);
xor_3  g26243(n13710, new_n24667, new_n24679);
not_3  g26244(new_n28593, new_n24204);
xor_3  g26245(n13722, new_n28593, new_n24183);
xnor_3 g26246(new_n28595, new_n17242, new_n17163_1);
xnor_3 g26247(n13754, new_n28595, new_n17334);
xor_3  g26248(n13764, new_n2973, new_n2935);
xor_3  g26249(new_n28598, new_n17542, new_n17537);
xor_3  g26250(n13798, new_n28598, new_n17547);
not_3  g26251(new_n28600, new_n21381);
xor_3  g26252(n13835, new_n28600, new_n21355);
not_3  g26253(new_n28602, new_n19340);
xor_3  g26254(n13850, new_n19343, new_n28602);
xor_3  g26255(n13922, new_n22039, new_n9218);
xnor_3 g26256(n13923, new_n23899_1, new_n23888_1);
not_3  g26257(new_n28606, new_n14142);
xor_3  g26258(n14004, new_n28606, new_n14141);
xor_3  g26259(n14036, new_n14397, new_n22953);
xnor_3 g26260(n14059, new_n26378, new_n26361);
xor_3  g26261(n14081, new_n21144, new_n21137);
not_3  g26262(new_n28611, new_n23215);
xor_3  g26263(n14095, new_n23219, new_n28611);
xor_3  g26264(n14107, new_n7914, new_n3613);
not_3  g26265(new_n28614, new_n10610);
xor_3  g26266(n14121, new_n10654, new_n28614);
xor_3  g26267(n14126, new_n14669, new_n14668);
xnor_3 g26268(n14136, new_n24208, new_n24174);
nor_4  g26269(new_n28618, new_n28483, new_n28478);
nor_4  g26270(new_n28619, new_n28618, new_n28477);
nor_4  g26271(new_n28620, new_n28476, new_n27284);
not_3  g26272(new_n28621, new_n28620);
nand_4 g26273(new_n28622, new_n28476, new_n27284);
nand_4 g26274(new_n28623, new_n28622, new_n28621);
xnor_3 g26275(n14147, new_n28623, new_n28619);
xnor_3 g26276(n14174, new_n26052, new_n26004);
xnor_3 g26277(n14190, new_n20241, new_n20210);
not_3  g26278(new_n28627, new_n6306);
xor_3  g26279(n14211, new_n28627, new_n6268);
not_3  g26280(new_n28629, new_n20471);
xor_3  g26281(n14222, new_n20476, new_n28629);
xnor_3 g26282(n14267, new_n16422, new_n16360);
not_3  g26283(new_n28632, new_n6701);
xor_3  g26284(n14271, new_n28632, new_n6686);
not_3  g26285(new_n28634, new_n11285);
xor_3  g26286(n14277, new_n28634, new_n11273_1);
not_3  g26287(new_n28636, new_n9976);
xor_3  g26288(n14294, new_n9979, new_n28636);
xnor_3 g26289(n14310, new_n28064, new_n28021);
not_3  g26290(new_n28639, new_n28085);
xor_3  g26291(n14326, new_n28088, new_n28639);
xnor_3 g26292(n14342, new_n15079, new_n15016);
not_3  g26293(new_n28642, new_n22646);
xor_3  g26294(n14353, new_n28642, new_n22630);
nor_4  g26295(new_n28644, new_n26357, new_n14164);
nor_4  g26296(new_n28645, new_n26356, new_n14166);
nor_4  g26297(new_n28646, new_n26380, new_n26358);
nor_4  g26298(new_n28647, new_n28646, new_n28645);
nor_4  g26299(new_n28648, new_n28647, new_n28644);
nor_4  g26300(new_n28649, new_n26356, new_n14171);
nor_4  g26301(new_n28650, new_n28649, new_n28646);
nor_4  g26302(n14364, new_n28650, new_n28648);
xor_3  g26303(n14375, new_n26940, new_n26937);
xnor_3 g26304(n14412, new_n27445, new_n27415);
nor_4  g26305(new_n28654, new_n21676, new_n7293);
not_3  g26306(new_n28655, new_n28654);
nor_4  g26307(new_n28656, new_n21731, new_n21730);
nor_4  g26308(new_n28657, new_n28656, new_n21711);
nor_4  g26309(new_n28658, new_n28657, new_n28655);
not_3  g26310(new_n28659, new_n28658);
nor_4  g26311(new_n28660, new_n28659, new_n14071_1);
not_3  g26312(new_n28661, new_n14071_1);
nor_4  g26313(new_n28662, new_n28658, new_n28661);
nor_4  g26314(new_n28663, new_n28662, new_n28660);
nor_4  g26315(new_n28664, new_n21716, new_n14072);
nor_4  g26316(new_n28665, new_n21755, new_n21717_1);
nor_4  g26317(new_n28666, new_n28665, new_n28664);
xnor_3 g26318(n14414, new_n28666, new_n28663);
xor_3  g26319(n14457, new_n19023, new_n19021);
xnor_3 g26320(n14464, new_n5738, new_n5691);
not_3  g26321(new_n28670, new_n13165);
xor_3  g26322(n14471, new_n13192, new_n28670);
not_3  g26323(new_n28672, new_n24240);
nand_4 g26324(new_n28673, new_n24251, new_n24243);
nand_4 g26325(new_n28674, new_n28673, new_n28672);
xnor_3 g26326(new_n28675, new_n28674, new_n28492);
nor_4  g26327(new_n28676, new_n28493, new_n24252);
nand_4 g26328(new_n28677, new_n28493, new_n24252);
nand_4 g26329(new_n28678, new_n28506, new_n28677);
not_3  g26330(new_n28679, new_n28678);
nor_4  g26331(new_n28680, new_n28679, new_n28676);
xnor_3 g26332(n14475, new_n28680, new_n28675);
not_3  g26333(new_n28682, new_n15064);
xor_3  g26334(n14541, new_n15067, new_n28682);
not_3  g26335(new_n28684, new_n26649);
nand_4 g26336(new_n28685, new_n26660_1, new_n26652);
nand_4 g26337(n14546, new_n28685, new_n28684);
xor_3  g26338(n14547, new_n13432, new_n13431);
not_3  g26339(new_n28688, new_n15482);
xor_3  g26340(n14593, new_n15502, new_n28688);
not_3  g26341(new_n28690, new_n11256);
xor_3  g26342(n14636, new_n11289, new_n28690);
not_3  g26343(new_n28692, new_n28241);
xor_3  g26344(n14701, new_n28256, new_n28692);
not_3  g26345(new_n28694, new_n14779);
xor_3  g26346(n14734, new_n14794, new_n28694);
xnor_3 g26347(n14746, new_n8457, new_n8404);
xor_3  g26348(n14763, new_n11694, new_n11691);
not_3  g26349(new_n28698, new_n27719);
xor_3  g26350(n14772, new_n28698, new_n27711);
xnor_3 g26351(n14801, new_n27656, new_n27655);
xnor_3 g26352(n14819, new_n26434, new_n26408_1);
xnor_3 g26353(n14827, new_n17879, new_n17833);
xnor_3 g26354(n14839, new_n25699, new_n25695);
not_3  g26355(new_n28704, new_n21371);
xor_3  g26356(n14849, new_n21373, new_n28704);
not_3  g26357(new_n28706, new_n25518_1);
not_3  g26358(new_n28707, new_n25522);
nor_4  g26359(new_n28708, new_n28707, new_n17816);
nor_4  g26360(new_n28709, new_n25590, new_n25523_1);
nor_4  g26361(new_n28710, new_n28709, new_n28708);
nor_4  g26362(n14891, new_n28710, new_n28706);
xor_3  g26363(n14931, new_n7662, new_n5397);
not_3  g26364(new_n28713, new_n28664);
xnor_3 g26365(new_n28714, new_n21716, new_n14073);
not_3  g26366(new_n28715, new_n21733);
xnor_3 g26367(new_n28716, new_n21732, new_n14078);
not_3  g26368(new_n28717, new_n21736);
nor_4  g26369(new_n28718, new_n21708, new_n21689);
nor_4  g26370(new_n28719, new_n28718, new_n21729);
nor_4  g26371(new_n28720, new_n28719, new_n14086);
nor_4  g26372(new_n28721, new_n28720, new_n21736);
nand_4 g26373(new_n28722, new_n21750_1, new_n28721);
nand_4 g26374(new_n28723, new_n28722, new_n28717);
nand_4 g26375(new_n28724, new_n28723, new_n28716);
nand_4 g26376(new_n28725, new_n28724, new_n28715);
nand_4 g26377(new_n28726, new_n28725, new_n28714);
nand_4 g26378(new_n28727, new_n28726, new_n28713);
nand_4 g26379(new_n28728, new_n28727, new_n28660);
nand_4 g26380(new_n28729, new_n28666, new_n28662);
nand_4 g26381(n14944, new_n28729, new_n28728);
xor_3  g26382(n14977, new_n22639, new_n10672);
not_3  g26383(new_n28732, new_n15465_1);
nand_4 g26384(new_n28733, new_n15508_1, new_n26901);
nand_4 g26385(new_n28734, new_n28733, new_n28732);
xor_3  g26386(n14989, new_n28734, new_n15462);
not_3  g26387(new_n28736, new_n13054_1);
xor_3  g26388(n15002, new_n28736, new_n13044_1);
xor_3  g26389(n15004, new_n27516, new_n21915_1);
xnor_3 g26390(n15011, new_n10857, new_n10806);
not_3  g26391(new_n28740, new_n27586);
nor_4  g26392(new_n28741, new_n23606, new_n23552);
nor_4  g26393(new_n28742, new_n27586, new_n28741);
nand_4 g26394(new_n28743, new_n23655, new_n28742);
nand_4 g26395(new_n28744, new_n28743, new_n28740);
nor_4  g26396(new_n28745, new_n28744, new_n27577);
nor_4  g26397(new_n28746, new_n27591, new_n27578);
nor_4  g26398(n15019, new_n28746, new_n28745);
nand_4 g26399(new_n28748, new_n18763, new_n18749);
nand_4 g26400(new_n28749, new_n18784, new_n18757);
nand_4 g26401(n15031, new_n28749, new_n28748);
xor_3  g26402(n15033, new_n22040, new_n22039);
xor_3  g26403(n15052, new_n14518, new_n8493);
xnor_3 g26404(n15082, new_n24091, new_n24081);
not_3  g26405(new_n28754, new_n9708);
xor_3  g26406(n15094, new_n9729, new_n28754);
not_3  g26407(new_n28756, new_n14200);
nor_4  g26408(new_n28757, new_n14199, new_n14196);
nor_4  g26409(n15118, new_n28757, new_n28756);
xnor_3 g26410(n15128, new_n28462, new_n28459);
xnor_3 g26411(n15139, new_n23105, new_n23062);
nor_4  g26412(new_n28761, new_n20601, new_n20590_1);
xnor_3 g26413(n15145, new_n28761, new_n20598);
xnor_3 g26414(n15165, new_n18145_1, new_n18101);
xor_3  g26415(n15176, new_n18683, new_n5850_1);
xor_3  g26416(n15180, new_n24933, new_n24932);
xnor_3 g26417(n15205, new_n19919, new_n19880);
xor_3  g26418(n15230, new_n6298, new_n20732);
xor_3  g26419(n15255, new_n20915_1, new_n20914);
not_3  g26420(new_n28769, new_n11656);
xor_3  g26421(n15275, new_n11706, new_n28769);
not_3  g26422(new_n28771, new_n17025);
xor_3  g26423(n15300, new_n17028, new_n28771);
not_3  g26424(new_n28773, new_n28169);
nor_4  g26425(new_n28774, new_n28773, new_n28164);
not_3  g26426(new_n28775, new_n28170);
nor_4  g26427(new_n28776, new_n28775, new_n28165);
nor_4  g26428(new_n28777, new_n28776, new_n28774);
xnor_3 g26429(new_n28778, new_n28777, new_n26644);
nor_4  g26430(new_n28779, new_n28172, new_n26592);
nor_4  g26431(new_n28780, new_n28185, new_n28173);
nor_4  g26432(new_n28781, new_n28780, new_n28779);
xnor_3 g26433(n15307, new_n28781, new_n28778);
xor_3  g26434(n15327, new_n24669, new_n24677);
not_3  g26435(new_n28784, new_n24641);
xor_3  g26436(n15345, new_n24654, new_n28784);
not_3  g26437(new_n28786, new_n15500);
xor_3  g26438(n15353, new_n28786, new_n15489);
not_3  g26439(new_n28788, new_n28271);
xnor_3 g26440(n15366, new_n28286, new_n28788);
xnor_3 g26441(n15382, new_n28450, new_n28447);
not_3  g26442(new_n28791, new_n11047);
xor_3  g26443(n15407, new_n11068, new_n28791);
not_3  g26444(new_n28793, new_n16515);
xor_3  g26445(n15428, new_n18302, new_n28793);
nor_4  g26446(new_n28795, new_n27998, new_n27994);
not_3  g26447(new_n28796, new_n28013);
nor_4  g26448(new_n28797, new_n28796, new_n27999);
nor_4  g26449(new_n28798, new_n28066, new_n28015);
nor_4  g26450(new_n28799, new_n28798, new_n28797);
nor_4  g26451(new_n28800, new_n28799, new_n28795);
nor_4  g26452(new_n28801, new_n28003, new_n13378);
nand_4 g26453(new_n28802, new_n28012, new_n28801);
nor_4  g26454(new_n28803, new_n28802, new_n28795);
nor_4  g26455(new_n28804, new_n28803, new_n28798);
nor_4  g26456(n15435, new_n28804, new_n28800);
nand_4 g26457(new_n28806, new_n27545, new_n27533);
nand_4 g26458(new_n28807, new_n27546, new_n27531);
nand_4 g26459(n15438, new_n28807, new_n28806);
xnor_3 g26460(n15465, new_n28059, new_n28030);
xor_3  g26461(n15467, new_n10208, new_n7841_1);
xnor_3 g26462(n15470, new_n9392, new_n9321);
xnor_3 g26463(n15477, new_n17883, new_n17827);
not_3  g26464(new_n28813, new_n28361);
xor_3  g26465(n15481, new_n28372, new_n28813);
not_3  g26466(new_n28815, new_n18417);
xor_3  g26467(n15496, new_n18420, new_n28815);
not_3  g26468(new_n28817, new_n14635);
xor_3  g26469(n15501, new_n14681, new_n28817);
xnor_3 g26470(n15555, new_n23221, new_n23212);
xnor_3 g26471(n15558, new_n26222, new_n26207);
not_3  g26472(new_n28821, new_n27383);
nand_4 g26473(new_n28822, new_n27388, new_n27385);
nand_4 g26474(n15559, new_n28822, new_n28821);
nand_4 g26475(new_n28824, new_n25037, new_n24971);
not_3  g26476(new_n28825, new_n28824);
nor_4  g26477(new_n28826, new_n25070, new_n28825);
nor_4  g26478(new_n28827, n23895, new_n19418);
nor_4  g26479(new_n28828, new_n24970, new_n24954);
nor_4  g26480(new_n28829, new_n28828, new_n28827);
nor_4  g26481(new_n28830, new_n28829, new_n26633);
nor_4  g26482(new_n28831, new_n28830, new_n28826);
nand_4 g26483(new_n28832, new_n28831, new_n27637);
nand_4 g26484(new_n28833, new_n28829, new_n27638);
nand_4 g26485(new_n28834, new_n28833, new_n28832);
not_3  g26486(new_n28835, new_n28829);
nor_4  g26487(new_n28836, new_n28835, new_n26633);
nor_4  g26488(new_n28837, new_n28836, new_n28831);
nor_4  g26489(n15570, new_n28837, new_n28834);
xnor_3 g26490(n15573, new_n15085, new_n14994);
nor_4  g26491(new_n28840, new_n14084, new_n14083);
xnor_3 g26492(n15588, new_n28840, new_n14152);
xnor_3 g26493(n15590, new_n26430, new_n26420);
xnor_3 g26494(n15598, new_n27132, new_n27120_1);
xnor_3 g26495(n15614, new_n11291, new_n11250);
xnor_3 g26496(n15662, new_n27723, new_n27697);
not_3  g26497(new_n28846, new_n3587);
xor_3  g26498(n15716, new_n3632, new_n28846);
xnor_3 g26499(n15749, new_n17735_1, new_n17683);
not_3  g26500(new_n28849, new_n23124);
xor_3  g26501(n15762, new_n23127, new_n28849);
xor_3  g26502(n15793, new_n9370, new_n9367);
not_3  g26503(new_n28852, new_n27423);
xor_3  g26504(n15812, new_n27439, new_n28852);
not_3  g26505(new_n28854, new_n15081);
xor_3  g26506(n15815, new_n28854, new_n15011_1);
not_3  g26507(new_n28856, new_n9971);
xor_3  g26508(n15816, new_n9974, new_n28856);
not_3  g26509(new_n28858, new_n14505);
xor_3  g26510(n15831, new_n14526, new_n28858);
not_3  g26511(new_n28860, new_n11542);
xor_3  g26512(n15846, new_n28860, new_n11539);
not_3  g26513(new_n28862, new_n10042);
xor_3  g26514(n15859, new_n10045, new_n28862);
nor_4  g26515(new_n28864, new_n9575, new_n4907);
nor_4  g26516(new_n28865, new_n24503, new_n28864);
nor_4  g26517(new_n28866, new_n28865, new_n9572);
xnor_3 g26518(new_n28867, new_n28866, new_n26711);
xnor_3 g26519(new_n28868, new_n28865, new_n9571);
nor_4  g26520(new_n28869, new_n28868, new_n24898);
nor_4  g26521(new_n28870, new_n24507, new_n24486);
nor_4  g26522(new_n28871, new_n24536, new_n24508);
nor_4  g26523(new_n28872, new_n28871, new_n28870);
xnor_3 g26524(new_n28873, new_n28868, new_n24898);
nor_4  g26525(new_n28874, new_n28873, new_n28872);
nor_4  g26526(new_n28875, new_n28874, new_n28869);
xnor_3 g26527(n15869, new_n28875, new_n28867);
xnor_3 g26528(n15885, new_n23277, new_n23247_1);
nor_4  g26529(new_n28878, new_n25998, new_n25915);
not_3  g26530(new_n28879, new_n26046);
nor_4  g26531(new_n28880, new_n28879, new_n26796);
nor_4  g26532(new_n28881, new_n28880, new_n26016);
nor_4  g26533(new_n28882, new_n28881, new_n26013);
nor_4  g26534(new_n28883, new_n28882, new_n26011);
nor_4  g26535(new_n28884, new_n28883, new_n26008);
nor_4  g26536(new_n28885, new_n28884, new_n26006);
nor_4  g26537(new_n28886, new_n28885, new_n26003);
nor_4  g26538(new_n28887, new_n28886, new_n26001);
nand_4 g26539(new_n28888, new_n28887, new_n28878);
nand_4 g26540(new_n28889, new_n28886, new_n25998);
nand_4 g26541(n15889, new_n28889, new_n28888);
xor_3  g26542(n15917, new_n23264, new_n27834);
xor_3  g26543(n15922, new_n16863, new_n16862);
xor_3  g26544(n15947, new_n8436, new_n8435);
not_3  g26545(new_n28894, new_n25598);
nand_4 g26546(new_n28895, new_n25610, new_n28894);
xor_3  g26547(new_n28896, new_n28895, new_n24031);
not_3  g26548(new_n28897, new_n25616);
nand_4 g26549(new_n28898, new_n25630, new_n25617);
nand_4 g26550(new_n28899, new_n28898, new_n28897);
not_3  g26551(new_n28900, new_n28899);
xnor_3 g26552(n15956, new_n28900, new_n28896);
not_3  g26553(new_n28902, new_n16534);
xnor_3 g26554(n15958, new_n16539, new_n28902);
not_3  g26555(new_n28904, new_n20950);
not_3  g26556(new_n28905, new_n20956);
nand_4 g26557(new_n28906, new_n28905, new_n14752);
nand_4 g26558(new_n28907, new_n28906, new_n28904);
nand_4 g26559(new_n28908, new_n20956, new_n14757);
nand_4 g26560(new_n28909, new_n28908, new_n20953);
nor_4  g26561(n15986, new_n28909, new_n28907);
xnor_3 g26562(n16013, new_n28183, new_n28179);
nor_4  g26563(new_n28912, new_n26897, new_n26884);
nor_4  g26564(new_n28913, new_n28912, new_n26882_1);
not_3  g26565(new_n28914, new_n26881);
nor_4  g26566(new_n28915, new_n28895, new_n28914);
not_3  g26567(new_n28916, new_n28895);
nor_4  g26568(new_n28917, new_n28916, new_n26881);
nor_4  g26569(new_n28918, new_n28917, new_n28915);
xnor_3 g26570(n16060, new_n28918, new_n28913);
not_3  g26571(new_n28920, new_n27888);
nor_4  g26572(new_n28921, new_n20153, new_n20945);
not_3  g26573(new_n28922, new_n28921);
nor_4  g26574(new_n28923, new_n20154, n25972);
nor_4  g26575(new_n28924, new_n28923, new_n28921);
nand_4 g26576(new_n28925, new_n20157, n21915);
nand_4 g26577(new_n28926, new_n27741, new_n27730);
nand_4 g26578(new_n28927, new_n28926, new_n28925);
nand_4 g26579(new_n28928, new_n28927, new_n28924);
nand_4 g26580(new_n28929, new_n28928, new_n28922);
xnor_3 g26581(new_n28930, new_n28929, new_n28920);
nand_4 g26582(new_n28931, new_n28930, new_n28013);
xnor_3 g26583(new_n28932, new_n28930, new_n28796);
xnor_3 g26584(new_n28933, new_n28927, new_n28924);
nand_4 g26585(new_n28934, new_n28933, new_n28020);
xnor_3 g26586(new_n28935, new_n28933, new_n28017);
nand_4 g26587(new_n28936, new_n28022, new_n27742);
nand_4 g26588(new_n28937, new_n27796, new_n27776);
nand_4 g26589(new_n28938, new_n28937, new_n28936);
nand_4 g26590(new_n28939, new_n28938, new_n28935);
nand_4 g26591(new_n28940, new_n28939, new_n28934);
nand_4 g26592(new_n28941, new_n28940, new_n28932);
nand_4 g26593(new_n28942, new_n28941, new_n28931);
not_3  g26594(new_n28943, new_n28942);
nand_4 g26595(new_n28944, new_n28929, new_n28920);
nor_4  g26596(new_n28945, new_n28944, new_n28802);
nand_4 g26597(new_n28946, new_n28944, new_n28802);
not_3  g26598(new_n28947, new_n28946);
nor_4  g26599(new_n28948, new_n28947, new_n28945);
xnor_3 g26600(n16062, new_n28948, new_n28943);
xnor_3 g26601(n16068, new_n28284, new_n28275);
xnor_3 g26602(n16080, new_n28557, new_n28554);
nand_4 g26603(new_n28952, new_n27895, new_n7429);
nand_4 g26604(new_n28953, new_n27901, new_n27897);
nand_4 g26605(new_n28954, new_n28953, new_n28952);
nor_4  g26606(new_n28955, new_n27888, new_n14468);
not_3  g26607(new_n28956, new_n27889);
nor_4  g26608(new_n28957, new_n27894, new_n28956);
nor_4  g26609(new_n28958, new_n28957, new_n28955);
not_3  g26610(new_n28959, new_n28958);
xnor_3 g26611(n16098, new_n28959, new_n28954);
not_3  g26612(new_n28961, new_n21642);
xor_3  g26613(n16110, new_n21658, new_n28961);
not_3  g26614(new_n28963, new_n18567);
xor_3  g26615(n16142, new_n18598, new_n28963);
not_3  g26616(new_n28965, new_n20394);
xor_3  g26617(n16185, new_n20407, new_n28965);
xnor_3 g26618(n16196, new_n15123, new_n15104);
xnor_3 g26619(n16206, new_n25651, new_n25650);
xor_3  g26620(n16215, new_n25746, new_n25741);
not_3  g26621(new_n28970, new_n23414_1);
xor_3  g26622(n16218, new_n28970, new_n23401_1);
xor_3  g26623(n16219, new_n4318, new_n4315);
not_3  g26624(new_n28973, new_n8181);
xor_3  g26625(n16230, new_n8184, new_n28973);
xor_3  g26626(n16243, new_n10040, new_n10030);
not_3  g26627(new_n28976, new_n21302_1);
xor_3  g26628(n16275, new_n21313, new_n28976);
xnor_3 g26629(n16279, new_n12303, new_n12302_1);
not_3  g26630(new_n28979, new_n25131);
nand_4 g26631(new_n28980, new_n25198, new_n25134);
nand_4 g26632(n16322, new_n28980, new_n28979);
xnor_3 g26633(n16327, new_n21321, new_n21276_1);
xnor_3 g26634(n16350, new_n26218, new_n26211);
xor_3  g26635(n16367, new_n7842, new_n7841_1);
xnor_3 g26636(n16379, new_n23541_1, new_n23540);
not_3  g26637(new_n28986, new_n24629_1);
xor_3  g26638(n16398, new_n24658, new_n28986);
not_3  g26639(new_n28988, new_n16522);
xor_3  g26640(n16406, new_n16524_1, new_n28988);
xnor_3 g26641(n16407, new_n27134_1, new_n27115);
xnor_3 g26642(n16419, new_n28940, new_n28932);
xnor_3 g26643(n16424, new_n9992, new_n9937);
nor_4  g26644(new_n28993, new_n16994_1, new_n16992);
xnor_3 g26645(n16428, new_n28993, new_n17041);
xnor_3 g26646(n16433, new_n14542, new_n14471_1);
xnor_3 g26647(n16440, new_n14538, new_n14477);
xor_3  g26648(n16445, new_n21660, new_n21638);
xnor_3 g26649(n16460, new_n17330, new_n17257);
xnor_3 g26650(n16481, new_n24531, new_n24519);
nor_4  g26651(new_n29000, new_n18090, new_n27665);
nand_4 g26652(new_n29001, new_n18153, new_n13381);
nand_4 g26653(new_n29002, new_n25265, new_n25246);
nand_4 g26654(new_n29003, new_n29002, new_n29001);
nor_4  g26655(new_n29004, new_n18153, new_n13375);
nor_4  g26656(new_n29005, new_n29004, new_n29000);
not_3  g26657(new_n29006, new_n29005);
nor_4  g26658(new_n29007, new_n29006, new_n29003);
nor_4  g26659(n16493, new_n29007, new_n29000);
not_3  g26660(new_n29009, new_n5413);
xor_3  g26661(n16506, new_n29009, new_n5383);
not_3  g26662(new_n29011, new_n15596);
xor_3  g26663(n16516, new_n15598_1, new_n29011);
xor_3  g26664(n16517, new_n27254, new_n27253);
not_3  g26665(new_n29014, new_n19220_1);
xor_3  g26666(n16527, new_n29014, new_n19219);
xor_3  g26667(n16554, new_n13046, new_n10998);
xor_3  g26668(n16583, new_n7179, new_n6771);
nor_4  g26669(new_n29018, new_n26559, new_n26553_1);
xnor_3 g26670(n16584, new_n29018, new_n26556);
not_3  g26671(new_n29020, new_n23623);
xor_3  g26672(n16589, new_n23648, new_n29020);
not_3  g26673(new_n29022, new_n24058);
xnor_3 g26674(n16596, new_n29022, new_n24057);
xnor_3 g26675(n16617, new_n27451, new_n27406);
xnor_3 g26676(n16630, new_n9018, new_n8971_1);
not_3  g26677(new_n29026, new_n5629);
xor_3  g26678(n16640, new_n27433, new_n29026);
xor_3  g26679(n16656, new_n2574, new_n2572);
xnor_3 g26680(n16674, new_n8196, new_n8140);
xor_3  g26681(n16682, new_n17327, new_n17262);
xnor_3 g26682(n16684, new_n27364, new_n27343);
not_3  g26683(new_n29032, new_n12735);
xor_3  g26684(n16688, new_n29032, new_n12732);
not_3  g26685(new_n29034, new_n7498);
xor_3  g26686(n16733, new_n29034, new_n7487);
xor_3  g26687(n16798, new_n9378, new_n9377);
xnor_3 g26688(n16834, new_n20526, new_n20525);
xnor_3 g26689(n16837, new_n3258, new_n3203);
xor_3  g26690(n16841, new_n26895, new_n26890);
not_3  g26691(new_n29040, new_n5852);
xor_3  g26692(n16885, new_n5855, new_n29040);
xnor_3 g26693(n16905, new_n9743, new_n9656);
nor_4  g26694(new_n29043, new_n26782, new_n26779);
xnor_3 g26695(n16951, new_n29043, new_n22345);
not_3  g26696(new_n29045, new_n19896);
xor_3  g26697(n16954, new_n19906, new_n29045);
xor_3  g26698(n16989, new_n9970, new_n4046);
xnor_3 g26699(n17006, new_n23543, new_n23503);
not_3  g26700(new_n29049, new_n16403);
xor_3  g26701(n17068, new_n16406_1, new_n29049);
xor_3  g26702(n17070, new_n18589, new_n18585);
xnor_3 g26703(n17075, new_n25194, new_n25140);
not_3  g26704(new_n29053, new_n20858);
xor_3  g26705(n17084, new_n20877, new_n29053);
xor_3  g26706(n17104, new_n5404, new_n13682);
xnor_3 g26707(n17106, new_n16134, new_n16099);
xor_3  g26708(n17119, new_n11698, new_n11684);
xnor_3 g26709(n17130, new_n15984, new_n15939);
xnor_3 g26710(n17138, new_n28055, new_n28039);
not_3  g26711(new_n29060, new_n27244);
xor_3  g26712(n17163, new_n27256, new_n29060);
xor_3  g26713(n17168, new_n24767, new_n24766);
not_3  g26714(new_n29063, new_n13887);
xor_3  g26715(n17202, new_n29063, new_n13878);
xnor_3 g26716(n17219, new_n23834, new_n23833);
xnor_3 g26717(n17232, new_n22910_1, new_n22868);
xor_3  g26718(n17236, new_n18728, new_n18725_1);
xor_3  g26719(n17243, new_n12635, new_n12633);
not_3  g26720(new_n29069, new_n13422);
xor_3  g26721(n17263, new_n13438, new_n29069);
not_3  g26722(new_n29071, new_n24034);
nor_4  g26723(new_n29072, new_n24062, new_n29071);
nor_4  g26724(n17285, new_n29072, new_n24033);
xnor_3 g26725(n17320, new_n14146, new_n14102);
xnor_3 g26726(n17337, new_n2977, new_n2923);
not_3  g26727(new_n29076, new_n27031_1);
xor_3  g26728(n17344, new_n27039, new_n29076);
xnor_3 g26729(n17359, new_n27047, new_n27011_1);
xor_3  g26730(n17387, new_n17307, new_n16214);
xor_3  g26731(n17391, new_n15768, new_n5849);
not_3  g26732(new_n29081, new_n23538);
xor_3  g26733(n17392, new_n29081, new_n23510);
xnor_3 g26734(n17421, new_n27366, new_n27339);
xor_3  g26735(n17432, new_n14720, new_n19054);
xnor_3 g26736(n17436, new_n26044, new_n26022);
xor_3  g26737(n17440, new_n8435, new_n5357);
not_3  g26738(new_n29087, new_n10083);
xor_3  g26739(n17450, new_n29087, new_n6771);
nand_4 g26740(new_n29089, new_n23232, new_n8703);
not_3  g26741(new_n29090, new_n8706);
not_3  g26742(new_n29091, new_n8705);
nand_4 g26743(new_n29092, new_n8787, new_n29091);
nand_4 g26744(new_n29093, new_n29092, new_n29090);
nand_4 g26745(new_n29094, new_n29093, new_n29089);
nand_4 g26746(new_n29095, new_n23233, new_n8704);
nand_4 g26747(new_n29096, new_n29095, new_n29092);
nand_4 g26748(new_n29097, new_n29096, new_n29094);
not_3  g26749(n17461, new_n29097);
not_3  g26750(new_n29099, new_n28501);
xnor_3 g26751(n17466, new_n28504, new_n29099);
not_3  g26752(new_n29101, new_n16420);
xor_3  g26753(n17493, new_n29101, new_n16366);
xor_3  g26754(n17500, new_n26607, new_n26604);
xnor_3 g26755(n17524, new_n27717, new_n27714);
xnor_3 g26756(n17529, new_n6709, new_n6657);
xor_3  g26757(new_n29106, new_n18335, new_n6763);
xor_3  g26758(n17557, new_n29106, new_n18339);
not_3  g26759(new_n29108, new_n20376);
xor_3  g26760(n17583, new_n20415, new_n29108);
not_3  g26761(new_n29110, new_n17319);
xor_3  g26762(n17592, new_n29110, new_n17285_1);
not_3  g26763(new_n29112, new_n9981);
xor_3  g26764(n17638, new_n29112, new_n9961);
xnor_3 g26765(n17687, new_n24534, new_n24512_1);
xnor_3 g26766(n17721, new_n16814, new_n16759);
xnor_3 g26767(n17735, new_n26856, new_n26831);
nor_4  g26768(new_n29117, new_n26131, new_n26128);
not_3  g26769(new_n29118, new_n26128);
nor_4  g26770(new_n29119, new_n26133, new_n29118);
nor_4  g26771(new_n29120, new_n29119, new_n29117);
nor_4  g26772(new_n29121, new_n29120, new_n26228);
xnor_3 g26773(new_n29122, new_n29120, new_n26228);
nor_4  g26774(new_n29123, new_n26135, new_n26118);
nor_4  g26775(new_n29124, new_n26146, new_n26136);
nor_4  g26776(new_n29125, new_n29124, new_n29123);
nor_4  g26777(new_n29126, new_n29125, new_n29122);
nor_4  g26778(new_n29127, new_n29126, new_n29121);
nor_4  g26779(n17738, new_n29127, new_n29117);
xor_3  g26780(n17746, new_n18827, new_n18824);
not_3  g26781(new_n29130, new_n28249);
xor_3  g26782(n17749, new_n28252, new_n29130);
xnor_3 g26783(n17820, new_n23096, new_n23075);
not_3  g26784(new_n29133, new_n17293);
xor_3  g26785(n17855, new_n17317, new_n29133);
not_3  g26786(new_n29135, new_n5591);
not_3  g26787(new_n29136, new_n5656);
nor_4  g26788(new_n29137, new_n29136, new_n29135);
not_3  g26789(new_n29138, new_n29137);
nand_4 g26790(new_n29139, new_n29136, new_n5593_1);
nand_4 g26791(new_n29140, new_n29139, new_n29138);
nor_4  g26792(new_n29141, new_n5749, new_n5750);
nor_4  g26793(new_n29142, new_n29141, new_n29140);
nor_4  g26794(n17877, new_n29142, new_n29137);
xnor_3 g26795(n17889, new_n19047, new_n19046);
nor_4  g26796(new_n29145, new_n28125, new_n28114);
nor_4  g26797(new_n29146, new_n28124, new_n28116);
nor_4  g26798(n17912, new_n29146, new_n29145);
xor_3  g26799(n17927, new_n27355, new_n27352);
not_3  g26800(new_n29149, new_n27417);
xor_3  g26801(n17931, new_n27443, new_n29149);
not_3  g26802(new_n29151, new_n9372_1);
xor_3  g26803(n17948, new_n29151, new_n9371_1);
xor_3  g26804(n17956, new_n19338, new_n19334);
xnor_3 g26805(new_n29154, new_n15435_1, new_n15431);
nor_4  g26806(new_n29155, new_n20942, new_n15446);
nor_4  g26807(new_n29156, new_n29155, new_n15444);
nor_4  g26808(new_n29157, new_n29156, new_n29154);
nor_4  g26809(new_n29158, new_n29157, new_n15436);
nor_4  g26810(new_n29159, new_n29158, new_n15249);
nor_4  g26811(new_n29160, new_n15429, new_n15249);
nor_4  g26812(new_n29161, new_n29157, new_n29160);
nor_4  g26813(n17963, new_n29161, new_n29159);
nor_4  g26814(new_n29163, n25494, new_n21610);
nor_4  g26815(new_n29164, new_n21628_1, new_n21612);
nor_4  g26816(new_n29165, new_n29164, new_n29163);
not_3  g26817(new_n29166, new_n29165);
nor_4  g26818(new_n29167, new_n29166, new_n15931);
nor_4  g26819(new_n29168, new_n29165, new_n15934);
xnor_3 g26820(new_n29169, new_n29165, new_n15934);
not_3  g26821(new_n29170, new_n21632);
nand_4 g26822(new_n29171, new_n21663, new_n29170);
nor_4  g26823(new_n29172, new_n29171, new_n29169);
nor_4  g26824(new_n29173, new_n29172, new_n29168);
nor_4  g26825(new_n29174, new_n29173, new_n29167);
not_3  g26826(new_n29175, new_n15931);
nor_4  g26827(new_n29176, new_n29165, new_n29175);
nor_4  g26828(new_n29177, new_n29176, new_n29172);
nor_4  g26829(n17976, new_n29177, new_n29174);
xnor_3 g26830(n17998, new_n8455, new_n8410);
xor_3  g26831(n18025, new_n17863, new_n2962);
xnor_3 g26832(n18043, new_n25583, new_n25582);
xnor_3 g26833(n18045, new_n27276, new_n27274);
not_3  g26834(new_n29183, new_n4324);
xor_3  g26835(n18059, new_n29183, new_n4310);
xnor_3 g26836(n18061, new_n25192, new_n25143);
xnor_3 g26837(n18071, new_n3641, new_n3561_1);
xnor_3 g26838(n18143, new_n12089, new_n12027);
xnor_3 g26839(n18152, new_n26609, new_n26602);
not_3  g26840(new_n29189, new_n8996);
xor_3  g26841(n18193, new_n9010, new_n29189);
nor_4  g26842(new_n29191, new_n14206, new_n14191);
xnor_3 g26843(n18232, new_n29191, new_n14203);
not_3  g26844(new_n29193, new_n20879_1);
xor_3  g26845(n18238, new_n29193, new_n20851);
not_3  g26846(new_n29195, new_n22899);
xor_3  g26847(n18241, new_n29195, new_n22896);
not_3  g26848(new_n29197, new_n26030);
xor_3  g26849(n18254, new_n26040, new_n29197);
xnor_3 g26850(n18288, new_n26854, new_n26836);
xnor_3 g26851(n18301, new_n14810, new_n14762);
not_3  g26852(new_n29201, new_n27258);
xor_3  g26853(n18304, new_n29201, new_n27240);
xnor_3 g26854(n18310, new_n16424_1, new_n16352);
not_3  g26855(new_n29204, new_n7845);
xor_3  g26856(n18311, new_n29204, new_n7844);
xnor_3 g26857(n18323, new_n21837, new_n21819);
not_3  g26858(new_n29207, new_n6260);
not_3  g26859(new_n29208, new_n6261);
nand_4 g26860(new_n29209, new_n28539, new_n29208);
nand_4 g26861(new_n29210, new_n29209, new_n29207);
xor_3  g26862(n18332, new_n29210, new_n6255);
xnor_3 g26863(n18343, new_n27454, new_n27453);
not_3  g26864(new_n29213, new_n23928);
xor_3  g26865(n18350, new_n23931, new_n29213);
not_3  g26866(new_n29215, new_n22414);
xor_3  g26867(n18362, new_n29215, new_n22413);
xnor_3 g26868(n18377, new_n5744, new_n5671);
not_3  g26869(new_n29218, new_n4549);
xor_3  g26870(n18405, new_n4587, new_n29218);
not_3  g26871(new_n29220, new_n20697);
xor_3  g26872(n18414, new_n29220, new_n20686);
not_3  g26873(new_n29222, new_n17943);
xor_3  g26874(n18418, new_n17954_1, new_n29222);
xnor_3 g26875(n18437, new_n9737, new_n9681);
xnor_3 g26876(n18439, new_n24948, new_n24902);
not_3  g26877(new_n29226, new_n13520);
xor_3  g26878(n18445, new_n29226, new_n13517);
xnor_3 g26879(n18467, new_n8194_1, new_n8145);
xnor_3 g26880(n18482, new_n22916, new_n22846);
xnor_3 g26881(n18509, new_n23275, new_n23249);
xor_3  g26882(n18513, new_n17081, new_n20964);
not_3  g26883(new_n29232, new_n18596);
xor_3  g26884(n18515, new_n29232, new_n18595);
not_3  g26885(new_n29234, new_n19686);
xor_3  g26886(n18572, new_n19715, new_n29234);
nand_4 g26887(new_n29236, new_n28945, new_n28943);
nand_4 g26888(new_n29237, new_n28947, new_n28942);
nand_4 g26889(n18574, new_n29237, new_n29236);
xnor_3 g26890(n18576, new_n26216, new_n26213);
xnor_3 g26891(n18582, new_n27879, new_n27867);
not_3  g26892(new_n29241, new_n24656);
xor_3  g26893(n18583, new_n29241, new_n24635);
not_3  g26894(new_n29243, new_n25175);
xor_3  g26895(n18610, new_n25178, new_n29243);
not_3  g26896(new_n29245, new_n18154);
nand_4 g26897(new_n29246, new_n18160, new_n18156);
nand_4 g26898(new_n29247, new_n29246, new_n29245);
xnor_3 g26899(n18635, new_n29247, new_n27286);
not_3  g26900(new_n29249, new_n7928);
xor_3  g26901(n18653, new_n29249, new_n7927);
xnor_3 g26902(n18679, new_n4070, new_n3994);
xnor_3 g26903(n18693, new_n25321, new_n25312);
not_3  g26904(new_n29253, new_n3209);
xor_3  g26905(n18708, new_n3256, new_n29253);
xnor_3 g26906(n18721, new_n28301, new_n28300);
xnor_3 g26907(n18725, new_n23103, new_n23065_1);
xnor_3 g26908(n18751, new_n25794, new_n25762);
xnor_3 g26909(n18780, new_n20409_1, new_n20391);
xnor_3 g26910(n18782, new_n24214, new_n24163);
nand_4 g26911(new_n29260, new_n9028, new_n8939);
nand_4 g26912(new_n29261, new_n9027, new_n8937);
nand_4 g26913(new_n29262, new_n29261, new_n29260);
not_3  g26914(n18802, new_n29262);
xor_3  g26915(n18830, new_n13188, new_n13186);
xor_3  g26916(n18831, new_n15636_1, new_n15631);
not_3  g26917(new_n29266, new_n14524);
xor_3  g26918(n18843, new_n29266, new_n14514);
not_3  g26919(new_n29268, new_n3222);
xor_3  g26920(n18858, new_n3252, new_n29268);
not_3  g26921(new_n29270, new_n12077);
xor_3  g26922(n18859, new_n29270, new_n12059);
xor_3  g26923(n18864, new_n21323, new_n21270);
xnor_3 g26924(n18865, new_n5225, new_n5138);
xnor_3 g26925(n18886, new_n26519, new_n26518);
not_3  g26926(new_n29275, new_n20405);
xor_3  g26927(n18887, new_n29275, new_n20404);
xnor_3 g26928(n18919, new_n10656, new_n10604);
not_3  g26929(new_n29278, new_n15069);
xor_3  g26930(n18940, new_n29278, new_n15055);
not_3  g26931(new_n29280, new_n28444);
not_3  g26932(new_n29281, new_n28445);
nor_4  g26933(new_n29282, new_n29281, new_n29280);
nor_4  g26934(n18945, new_n29282, new_n28446);
xnor_3 g26935(n18970, new_n28092, new_n28080);
nand_4 g26936(new_n29285, new_n20954, new_n20953);
xnor_3 g26937(n18977, new_n29285, new_n28905);
xor_3  g26938(n18982, new_n18731, new_n19950);
xor_3  g26939(n18999, new_n25902, new_n25900);
xnor_3 g26940(n19044, new_n11752, new_n11747);
xor_3  g26941(n19125, new_n18341, new_n18330);
xor_3  g26942(n19141, new_n6714, new_n6643);
not_3  g26943(new_n29292, new_n17251_1);
nor_4  g26944(new_n29293, new_n21462, new_n29292);
nor_4  g26945(new_n29294, new_n21463, new_n17251_1);
nor_4  g26946(new_n29295, new_n29294, new_n29293);
nor_4  g26947(new_n29296, new_n21470, new_n17260);
not_3  g26948(new_n29297, new_n29296);
not_3  g26949(new_n29298, new_n17260);
nor_4  g26950(new_n29299, new_n21483, new_n29298);
nor_4  g26951(new_n29300, new_n29299, new_n29296);
not_3  g26952(new_n29301, new_n21473);
nand_4 g26953(new_n29302, new_n29301, new_n17265);
nand_4 g26954(new_n29303, new_n23133, new_n23115);
nand_4 g26955(new_n29304, new_n29303, new_n29302);
nand_4 g26956(new_n29305, new_n29304, new_n29300);
nand_4 g26957(new_n29306, new_n29305, new_n29297);
xnor_3 g26958(n19164, new_n29306, new_n29295);
not_3  g26959(new_n29308, new_n9988);
xor_3  g26960(n19174, new_n29308, new_n9987);
xnor_3 g26961(n19176, new_n26105, new_n26102);
not_3  g26962(new_n29311, new_n27260);
xor_3  g26963(n19202, new_n29311, new_n27236);
not_3  g26964(new_n29313, new_n25065);
xor_3  g26965(n19220, new_n29313, new_n25053);
xor_3  g26966(n19221, new_n9390, new_n9327);
not_3  g26967(new_n29316, new_n13689);
xor_3  g26968(n19223, new_n13692, new_n29316);
xor_3  g26969(n19224, new_n21309, new_n21308);
xnor_3 g26970(n19233, new_n19257, new_n19248);
xnor_3 g26971(n19244, new_n15612, new_n15568);
xnor_3 g26972(n19314, new_n10658, new_n10599);
not_3  g26973(new_n29322, new_n13056);
xor_3  g26974(n19315, new_n13059, new_n29322);
xnor_3 g26975(n19323, new_n16416, new_n16374);
not_3  g26976(new_n29325, new_n27034);
xor_3  g26977(n19333, new_n27037_1, new_n29325);
nand_4 g26978(new_n29327, new_n21451, new_n12015);
not_3  g26979(new_n29328, new_n21457);
nand_4 g26980(new_n29329, new_n21489_1, new_n21458);
nand_4 g26981(new_n29330, new_n29329, new_n29328);
not_3  g26982(new_n29331, new_n21451);
xnor_3 g26983(new_n29332, new_n29331, new_n12014);
not_3  g26984(new_n29333, new_n29332);
nand_4 g26985(new_n29334, new_n29333, new_n29330);
nand_4 g26986(n19348, new_n29334, new_n29327);
xnor_3 g26987(n19354, new_n20891, new_n20814);
xnor_3 g26988(n19367, new_n13448, new_n13405);
xnor_3 g26989(n19385, new_n23729, new_n23701);
xnor_3 g26990(new_n29339, new_n21045, new_n26528);
xnor_3 g26991(n19389, new_n29339, new_n21089);
xnor_3 g26992(n19401, new_n20243, new_n20206);
nor_4  g26993(new_n29342, new_n28745, new_n27575);
nor_4  g26994(new_n29343, new_n27572, new_n27570);
xnor_3 g26995(n19414, new_n29343, new_n29342);
xor_3  g26996(n19424, new_n23953, new_n28145);
xnor_3 g26997(n19450, new_n26523, new_n26503);
nand_4 g26998(new_n29347, new_n21451, new_n17163_1);
xnor_3 g26999(new_n29348, new_n29331, new_n17163_1);
nor_4  g27000(new_n29349, new_n21456, new_n17246);
not_3  g27001(new_n29350, new_n29349);
not_3  g27002(new_n29351, new_n17246);
nor_4  g27003(new_n29352, new_n21454, new_n29351);
nor_4  g27004(new_n29353, new_n29352, new_n29349);
not_3  g27005(new_n29354, new_n29294);
nand_4 g27006(new_n29355, new_n29306, new_n29295);
nand_4 g27007(new_n29356, new_n29355, new_n29354);
nand_4 g27008(new_n29357, new_n29356, new_n29353);
nand_4 g27009(new_n29358, new_n29357, new_n29350);
nand_4 g27010(new_n29359, new_n29358, new_n29348);
nand_4 g27011(n19458, new_n29359, new_n29347);
not_3  g27012(new_n29361, new_n18821);
xor_3  g27013(n19467, new_n18829, new_n29361);
not_3  g27014(new_n29363, new_n9672);
xor_3  g27015(n19496, new_n9739, new_n29363);
not_3  g27016(new_n29365, new_n18771);
not_3  g27017(new_n29366, new_n18780_1);
nor_4  g27018(new_n29367, new_n29366, new_n29365);
nor_4  g27019(n19523, new_n29367, new_n18781);
xnor_3 g27020(n19570, new_n5216, new_n5163);
not_3  g27021(new_n29370, new_n14675);
xor_3  g27022(n19602, new_n29370, new_n14658);
not_3  g27023(new_n29372, new_n15110);
xor_3  g27024(n19617, new_n15116, new_n29372);
xnor_3 g27025(n19623, new_n16812_1, new_n16764);
not_3  g27026(new_n29375, new_n27642);
xnor_3 g27027(n19641, new_n27643, new_n29375);
xnor_3 g27028(n19648, new_n27368, new_n27335);
not_3  g27029(new_n29378, new_n19691);
xor_3  g27030(n19664, new_n19713, new_n29378);
xor_3  g27031(n19736, new_n24764, new_n24748);
nand_4 g27032(new_n29381, new_n27595, new_n27566);
nor_4  g27033(new_n29382, new_n27566, new_n3650);
nor_4  g27034(new_n29383, new_n29342, new_n27572);
nor_4  g27035(new_n29384, new_n29383, new_n27570);
nand_4 g27036(new_n29385, new_n29384, new_n29382);
nand_4 g27037(n19749, new_n29385, new_n29381);
xnor_3 g27038(n19756, new_n18424, new_n18410);
not_3  g27039(new_n29388, new_n14673);
xor_3  g27040(n19767, new_n29388, new_n14670);
not_3  g27041(new_n29390, new_n3645);
xnor_3 g27042(n19780, new_n29390, new_n3643);
xnor_3 g27043(n19792, new_n28324, new_n28320);
not_3  g27044(new_n29393, new_n25550_1);
xor_3  g27045(n19798, new_n25572, new_n29393);
xor_3  g27046(n19873, new_n20523, new_n20520);
nor_4  g27047(new_n29396, new_n14399, new_n14346);
nor_4  g27048(new_n29397, new_n29396, new_n22947);
nor_4  g27049(new_n29398, new_n29397, new_n22945);
nor_4  g27050(new_n29399, new_n29398, new_n22943);
nor_4  g27051(new_n29400, new_n29399, new_n22928);
nor_4  g27052(new_n29401, new_n22938, new_n22928);
nor_4  g27053(new_n29402, new_n29398, new_n29401);
nor_4  g27054(n19909, new_n29402, new_n29400);
xor_3  g27055(n19916, new_n24762, new_n24753);
not_3  g27056(new_n29405, new_n25544);
xor_3  g27057(n19923, new_n25576, new_n29405);
xnor_3 g27058(n19930, new_n23545, new_n23499);
xnor_3 g27059(n19968, new_n7517, new_n7387);
not_3  g27060(new_n29409, new_n24187);
xor_3  g27061(n19988, new_n24202, new_n29409);
not_3  g27062(new_n29411, new_n25664);
nor_4  g27063(new_n29412, new_n26552, new_n29411);
nor_4  g27064(new_n29413, new_n25664, new_n12233);
nor_4  g27065(new_n29414, new_n25668, new_n25665_1);
nor_4  g27066(new_n29415, new_n29414, new_n29413);
nor_4  g27067(new_n29416, new_n29415, new_n29412);
nor_4  g27068(new_n29417, new_n26558, new_n25664);
nor_4  g27069(new_n29418, new_n29417, new_n29414);
nor_4  g27070(n20004, new_n29418, new_n29416);
not_3  g27071(new_n29420, new_n25771);
xor_3  g27072(n20017, new_n25790, new_n29420);
xnor_3 g27073(n20033, new_n22912, new_n22861);
xnor_3 g27074(n20061, new_n17033, new_n17032);
xnor_3 g27075(n20069, new_n22360, new_n22355);
nand_4 g27076(new_n29425, new_n17816, new_n17808);
nand_4 g27077(new_n29426, new_n17887, new_n17818);
nand_4 g27078(n20086, new_n29426, new_n29425);
xnor_3 g27079(n20096, new_n24055, new_n24052_1);
not_3  g27080(new_n29429, new_n16408);
xor_3  g27081(n20103, new_n29429, new_n16398_1);
xnor_3 g27082(n20126, new_n14148_1, new_n14096);
xnor_3 g27083(n20149, new_n26294, new_n26263);
xnor_3 g27084(n20187, new_n14536, new_n14480);
xnor_3 g27085(n20279, new_n21606, new_n21569);
nand_4 g27086(new_n29435, new_n27860, new_n27854);
nand_4 g27087(new_n29436, new_n27864, new_n29435);
not_3  g27088(new_n29437, new_n27860);
nand_4 g27089(new_n29438, new_n27881, new_n29437);
not_3  g27090(new_n29439, new_n27881);
nand_4 g27091(new_n29440, new_n29439, new_n21807);
nand_4 g27092(new_n29441, new_n29440, new_n29438);
nor_4  g27093(n20287, new_n29441, new_n29436);
xnor_3 g27094(n20301, new_n25368, new_n25363);
not_3  g27095(new_n29444, new_n9745);
nor_4  g27096(new_n29445, new_n29444, new_n9649);
nor_4  g27097(n20330, new_n29445, new_n9525);
xnor_3 g27098(n20333, new_n14532, new_n14486);
not_3  g27099(new_n29448, new_n12562_1);
not_3  g27100(new_n29449, new_n12563);
nor_4  g27101(new_n29450, new_n23286, new_n12567);
nand_4 g27102(new_n29451, new_n29450, new_n29449);
nand_4 g27103(new_n29452, new_n29451, new_n29448);
nand_4 g27104(new_n29453, new_n29452, new_n12557);
nand_4 g27105(new_n29454, new_n12642, new_n12555);
nand_4 g27106(n20355, new_n29454, new_n29453);
xor_3  g27107(n20366, new_n10031, new_n5986);
xnor_3 g27108(n20388, new_n23774, new_n23771);
not_3  g27109(new_n29458, new_n27419);
xor_3  g27110(n20402, new_n27441, new_n29458);
not_3  g27111(new_n29460, new_n19003);
xor_3  g27112(n20403, new_n19034, new_n29460);
xor_3  g27113(n20424, new_n3237, new_n3234);
not_3  g27114(new_n29463, new_n25182);
xor_3  g27115(n20436, new_n29463, new_n25163);
xor_3  g27116(n20441, new_n9725, new_n9724);
xnor_3 g27117(n20445, new_n9026, new_n8945);
xnor_3 g27118(n20450, new_n5746, new_n5664);
xor_3  g27119(n20490, new_n20424_1, new_n7843);
xor_3  g27120(n20495, new_n25063, new_n25059);
nor_4  g27121(new_n29470, new_n19049, new_n19050);
nand_4 g27122(new_n29471, new_n25915, new_n19050);
nand_4 g27123(new_n29472, new_n19049, new_n19051);
nand_4 g27124(new_n29473, new_n29472, new_n29471);
nor_4  g27125(n20515, new_n29473, new_n29470);
nor_4  g27126(new_n29475, new_n28326, new_n28314);
nor_4  g27127(n20533, new_n29475, new_n28310);
not_3  g27128(new_n29477, new_n22195);
xor_3  g27129(n20582, new_n29477, new_n22185);
not_3  g27130(new_n29479, new_n24357);
xor_3  g27131(n20590, new_n24394, new_n29479);
not_3  g27132(new_n29481, new_n3624);
xor_3  g27133(n20602, new_n29481, new_n3620);
not_3  g27134(new_n29483, new_n20402_1);
xor_3  g27135(n20609, new_n29483, new_n20400);
not_3  g27136(new_n29485, new_n7719);
xor_3  g27137(n20623, new_n29485, new_n7710);
xnor_3 g27138(n20629, new_n25588, new_n25528);
not_3  g27139(new_n29488, new_n17021);
xor_3  g27140(n20661, new_n17030, new_n29488);
not_3  g27141(new_n29490, new_n10085);
xor_3  g27142(n20673, new_n10088, new_n29490);
xnor_3 g27143(n20678, new_n25580, new_n25536);
nor_4  g27144(new_n29493, new_n18394, new_n13774);
nor_4  g27145(new_n29494, new_n18431, new_n18395);
nor_4  g27146(new_n29495, new_n29494, new_n29493);
nor_4  g27147(n20680, new_n29495, new_n18391);
xor_3  g27148(n20685, new_n7493, new_n4657);
nor_4  g27149(new_n29498, new_n29176, new_n29167);
xnor_3 g27150(n20691, new_n29498, new_n29173);
not_3  g27151(new_n29500, new_n19697);
xor_3  g27152(n20696, new_n19711, new_n29500);
not_3  g27153(new_n29502, new_n28043);
xor_3  g27154(n20704, new_n28053, new_n29502);
xor_3  g27155(n20705, new_n26848, new_n26847_1);
not_3  g27156(new_n29505, new_n12087);
xor_3  g27157(n20709, new_n29505, new_n12032);
xnor_3 g27158(n20713, new_n18290_1, new_n18261);
not_3  g27159(new_n29508, new_n10310);
nor_4  g27160(new_n29509, new_n10308, new_n10307);
xor_3  g27161(n20722, new_n29509, new_n29508);
not_3  g27162(new_n29511, new_n28674);
nor_4  g27163(new_n29512, new_n29511, new_n24263);
nor_4  g27164(new_n29513, new_n24282, new_n24264);
nor_4  g27165(new_n29514, new_n29513, new_n24266);
nor_4  g27166(new_n29515, new_n29514, new_n29512);
nor_4  g27167(new_n29516, new_n28674, new_n24262);
nor_4  g27168(new_n29517, new_n29516, new_n29513);
nor_4  g27169(n20723, new_n29517, new_n29515);
nand_4 g27170(new_n29519, new_n27864, new_n27862);
xnor_3 g27171(n20748, new_n29519, new_n27881);
xor_3  g27172(n20761, new_n6302, new_n6285);
xnor_3 g27173(n20774, new_n25190, new_n25146);
xnor_3 g27174(n20788, new_n29358, new_n29348);
not_3  g27175(new_n29524, new_n28622);
nor_4  g27176(new_n29525, new_n29524, new_n28619);
nor_4  g27177(new_n29526, new_n28620, new_n28618);
nor_4  g27178(n20795, new_n29526, new_n29525);
nand_4 g27179(new_n29528, new_n27396, new_n25228);
xnor_3 g27180(new_n29529, new_n25232, new_n25226);
xnor_3 g27181(n20803, new_n29529, new_n29528);
not_3  g27182(new_n29531, new_n5750);
nand_4 g27183(new_n29532, new_n5754, new_n5753);
nand_4 g27184(new_n29533, new_n29532, new_n29531);
xnor_3 g27185(n20869, new_n29533, new_n29140);
xnor_3 g27186(n20879, new_n28254, new_n28245);
xnor_3 g27187(n20915, new_n7504, new_n7462);
xor_3  g27188(new_n29537, n19282, new_n14210);
not_3  g27189(new_n29538, new_n29537);
nor_4  g27190(new_n29539, n12657, new_n20487);
nand_4 g27191(new_n29540, new_n26865, new_n26861);
not_3  g27192(new_n29541, new_n29540);
nor_4  g27193(new_n29542, new_n29541, new_n29539);
xor_3  g27194(new_n29543, new_n29542, new_n29538);
not_3  g27195(new_n29544, new_n29543);
nand_4 g27196(new_n29545, new_n29544, new_n26689);
nand_4 g27197(new_n29546, new_n26866, new_n24701);
nand_4 g27198(new_n29547, new_n26870, new_n26867);
nand_4 g27199(new_n29548, new_n29547, new_n29546);
xnor_3 g27200(new_n29549, new_n29543, new_n26689);
nand_4 g27201(new_n29550, new_n29549, new_n29548);
nand_4 g27202(new_n29551, new_n29550, new_n29545);
nor_4  g27203(new_n29552, n19282, new_n14210);
nor_4  g27204(new_n29553, new_n29542, new_n29538);
nor_4  g27205(new_n29554, new_n29553, new_n29552);
not_3  g27206(new_n29555, new_n29554);
nand_4 g27207(new_n29556, new_n29555, new_n28118);
nor_4  g27208(new_n29557, new_n29556, new_n29551);
nor_4  g27209(new_n29558, new_n29557, new_n28112);
not_3  g27210(new_n29559, new_n29551);
not_3  g27211(new_n29560, new_n28118);
nand_4 g27212(new_n29561, new_n29554, new_n29560);
nor_4  g27213(new_n29562, new_n29561, new_n29559);
nor_4  g27214(new_n29563, new_n29562, new_n28113);
nor_4  g27215(n20935, new_n29563, new_n29558);
not_3  g27216(new_n29565, new_n27346);
xor_3  g27217(n20936, new_n27362, new_n29565);
not_3  g27218(new_n29567, new_n20933);
xor_3  g27219(n21008, new_n29567, new_n20932);
not_3  g27220(new_n29569, new_n24212);
xor_3  g27221(n21017, new_n29569, new_n24166);
nor_4  g27222(new_n29571, new_n28777, new_n26644);
nor_4  g27223(new_n29572, new_n28781, new_n28778);
nor_4  g27224(new_n29573, new_n29572, new_n29571);
nor_4  g27225(n21034, new_n29573, new_n28774);
xnor_3 g27226(n21046, new_n27543, new_n27541);
not_3  g27227(new_n29576, new_n10218);
xor_3  g27228(n21062, new_n29576, new_n10193);
not_3  g27229(new_n29578, new_n28310);
not_3  g27230(new_n29579, new_n28416);
xnor_3 g27231(new_n29580, new_n28425, new_n29579);
nand_4 g27232(new_n29581, new_n29580, new_n29578);
xnor_3 g27233(new_n29582, new_n28425, new_n28416);
nand_4 g27234(new_n29583, new_n29582, new_n28310);
nand_4 g27235(n21093, new_n29583, new_n29581);
xor_3  g27236(n21094, new_n11738, new_n9361);
xnor_3 g27237(n21123, new_n18143_1, new_n18106);
xor_3  g27238(n21154, new_n23412, new_n22442_1);
xnor_3 g27239(n21157, new_n19229, new_n19189);
xnor_3 g27240(n21168, new_n26286, new_n26278);
xor_3  g27241(n21173, new_n8758, new_n8757);
not_3  g27242(new_n29591, new_n5178);
xor_3  g27243(n21176, new_n5212, new_n29591);
not_3  g27244(new_n29593, new_n17723);
xor_3  g27245(n21182, new_n29593, new_n17716);
nand_4 g27246(new_n29595, new_n27327, new_n26315);
nand_4 g27247(new_n29596, new_n27370, new_n26323);
nand_4 g27248(new_n29597, new_n29596, new_n29595);
not_3  g27249(new_n29598, new_n26315);
nand_4 g27250(new_n29599, new_n27371, new_n29598);
nand_4 g27251(new_n29600, new_n29599, new_n27332);
nor_4  g27252(n21193, new_n29600, new_n29597);
not_3  g27253(new_n29602, new_n11408);
xor_3  g27254(n21203, new_n11411, new_n29602);
xor_3  g27255(n21225, new_n20399, new_n2595);
xnor_3 g27256(n21238, new_n24671, new_n24607);
xnor_3 g27257(n21254, new_n17035_1, new_n17014);
xnor_3 g27258(n21298, new_n24943, new_n24908);
xor_3  g27259(n21302, new_n24648, new_n11277);
not_3  g27260(new_n29609, new_n24757);
xor_3  g27261(n21349, new_n24760, new_n29609);
xor_3  g27262(n21365, new_n19908, new_n19892);
xnor_3 g27263(n21367, new_n18782_1, new_n18767);
xnor_3 g27264(n21396, new_n14392, new_n14361);
xnor_3 g27265(n21399, new_n9024, new_n8954);
not_3  g27266(new_n29615, new_n3655);
xnor_3 g27267(n21404, new_n29615, new_n3647);
not_3  g27268(new_n29617, new_n10090);
xor_3  g27269(n21446, new_n29617, new_n10078);
xnor_3 g27270(n21472, new_n14201, new_n14193);
xnor_3 g27271(n21525, new_n8781, new_n8727);
not_3  g27272(new_n29621, new_n21383);
xor_3  g27273(n21549, new_n29621, new_n21349_1);
xnor_3 g27274(n21615, new_n24529, new_n24525);
nor_4  g27275(new_n29624, new_n27860, new_n9313);
xnor_3 g27276(new_n29625, new_n27860, new_n9313);
nor_4  g27277(new_n29626, new_n21843, new_n21848);
nor_4  g27278(new_n29627, new_n29626, new_n29625);
nor_4  g27279(n21628, new_n29627, new_n29624);
nor_4  g27280(new_n29629, new_n26926, new_n26319);
xnor_3 g27281(new_n29630, new_n26926, new_n26322);
not_3  g27282(new_n29631, new_n29630);
nor_4  g27283(new_n29632, new_n26929_1, new_n26322);
nor_4  g27284(new_n29633, new_n28576, new_n28572);
nor_4  g27285(new_n29634, new_n29633, new_n29632);
nor_4  g27286(new_n29635, new_n29634, new_n29631);
nor_4  g27287(n21637, new_n29635, new_n29629);
not_3  g27288(new_n29637, new_n26850);
xor_3  g27289(n21645, new_n29637, new_n26842);
xor_3  g27290(n21665, new_n14711, new_n7711);
xnor_3 g27291(n21680, new_n18429, new_n18399);
xnor_3 g27292(n21685, new_n27449, new_n27409);
xor_3  g27293(n21717, new_n23098, new_n23071);
not_3  g27294(new_n29643, new_n20917);
xor_3  g27295(n21719, new_n29643, new_n20911);
not_3  g27296(new_n29645, new_n23087);
xor_3  g27297(n21750, new_n23090, new_n29645);
xnor_3 g27298(n21765, new_n27159, new_n27156);
xnor_3 g27299(n21800, new_n29549, new_n29548);
xor_3  g27300(new_n29649, new_n4837, new_n4833);
xor_3  g27301(n21820, new_n29649, new_n4843);
not_3  g27302(new_n29651, new_n24178);
xor_3  g27303(n21874, new_n24206, new_n29651);
not_3  g27304(new_n29653, new_n16393);
xor_3  g27305(n21943, new_n16410, new_n29653);
xnor_3 g27306(n21960, new_n19912, new_n19887);
xor_3  g27307(n21976, new_n8444, new_n8443);
xnor_3 g27308(n21986, new_n13702, new_n13658);
xnor_3 g27309(n22016, new_n13450, new_n13401);
not_3  g27310(new_n29659, new_n23083);
xor_3  g27311(n22027, new_n23092, new_n29659);
xor_3  g27312(n22050, new_n16130, new_n16118);
xor_3  g27313(n22063, new_n4660, new_n4657);
xnor_3 g27314(n22076, new_n26284, new_n26281);
not_3  g27315(new_n29664, new_n25636);
nor_4  g27316(new_n29665, new_n25659, new_n29664);
nor_4  g27317(n22090, new_n29665, new_n25635);
xnor_3 g27318(n22107, new_n28090, new_n28082);
xor_3  g27319(n22113, new_n22054, new_n22021);
nor_4  g27320(new_n29669, new_n17043, new_n16984);
nor_4  g27321(new_n29670, new_n17042, new_n16987);
nor_4  g27322(n22124, new_n29670, new_n29669);
nor_4  g27323(new_n29672, new_n28895, new_n24030);
nor_4  g27324(new_n29673, new_n28899, new_n28896);
nor_4  g27325(n22126, new_n29673, new_n29672);
nor_4  g27326(new_n29675, new_n29562, new_n29557);
xnor_3 g27327(n22130, new_n29675, new_n28113);
xor_3  g27328(n22144, new_n22300, new_n22296);
xnor_3 g27329(n22150, new_n28565, new_n28559);
not_3  g27330(new_n29679, new_n24447);
xor_3  g27331(n22157, new_n29679, new_n24436);
not_3  g27332(new_n29681, new_n29304);
xor_3  g27333(n22213, new_n29681, new_n29300);
xor_3  g27334(n22283, new_n12618, new_n12615);
xor_3  g27335(n22311, new_n25258, new_n25254_1);
xor_3  g27336(n22317, new_n10660, new_n10590);
xor_3  g27337(n22341, new_n21750_1, new_n21737);
nand_4 g27338(new_n29687, new_n8487, new_n8464);
not_3  g27339(new_n29688, new_n8390);
xnor_3 g27340(new_n29689, new_n22543, new_n8252);
not_3  g27341(new_n29690, new_n8396);
nor_4  g27342(new_n29691, new_n8398, new_n8397);
nor_4  g27343(new_n29692, new_n29691, new_n8396);
nand_4 g27344(new_n29693, new_n8459, new_n29692);
nand_4 g27345(new_n29694, new_n29693, new_n29690);
nand_4 g27346(new_n29695, new_n29694, new_n29689);
nand_4 g27347(new_n29696, new_n29695, new_n29688);
nand_4 g27348(new_n29697, new_n8485, new_n29696);
nand_4 g27349(new_n29698, new_n29697, new_n29687);
xnor_3 g27350(n22353, new_n29698, new_n22657);
xnor_3 g27351(n22444, new_n21748, new_n21740);
xor_3  g27352(n22467, new_n12291, new_n12289);
xor_3  g27353(n22484, new_n10635, new_n10633);
xnor_3 g27354(n22489, new_n22524, new_n22519);
xnor_3 g27355(n22494, new_n9994, new_n9933);
xor_3  g27356(n22533, new_n12626_1, new_n12592);
not_3  g27357(new_n29706, new_n28048);
xor_3  g27358(n22584, new_n28051, new_n29706);
nor_4  g27359(new_n29708, new_n22306, new_n22269);
nor_4  g27360(n22589, new_n29708, new_n22270_1);
xnor_3 g27361(n22620, new_n29356, new_n29353);
xor_3  g27362(n22623, new_n10084, new_n29087);
xnor_3 g27363(n22697, new_n21085, new_n21068);
not_3  g27364(new_n29713, new_n10623);
xor_3  g27365(n22714, new_n10650_1, new_n29713);
xnor_3 g27366(n22761, new_n14540, new_n14474);
not_3  g27367(new_n29716, new_n23626);
xor_3  g27368(n22779, new_n23646, new_n29716);
xnor_3 g27369(n22787, new_n28061, new_n28026);
xnor_3 g27370(n22819, new_n2589, new_n2546);
xor_3  g27371(n22858, new_n11060, new_n5198);
nor_4  g27372(new_n29721, new_n28649, new_n28644);
xnor_3 g27373(n22870, new_n29721, new_n28647);
xor_3  g27374(n22891, new_n11700, new_n11679);
xor_3  g27375(n22897, new_n24387, new_n24370);
xnor_3 g27376(n22903, new_n12312, new_n12238);
xnor_3 g27377(n22907, new_n17737, new_n17676);
not_3  g27378(new_n29727, new_n8448);
xor_3  g27379(n22910, new_n8449, new_n29727);
xnor_3 g27380(n22914, new_n15094_1, new_n15087);
xor_3  g27381(n22939, new_n6725, new_n6687);
not_3  g27382(new_n29731, new_n23776);
xnor_3 g27383(new_n29732, new_n23767, new_n5129);
xnor_3 g27384(n22998, new_n29732, new_n29731);
xor_3  g27385(n23006, new_n10646, new_n20079);
not_3  g27386(new_n29735, new_n15627);
xor_3  g27387(n23007, new_n15638, new_n29735);
xnor_3 g27388(n23009, new_n22548, new_n22545);
xnor_3 g27389(n23014, new_n20889, new_n20821);
xnor_3 g27390(n23047, new_n29634, new_n29630);
xnor_3 g27391(n23058, new_n21835, new_n21822);
nor_4  g27392(n23066, new_n23111, new_n23107);
nor_4  g27393(new_n29742, new_n22983, new_n12369);
nor_4  g27394(new_n29743, new_n29742, new_n22985);
xnor_3 g27395(n23067, new_n29743, new_n22982);
xor_3  g27396(n23238, new_n19904, new_n19898);
xnor_3 g27397(n23247, new_n21487, new_n21467);
xor_3  g27398(n23248, new_n18591, new_n18580);
not_3  g27399(new_n29748, new_n21582);
xor_3  g27400(n23270, new_n21599_1, new_n29748);
xnor_3 g27401(n23289, new_n28123, new_n28120);
xnor_3 g27402(n23305, new_n6312, new_n6244);
not_3  g27403(new_n29752, new_n26034);
xor_3  g27404(n23341, new_n26038, new_n29752);
xor_3  g27405(n23342, new_n11278, new_n5631);
nand_4 g27406(new_n29755, new_n26404, new_n8938);
nand_4 g27407(new_n29756, new_n26436, new_n29755);
not_3  g27408(new_n29757, new_n29756);
nor_4  g27409(new_n29758, new_n26404, new_n8938);
not_3  g27410(new_n29759, new_n26435);
nor_4  g27411(new_n29760, new_n29759, new_n29758);
nor_4  g27412(n23355, new_n29760, new_n29757);
xnor_3 g27413(n23371, new_n23897, new_n23894);
xnor_3 g27414(n23401, new_n19038, new_n18993);
xor_3  g27415(n23414, new_n16127, new_n16125);
not_3  g27416(new_n29765, new_n21575);
xor_3  g27417(n23429, new_n21604, new_n29765);
nor_4  g27418(new_n29767, new_n26715, new_n26708);
not_3  g27419(new_n29768, new_n26711);
nor_4  g27420(new_n29769, new_n29768, new_n26708);
nor_4  g27421(new_n29770, new_n29769, new_n26714);
nor_4  g27422(n23433, new_n29770, new_n29767);
not_3  g27423(new_n29772, new_n22888);
xor_3  g27424(n23434, new_n22904, new_n29772);
nor_4  g27425(new_n29774, new_n28915, new_n28913);
nor_4  g27426(new_n29775, new_n28917, new_n28912);
nor_4  g27427(n23450, new_n29775, new_n29774);
not_3  g27428(new_n29777, new_n20887);
xor_3  g27429(n23471, new_n29777, new_n20828);
xor_3  g27430(n23480, new_n26048, new_n26013);
xnor_3 g27431(n23546, new_n22092, new_n22086);
not_3  g27432(new_n29781, new_n25557);
xor_3  g27433(n23550, new_n25570, new_n29781);
not_3  g27434(new_n29783, new_n8745_1);
xor_3  g27435(n23585, new_n8775, new_n29783);
xor_3  g27436(n23588, new_n24385, new_n24374_1);
xor_3  g27437(n23619, new_n25898, new_n25897);
not_3  g27438(new_n29787, new_n3233);
xor_3  g27439(n23624, new_n3250, new_n29787);
not_3  g27440(new_n29789, new_n14377);
xor_3  g27441(n23628, new_n14384, new_n29789);
xnor_3 g27442(n23637, new_n27041, new_n27027);
xnor_3 g27443(n23663, new_n27792, new_n27789);
not_3  g27444(new_n29793, new_n14386);
xor_3  g27445(n23669, new_n29793, new_n14373);
xnor_3 g27446(n23684, new_n15982, new_n15947_1);
not_3  g27447(new_n29796, new_n23531);
xor_3  g27448(n23690, new_n29796, new_n23521);
not_3  g27449(new_n29798, new_n27447);
xor_3  g27450(n23714, new_n29798, new_n27413);
not_3  g27451(new_n29800, new_n28954);
nor_4  g27452(n23719, new_n28958, new_n29800);
xnor_3 g27453(n23748, new_n26373, new_n26370);
xor_3  g27454(n23856, new_n13177, new_n8490);
not_3  g27455(new_n29804, new_n8773);
xor_3  g27456(n23883, new_n29804, new_n8772);
xor_3  g27457(new_n29806, new_n17717, new_n6793);
xor_3  g27458(n23888, new_n29806, new_n17720);
not_3  g27459(new_n29808, new_n3593);
xor_3  g27460(n23899, new_n3630, new_n29808);
xor_3  g27461(n23903, new_n21306, new_n11401);
xnor_3 g27462(n23924, new_n15610, new_n15573_1);
not_3  g27463(new_n29812, new_n20479);
xor_3  g27464(n23935, new_n29812, new_n20478_1);
not_3  g27465(new_n29814, new_n15978);
xor_3  g27466(n23942, new_n29814, new_n15958_1);
xor_3  g27467(n23954, new_n21883, new_n21870);
not_3  g27468(new_n29817, new_n23168);
xor_3  g27469(n23958, new_n23191, new_n29817);
xor_3  g27470(n23986, new_n27629, new_n27628);
xor_3  g27471(n24002, new_n20935_1, new_n20929_1);
not_3  g27472(new_n29821, new_n15845);
xor_3  g27473(n24039, new_n29821, new_n15832);
xnor_3 g27474(n24052, new_n28873, new_n28872);
not_3  g27475(new_n29824, new_n25156);
xor_3  g27476(n24092, new_n25184, new_n29824);
not_3  g27477(new_n29826, new_n19225);
xor_3  g27478(n24096, new_n29826, new_n19224_1);
xnor_3 g27479(n24097, new_n14802, new_n14771);
xnor_3 g27480(n24105, new_n14390, new_n14365);
not_3  g27481(new_n29830, new_n22484_1);
xor_3  g27482(n24119, new_n22511, new_n29830);
xnor_3 g27483(n24133, new_n18426, new_n18404);
xnor_3 g27484(n24141, new_n24662, new_n24621);
xnor_3 g27485(n24145, new_n26298, new_n26296);
xnor_3 g27486(n24146, new_n27130_1, new_n27126);
not_3  g27487(new_n29836, new_n15456);
xor_3  g27488(n24155, new_n15513, new_n29836);
xnor_3 g27489(n24160, new_n29171, new_n29169);
xnor_3 g27490(n24167, new_n11074, new_n11033);
nand_4 g27491(new_n29840, new_n25327, new_n25323);
not_3  g27492(n24172, new_n29840);
not_3  g27493(new_n29842, new_n17709);
xor_3  g27494(n24177, new_n17725, new_n29842);
xnor_3 g27495(n24228, new_n29005, new_n29003);
xnor_3 g27496(n24258, new_n21753_1, new_n21734);
nor_4  g27497(new_n29846, new_n22654, new_n8467);
not_3  g27498(new_n29847, new_n29687);
nor_4  g27499(new_n29848, new_n29697, new_n22654);
nor_4  g27500(new_n29849, new_n29848, new_n29847);
nor_4  g27501(n24260, new_n29849, new_n29846);
xor_3  g27502(n24289, new_n23650, new_n23619_1);
not_3  g27503(new_n29852, new_n5406);
xor_3  g27504(n24297, new_n29852, new_n5393);
xor_3  g27505(n24307, new_n14382, new_n4311);
not_3  g27506(new_n29855, new_n2582_1);
xor_3  g27507(n24342, new_n29855, new_n2570_1);
xnor_3 g27508(n24345, new_n19910, new_n19890);
not_3  g27509(new_n29858, new_n11413);
xor_3  g27510(n24347, new_n29858, new_n11399);
xnor_3 g27511(n24373, new_n5742_1, new_n5677);
xor_3  g27512(n24406, new_n22429, new_n22428);
not_3  g27513(new_n29862, new_n16875);
xor_3  g27514(n24415, new_n29862, new_n16861);
not_3  g27515(new_n29864, new_n13052);
xor_3  g27516(n24421, new_n29864, new_n13051);
not_3  g27517(new_n29866, new_n16616);
xor_3  g27518(n24431, new_n16653, new_n29866);
xnor_3 g27519(n24472, new_n14530, new_n14490);
nor_4  g27520(new_n29869, new_n28129, new_n27524);
nor_4  g27521(new_n29870, new_n29869, new_n28131);
xnor_3 g27522(n24476, new_n29870, new_n28128);
xnor_3 g27523(n24483, new_n12305, new_n12254);
xor_3  g27524(n24501, new_n16515, new_n16513);
xnor_3 g27525(n24512, new_n22571, new_n22567);
xor_3  g27526(n24558, new_n5411, new_n5408);
xor_3  g27527(n24576, new_n2963, new_n2962);
not_3  g27528(new_n29877, new_n2965);
xor_3  g27529(n24579, new_n29877, new_n2964);
xnor_3 g27530(n24602, new_n25263, new_n25250);
not_3  g27531(new_n29880, new_n17556);
xor_3  g27532(n24604, new_n29880, new_n17510);
xnor_3 g27533(n24626, new_n28282, new_n28279);
nand_4 g27534(new_n29883, new_n27142, new_n27081);
xnor_3 g27535(n24629, new_n29883, new_n27141);
not_3  g27536(new_n29885, new_n26852);
xor_3  g27537(n24636, new_n29885, new_n26838);
xnor_3 g27538(n24715, new_n26516, new_n26513);
xnor_3 g27539(n24723, new_n25196, new_n25137);
nand_4 g27540(new_n29889, new_n20895, new_n20808);
xnor_3 g27541(n24749, new_n29889, new_n20893);
xnor_3 g27542(n24758, new_n25186, new_n25152);
xnor_3 g27543(n24784, new_n28369, new_n28366);
not_3  g27544(new_n29893, new_n20114);
xor_3  g27545(n24807, new_n29893, new_n20113);
xor_3  g27546(n24826, new_n11729, new_n9369);
xnor_3 g27547(n24840, new_n9020, new_n8966);
not_3  g27548(new_n29897, new_n12064);
xor_3  g27549(n24841, new_n12075, new_n29897);
xor_3  g27550(n24853, new_n5997, new_n5982);
not_3  g27551(new_n29900, new_n3254);
xor_3  g27552(n24857, new_n29900, new_n3214);
not_3  g27553(new_n29902, new_n7478);
xor_3  g27554(n24887, new_n7500, new_n29902);
xor_3  g27555(n24934, new_n11064, new_n11055);
xnor_3 g27556(n24998, new_n8785, new_n8712);
not_3  g27557(new_n29906, new_n14139);
xor_3  g27558(n25006, new_n29906, new_n14120);
xnor_3 g27559(n25032, new_n25655, new_n25642);
xnor_3 g27560(n25062, new_n20045, new_n20023);
nand_4 g27561(new_n29910, new_n24220, new_n24152);
xnor_3 g27562(n25083, new_n29910, new_n24218);
xor_3  g27563(n25097, new_n15974, new_n15971);
xnor_3 g27564(n25133, new_n22084, new_n22081);
xnor_3 g27565(n25155, new_n22906, new_n22882);
nand_4 g27566(new_n29915, new_n29561, new_n29556);
xnor_3 g27567(n25181, new_n29915, new_n29551);
xnor_3 g27568(n25200, new_n25657, new_n25640);
nor_4  g27569(new_n29918, new_n26533, new_n26497);
nand_4 g27570(new_n29919, new_n26529, new_n26527);
xnor_3 g27571(n25209, new_n29919, new_n29918);
not_3  g27572(new_n29921, new_n18688);
xor_3  g27573(n25215, new_n29921, new_n18687);
xnor_3 g27574(n25244, new_n22663, new_n22659);
not_3  g27575(new_n29924, new_n22171);
xor_3  g27576(n25254, new_n22199, new_n29924);
xor_3  g27577(n25256, new_n25904, new_n25871);
nand_4 g27578(new_n29927, new_n25072, new_n25071);
nand_4 g27579(new_n29928, new_n29927, new_n28824);
not_3  g27580(new_n29929, new_n28830);
nand_4 g27581(new_n29930, new_n29929, new_n29928);
nor_4  g27582(new_n29931, new_n28835, new_n26636);
not_3  g27583(new_n29932, new_n29931);
nand_4 g27584(new_n29933, new_n29932, new_n29930);
xnor_3 g27585(new_n29934, new_n28835, new_n27637);
xnor_3 g27586(n25293, new_n29934, new_n29933);
xor_3  g27587(n25328, new_n25893, new_n25885);
xor_3  g27588(n25332, new_n13426, new_n4840);
nor_4  g27589(new_n29938, new_n28378, new_n28350);
nor_4  g27590(new_n29939, new_n28377, new_n28348);
nor_4  g27591(n25337, new_n29939, new_n29938);
not_3  g27592(new_n29941, new_n13885);
nor_4  g27593(new_n29942, new_n13882, new_n13881);
xor_3  g27594(n25356, new_n29942, new_n29941);
not_3  g27595(new_n29944, new_n10848);
xor_3  g27596(n25362, new_n29944, new_n10832);
not_3  g27597(new_n29946, new_n17847);
xor_3  g27598(n25412, new_n17873, new_n29946);
xor_3  g27599(n25460, new_n19025, new_n19024);
not_3  g27600(new_n29949, new_n8739);
xor_3  g27601(n25468, new_n8777, new_n29949);
xnor_3 g27602(n25499, new_n17875, new_n17839);
not_3  g27603(new_n29952, new_n24652);
xor_3  g27604(n25513, new_n29952, new_n24649);
xnor_3 g27605(n25518, new_n14800, new_n14773);
xnor_3 g27606(n25532, new_n16418, new_n16370);
xor_3  g27607(n25539, new_n25067, new_n25044);
not_3  g27608(new_n29957, new_n21083);
xor_3  g27609(n25550, new_n29957, new_n21073);
not_3  g27610(new_n29959, new_n26026);
xor_3  g27611(n25611, new_n26042, new_n29959);
xor_3  g27612(new_n29961, new_n6292, new_n6289);
xor_3  g27613(n25614, new_n29961, new_n6300);
xnor_3 g27614(n25619, new_n15608, new_n15578);
nor_4  g27615(new_n29964, new_n28674, new_n28492);
nor_4  g27616(new_n29965, new_n28680, new_n29964);
nor_4  g27617(new_n29966, new_n29511, new_n28493);
nor_4  g27618(new_n29967, new_n28679, new_n29966);
nor_4  g27619(n25665, new_n29967, new_n29965);
not_3  g27620(new_n29969, new_n11041);
xor_3  g27621(n25706, new_n11070, new_n29969);
nor_4  g27622(new_n29971, new_n29516, new_n29512);
xnor_3 g27623(n25719, new_n29971, new_n29514);
xor_3  g27624(n25756, new_n11708, new_n11652);
nor_4  g27625(new_n29974, new_n15931, new_n15882);
not_3  g27626(new_n29975, new_n15986_1);
nor_4  g27627(new_n29976, new_n29975, new_n29974);
nand_4 g27628(new_n29977, new_n15931, new_n15882);
nand_4 g27629(new_n29978, new_n15985, new_n29977);
not_3  g27630(new_n29979, new_n29978);
nor_4  g27631(n25758, new_n29979, new_n29976);
xor_3  g27632(n25773, new_n21306, new_n15619);
xor_3  g27633(n25784, new_n25784_1, new_n22046);
not_3  g27634(new_n29983, new_n9985);
xor_3  g27635(n25792, new_n29983, new_n9949);
xnor_3 g27636(n25816, new_n8192, new_n8151);
xnor_3 g27637(n25826, new_n7506, new_n7456);
xor_3  g27638(n25839, new_n15057, new_n15056);
xnor_3 g27639(n25840, new_n17325, new_n17269);
not_3  g27640(new_n29989, new_n9695_1);
xor_3  g27641(n25873, new_n9733, new_n29989);
not_3  g27642(new_n29991, new_n21848);
nand_4 g27643(new_n29992, new_n21850, new_n21849);
nand_4 g27644(new_n29993, new_n29992, new_n29991);
xnor_3 g27645(n25934, new_n29993, new_n29625);
xnor_3 g27646(n25938, new_n26288, new_n26274_1);
xnor_3 g27647(n25985, new_n26658, new_n26655);
xor_3  g27648(n25994, new_n17072, new_n10834_1);
not_3  g27649(new_n29998, new_n22838);
nand_4 g27650(new_n29999, new_n22918_1, new_n22841);
nand_4 g27651(n26084, new_n29999, new_n29998);
xnor_3 g27652(n26096, new_n28374, new_n28357);
nand_4 g27653(new_n30002, new_n14156, new_n28661);
nor_4  g27654(n26111, new_n30002, new_n14040);
not_3  g27655(new_n30004, new_n14113);
xor_3  g27656(n26113, new_n14144, new_n30004);
xor_3  g27657(n26156, new_n25208, new_n25205);
not_3  g27658(new_n30007, new_n21290);
xor_3  g27659(n26159, new_n21317_1, new_n30007);
not_3  g27660(new_n30009, new_n4068);
xor_3  g27661(n26179, new_n30009, new_n4000_1);
xor_3  g27662(n26220, new_n17309, new_n17307);
xnor_3 g27663(n26229, new_n28423, new_n28421);
not_3  g27664(new_n30013, new_n15471);
xor_3  g27665(n26237, new_n15506_1, new_n30013);
not_3  g27666(new_n30015, new_n19552);
xor_3  g27667(n26250, new_n19570_1, new_n30015);
nor_4  g27668(new_n30017, new_n26790, new_n26787);
nor_4  g27669(n26274, new_n30017, new_n26330);
xnor_3 g27670(n26287, new_n19574, new_n19538);
nor_4  g27671(new_n30020, new_n29417, new_n29412);
xnor_3 g27672(n26317, new_n30020, new_n29415);
nor_4  g27673(new_n30022, new_n23234, new_n23226);
nor_4  g27674(new_n30023, new_n23235, new_n23225);
nor_4  g27675(n26353, new_n30023, new_n30022);
not_3  g27676(new_n30025, new_n25252);
xor_3  g27677(n26375, new_n25261, new_n30025);
nor_4  g27678(new_n30027, new_n28866, new_n26711);
nor_4  g27679(new_n30028, new_n28875, new_n28867);
nor_4  g27680(n26396, new_n30028, new_n30027);
xor_3  g27681(n26429, new_n6298, new_n6295);
not_3  g27682(new_n30031, new_n17938);
xor_3  g27683(n26431, new_n17956_1, new_n30031);
xnor_3 g27684(n26439, new_n8462, new_n8391);
not_3  g27685(new_n30034, new_n25568);
xor_3  g27686(n26492, new_n30034, new_n25565_1);
not_3  g27687(new_n30036, new_n12295);
xor_3  g27688(n26515, new_n12298, new_n30036);
xnor_3 g27689(n26538, new_n2587, new_n2553_1);
not_3  g27690(new_n30039, new_n18576_1);
xor_3  g27691(n26590, new_n18593, new_n30039);
xor_3  g27692(n26598, new_n24197, new_n20872);
nor_4  g27693(new_n30042, new_n29931, new_n28830);
xnor_3 g27694(n26605, new_n30042, new_n28826);
not_3  g27695(new_n30044, new_n28797);
not_3  g27696(new_n30045, new_n28018);
not_3  g27697(new_n30046, new_n28021);
nand_4 g27698(new_n30047, new_n28063, new_n30046);
nand_4 g27699(new_n30048, new_n30047, new_n30045);
nand_4 g27700(new_n30049, new_n30048, new_n28014);
nand_4 g27701(new_n30050, new_n30049, new_n30044);
xnor_3 g27702(new_n30051, new_n28802, new_n28795);
xnor_3 g27703(n26656, new_n30051, new_n30050);
not_3  g27704(new_n30053, new_n14132);
xor_3  g27705(n26674, new_n30053, new_n14129);
not_3  g27706(new_n30055, new_n11525);
xor_3  g27707(n26675, new_n11546, new_n30055);
not_3  g27708(new_n30057, new_n25578);
xor_3  g27709(n26681, new_n30057, new_n25539_1);
nor_4  g27710(new_n30059, new_n11754, new_n6631_1);
nor_4  g27711(new_n30060, new_n30059, new_n6628_1);
nor_4  g27712(new_n30061, new_n30060, new_n6621);
nor_4  g27713(new_n30062, new_n30059, new_n6624);
nor_4  g27714(n26696, new_n30062, new_n30061);
xnor_3 g27715(n26698, new_n18288_1, new_n18267);
xor_3  g27716(n26707, new_n19218, new_n19216);
xnor_3 g27717(n26719, new_n29333, new_n29330);
not_3  g27718(new_n30067, new_n11051);
xor_3  g27719(n26727, new_n11066, new_n30067);
not_3  g27720(new_n30069, new_n26732);
nor_4  g27721(new_n30070, new_n26735, new_n30069);
nor_4  g27722(n26729, new_n30070, new_n26729_1);
not_3  g27723(new_n30072, new_n23165);
not_3  g27724(new_n30073, new_n23167);
not_3  g27725(new_n30074, new_n23189);
nand_4 g27726(new_n30075, new_n30074, new_n26798);
nand_4 g27727(new_n30076, new_n30075, new_n23171);
nand_4 g27728(new_n30077, new_n30076, new_n29817);
nand_4 g27729(new_n30078, new_n30077, new_n30073);
nor_4  g27730(new_n30079, new_n30078, new_n30072);
nor_4  g27731(new_n30080, new_n30079, new_n23162);
xnor_3 g27732(n26745, new_n30080, new_n26759);
not_3  g27733(new_n30082, new_n9347);
xor_3  g27734(n26775, new_n9384, new_n30082);
xnor_3 g27735(n26780, new_n12739, new_n12719);
not_3  g27736(new_n30085, new_n27269);
xnor_3 g27737(n26794, new_n27278, new_n30085);
not_3  g27738(new_n30087, new_n3567);
xor_3  g27739(n26795, new_n3639, new_n30087);
xnor_3 g27740(n26801, new_n13069, new_n13017);
xnor_3 g27741(n26815, new_n13526, new_n13503);
xnor_3 g27742(n26847, new_n28938, new_n28935);
nand_4 g27743(new_n30092, new_n29095, new_n29089);
xnor_3 g27744(n26900, new_n30092, new_n29093);
xor_3  g27745(n26902, new_n23419, new_n23418);
xor_3  g27746(n26905, new_n21656, new_n21648);
xnor_3 g27747(n26921, new_n9735, new_n9689_1);
not_3  g27748(new_n30097, new_n27703);
xor_3  g27749(n26923, new_n27721, new_n30097);
xor_3  g27750(n26929, new_n13182, new_n13179);
xnor_3 g27751(n26930, new_n29156, new_n29154);
xnor_3 g27752(n26943, new_n19572, new_n19543);
xnor_3 g27753(n26970, new_n17877_1, new_n17836);
xnor_3 g27754(n27004, new_n26220_1, new_n26209);
xnor_3 g27755(n27011, new_n12640, new_n12563);
xnor_3 g27756(n27019, new_n24216, new_n24156);
not_3  g27757(new_n30106, new_n5732_1);
xor_3  g27758(n27031, new_n30106, new_n5716);
not_3  g27759(new_n30108, new_n27332);
nor_4  g27760(new_n30109, new_n30108, new_n27330);
xnor_3 g27761(n27051, new_n30109, new_n27370);
xor_3  g27762(n27072, new_n21479, new_n21476);
xnor_3 g27763(n27079, new_n19042_1, new_n18980);
xor_3  g27764(n27096, new_n4842, new_n4840);
xor_3  g27765(n27110, new_n17549, new_n17536);
not_3  g27766(new_n30115, new_n16798_1);
xor_3  g27767(n27112, new_n16802, new_n30115);
xnor_3 g27768(n27130, new_n27727, new_n29883);
xnor_3 g27769(n27145, new_n20040_1, new_n20031);
not_3  g27770(new_n30119, new_n26958);
nor_4  g27771(new_n30120, new_n26961, new_n30119);
nor_4  g27772(n27158, new_n30120, new_n26957);
not_3  g27773(new_n30122, new_n26455);
xor_3  g27774(n27163, new_n26458, new_n30122);
xnor_3 g27775(n27194, new_n29125, new_n29122);
endmodule


