// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Sun Jun 23 19:34:26 2024

module top_810026173_826291639_946996917_1246901 ( 
    n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213, n223,
    n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414, n424,
    n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649, n653,
    n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788, n801,
    n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764,
    n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156, n174,
    n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299, n317,
    n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457, n460,
    n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547, n549,
    n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648, n665,
    n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773, n790,
    n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888, n891,
    n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989, n991,
    n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103, n1113,
    n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183, n1191,
    n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255, n1260,
    n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347, n1348,
    n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426, n1440,
    n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502, n1507,
    n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633, n1635,
    n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690, n1721,
    n1727, n1729, n1731, n1737, n1746  );
  input  n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213,
    n223, n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414,
    n424, n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649,
    n653, n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788,
    n801, n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764;
  output n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156,
    n174, n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299,
    n317, n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457,
    n460, n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547,
    n549, n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648,
    n665, n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773,
    n790, n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888,
    n891, n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989,
    n991, n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103,
    n1113, n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183,
    n1191, n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255,
    n1260, n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347,
    n1348, n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426,
    n1440, n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502,
    n1507, n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633,
    n1635, n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690,
    n1721, n1727, n1729, n1731, n1737, n1746;
  wire new_n276_1, new_n277_1, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290_1, new_n291, new_n292_1, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299_1, new_n300, new_n301,
    new_n302, new_n303_1, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317_1, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329_1,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347_1, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353_1, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372_1, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378_1, new_n379_1, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387_1, new_n388, new_n389, new_n390,
    new_n391_1, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401_1, new_n402_1, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414_1, new_n415, new_n416_1,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423_1,
    new_n424_1, new_n425, new_n426_1, new_n427, new_n428, new_n429_1,
    new_n430, new_n431, new_n432_1, new_n433_1, new_n434, new_n435,
    new_n436, new_n437, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444_1, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452_1, new_n453, new_n454, new_n455, new_n456,
    new_n457_1, new_n458, new_n459, new_n460_1, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469_1,
    new_n470, new_n471, new_n472_1, new_n473, new_n474, new_n475,
    new_n476_1, new_n477, new_n478, new_n480, new_n481, new_n482_1,
    new_n483, new_n484, new_n485, new_n486, new_n487, new_n488_1, new_n489,
    new_n490, new_n491, new_n492, new_n493_1, new_n494, new_n495, new_n496,
    new_n497, new_n498_1, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510_1,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517_1,
    new_n518, new_n519, new_n520, new_n521, new_n522_1, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532_1, new_n533, new_n534_1, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541_1, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547_1, new_n548, new_n549_1, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555_1, new_n556,
    new_n557_1, new_n558, new_n560, new_n564, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585_1, new_n586,
    new_n587, new_n588_1, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599_1, new_n600_1, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607_1, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627_1, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638_1, new_n639, new_n640, new_n641, new_n642,
    new_n643_1, new_n644, new_n645, new_n646_1, new_n647_1, new_n648_1,
    new_n649_1, new_n650, new_n651, new_n652, new_n653_1, new_n654,
    new_n655_1, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665_1, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675_1,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682_1,
    new_n683_1, new_n684_1, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693_1, new_n694,
    new_n695_1, new_n696, new_n697, new_n698, new_n699_1, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712_1, new_n713, new_n714,
    new_n715_1, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724_1, new_n725_1, new_n726, new_n727,
    new_n728, new_n729_1, new_n730, new_n731_1, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738_1, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747_1,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759_1, new_n760, new_n761_1,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770_1, new_n771, new_n772, new_n773_1, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788_1,
    new_n789, new_n790_1, new_n791, new_n792_1, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801_1,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813_1, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823_1,
    new_n824_1, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836_1, new_n837,
    new_n838, new_n839_1, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846_1, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858_1,
    new_n859, new_n860, new_n861, new_n862_1, new_n863, new_n864,
    new_n865_1, new_n866, new_n867_1, new_n868, new_n870_1, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882_1, new_n883_1, new_n884,
    new_n885, new_n886, new_n887, new_n888_1, new_n889, new_n890,
    new_n891_1, new_n892_1, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902_1, new_n903,
    new_n904, new_n906_1, new_n907, new_n909, new_n910, new_n911,
    new_n912_1, new_n913, new_n916, new_n917, new_n918, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927_1, new_n928, new_n929,
    new_n930, new_n931_1, new_n932, new_n933, new_n934, new_n935_1,
    new_n936, new_n937, new_n938, new_n941, new_n942_1, new_n943,
    new_n944_1, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952_1, new_n953_1, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961_1, new_n965, new_n966,
    new_n967, new_n968_1, new_n970, new_n972, new_n973, new_n974_1,
    new_n975, new_n976, new_n977, new_n978, new_n979_1, new_n980_1,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989_1, new_n990, new_n991_1, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000_1, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005_1,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012_1, new_n1013, new_n1014, new_n1015_1, new_n1016_1, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025_1, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030_1, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1059, new_n1060, new_n1061, new_n1062_1,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067_1, new_n1068_1,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103_1, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113_1, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119_1, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1133, new_n1134, new_n1135_1, new_n1136,
    new_n1137, new_n1138_1, new_n1139, new_n1140_1, new_n1141, new_n1142_1,
    new_n1143, new_n1144, new_n1145_1, new_n1146, new_n1147, new_n1148,
    new_n1149_1, new_n1150, new_n1152, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161_1, new_n1162_1, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172_1, new_n1173, new_n1174, new_n1175_1,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183_1, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191_1, new_n1192, new_n1193, new_n1194_1,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199_1, new_n1200,
    new_n1201_1, new_n1202_1, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222_1, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234_1, new_n1235_1, new_n1236,
    new_n1237_1, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249_1, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255_1, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260_1,
    new_n1262, new_n1264, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277_1, new_n1284, new_n1285, new_n1286, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1294, new_n1295, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305_1, new_n1306, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315_1, new_n1316,
    new_n1317, new_n1320, new_n1321_1, new_n1322, new_n1323, new_n1326,
    new_n1327, new_n1328, new_n1331, new_n1332_1, new_n1333, new_n1334,
    new_n1338_1, new_n1341_1, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1346, new_n1347_1, new_n1348_1, new_n1349_1, new_n1350,
    new_n1351_1, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363_1, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369_1, new_n1370, new_n1371, new_n1372, new_n1373, new_n1375,
    new_n1376, new_n1377, new_n1378, new_n1379, new_n1380, new_n1381_1,
    new_n1382, new_n1383_1, new_n1384, new_n1385_1, new_n1386, new_n1387,
    new_n1388, new_n1389, new_n1390, new_n1391, new_n1392, new_n1393_1,
    new_n1394, new_n1395, new_n1396, new_n1397, new_n1398, new_n1399_1,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407_1, new_n1408, new_n1409, new_n1411, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422_1, new_n1423, new_n1424,
    new_n1425_1, new_n1426_1, new_n1427, new_n1428, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435_1, new_n1436, new_n1437,
    new_n1439, new_n1440_1, new_n1441, new_n1442, new_n1443, new_n1444,
    new_n1445, new_n1446, new_n1447, new_n1448, new_n1449, new_n1450,
    new_n1451, new_n1452, new_n1453_1, new_n1454, new_n1455, new_n1456,
    new_n1457_1, new_n1458, new_n1459, new_n1460_1, new_n1461_1, new_n1462,
    new_n1463_1, new_n1464, new_n1465, new_n1466, new_n1467, new_n1468,
    new_n1469, new_n1470_1, new_n1471, new_n1472, new_n1473, new_n1474,
    new_n1475, new_n1476, new_n1477, new_n1478, new_n1479, new_n1480,
    new_n1481_1, new_n1482, new_n1483, new_n1484, new_n1485, new_n1486,
    new_n1487, new_n1488, new_n1489, new_n1490, new_n1491, new_n1492,
    new_n1493, new_n1494, new_n1495_1, new_n1496, new_n1497, new_n1498_1,
    new_n1499, new_n1500, new_n1501_1, new_n1502_1, new_n1503, new_n1504,
    new_n1505, new_n1506, new_n1507_1, new_n1508, new_n1509, new_n1510,
    new_n1511, new_n1512, new_n1513, new_n1514, new_n1515, new_n1516,
    new_n1517, new_n1518, new_n1519, new_n1520, new_n1521, new_n1522,
    new_n1523, new_n1524, new_n1525_1, new_n1526, new_n1527_1, new_n1528,
    new_n1529, new_n1530_1, new_n1531, new_n1532, new_n1533, new_n1534,
    new_n1535_1, new_n1536, new_n1537_1, new_n1538, new_n1539, new_n1540,
    new_n1541, new_n1542, new_n1543, new_n1544_1, new_n1545, new_n1546,
    new_n1547, new_n1548, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1554, new_n1555, new_n1556_1, new_n1557, new_n1558,
    new_n1559, new_n1560, new_n1561, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1566, new_n1567, new_n1568, new_n1569, new_n1570,
    new_n1571, new_n1572, new_n1575, new_n1576, new_n1577, new_n1578,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1589, new_n1591,
    new_n1593, new_n1594, new_n1595_1, new_n1596, new_n1597_1, new_n1598,
    new_n1599, new_n1600_1, new_n1601_1, new_n1606, new_n1607, new_n1608,
    new_n1609, new_n1610, new_n1611, new_n1612, new_n1613_1, new_n1614,
    new_n1615, new_n1616, new_n1617, new_n1618, new_n1619, new_n1620,
    new_n1621, new_n1622_1, new_n1623, new_n1624, new_n1625, new_n1626,
    new_n1627, new_n1628, new_n1629_1, new_n1630, new_n1631, new_n1632,
    new_n1633_1, new_n1634, new_n1635_1, new_n1636, new_n1637, new_n1638,
    new_n1639, new_n1641, new_n1643_1, new_n1644, new_n1645, new_n1650,
    new_n1652, new_n1653, new_n1654_1, new_n1655, new_n1656, new_n1657_1,
    new_n1658, new_n1659, new_n1660_1, new_n1661, new_n1662, new_n1664,
    new_n1666, new_n1667, new_n1668, new_n1669, new_n1673, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683_1, new_n1684, new_n1685,
    new_n1688_1, new_n1689, new_n1690_1, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1706,
    new_n1707_1, new_n1708, new_n1709, new_n1710, new_n1711, new_n1712,
    new_n1715, new_n1721_1, new_n1723, new_n1725, new_n1726, new_n1727_1,
    new_n1728, new_n1729_1, new_n1730, new_n1731_1, new_n1732, new_n1733,
    new_n1734, new_n1741, new_n1742, new_n1743_1, new_n1744, new_n1745,
    new_n1749, new_n1753, new_n1754, new_n1755, new_n1756, new_n1758,
    new_n1759, new_n1760, new_n1762, new_n1765, new_n1766, new_n1767,
    new_n1769, new_n1770, new_n1771, new_n1772, new_n1773, new_n1774,
    new_n1775, new_n1776, new_n1777, new_n1782, new_n1783, new_n1784,
    new_n1785, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1797, new_n1798, new_n1799, new_n1800, new_n1801,
    new_n1803, new_n1804, new_n1805, new_n1806, new_n1807, new_n1808,
    new_n1810, new_n1811, new_n1815, new_n1819, new_n1822, new_n1825,
    new_n1828, new_n1830, new_n1834, new_n1842, new_n1846, new_n1849,
    new_n1850, new_n1851, new_n1854, new_n1855, new_n1856, new_n1857,
    new_n1858, new_n1859, new_n1860, new_n1861, new_n1862, new_n1873,
    new_n1874, new_n1875, new_n1876;
not_8  g0000(n1501, new_n276_1);
not_8  g0001(n36, new_n277_1);
not_8  g0002(n1643, new_n278);
nand_5 g0003(new_n278, new_n277_1, new_n279);
xnor_4 g0004(n1643, new_n277_1, new_n280);
not_8  g0005(n555, new_n281);
not_8  g0006(n788, new_n282);
nand_5 g0007(new_n282, new_n281, new_n283);
xnor_4 g0008(n788, new_n281, new_n284);
not_8  g0009(n353, new_n285);
not_8  g0010(n747, new_n286);
nand_5 g0011(new_n286, new_n285, new_n287);
xnor_4 g0012(n747, new_n285, new_n288);
not_8  g0013(n329, new_n289);
not_8  g0014(n952, new_n290_1);
nand_5 g0015(new_n290_1, new_n289, new_n291);
nand_5 g0016(n1145, n931, new_n292_1);
xnor_4 g0017(n952, new_n289, new_n293);
nand_5 g0018(new_n293, new_n292_1, new_n294);
nand_5 g0019(new_n294, new_n291, new_n295);
nand_5 g0020(new_n295, new_n288, new_n296);
nand_5 g0021(new_n296, new_n287, new_n297);
nand_5 g0022(new_n297, new_n284, new_n298);
nand_5 g0023(new_n298, new_n283, new_n299_1);
nand_5 g0024(new_n299_1, new_n280, new_n300);
nand_5 g0025(new_n300, new_n279, new_n301);
nor_7  g0026(new_n301, new_n276_1, new_n302);
xnor_4 g0027(new_n302, n433, new_n303_1);
nand_5 g0028(n1000, n870, new_n304);
not_8  g0029(n1000, new_n305);
nand_5 g0030(new_n305, n66, new_n306);
nand_5 g0031(new_n306, new_n304, new_n307);
not_8  g0032(new_n307, new_n308);
nand_5 g0033(n1000, n585, new_n309);
nand_5 g0034(new_n305, n968, new_n310);
nand_5 g0035(new_n310, new_n309, new_n311);
not_8  g0036(new_n311, new_n312);
nand_5 g0037(new_n312, new_n308, new_n313);
not_8  g0038(new_n313, new_n314);
nand_5 g0039(n1000, n155, new_n315);
nand_5 g0040(n1435, new_n305, new_n316);
nand_5 g0041(new_n316, new_n315, new_n317_1);
not_8  g0042(new_n317_1, new_n318);
nand_5 g0043(new_n318, new_n314, new_n319);
not_8  g0044(new_n319, new_n320);
not_8  g0045(n682, new_n321);
nand_5 g0046(new_n305, new_n321, new_n322);
not_8  g0047(n1678, new_n323);
nand_5 g0048(new_n323, n1000, new_n324);
nand_5 g0049(new_n324, new_n322, new_n325);
not_8  g0050(new_n325, new_n326);
nand_5 g0051(new_n326, new_n320, new_n327);
xnor_4 g0052(n1597, n682, new_n328);
nand_5 g0053(new_n328, new_n305, new_n329_1);
not_8  g0054(n607, new_n330);
xnor_4 g0055(n1678, new_n330, new_n331);
nand_5 g0056(new_n331, n1000, new_n332);
nand_5 g0057(new_n332, new_n329_1, new_n333);
not_8  g0058(new_n333, new_n334);
xnor_4 g0059(new_n334, new_n327, new_n335);
not_8  g0060(new_n335, new_n336);
xnor_4 g0061(new_n326, new_n319, new_n337);
not_8  g0062(new_n337, new_n338);
xnor_4 g0063(new_n318, new_n313, new_n339);
not_8  g0064(new_n339, new_n340);
not_8  g0065(n693, new_n341);
xnor_4 g0066(new_n311, new_n307, new_n342);
not_8  g0067(new_n342, new_n343);
nand_5 g0068(new_n343, new_n341, new_n344);
nand_5 g0069(new_n342, n693, new_n345);
nand_5 g0070(new_n312, n1763, new_n346);
not_8  g0071(n1763, new_n347_1);
nand_5 g0072(new_n311, new_n347_1, new_n348);
nand_5 g0073(n1461, n1000, new_n349);
nand_5 g0074(new_n305, n347, new_n350);
nand_5 g0075(new_n350, new_n349, new_n351);
nand_5 g0076(new_n351, n1530, new_n352);
not_8  g0077(new_n352, new_n353_1);
nand_5 g0078(new_n353_1, new_n348, new_n354);
nand_5 g0079(new_n354, new_n346, new_n355);
not_8  g0080(new_n355, new_n356);
nand_5 g0081(new_n356, new_n345, new_n357);
nand_5 g0082(new_n357, new_n344, new_n358);
not_8  g0083(new_n358, new_n359);
nand_5 g0084(new_n359, new_n340, new_n360);
not_8  g0085(new_n360, new_n361);
nand_5 g0086(new_n361, new_n338, new_n362);
not_8  g0087(new_n362, new_n363);
nand_5 g0088(new_n363, new_n336, new_n364);
not_8  g0089(new_n327, new_n365);
nand_5 g0090(new_n334, new_n365, new_n366);
not_8  g0091(n26, new_n367);
nand_5 g0092(n1678, n607, new_n368);
nand_5 g0093(new_n368, new_n367, new_n369);
nand_5 g0094(n607, n26, new_n370);
not_8  g0095(new_n370, new_n371);
nand_5 g0096(new_n371, n1678, new_n372_1);
nand_5 g0097(new_n372_1, new_n369, new_n373);
nand_5 g0098(new_n373, n1000, new_n374);
not_8  g0099(n46, new_n375);
not_8  g0100(n1597, new_n376);
nand_5 g0101(new_n376, new_n375, new_n377);
not_8  g0102(new_n377, new_n378_1);
nand_5 g0103(new_n378_1, new_n321, new_n379_1);
nand_5 g0104(new_n376, new_n321, new_n380);
nand_5 g0105(new_n380, n46, new_n381);
nand_5 g0106(new_n381, new_n379_1, new_n382);
not_8  g0107(new_n382, new_n383);
nand_5 g0108(new_n383, new_n305, new_n384);
nand_5 g0109(new_n384, new_n374, new_n385);
xnor_4 g0110(new_n385, new_n366, new_n386);
not_8  g0111(new_n386, new_n387_1);
xnor_4 g0112(new_n387_1, new_n364, new_n388);
xnor_4 g0113(new_n388, new_n303_1, new_n389);
xnor_4 g0114(new_n362, new_n336, new_n390);
not_8  g0115(new_n390, new_n391_1);
xnor_4 g0116(new_n301, n1501, new_n392);
not_8  g0117(new_n392, new_n393);
nand_5 g0118(new_n393, new_n391_1, new_n394);
xnor_4 g0119(new_n392, new_n391_1, new_n395);
xnor_4 g0120(new_n360, new_n338, new_n396);
xnor_4 g0121(new_n299_1, new_n280, new_n397);
nand_5 g0122(new_n397, new_n396, new_n398);
xnor_4 g0123(new_n358, new_n340, new_n399);
not_8  g0124(new_n399, new_n400);
xnor_4 g0125(new_n297, new_n284, new_n401_1);
not_8  g0126(new_n401_1, new_n402_1);
nand_5 g0127(new_n402_1, new_n400, new_n403);
xnor_4 g0128(new_n402_1, new_n399, new_n404);
xnor_4 g0129(new_n295, new_n288, new_n405);
not_8  g0130(new_n405, new_n406);
xnor_4 g0131(n1145, n931, new_n407);
not_8  g0132(new_n407, new_n408);
not_8  g0133(n1530, new_n409);
xnor_4 g0134(new_n351, new_n409, new_n410);
nand_5 g0135(new_n410, new_n408, new_n411);
xnor_4 g0136(new_n293, new_n292_1, new_n412);
not_8  g0137(new_n412, new_n413);
nand_5 g0138(new_n413, new_n411, new_n414_1);
not_8  g0139(new_n411, new_n415);
nand_5 g0140(new_n415, new_n293, new_n416_1);
xnor_4 g0141(new_n311, new_n347_1, new_n417);
xnor_4 g0142(new_n417, new_n352, new_n418);
nand_5 g0143(new_n418, new_n416_1, new_n419);
nand_5 g0144(new_n419, new_n414_1, new_n420);
nand_5 g0145(new_n420, new_n406, new_n421);
not_8  g0146(new_n420, new_n422);
nand_5 g0147(new_n422, new_n405, new_n423_1);
xnor_4 g0148(new_n342, new_n341, new_n424_1);
xnor_4 g0149(new_n424_1, new_n355, new_n425);
nand_5 g0150(new_n425, new_n423_1, new_n426_1);
nand_5 g0151(new_n426_1, new_n421, new_n427);
nand_5 g0152(new_n427, new_n404, new_n428);
nand_5 g0153(new_n428, new_n403, new_n429_1);
not_8  g0154(new_n429_1, new_n430);
not_8  g0155(new_n397, new_n431);
xnor_4 g0156(new_n431, new_n396, new_n432_1);
nand_5 g0157(new_n432_1, new_n430, new_n433_1);
nand_5 g0158(new_n433_1, new_n398, new_n434);
not_8  g0159(new_n434, new_n435);
nand_5 g0160(new_n435, new_n395, new_n436);
nand_5 g0161(new_n436, new_n394, new_n437);
xnor_4 g0162(new_n437, new_n389, n19);
not_8  g0163(n870, new_n439);
not_8  g0164(n1381, new_n440);
nand_5 g0165(new_n440, n402, new_n441);
nand_5 g0166(new_n441, new_n439, new_n442);
not_8  g0167(n66, new_n443);
not_8  g0168(new_n441, new_n444_1);
nand_5 g0169(new_n444_1, new_n443, new_n445);
nand_5 g0170(new_n445, new_n442, new_n446);
xnor_4 g0171(new_n446, n69, new_n447);
not_8  g0172(n585, new_n448);
nand_5 g0173(new_n441, new_n448, new_n449);
not_8  g0174(n968, new_n450);
nand_5 g0175(new_n444_1, new_n450, new_n451);
nand_5 g0176(new_n451, new_n449, new_n452_1);
not_8  g0177(new_n452_1, new_n453);
nand_5 g0178(new_n453, n953, new_n454);
not_8  g0179(n1461, new_n455);
nand_5 g0180(new_n441, new_n455, new_n456);
not_8  g0181(n347, new_n457_1);
nand_5 g0182(new_n444_1, new_n457_1, new_n458);
nand_5 g0183(new_n458, new_n456, new_n459);
not_8  g0184(new_n459, new_n460_1);
nand_5 g0185(new_n460_1, n303, new_n461);
not_8  g0186(new_n461, new_n462);
xnor_4 g0187(new_n452_1, n953, new_n463);
nand_5 g0188(new_n463, new_n462, new_n464);
nand_5 g0189(new_n464, new_n454, new_n465);
xnor_4 g0190(new_n465, new_n447, new_n466);
xnor_4 g0191(new_n466, new_n405, new_n467);
xnor_4 g0192(new_n459, n303, new_n468);
nand_5 g0193(new_n468, new_n408, new_n469_1);
nand_5 g0194(new_n469_1, new_n413, new_n470);
not_8  g0195(new_n463, new_n471);
xnor_4 g0196(new_n471, new_n461, new_n472_1);
not_8  g0197(new_n469_1, new_n473);
nand_5 g0198(new_n473, new_n293, new_n474);
nand_5 g0199(new_n474, new_n470, new_n475);
not_8  g0200(new_n475, new_n476_1);
nand_5 g0201(new_n476_1, new_n472_1, new_n477);
nand_5 g0202(new_n477, new_n470, new_n478);
xnor_4 g0203(new_n478, new_n467, n33);
not_8  g0204(n247, new_n480);
nand_5 g0205(new_n330, new_n367, new_n481);
not_8  g0206(new_n481, new_n482_1);
nand_5 g0207(new_n482_1, new_n480, new_n483);
xnor_4 g0208(new_n483, n1642, new_n484);
nand_5 g0209(new_n484, n1381, new_n485);
not_8  g0210(n379, new_n486);
not_8  g0211(n1527, new_n487);
nand_5 g0212(new_n487, new_n375, new_n488_1);
not_8  g0213(new_n488_1, new_n489);
nand_5 g0214(new_n489, new_n486, new_n490);
nand_5 g0215(new_n488_1, n379, new_n491);
nand_5 g0216(new_n491, n402, new_n492);
not_8  g0217(new_n492, new_n493_1);
nand_5 g0218(new_n493_1, new_n490, new_n494);
nand_5 g0219(n1642, new_n440, new_n495);
nand_5 g0220(new_n495, new_n441, new_n496);
nand_5 g0221(new_n496, new_n494, new_n497);
nand_5 g0222(new_n497, new_n485, new_n498_1);
xnor_4 g0223(new_n481, n247, new_n499);
nand_5 g0224(new_n499, n1381, new_n500);
nand_5 g0225(n1527, n46, new_n501);
nand_5 g0226(new_n501, n402, new_n502);
not_8  g0227(new_n502, new_n503);
nand_5 g0228(new_n503, new_n488_1, new_n504);
nand_5 g0229(new_n440, n247, new_n505);
nand_5 g0230(new_n505, new_n441, new_n506);
nand_5 g0231(new_n506, new_n504, new_n507);
nand_5 g0232(new_n507, new_n500, new_n508);
nand_5 g0233(new_n441, new_n323, new_n509);
nand_5 g0234(new_n444_1, new_n321, new_n510_1);
nand_5 g0235(new_n510_1, new_n509, new_n511);
nand_5 g0236(new_n511, new_n278, new_n512);
xnor_4 g0237(new_n511, n1643, new_n513);
not_8  g0238(n155, new_n514);
nand_5 g0239(new_n441, new_n514, new_n515);
not_8  g0240(n1435, new_n516);
nand_5 g0241(new_n444_1, new_n516, new_n517_1);
nand_5 g0242(new_n517_1, new_n515, new_n518);
not_8  g0243(new_n518, new_n519);
nand_5 g0244(new_n519, n555, new_n520);
nand_5 g0245(new_n446, new_n285, new_n521);
xnor_4 g0246(new_n446, n353, new_n522_1);
nand_5 g0247(new_n452_1, new_n290_1, new_n523);
nand_5 g0248(new_n460_1, n1145, new_n524);
xnor_4 g0249(new_n452_1, n952, new_n525);
nand_5 g0250(new_n525, new_n524, new_n526);
nand_5 g0251(new_n526, new_n523, new_n527);
nand_5 g0252(new_n527, new_n522_1, new_n528);
nand_5 g0253(new_n528, new_n521, new_n529);
not_8  g0254(new_n529, new_n530);
xnor_4 g0255(new_n518, n555, new_n531);
nand_5 g0256(new_n531, new_n530, new_n532_1);
nand_5 g0257(new_n532_1, new_n520, new_n533);
not_8  g0258(new_n533, new_n534_1);
nand_5 g0259(new_n534_1, new_n513, new_n535);
nand_5 g0260(new_n535, new_n512, new_n536);
not_8  g0261(new_n536, new_n537);
nand_5 g0262(n1381, n607, new_n538);
nand_5 g0263(new_n376, n402, new_n539);
not_8  g0264(n402, new_n540);
nand_5 g0265(new_n330, new_n540, new_n541_1);
nand_5 g0266(new_n541_1, new_n539, new_n542);
nand_5 g0267(new_n542, new_n440, new_n543);
nand_5 g0268(new_n543, new_n538, new_n544);
not_8  g0269(new_n544, new_n545);
nand_5 g0270(new_n545, new_n537, new_n546);
not_8  g0271(new_n546, new_n547_1);
nand_5 g0272(n402, n46, new_n548);
nand_5 g0273(new_n540, new_n367, new_n549_1);
nand_5 g0274(new_n549_1, new_n548, new_n550);
nand_5 g0275(new_n550, new_n440, new_n551);
xnor_4 g0276(n607, new_n367, new_n552);
nand_5 g0277(new_n552, n1381, new_n553);
nand_5 g0278(new_n553, new_n551, new_n554);
not_8  g0279(new_n554, new_n555_1);
nand_5 g0280(new_n555_1, new_n547_1, new_n556);
not_8  g0281(new_n556, new_n557_1);
nand_5 g0282(new_n557_1, new_n508, new_n558);
xnor_4 g0283(new_n558, new_n498_1, n1731);
not_8  g0284(n1731, new_n560);
xnor_4 g0285(new_n556, new_n508, n1138);
xnor_4 g0286(new_n545, new_n536, n1727);
xnor_4 g0287(new_n525, new_n524, n1457);
not_8  g0288(n1457, new_n564);
xnor_4 g0289(new_n459, n1145, n1183);
not_8  g0290(n1183, n1237);
nand_5 g0291(n1237, new_n564, new_n567);
not_8  g0292(new_n567, new_n568);
xnor_4 g0293(new_n527, new_n522_1, n416);
not_8  g0294(n416, new_n570);
nand_5 g0295(new_n570, new_n568, new_n571);
not_8  g0296(new_n571, new_n572);
xnor_4 g0297(new_n531, new_n529, n1721);
not_8  g0298(n1721, new_n574);
nand_5 g0299(new_n574, new_n572, new_n575);
xnor_4 g0300(new_n533, new_n513, new_n576);
not_8  g0301(new_n576, n715);
nand_5 g0302(n715, new_n575, new_n578);
not_8  g0303(new_n578, new_n579);
nand_5 g0304(new_n579, n1727, new_n580);
not_8  g0305(new_n580, new_n581);
nand_5 g0306(new_n581, new_n555_1, new_n582);
not_8  g0307(new_n582, new_n583);
nand_5 g0308(new_n583, n1138, new_n584);
nand_5 g0309(new_n584, new_n560, new_n585_1);
not_8  g0310(new_n584, new_n586);
nand_5 g0311(new_n586, new_n498_1, new_n587);
nand_5 g0312(new_n587, new_n585_1, new_n588_1);
not_8  g0313(new_n588_1, n44);
xnor_4 g0314(new_n410, new_n407, n55);
not_8  g0315(n1544, new_n591);
not_8  g0316(n1332, new_n592);
not_8  g0317(n1707, new_n593);
nand_5 g0318(new_n593, new_n278, new_n594);
xnor_4 g0319(n1707, new_n278, new_n595);
not_8  g0320(n1140, new_n596);
nand_5 g0321(new_n596, new_n281, new_n597);
xnor_4 g0322(n1140, new_n281, new_n598);
not_8  g0323(n1351, new_n599_1);
nand_5 g0324(new_n599_1, new_n285, new_n600_1);
xnor_4 g0325(n1351, new_n285, new_n601);
not_8  g0326(n729, new_n602);
nand_5 g0327(new_n290_1, new_n602, new_n603);
nand_5 g0328(n1145, n684, new_n604);
xnor_4 g0329(n952, new_n602, new_n605);
nand_5 g0330(new_n605, new_n604, new_n606);
nand_5 g0331(new_n606, new_n603, new_n607_1);
nand_5 g0332(new_n607_1, new_n601, new_n608);
nand_5 g0333(new_n608, new_n600_1, new_n609);
nand_5 g0334(new_n609, new_n598, new_n610);
nand_5 g0335(new_n610, new_n597, new_n611);
nand_5 g0336(new_n611, new_n595, new_n612);
nand_5 g0337(new_n612, new_n594, new_n613);
nor_7  g0338(new_n613, new_n592, new_n614);
nand_5 g0339(new_n614, n391, new_n615);
xnor_4 g0340(new_n615, new_n591, new_n616);
nand_5 g0341(n266, n155, new_n617);
not_8  g0342(n266, new_n618);
nand_5 g0343(n1435, new_n618, new_n619);
nand_5 g0344(new_n619, new_n617, new_n620);
not_8  g0345(new_n620, new_n621);
nand_5 g0346(n870, n266, new_n622);
nand_5 g0347(new_n618, n66, new_n623);
nand_5 g0348(new_n623, new_n622, new_n624);
not_8  g0349(new_n624, new_n625);
nand_5 g0350(new_n625, new_n621, new_n626);
not_8  g0351(new_n626, new_n627_1);
nand_5 g0352(n1678, n266, new_n628);
nand_5 g0353(n682, new_n618, new_n629);
nand_5 g0354(new_n629, new_n628, new_n630);
not_8  g0355(new_n630, new_n631);
nand_5 g0356(new_n631, new_n627_1, new_n632);
not_8  g0357(new_n632, new_n633);
nand_5 g0358(n1597, new_n618, new_n634);
nand_5 g0359(new_n330, n266, new_n635);
nand_5 g0360(new_n635, new_n634, new_n636);
nand_5 g0361(new_n636, new_n633, new_n637);
nand_5 g0362(n266, new_n367, new_n638_1);
xnor_4 g0363(n1597, new_n375, new_n639);
nand_5 g0364(new_n639, new_n618, new_n640);
nand_5 g0365(new_n640, new_n638_1, new_n641);
xnor_4 g0366(new_n641, new_n637, new_n642);
not_8  g0367(new_n642, new_n643_1);
xnor_4 g0368(new_n636, new_n632, new_n644);
not_8  g0369(new_n644, new_n645);
xnor_4 g0370(new_n631, new_n626, new_n646_1);
not_8  g0371(new_n646_1, new_n647_1);
xnor_4 g0372(new_n624, new_n620, new_n648_1);
nand_5 g0373(new_n648_1, n223, new_n649_1);
xnor_4 g0374(new_n648_1, n223, new_n650);
not_8  g0375(new_n650, new_n651);
nand_5 g0376(new_n625, n444, new_n652);
not_8  g0377(n472, new_n653_1);
nand_5 g0378(n585, n266, new_n654);
nand_5 g0379(n968, new_n618, new_n655_1);
nand_5 g0380(new_n655_1, new_n654, new_n656);
not_8  g0381(new_n656, new_n657);
nand_5 g0382(new_n657, new_n653_1, new_n658);
nand_5 g0383(n1461, n266, new_n659);
nand_5 g0384(n347, new_n618, new_n660);
nand_5 g0385(new_n660, new_n659, new_n661);
nand_5 g0386(new_n661, n801, new_n662);
xnor_4 g0387(new_n656, new_n653_1, new_n663);
nand_5 g0388(new_n663, new_n662, new_n664);
nand_5 g0389(new_n664, new_n658, new_n665_1);
not_8  g0390(new_n665_1, new_n666);
xnor_4 g0391(new_n624, n444, new_n667);
nand_5 g0392(new_n667, new_n666, new_n668);
nand_5 g0393(new_n668, new_n652, new_n669);
nand_5 g0394(new_n669, new_n651, new_n670);
nand_5 g0395(new_n670, new_n649_1, new_n671);
nand_5 g0396(new_n671, new_n647_1, new_n672);
not_8  g0397(new_n672, new_n673);
nand_5 g0398(new_n673, new_n645, new_n674);
not_8  g0399(new_n674, new_n675_1);
nand_5 g0400(new_n675_1, new_n643_1, new_n676);
not_8  g0401(new_n637, new_n677);
nand_5 g0402(new_n641, new_n677, new_n678);
nand_5 g0403(new_n489, new_n376, new_n679);
nand_5 g0404(new_n377, n1527, new_n680);
nand_5 g0405(new_n680, new_n679, new_n681);
not_8  g0406(new_n681, new_n682_1);
nand_5 g0407(new_n682_1, new_n618, new_n683_1);
nand_5 g0408(n266, new_n480, new_n684_1);
nand_5 g0409(new_n684_1, new_n683_1, new_n685);
not_8  g0410(new_n685, new_n686);
xnor_4 g0411(new_n686, new_n678, new_n687);
xnor_4 g0412(new_n687, new_n676, new_n688);
xnor_4 g0413(new_n688, new_n616, new_n689);
xnor_4 g0414(new_n614, n391, new_n690);
xnor_4 g0415(new_n674, new_n643_1, new_n691);
not_8  g0416(new_n691, new_n692);
nand_5 g0417(new_n692, new_n690, new_n693_1);
xnor_4 g0418(new_n672, new_n645, new_n694);
not_8  g0419(new_n694, new_n695_1);
xnor_4 g0420(new_n613, n1332, new_n696);
not_8  g0421(new_n696, new_n697);
nand_5 g0422(new_n697, new_n695_1, new_n698);
xnor_4 g0423(new_n696, new_n695_1, new_n699_1);
xnor_4 g0424(new_n671, new_n646_1, new_n700);
not_8  g0425(new_n700, new_n701);
not_8  g0426(new_n595, new_n702);
xnor_4 g0427(new_n611, new_n702, new_n703);
nand_5 g0428(new_n703, new_n701, new_n704);
xnor_4 g0429(new_n703, new_n700, new_n705);
xnor_4 g0430(new_n669, new_n650, new_n706);
not_8  g0431(new_n706, new_n707);
not_8  g0432(new_n598, new_n708);
xnor_4 g0433(new_n609, new_n708, new_n709);
nand_5 g0434(new_n709, new_n707, new_n710);
xnor_4 g0435(new_n709, new_n706, new_n711);
xnor_4 g0436(new_n667, new_n665_1, new_n712_1);
not_8  g0437(new_n712_1, new_n713);
not_8  g0438(new_n601, new_n714);
xnor_4 g0439(new_n607_1, new_n714, new_n715_1);
nand_5 g0440(new_n715_1, new_n713, new_n716);
not_8  g0441(new_n604, new_n717);
not_8  g0442(new_n605, new_n718);
nand_5 g0443(new_n718, new_n717, new_n719);
not_8  g0444(n684, new_n720);
xnor_4 g0445(n1145, new_n720, new_n721);
not_8  g0446(n801, new_n722);
xnor_4 g0447(new_n661, new_n722, new_n723);
nand_5 g0448(new_n723, new_n721, new_n724_1);
nand_5 g0449(new_n724_1, new_n606, new_n725_1);
not_8  g0450(new_n725_1, new_n726);
nand_5 g0451(new_n726, new_n719, new_n727);
xnor_4 g0452(new_n663, new_n662, new_n728);
not_8  g0453(new_n728, new_n729_1);
not_8  g0454(new_n724_1, new_n730);
nand_5 g0455(new_n730, new_n605, new_n731_1);
nand_5 g0456(new_n731_1, new_n727, new_n732);
not_8  g0457(new_n732, new_n733);
nand_5 g0458(new_n733, new_n729_1, new_n734);
nand_5 g0459(new_n734, new_n727, new_n735);
xnor_4 g0460(new_n715_1, new_n712_1, new_n736);
nand_5 g0461(new_n736, new_n735, new_n737);
nand_5 g0462(new_n737, new_n716, new_n738_1);
nand_5 g0463(new_n738_1, new_n711, new_n739);
nand_5 g0464(new_n739, new_n710, new_n740);
nand_5 g0465(new_n740, new_n705, new_n741);
nand_5 g0466(new_n741, new_n704, new_n742);
nand_5 g0467(new_n742, new_n699_1, new_n743);
nand_5 g0468(new_n743, new_n698, new_n744);
xnor_4 g0469(new_n691, new_n690, new_n745);
nand_5 g0470(new_n745, new_n744, new_n746);
nand_5 g0471(new_n746, new_n693_1, new_n747_1);
xnor_4 g0472(new_n747_1, new_n689, n56);
not_8  g0473(new_n676, new_n749);
nand_5 g0474(new_n687, new_n749, new_n750);
not_8  g0475(new_n750, new_n751);
not_8  g0476(new_n678, new_n752);
nand_5 g0477(new_n685, new_n752, new_n753);
not_8  g0478(n1642, new_n754);
nand_5 g0479(new_n754, n266, new_n755);
xnor_4 g0480(new_n679, new_n486, new_n756);
nand_5 g0481(new_n756, new_n618, new_n757);
nand_5 g0482(new_n757, new_n755, new_n758);
xnor_4 g0483(new_n758, new_n753, new_n759_1);
not_8  g0484(new_n759_1, new_n760);
nand_5 g0485(new_n760, new_n751, new_n761_1);
not_8  g0486(new_n761_1, new_n762);
not_8  g0487(new_n753, new_n763);
nand_5 g0488(new_n758, new_n763, new_n764);
not_8  g0489(n171, new_n765);
nand_5 g0490(n266, new_n765, new_n766);
not_8  g0491(new_n679, new_n767);
nand_5 g0492(new_n767, new_n486, new_n768);
nand_5 g0493(new_n768, n1263, new_n769);
not_8  g0494(n1263, new_n770_1);
not_8  g0495(new_n768, new_n771);
nand_5 g0496(new_n771, new_n770_1, new_n772);
nand_5 g0497(new_n772, new_n618, new_n773_1);
not_8  g0498(new_n773_1, new_n774);
nand_5 g0499(new_n774, new_n769, new_n775);
nand_5 g0500(new_n775, new_n766, new_n776);
xnor_4 g0501(new_n776, new_n764, new_n777);
not_8  g0502(new_n777, new_n778);
nand_5 g0503(new_n778, new_n762, new_n779);
not_8  g0504(new_n764, new_n780);
nand_5 g0505(new_n776, new_n780, new_n781);
nand_5 g0506(n557, n266, new_n782);
not_8  g0507(n1422, new_n783);
not_8  g0508(new_n772, new_n784);
nand_5 g0509(new_n784, new_n783, new_n785);
not_8  g0510(new_n785, new_n786);
nand_5 g0511(new_n786, new_n618, new_n787);
nand_5 g0512(new_n774, n1422, new_n788_1);
nand_5 g0513(new_n788_1, new_n787, new_n789);
not_8  g0514(new_n789, new_n790_1);
nand_5 g0515(new_n790_1, new_n782, new_n791);
not_8  g0516(new_n791, new_n792_1);
xnor_4 g0517(new_n792_1, new_n781, new_n793);
not_8  g0518(new_n793, new_n794);
xnor_4 g0519(new_n794, new_n779, new_n795);
not_8  g0520(new_n615, new_n796);
nand_5 g0521(new_n796, n1544, new_n797);
not_8  g0522(new_n797, new_n798);
nand_5 g0523(new_n798, n649, new_n799);
xnor_4 g0524(new_n778, new_n761_1, new_n800);
not_8  g0525(new_n800, new_n801_1);
nand_5 g0526(new_n801_1, new_n799, new_n802);
xnor_4 g0527(new_n800, new_n799, new_n803);
not_8  g0528(n649, new_n804);
xnor_4 g0529(new_n797, new_n804, new_n805);
xnor_4 g0530(new_n760, new_n750, new_n806);
not_8  g0531(new_n806, new_n807);
nand_5 g0532(new_n807, new_n805, new_n808);
xnor_4 g0533(new_n806, new_n805, new_n809);
not_8  g0534(new_n688, new_n810);
nand_5 g0535(new_n810, new_n616, new_n811);
nand_5 g0536(new_n747_1, new_n689, new_n812);
nand_5 g0537(new_n812, new_n811, new_n813_1);
nand_5 g0538(new_n813_1, new_n809, new_n814);
nand_5 g0539(new_n814, new_n808, new_n815);
nand_5 g0540(new_n815, new_n803, new_n816);
nand_5 g0541(new_n816, new_n802, new_n817);
xnor_4 g0542(new_n817, new_n795, n67);
not_8  g0543(n469, new_n819);
xnor_4 g0544(n1643, new_n819, new_n820);
not_8  g0545(n927, new_n821);
nand_5 g0546(new_n821, new_n281, new_n822);
xnor_4 g0547(n927, new_n281, new_n823_1);
not_8  g0548(n655, new_n824_1);
nand_5 g0549(new_n824_1, new_n285, new_n825);
xnor_4 g0550(n655, new_n285, new_n826);
not_8  g0551(n653, new_n827);
nand_5 g0552(new_n290_1, new_n827, new_n828);
nand_5 g0553(n1764, n1145, new_n829);
xnor_4 g0554(n952, new_n827, new_n830);
nand_5 g0555(new_n830, new_n829, new_n831);
nand_5 g0556(new_n831, new_n828, new_n832);
nand_5 g0557(new_n832, new_n826, new_n833);
nand_5 g0558(new_n833, new_n825, new_n834);
nand_5 g0559(new_n834, new_n823_1, new_n835);
nand_5 g0560(new_n835, new_n822, new_n836_1);
xnor_4 g0561(new_n836_1, new_n820, new_n837);
not_8  g0562(new_n837, new_n838);
xnor_4 g0563(new_n838, new_n396, new_n839_1);
not_8  g0564(new_n823_1, new_n840);
xnor_4 g0565(new_n834, new_n840, new_n841);
nand_5 g0566(new_n841, new_n400, new_n842);
xnor_4 g0567(new_n841, new_n399, new_n843);
not_8  g0568(new_n829, new_n844);
not_8  g0569(new_n830, new_n845);
nand_5 g0570(new_n845, new_n844, new_n846_1);
not_8  g0571(n1145, new_n847);
xnor_4 g0572(n1764, new_n847, new_n848);
nand_5 g0573(new_n848, new_n410, new_n849);
nand_5 g0574(new_n849, new_n831, new_n850);
not_8  g0575(new_n850, new_n851);
nand_5 g0576(new_n851, new_n846_1, new_n852);
not_8  g0577(new_n849, new_n853);
nand_5 g0578(new_n853, new_n830, new_n854);
nand_5 g0579(new_n854, new_n852, new_n855);
not_8  g0580(new_n855, new_n856);
nand_5 g0581(new_n856, new_n418, new_n857);
nand_5 g0582(new_n857, new_n852, new_n858_1);
not_8  g0583(new_n858_1, new_n859);
xnor_4 g0584(new_n832, new_n826, new_n860);
nand_5 g0585(new_n860, new_n859, new_n861);
not_8  g0586(new_n425, new_n862_1);
xnor_4 g0587(new_n860, new_n858_1, new_n863);
nand_5 g0588(new_n863, new_n862_1, new_n864);
nand_5 g0589(new_n864, new_n861, new_n865_1);
not_8  g0590(new_n865_1, new_n866);
nand_5 g0591(new_n866, new_n843, new_n867_1);
nand_5 g0592(new_n867_1, new_n842, new_n868);
xnor_4 g0593(new_n868, new_n839_1, n74);
not_8  g0594(new_n558, new_n870_1);
nand_5 g0595(new_n870_1, new_n498_1, new_n871);
not_8  g0596(new_n871, new_n872);
not_8  g0597(new_n483, new_n873);
nand_5 g0598(new_n873, new_n754, new_n874);
xnor_4 g0599(new_n874, n171, new_n875);
nand_5 g0600(new_n875, n1381, new_n876);
not_8  g0601(new_n490, new_n877);
nand_5 g0602(new_n877, new_n770_1, new_n878);
nand_5 g0603(new_n490, n1263, new_n879);
nand_5 g0604(new_n879, n402, new_n880);
not_8  g0605(new_n880, new_n881);
nand_5 g0606(new_n881, new_n878, new_n882_1);
nand_5 g0607(new_n440, n171, new_n883_1);
nand_5 g0608(new_n883_1, new_n441, new_n884);
nand_5 g0609(new_n884, new_n882_1, new_n885);
nand_5 g0610(new_n885, new_n876, new_n886);
nand_5 g0611(new_n886, new_n872, new_n887);
not_8  g0612(new_n874, new_n888_1);
nand_5 g0613(new_n888_1, new_n765, new_n889);
nand_5 g0614(new_n889, n557, new_n890);
not_8  g0615(n557, new_n891_1);
not_8  g0616(new_n889, new_n892_1);
nand_5 g0617(new_n892_1, new_n891_1, new_n893);
nand_5 g0618(new_n893, n1381, new_n894);
not_8  g0619(new_n894, new_n895);
nand_5 g0620(new_n895, new_n890, new_n896);
nand_5 g0621(n557, new_n540, new_n897);
xnor_4 g0622(new_n878, n1422, new_n898);
nand_5 g0623(new_n898, n402, new_n899);
nand_5 g0624(new_n899, new_n897, new_n900);
not_8  g0625(new_n900, new_n901);
nand_5 g0626(new_n901, new_n440, new_n902_1);
nand_5 g0627(new_n902_1, new_n896, new_n903);
not_8  g0628(new_n903, new_n904);
xnor_4 g0629(new_n904, new_n887, n156);
not_8  g0630(n156, new_n906_1);
not_8  g0631(new_n587, new_n907);
xnor_4 g0632(new_n886, new_n871, n1149);
nand_5 g0633(n1149, new_n907, new_n909);
nand_5 g0634(new_n909, new_n906_1, new_n910);
not_8  g0635(new_n909, new_n911);
nand_5 g0636(new_n911, new_n904, new_n912_1);
nand_5 g0637(new_n912_1, new_n910, new_n913);
not_8  g0638(new_n913, n106);
xnor_4 g0639(new_n555_1, new_n546, n1385);
not_8  g0640(n1385, new_n916);
nand_5 g0641(new_n916, new_n580, new_n917);
nand_5 g0642(new_n917, new_n582, new_n918);
not_8  g0643(new_n918, n126);
xnor_4 g0644(new_n740, new_n705, n135);
nand_5 g0645(new_n631, new_n278, new_n921);
xnor_4 g0646(new_n630, new_n278, new_n922);
nand_5 g0647(new_n621, new_n281, new_n923);
nand_5 g0648(new_n625, new_n285, new_n924);
xnor_4 g0649(new_n624, new_n285, new_n925);
nand_5 g0650(new_n657, new_n290_1, new_n926);
nand_5 g0651(new_n661, n1145, new_n927_1);
xnor_4 g0652(new_n656, new_n290_1, new_n928);
nand_5 g0653(new_n928, new_n927_1, new_n929);
nand_5 g0654(new_n929, new_n926, new_n930);
nand_5 g0655(new_n930, new_n925, new_n931_1);
nand_5 g0656(new_n931_1, new_n924, new_n932);
xnor_4 g0657(new_n620, new_n281, new_n933);
nand_5 g0658(new_n933, new_n932, new_n934);
nand_5 g0659(new_n934, new_n923, new_n935_1);
nand_5 g0660(new_n935_1, new_n922, new_n936);
nand_5 g0661(new_n936, new_n921, new_n937);
nor_7  g0662(new_n937, new_n636, new_n938);
xnor_4 g0663(new_n938, new_n641, n145);
xnor_4 g0664(new_n407, n347, n174);
xnor_4 g0665(new_n392, new_n376, new_n941);
nand_5 g0666(new_n397, n682, new_n942_1);
xnor_4 g0667(new_n397, new_n321, new_n943);
nand_5 g0668(new_n401_1, n1435, new_n944_1);
xnor_4 g0669(new_n401_1, new_n516, new_n945);
nand_5 g0670(new_n405, n66, new_n946);
xnor_4 g0671(new_n405, new_n443, new_n947);
nand_5 g0672(new_n413, new_n450, new_n948);
nand_5 g0673(new_n408, n347, new_n949);
xnor_4 g0674(new_n412, new_n450, new_n950);
nand_5 g0675(new_n950, new_n949, new_n951);
nand_5 g0676(new_n951, new_n948, new_n952_1);
not_8  g0677(new_n952_1, new_n953_1);
nand_5 g0678(new_n953_1, new_n947, new_n954);
nand_5 g0679(new_n954, new_n946, new_n955);
nand_5 g0680(new_n955, new_n945, new_n956);
nand_5 g0681(new_n956, new_n944_1, new_n957);
nand_5 g0682(new_n957, new_n943, new_n958);
nand_5 g0683(new_n958, new_n942_1, new_n959);
xnor_4 g0684(new_n959, new_n941, new_n960);
xnor_4 g0685(new_n957, new_n943, new_n961_1);
xnor_4 g0686(new_n952_1, new_n947, n1426);
not_8  g0687(n1426, n547);
xnor_4 g0688(new_n955, new_n945, n1601);
nand_5 g0689(n1601, n547, new_n965);
not_8  g0690(new_n965, new_n966);
nand_5 g0691(new_n966, new_n961_1, new_n967);
not_8  g0692(new_n967, new_n968_1);
xnor_4 g0693(new_n968_1, new_n960, n181);
xnor_4 g0694(new_n420, new_n405, new_n970);
xnor_4 g0695(new_n970, new_n425, n208);
not_8  g0696(new_n636, new_n972);
not_8  g0697(n213, new_n973);
nand_5 g0698(new_n625, new_n973, new_n974_1);
xnor_4 g0699(new_n624, new_n973, new_n975);
not_8  g0700(n1743, new_n976);
nand_5 g0701(new_n657, new_n976, new_n977);
nand_5 g0702(new_n661, n600, new_n978);
xnor_4 g0703(new_n656, new_n976, new_n979_1);
nand_5 g0704(new_n979_1, new_n978, new_n980_1);
nand_5 g0705(new_n980_1, new_n977, new_n981);
nand_5 g0706(new_n981, new_n975, new_n982);
nand_5 g0707(new_n982, new_n974_1, new_n983);
not_8  g0708(new_n983, new_n984);
nand_5 g0709(new_n984, new_n620, new_n985);
not_8  g0710(new_n985, new_n986);
nand_5 g0711(new_n986, new_n630, new_n987);
xnor_4 g0712(new_n987, new_n972, new_n988);
not_8  g0713(n424, new_n989_1);
nand_5 g0714(new_n278, new_n989_1, new_n990);
xnor_4 g0715(n1643, new_n989_1, new_n991_1);
not_8  g0716(n1363, new_n992);
nand_5 g0717(new_n992, new_n281, new_n993);
xnor_4 g0718(n1363, new_n281, new_n994);
not_8  g0719(n498, new_n995);
nand_5 g0720(new_n995, new_n285, new_n996);
xnor_4 g0721(n498, new_n285, new_n997);
not_8  g0722(n414, new_n998);
nand_5 g0723(new_n290_1, new_n998, new_n999);
nand_5 g0724(n1145, n183, new_n1000_1);
xnor_4 g0725(n952, new_n998, new_n1001);
nand_5 g0726(new_n1001, new_n1000_1, new_n1002);
nand_5 g0727(new_n1002, new_n999, new_n1003);
nand_5 g0728(new_n1003, new_n997, new_n1004);
nand_5 g0729(new_n1004, new_n996, new_n1005_1);
nand_5 g0730(new_n1005_1, new_n994, new_n1006);
nand_5 g0731(new_n1006, new_n993, new_n1007);
nand_5 g0732(new_n1007, new_n991_1, new_n1008);
nand_5 g0733(new_n1008, new_n990, new_n1009);
xnor_4 g0734(new_n1009, n17, new_n1010);
not_8  g0735(new_n1010, new_n1011);
xnor_4 g0736(new_n1011, new_n988, new_n1012_1);
xnor_4 g0737(new_n985, new_n630, new_n1013);
not_8  g0738(new_n1013, new_n1014);
not_8  g0739(new_n991_1, new_n1015_1);
xnor_4 g0740(new_n1007, new_n1015_1, new_n1016_1);
nand_5 g0741(new_n1016_1, new_n1014, new_n1017);
xnor_4 g0742(new_n983, new_n620, new_n1018);
not_8  g0743(new_n1018, new_n1019);
not_8  g0744(new_n994, new_n1020);
xnor_4 g0745(new_n1005_1, new_n1020, new_n1021);
nand_5 g0746(new_n1021, new_n1019, new_n1022);
xnor_4 g0747(new_n1021, new_n1018, new_n1023);
xnor_4 g0748(new_n981, new_n975, new_n1024);
not_8  g0749(new_n1024, new_n1025_1);
not_8  g0750(new_n997, new_n1026);
xnor_4 g0751(new_n1003, new_n1026, new_n1027);
nand_5 g0752(new_n1027, new_n1025_1, new_n1028);
not_8  g0753(new_n1000_1, new_n1029);
not_8  g0754(new_n1001, new_n1030_1);
nand_5 g0755(new_n1030_1, new_n1029, new_n1031);
xnor_4 g0756(n1145, n183, new_n1032);
not_8  g0757(new_n1032, new_n1033);
not_8  g0758(n600, new_n1034);
xnor_4 g0759(new_n661, new_n1034, new_n1035);
nand_5 g0760(new_n1035, new_n1033, new_n1036);
nand_5 g0761(new_n1036, new_n1002, new_n1037);
not_8  g0762(new_n1037, new_n1038);
nand_5 g0763(new_n1038, new_n1031, new_n1039);
xnor_4 g0764(new_n979_1, new_n978, new_n1040);
not_8  g0765(new_n1040, new_n1041);
not_8  g0766(new_n1036, new_n1042);
nand_5 g0767(new_n1042, new_n1001, new_n1043);
nand_5 g0768(new_n1043, new_n1039, new_n1044);
not_8  g0769(new_n1044, new_n1045);
nand_5 g0770(new_n1045, new_n1041, new_n1046);
nand_5 g0771(new_n1046, new_n1039, new_n1047);
xnor_4 g0772(new_n1027, new_n1024, new_n1048);
nand_5 g0773(new_n1048, new_n1047, new_n1049);
nand_5 g0774(new_n1049, new_n1028, new_n1050);
nand_5 g0775(new_n1050, new_n1023, new_n1051);
nand_5 g0776(new_n1051, new_n1022, new_n1052);
xnor_4 g0777(new_n1016_1, new_n1013, new_n1053);
nand_5 g0778(new_n1053, new_n1052, new_n1054);
nand_5 g0779(new_n1054, new_n1017, new_n1055);
xnor_4 g0780(new_n1055, new_n1012_1, n216);
xnor_4 g0781(new_n1048, new_n1047, n218);
xnor_4 g0782(new_n815, new_n803, n231);
not_8  g0783(n1747, new_n1059);
not_8  g0784(n17, new_n1060);
nor_7  g0785(new_n1009, new_n1060, new_n1061);
nand_5 g0786(new_n1061, n961, new_n1062_1);
not_8  g0787(new_n1062_1, new_n1063);
nand_5 g0788(new_n1063, n738, new_n1064);
xnor_4 g0789(new_n1064, new_n1059, new_n1065);
not_8  g0790(new_n758, new_n1066);
not_8  g0791(new_n641, new_n1067_1);
not_8  g0792(new_n987, new_n1068_1);
nand_5 g0793(new_n1068_1, new_n972, new_n1069);
not_8  g0794(new_n1069, new_n1070);
nand_5 g0795(new_n1070, new_n1067_1, new_n1071);
not_8  g0796(new_n1071, new_n1072);
nand_5 g0797(new_n1072, new_n686, new_n1073);
xnor_4 g0798(new_n1073, new_n1066, new_n1074);
xnor_4 g0799(new_n1074, new_n1065, new_n1075);
not_8  g0800(n738, new_n1076);
xnor_4 g0801(new_n1062_1, new_n1076, new_n1077);
xnor_4 g0802(new_n1071, new_n686, new_n1078);
not_8  g0803(new_n1078, new_n1079);
nand_5 g0804(new_n1079, new_n1077, new_n1080);
xnor_4 g0805(new_n1078, new_n1077, new_n1081);
xnor_4 g0806(new_n1061, n961, new_n1082);
xnor_4 g0807(new_n1069, new_n1067_1, new_n1083);
not_8  g0808(new_n1083, new_n1084);
nand_5 g0809(new_n1084, new_n1082, new_n1085);
xnor_4 g0810(new_n1083, new_n1082, new_n1086);
not_8  g0811(new_n988, new_n1087);
nand_5 g0812(new_n1011, new_n1087, new_n1088);
nand_5 g0813(new_n1055, new_n1012_1, new_n1089);
nand_5 g0814(new_n1089, new_n1088, new_n1090);
nand_5 g0815(new_n1090, new_n1086, new_n1091);
nand_5 g0816(new_n1091, new_n1085, new_n1092);
nand_5 g0817(new_n1092, new_n1081, new_n1093);
nand_5 g0818(new_n1093, new_n1080, new_n1094);
xnor_4 g0819(new_n1094, new_n1075, n238);
nand_5 g0820(new_n302, n433, new_n1096);
not_8  g0821(new_n1096, new_n1097);
nand_5 g0822(new_n1097, n1537, new_n1098);
not_8  g0823(new_n1098, new_n1099);
nand_5 g0824(new_n1099, n675, new_n1100);
xnor_4 g0825(new_n1100, n1263, new_n1101);
xnor_4 g0826(new_n1098, n675, new_n1102);
nand_5 g0827(new_n1102, n379, new_n1103_1);
xnor_4 g0828(new_n1102, new_n486, new_n1104);
xnor_4 g0829(new_n1096, n1537, new_n1105);
nand_5 g0830(new_n1105, n1527, new_n1106);
xnor_4 g0831(new_n1105, new_n487, new_n1107);
not_8  g0832(new_n303_1, new_n1108);
nand_5 g0833(new_n1108, n46, new_n1109);
nand_5 g0834(new_n392, n1597, new_n1110);
nand_5 g0835(new_n959, new_n941, new_n1111);
nand_5 g0836(new_n1111, new_n1110, new_n1112);
xnor_4 g0837(new_n303_1, n46, new_n1113_1);
nand_5 g0838(new_n1113_1, new_n1112, new_n1114);
nand_5 g0839(new_n1114, new_n1109, new_n1115);
nand_5 g0840(new_n1115, new_n1107, new_n1116);
nand_5 g0841(new_n1116, new_n1106, new_n1117);
nand_5 g0842(new_n1117, new_n1104, new_n1118);
nand_5 g0843(new_n1118, new_n1103_1, new_n1119_1);
xnor_4 g0844(new_n1119_1, new_n1101, new_n1120);
xnor_4 g0845(new_n1117, new_n1104, new_n1121);
xnor_4 g0846(new_n1115, new_n1107, new_n1122);
nand_5 g0847(new_n968_1, new_n960, new_n1123);
not_8  g0848(new_n1123, new_n1124);
xnor_4 g0849(new_n1113_1, new_n1112, new_n1125);
nand_5 g0850(new_n1125, new_n1124, new_n1126);
not_8  g0851(new_n1126, new_n1127);
nand_5 g0852(new_n1127, new_n1122, new_n1128);
not_8  g0853(new_n1128, new_n1129);
nand_5 g0854(new_n1129, new_n1121, new_n1130);
not_8  g0855(new_n1130, new_n1131);
xnor_4 g0856(new_n1131, new_n1120, n270);
xnor_4 g0857(new_n700, new_n397, new_n1133);
nand_5 g0858(new_n706, new_n401_1, new_n1134);
nand_5 g0859(new_n707, new_n402_1, new_n1135_1);
nand_5 g0860(new_n712_1, new_n405, new_n1136);
nand_5 g0861(new_n713, new_n406, new_n1137);
nand_5 g0862(new_n723, new_n408, new_n1138_1);
nand_5 g0863(new_n1138_1, new_n413, new_n1139);
not_8  g0864(new_n1138_1, new_n1140_1);
nand_5 g0865(new_n1140_1, new_n293, new_n1141);
nand_5 g0866(new_n1141, new_n1139, new_n1142_1);
not_8  g0867(new_n1142_1, new_n1143);
nand_5 g0868(new_n1143, new_n729_1, new_n1144);
nand_5 g0869(new_n1144, new_n1139, new_n1145_1);
not_8  g0870(new_n1145_1, new_n1146);
nand_5 g0871(new_n1146, new_n1137, new_n1147);
nand_5 g0872(new_n1147, new_n1136, new_n1148);
nand_5 g0873(new_n1148, new_n1135_1, new_n1149_1);
nand_5 g0874(new_n1149_1, new_n1134, new_n1150);
xnor_4 g0875(new_n1150, new_n1133, n276);
not_8  g0876(new_n848, new_n1152);
xnor_4 g0877(new_n1152, new_n410, n290);
xnor_4 g0878(new_n950, new_n949, n292);
not_8  g0879(new_n1064, new_n1155);
nand_5 g0880(new_n1155, n1747, new_n1156);
not_8  g0881(new_n776, new_n1157);
not_8  g0882(new_n1073, new_n1158);
nand_5 g0883(new_n1158, new_n1066, new_n1159);
xnor_4 g0884(new_n1159, new_n1157, new_n1160);
not_8  g0885(new_n1160, new_n1161_1);
nand_5 g0886(new_n1161_1, new_n1156, new_n1162_1);
xnor_4 g0887(new_n1160, new_n1156, new_n1163);
not_8  g0888(new_n1074, new_n1164);
nand_5 g0889(new_n1164, new_n1065, new_n1165);
nand_5 g0890(new_n1094, new_n1075, new_n1166);
nand_5 g0891(new_n1166, new_n1165, new_n1167);
nand_5 g0892(new_n1167, new_n1163, new_n1168);
nand_5 g0893(new_n1168, new_n1162_1, new_n1169);
not_8  g0894(new_n787, new_n1170);
not_8  g0895(new_n1159, new_n1171);
nand_5 g0896(new_n1171, new_n1157, new_n1172_1);
nand_5 g0897(new_n1172_1, new_n1170, new_n1173);
not_8  g0898(new_n1173, new_n1174);
nand_5 g0899(new_n1174, new_n1169, new_n1175_1);
not_8  g0900(new_n1175_1, n299);
not_8  g0901(new_n511, new_n1177);
nand_5 g0902(new_n519, n1341, new_n1178);
xnor_4 g0903(new_n518, n1341, new_n1179);
not_8  g0904(new_n446, new_n1180);
nand_5 g0905(new_n1180, n69, new_n1181);
nand_5 g0906(new_n465, new_n447, new_n1182);
nand_5 g0907(new_n1182, new_n1181, new_n1183_1);
nand_5 g0908(new_n1183_1, new_n1179, new_n1184);
nand_5 g0909(new_n1184, new_n1178, new_n1185);
nand_5 g0910(new_n1185, new_n1177, new_n1186);
nor_7  g0911(new_n1186, new_n544, new_n1187);
xnor_4 g0912(new_n1187, new_n555_1, new_n1188);
not_8  g0913(n862, new_n1189);
not_8  g0914(n761, new_n1190);
nand_5 g0915(new_n278, new_n1190, new_n1191_1);
xnor_4 g0916(n1643, new_n1190, new_n1192);
not_8  g0917(n1172, new_n1193);
nand_5 g0918(new_n1193, new_n281, new_n1194_1);
xnor_4 g0919(n1172, new_n281, new_n1195);
not_8  g0920(n695, new_n1196);
nand_5 g0921(new_n1196, new_n285, new_n1197);
xnor_4 g0922(n695, new_n285, new_n1198);
not_8  g0923(n1296, new_n1199_1);
nand_5 g0924(new_n1199_1, new_n290_1, new_n1200);
nand_5 g0925(n1145, n1062, new_n1201_1);
xnor_4 g0926(n1296, new_n290_1, new_n1202_1);
nand_5 g0927(new_n1202_1, new_n1201_1, new_n1203);
nand_5 g0928(new_n1203, new_n1200, new_n1204);
nand_5 g0929(new_n1204, new_n1198, new_n1205);
nand_5 g0930(new_n1205, new_n1197, new_n1206);
nand_5 g0931(new_n1206, new_n1195, new_n1207);
nand_5 g0932(new_n1207, new_n1194_1, new_n1208);
nand_5 g0933(new_n1208, new_n1192, new_n1209);
nand_5 g0934(new_n1209, new_n1191_1, new_n1210);
nor_7  g0935(new_n1210, new_n1189, new_n1211);
xnor_4 g0936(new_n1211, n1222, new_n1212);
not_8  g0937(new_n1212, new_n1213);
xnor_4 g0938(new_n1213, new_n1188, new_n1214);
xnor_4 g0939(new_n1186, new_n545, new_n1215);
not_8  g0940(new_n1215, new_n1216);
xnor_4 g0941(new_n1210, n862, new_n1217);
not_8  g0942(new_n1217, new_n1218);
nand_5 g0943(new_n1218, new_n1216, new_n1219);
xnor_4 g0944(new_n1218, new_n1215, new_n1220);
xnor_4 g0945(new_n1185, new_n511, new_n1221);
not_8  g0946(new_n1221, new_n1222_1);
not_8  g0947(new_n1192, new_n1223);
xnor_4 g0948(new_n1208, new_n1223, new_n1224);
nand_5 g0949(new_n1224, new_n1222_1, new_n1225);
xnor_4 g0950(new_n1224, new_n1221, new_n1226);
xnor_4 g0951(new_n1183_1, new_n1179, new_n1227);
not_8  g0952(new_n1195, new_n1228);
xnor_4 g0953(new_n1206, new_n1228, new_n1229);
nand_5 g0954(new_n1229, new_n1227, new_n1230);
xnor_4 g0955(new_n1206, new_n1195, new_n1231);
xnor_4 g0956(new_n1231, new_n1227, new_n1232);
not_8  g0957(new_n1198, new_n1233);
xnor_4 g0958(new_n1204, new_n1233, new_n1234_1);
nand_5 g0959(new_n1234_1, new_n466, new_n1235_1);
xnor_4 g0960(new_n1204, new_n1198, new_n1236);
xnor_4 g0961(new_n1236, new_n466, new_n1237_1);
not_8  g0962(new_n1201_1, new_n1238);
not_8  g0963(new_n1202_1, new_n1239);
nand_5 g0964(new_n1239, new_n1238, new_n1240);
not_8  g0965(n1062, new_n1241);
xnor_4 g0966(n1145, new_n1241, new_n1242);
nand_5 g0967(new_n1242, new_n468, new_n1243);
nand_5 g0968(new_n1243, new_n1203, new_n1244);
not_8  g0969(new_n1244, new_n1245);
nand_5 g0970(new_n1245, new_n1240, new_n1246);
not_8  g0971(new_n1243, new_n1247);
nand_5 g0972(new_n1247, new_n1202_1, new_n1248);
nand_5 g0973(new_n1248, new_n1246, new_n1249_1);
not_8  g0974(new_n1249_1, new_n1250);
nand_5 g0975(new_n1250, new_n472_1, new_n1251);
nand_5 g0976(new_n1251, new_n1246, new_n1252);
nand_5 g0977(new_n1252, new_n1237_1, new_n1253);
nand_5 g0978(new_n1253, new_n1235_1, new_n1254);
nand_5 g0979(new_n1254, new_n1232, new_n1255_1);
nand_5 g0980(new_n1255_1, new_n1230, new_n1256);
nand_5 g0981(new_n1256, new_n1226, new_n1257);
nand_5 g0982(new_n1257, new_n1225, new_n1258);
nand_5 g0983(new_n1258, new_n1220, new_n1259);
nand_5 g0984(new_n1259, new_n1219, new_n1260_1);
xnor_4 g0985(new_n1260_1, new_n1214, n317);
not_8  g0986(new_n1242, new_n1262);
xnor_4 g0987(new_n1262, new_n468, n372);
not_8  g0988(new_n843, new_n1264);
xnor_4 g0989(new_n865_1, new_n1264, n378);
nand_5 g0990(new_n938, new_n1067_1, new_n1266);
not_8  g0991(new_n1266, new_n1267);
nand_5 g0992(new_n1267, new_n686, new_n1268);
not_8  g0993(new_n1268, new_n1269);
nand_5 g0994(new_n1269, new_n1066, new_n1270);
not_8  g0995(new_n1270, new_n1271);
nand_5 g0996(new_n1271, new_n1157, new_n1272);
not_8  g0997(new_n1272, new_n1273);
nand_5 g0998(new_n1273, new_n791, new_n1274);
not_8  g0999(new_n1274, new_n1275);
nand_5 g1000(new_n1275, new_n787, new_n1276);
nand_5 g1001(new_n1272, new_n1170, new_n1277_1);
nand_5 g1002(new_n1277_1, new_n1276, n1425);
xnor_4 g1003(new_n1270, new_n1157, n1249);
xnor_4 g1004(new_n1266, new_n686, n1119);
xnor_4 g1005(new_n661, new_n847, n647);
not_8  g1006(n647, n1255);
xnor_4 g1007(new_n928, new_n927_1, n646);
not_8  g1008(n646, new_n1284);
nand_5 g1009(new_n1284, n1255, new_n1285);
not_8  g1010(new_n1285, new_n1286);
xnor_4 g1011(new_n930, new_n925, n1016);
not_8  g1012(n1016, new_n1288);
nand_5 g1013(new_n1288, new_n1286, new_n1289);
xnor_4 g1014(new_n933, new_n932, n1683);
nand_5 g1015(n1683, new_n1289, new_n1291);
not_8  g1016(new_n1291, new_n1292);
xnor_4 g1017(new_n935_1, new_n922, n569);
nand_5 g1018(n569, new_n1292, new_n1294);
not_8  g1019(new_n1294, new_n1295);
xnor_4 g1020(new_n937, new_n972, n773);
nand_5 g1021(n773, new_n1295, new_n1297);
not_8  g1022(new_n1297, new_n1298);
nand_5 g1023(new_n1298, new_n1067_1, new_n1299);
not_8  g1024(new_n1299, new_n1300);
nand_5 g1025(new_n1300, n1119, new_n1301);
not_8  g1026(new_n1301, new_n1302);
nand_5 g1027(new_n1302, new_n1066, new_n1303);
not_8  g1028(new_n1303, new_n1304);
nand_5 g1029(new_n1304, n1249, new_n1305_1);
not_8  g1030(new_n1305_1, new_n1306);
nand_5 g1031(new_n1306, new_n791, new_n1307);
xnor_4 g1032(new_n1307, n1425, n387);
nand_5 g1033(new_n1187, new_n555_1, new_n1309);
xnor_4 g1034(new_n1309, new_n508, new_n1310);
nand_5 g1035(new_n1211, n1222, new_n1311);
xnor_4 g1036(new_n1311, n1757, new_n1312);
not_8  g1037(new_n1312, new_n1313);
xnor_4 g1038(new_n1313, new_n1310, new_n1314);
nand_5 g1039(new_n1212, new_n1188, new_n1315_1);
nand_5 g1040(new_n1260_1, new_n1214, new_n1316);
nand_5 g1041(new_n1316, new_n1315_1, new_n1317);
xnor_4 g1042(new_n1317, new_n1314, n401);
xnor_4 g1043(new_n863, new_n425, n423);
xnor_4 g1044(new_n1227, new_n401_1, new_n1320);
nand_5 g1045(new_n466, new_n406, new_n1321_1);
nand_5 g1046(new_n478, new_n467, new_n1322);
nand_5 g1047(new_n1322, new_n1321_1, new_n1323);
xnor_4 g1048(new_n1323, new_n1320, n426);
xnor_4 g1049(new_n1272, new_n791, n493);
not_8  g1050(n493, new_n1326);
nand_5 g1051(new_n1326, new_n1305_1, new_n1327);
nand_5 g1052(new_n1327, new_n1307, new_n1328);
not_8  g1053(new_n1328, n429);
xnor_4 g1054(n773, new_n1294, n432);
xnor_4 g1055(new_n1221, new_n431, new_n1331);
nand_5 g1056(new_n1227, new_n402_1, new_n1332_1);
nand_5 g1057(new_n1323, new_n1320, new_n1333);
nand_5 g1058(new_n1333, new_n1332_1, new_n1334);
xnor_4 g1059(new_n1334, new_n1331, n452);
xnor_4 g1060(new_n1125, new_n1124, n457);
xnor_4 g1061(new_n1167, new_n1163, n460);
not_8  g1062(new_n721, new_n1338_1);
xnor_4 g1063(new_n723, new_n1338_1, n476);
xnor_4 g1064(new_n427, new_n404, n482);
not_8  g1065(new_n1309, new_n1341_1);
nand_5 g1066(new_n1341_1, new_n508, new_n1342);
not_8  g1067(new_n1342, new_n1343);
nand_5 g1068(new_n1343, new_n498_1, new_n1344);
xnor_4 g1069(new_n1344, new_n886, new_n1345);
xnor_4 g1070(new_n1345, new_n1100, new_n1346);
not_8  g1071(new_n1102, new_n1347_1);
xnor_4 g1072(new_n1342, new_n498_1, new_n1348_1);
not_8  g1073(new_n1348_1, new_n1349_1);
nand_5 g1074(new_n1349_1, new_n1347_1, new_n1350);
xnor_4 g1075(new_n1348_1, new_n1347_1, new_n1351_1);
not_8  g1076(new_n1105, new_n1352);
not_8  g1077(new_n1310, new_n1353);
nand_5 g1078(new_n1353, new_n1352, new_n1354);
xnor_4 g1079(new_n1310, new_n1352, new_n1355);
not_8  g1080(new_n1188, new_n1356);
nand_5 g1081(new_n1356, new_n1108, new_n1357);
nand_5 g1082(new_n1216, new_n393, new_n1358);
xnor_4 g1083(new_n1215, new_n393, new_n1359);
nand_5 g1084(new_n1222_1, new_n431, new_n1360);
nand_5 g1085(new_n1334, new_n1331, new_n1361);
nand_5 g1086(new_n1361, new_n1360, new_n1362);
nand_5 g1087(new_n1362, new_n1359, new_n1363_1);
nand_5 g1088(new_n1363_1, new_n1358, new_n1364);
not_8  g1089(new_n1364, new_n1365);
xnor_4 g1090(new_n1188, new_n1108, new_n1366);
nand_5 g1091(new_n1366, new_n1365, new_n1367);
nand_5 g1092(new_n1367, new_n1357, new_n1368);
not_8  g1093(new_n1368, new_n1369_1);
nand_5 g1094(new_n1369_1, new_n1355, new_n1370);
nand_5 g1095(new_n1370, new_n1354, new_n1371);
nand_5 g1096(new_n1371, new_n1351_1, new_n1372);
nand_5 g1097(new_n1372, new_n1350, new_n1373);
xnor_4 g1098(new_n1373, new_n1346, n510);
xnor_4 g1099(new_n1347_1, new_n1074, new_n1375);
nand_5 g1100(new_n1352, new_n1079, new_n1376);
xnor_4 g1101(new_n1352, new_n1078, new_n1377);
nand_5 g1102(new_n1084, new_n303_1, new_n1378);
xnor_4 g1103(new_n1083, new_n303_1, new_n1379);
nand_5 g1104(new_n1087, new_n393, new_n1380);
xnor_4 g1105(new_n988, new_n393, new_n1381_1);
nand_5 g1106(new_n1013, new_n397, new_n1382);
nand_5 g1107(new_n1019, new_n402_1, new_n1383_1);
xnor_4 g1108(new_n1018, new_n402_1, new_n1384);
nand_5 g1109(new_n1025_1, new_n406, new_n1385_1);
xnor_4 g1110(new_n1024, new_n406, new_n1386);
nand_5 g1111(new_n1035, new_n408, new_n1387);
nand_5 g1112(new_n1387, new_n413, new_n1388);
not_8  g1113(new_n1387, new_n1389);
nand_5 g1114(new_n1389, new_n293, new_n1390);
nand_5 g1115(new_n1390, new_n1388, new_n1391);
not_8  g1116(new_n1391, new_n1392);
nand_5 g1117(new_n1392, new_n1041, new_n1393_1);
nand_5 g1118(new_n1393_1, new_n1388, new_n1394);
nand_5 g1119(new_n1394, new_n1386, new_n1395);
nand_5 g1120(new_n1395, new_n1385_1, new_n1396);
nand_5 g1121(new_n1396, new_n1384, new_n1397);
nand_5 g1122(new_n1397, new_n1383_1, new_n1398);
not_8  g1123(new_n1398, new_n1399_1);
xnor_4 g1124(new_n1013, new_n431, new_n1400);
nand_5 g1125(new_n1400, new_n1399_1, new_n1401);
nand_5 g1126(new_n1401, new_n1382, new_n1402);
not_8  g1127(new_n1402, new_n1403);
nand_5 g1128(new_n1403, new_n1381_1, new_n1404);
nand_5 g1129(new_n1404, new_n1380, new_n1405);
nand_5 g1130(new_n1405, new_n1379, new_n1406);
nand_5 g1131(new_n1406, new_n1378, new_n1407_1);
nand_5 g1132(new_n1407_1, new_n1377, new_n1408);
nand_5 g1133(new_n1408, new_n1376, new_n1409);
xnor_4 g1134(new_n1409, new_n1375, n517);
xnor_4 g1135(new_n1347_1, new_n806, new_n1411);
nand_5 g1136(new_n1352, new_n810, new_n1412);
xnor_4 g1137(new_n1352, new_n688, new_n1413);
nand_5 g1138(new_n692, new_n303_1, new_n1414);
nand_5 g1139(new_n695_1, new_n393, new_n1415);
xnor_4 g1140(new_n695_1, new_n392, new_n1416);
nand_5 g1141(new_n700, new_n397, new_n1417);
nand_5 g1142(new_n701, new_n431, new_n1418);
nand_5 g1143(new_n1150, new_n1418, new_n1419);
nand_5 g1144(new_n1419, new_n1417, new_n1420);
not_8  g1145(new_n1420, new_n1421);
nand_5 g1146(new_n1421, new_n1416, new_n1422_1);
nand_5 g1147(new_n1422_1, new_n1415, new_n1423);
xnor_4 g1148(new_n691, new_n303_1, new_n1424);
nand_5 g1149(new_n1424, new_n1423, new_n1425_1);
nand_5 g1150(new_n1425_1, new_n1414, new_n1426_1);
nand_5 g1151(new_n1426_1, new_n1413, new_n1427);
nand_5 g1152(new_n1427, new_n1412, new_n1428);
xnor_4 g1153(new_n1428, new_n1411, n522);
nand_5 g1154(n1601, new_n961_1, new_n1430);
not_8  g1155(new_n1430, new_n1431);
nand_5 g1156(new_n1431, new_n960, new_n1432);
not_8  g1157(new_n1432, new_n1433);
nand_5 g1158(new_n1433, new_n1125, new_n1434);
not_8  g1159(new_n1434, new_n1435_1);
nand_5 g1160(new_n1435_1, new_n1122, new_n1436);
not_8  g1161(new_n1436, new_n1437);
xnor_4 g1162(new_n1437, new_n1121, n532);
not_8  g1163(new_n322, new_n1439);
nand_5 g1164(new_n786, new_n1439, new_n1440_1);
not_8  g1165(new_n372_1, new_n1441);
nand_5 g1166(new_n1441, n247, new_n1442);
not_8  g1167(new_n1442, new_n1443);
nand_5 g1168(new_n1443, n1642, new_n1444);
not_8  g1169(new_n1444, new_n1445);
nand_5 g1170(new_n1445, n171, new_n1446);
not_8  g1171(new_n1446, new_n1447);
nand_5 g1172(new_n1447, n557, new_n1448);
not_8  g1173(new_n1448, new_n1449);
nand_5 g1174(new_n1449, n1000, new_n1450);
not_8  g1175(new_n366, new_n1451);
nand_5 g1176(new_n385, new_n1451, new_n1452);
not_8  g1177(new_n1452, new_n1453_1);
xnor_4 g1178(new_n372_1, new_n480, new_n1454);
nand_5 g1179(new_n1454, n1000, new_n1455);
nand_5 g1180(new_n767, new_n321, new_n1456);
nand_5 g1181(new_n379_1, n1527, new_n1457_1);
nand_5 g1182(new_n1457_1, new_n1456, new_n1458);
not_8  g1183(new_n1458, new_n1459);
nand_5 g1184(new_n1459, new_n305, new_n1460_1);
nand_5 g1185(new_n1460_1, new_n1455, new_n1461_1);
nand_5 g1186(new_n1461_1, new_n1453_1, new_n1462);
not_8  g1187(new_n1462, new_n1463_1);
xnor_4 g1188(new_n1456, n379, new_n1464);
nand_5 g1189(new_n1464, new_n305, new_n1465);
xnor_4 g1190(new_n1442, n1642, new_n1466);
nand_5 g1191(new_n1466, n1000, new_n1467);
nand_5 g1192(new_n1467, new_n1465, new_n1468);
not_8  g1193(new_n1468, new_n1469);
nand_5 g1194(new_n1469, new_n1463_1, new_n1470_1);
not_8  g1195(new_n1470_1, new_n1471);
not_8  g1196(new_n1456, new_n1472);
nand_5 g1197(new_n1472, new_n486, new_n1473);
nand_5 g1198(new_n1473, n1263, new_n1474);
not_8  g1199(new_n380, new_n1475);
not_8  g1200(new_n878, new_n1476);
nand_5 g1201(new_n1476, new_n1475, new_n1477);
nand_5 g1202(new_n1477, new_n1474, new_n1478);
nand_5 g1203(new_n1478, new_n305, new_n1479);
nand_5 g1204(new_n1444, new_n765, new_n1480);
nand_5 g1205(new_n1446, n1000, new_n1481_1);
not_8  g1206(new_n1481_1, new_n1482);
nand_5 g1207(new_n1482, new_n1480, new_n1483);
nand_5 g1208(new_n1483, new_n1479, new_n1484);
not_8  g1209(new_n1484, new_n1485);
nand_5 g1210(new_n1485, new_n1471, new_n1486);
not_8  g1211(new_n1486, new_n1487);
nand_5 g1212(new_n1482, new_n891_1, new_n1488);
nand_5 g1213(new_n1477, n1422, new_n1489);
nand_5 g1214(new_n1489, new_n305, new_n1490);
nand_5 g1215(new_n1490, new_n1450, new_n1491);
not_8  g1216(new_n1491, new_n1492);
nand_5 g1217(new_n1492, new_n1488, new_n1493);
nand_5 g1218(new_n1493, new_n1440_1, new_n1494);
not_8  g1219(new_n1494, new_n1495_1);
nand_5 g1220(new_n1495_1, new_n1487, new_n1496);
not_8  g1221(new_n1496, new_n1497);
nand_5 g1222(new_n1497, new_n1450, new_n1498_1);
nand_5 g1223(new_n1498_1, new_n1440_1, new_n1499);
xnor_4 g1224(new_n1495_1, new_n1486, new_n1500);
not_8  g1225(new_n1500, new_n1501_1);
xnor_4 g1226(new_n1469, new_n1462, new_n1502_1);
not_8  g1227(new_n1502_1, new_n1503);
not_8  g1228(new_n364, new_n1504);
nand_5 g1229(new_n387_1, new_n1504, new_n1505);
not_8  g1230(new_n1505, new_n1506);
xnor_4 g1231(new_n1461_1, new_n1452, new_n1507_1);
not_8  g1232(new_n1507_1, new_n1508);
nand_5 g1233(new_n1508, new_n1506, new_n1509);
not_8  g1234(new_n1509, new_n1510);
nand_5 g1235(new_n1510, new_n1503, new_n1511);
not_8  g1236(new_n1511, new_n1512);
xnor_4 g1237(new_n1485, new_n1470_1, new_n1513);
not_8  g1238(new_n1513, new_n1514);
nand_5 g1239(new_n1514, new_n1512, new_n1515);
not_8  g1240(new_n1515, new_n1516);
nand_5 g1241(new_n1516, new_n1501_1, new_n1517);
nand_5 g1242(new_n1517, new_n1499, new_n1518);
not_8  g1243(new_n1518, new_n1519);
xnor_4 g1244(new_n1515, new_n1501_1, new_n1520);
not_8  g1245(n49, new_n1521);
nand_5 g1246(new_n278, new_n819, new_n1522);
nand_5 g1247(new_n836_1, new_n820, new_n1523);
nand_5 g1248(new_n1523, new_n1522, new_n1524);
nor_7  g1249(new_n1524, new_n1521, new_n1525_1);
nand_5 g1250(new_n1525_1, n1622, new_n1526);
not_8  g1251(new_n1526, new_n1527_1);
nand_5 g1252(new_n1527_1, n906, new_n1528);
not_8  g1253(new_n1528, new_n1529);
nand_5 g1254(new_n1529, n277, new_n1530_1);
xnor_4 g1255(new_n1514, new_n1511, new_n1531);
not_8  g1256(new_n1531, new_n1532);
nand_5 g1257(new_n1532, new_n1530_1, new_n1533);
xnor_4 g1258(new_n1531, new_n1530_1, new_n1534);
not_8  g1259(n277, new_n1535_1);
xnor_4 g1260(new_n1528, new_n1535_1, new_n1536);
xnor_4 g1261(new_n1509, new_n1503, new_n1537_1);
not_8  g1262(new_n1537_1, new_n1538);
nand_5 g1263(new_n1538, new_n1536, new_n1539);
xnor_4 g1264(new_n1537_1, new_n1536, new_n1540);
not_8  g1265(n906, new_n1541);
xnor_4 g1266(new_n1526, new_n1541, new_n1542);
xnor_4 g1267(new_n1508, new_n1505, new_n1543);
not_8  g1268(new_n1543, new_n1544_1);
nand_5 g1269(new_n1544_1, new_n1542, new_n1545);
xnor_4 g1270(new_n1543, new_n1542, new_n1546);
not_8  g1271(new_n388, new_n1547);
xnor_4 g1272(new_n1525_1, n1622, new_n1548);
nand_5 g1273(new_n1548, new_n1547, new_n1549);
xnor_4 g1274(new_n1548, new_n388, new_n1550);
xnor_4 g1275(new_n1524, n49, new_n1551);
nand_5 g1276(new_n1551, new_n390, new_n1552);
xnor_4 g1277(new_n1551, new_n390, new_n1553);
not_8  g1278(new_n1553, new_n1554);
nand_5 g1279(new_n837, new_n396, new_n1555);
not_8  g1280(new_n868, new_n1556_1);
nand_5 g1281(new_n1556_1, new_n839_1, new_n1557);
nand_5 g1282(new_n1557, new_n1555, new_n1558);
nand_5 g1283(new_n1558, new_n1554, new_n1559);
nand_5 g1284(new_n1559, new_n1552, new_n1560);
not_8  g1285(new_n1560, new_n1561);
nand_5 g1286(new_n1561, new_n1550, new_n1562);
nand_5 g1287(new_n1562, new_n1549, new_n1563);
nand_5 g1288(new_n1563, new_n1546, new_n1564);
nand_5 g1289(new_n1564, new_n1545, new_n1565);
nand_5 g1290(new_n1565, new_n1540, new_n1566);
nand_5 g1291(new_n1566, new_n1539, new_n1567);
nand_5 g1292(new_n1567, new_n1534, new_n1568);
nand_5 g1293(new_n1568, new_n1533, new_n1569);
not_8  g1294(new_n1569, new_n1570);
nand_5 g1295(new_n1570, new_n1520, new_n1571);
nand_5 g1296(new_n1571, new_n1519, new_n1572);
not_8  g1297(new_n1572, n534);
xnor_4 g1298(n1721, new_n571, n541);
nand_5 g1299(new_n1161_1, new_n1100, new_n1575);
xnor_4 g1300(new_n1160, new_n1100, new_n1576);
nand_5 g1301(new_n1347_1, new_n1164, new_n1577);
nand_5 g1302(new_n1409, new_n1375, new_n1578);
nand_5 g1303(new_n1578, new_n1577, new_n1579);
nand_5 g1304(new_n1579, new_n1576, new_n1580);
nand_5 g1305(new_n1580, new_n1575, new_n1581);
nand_5 g1306(new_n1581, new_n1174, new_n1582);
not_8  g1307(new_n1582, n549);
xnor_4 g1308(new_n1424, new_n1423, n559);
xnor_4 g1309(new_n1400, new_n1398, n573);
xnor_4 g1310(new_n1579, new_n1576, n588);
xnor_4 g1311(n416, new_n567, n599);
not_8  g1312(new_n1277_1, n824);
nand_5 g1313(new_n1305_1, n824, new_n1589);
not_8  g1314(new_n1589, n627);
xnor_4 g1315(new_n1172_1, new_n791, new_n1591);
xnor_4 g1316(new_n1591, new_n1169, n638);
not_8  g1317(new_n887, new_n1593);
nand_5 g1318(new_n904, new_n1593, new_n1594);
nand_5 g1319(new_n1476, new_n783, new_n1595_1);
not_8  g1320(new_n1595_1, new_n1596);
nand_5 g1321(new_n1596, new_n444_1, new_n1597_1);
not_8  g1322(new_n893, new_n1598);
nand_5 g1323(new_n1598, n1381, new_n1599);
nand_5 g1324(new_n1599, new_n1597_1, new_n1600_1);
nand_5 g1325(new_n1600_1, new_n1594, new_n1601_1);
not_8  g1326(new_n1601_1, n643);
xnor_4 g1327(new_n1558, new_n1553, n648);
xnor_4 g1328(new_n742, new_n699_1, n665);
xnor_4 g1329(new_n1092, new_n1081, n683);
not_8  g1330(new_n1520, new_n1606);
nand_5 g1331(new_n1606, new_n1100, new_n1607);
xnor_4 g1332(new_n1520, new_n1100, new_n1608);
nand_5 g1333(new_n1532, new_n1100, new_n1609);
xnor_4 g1334(new_n1531, new_n1100, new_n1610);
nand_5 g1335(new_n1538, new_n1347_1, new_n1611);
xnor_4 g1336(new_n1537_1, new_n1347_1, new_n1612);
nand_5 g1337(new_n1544_1, new_n1352, new_n1613_1);
xnor_4 g1338(new_n1543, new_n1352, new_n1614);
nand_5 g1339(new_n1547, new_n303_1, new_n1615);
nand_5 g1340(new_n437, new_n389, new_n1616);
nand_5 g1341(new_n1616, new_n1615, new_n1617);
nand_5 g1342(new_n1617, new_n1614, new_n1618);
nand_5 g1343(new_n1618, new_n1613_1, new_n1619);
nand_5 g1344(new_n1619, new_n1612, new_n1620);
nand_5 g1345(new_n1620, new_n1611, new_n1621);
nand_5 g1346(new_n1621, new_n1610, new_n1622_1);
nand_5 g1347(new_n1622_1, new_n1609, new_n1623);
nand_5 g1348(new_n1623, new_n1608, new_n1624);
nand_5 g1349(new_n1624, new_n1607, new_n1625);
not_8  g1350(new_n1499, new_n1626);
not_8  g1351(new_n1450, new_n1627);
nand_5 g1352(new_n1486, new_n1627, new_n1628);
nand_5 g1353(new_n1628, new_n1626, new_n1629_1);
not_8  g1354(new_n1629_1, new_n1630);
xnor_4 g1355(new_n1630, new_n1517, new_n1631);
not_8  g1356(new_n1631, new_n1632);
nand_5 g1357(new_n1632, new_n1625, new_n1633_1);
nand_5 g1358(new_n1631, new_n1100, new_n1634);
not_8  g1359(new_n1100, new_n1635_1);
nand_5 g1360(new_n1624, new_n1635_1, new_n1636);
nand_5 g1361(new_n1636, new_n1634, new_n1637);
not_8  g1362(new_n1637, new_n1638);
nand_5 g1363(new_n1638, new_n1633_1, new_n1639);
xnor_4 g1364(new_n1639, new_n1519, n699);
not_8  g1365(new_n418, new_n1641);
xnor_4 g1366(new_n855, new_n1641, n712);
not_8  g1367(n145, new_n1643_1);
nand_5 g1368(new_n1297, new_n1643_1, new_n1644);
nand_5 g1369(new_n1644, new_n1299, new_n1645);
not_8  g1370(new_n1645, n724);
xnor_4 g1371(n1016, new_n1285, n725);
xnor_4 g1372(new_n1426_1, new_n1413, n731);
xnor_4 g1373(new_n1617, new_n1614, n748);
not_8  g1374(new_n1355, new_n1650);
xnor_4 g1375(new_n1368, new_n1650, n759);
nand_5 g1376(new_n1437, new_n1121, new_n1652);
not_8  g1377(new_n1652, new_n1653);
nand_5 g1378(new_n1653, new_n1120, new_n1654_1);
not_8  g1379(new_n1654_1, new_n1655);
nand_5 g1380(new_n1100, new_n770_1, new_n1656);
not_8  g1381(new_n1119_1, new_n1657_1);
nand_5 g1382(new_n1657_1, new_n1101, new_n1658);
nand_5 g1383(new_n1658, new_n1656, new_n1659);
nand_5 g1384(new_n1659, new_n783, new_n1660_1);
not_8  g1385(new_n1660_1, new_n1661);
nand_5 g1386(new_n1661, new_n1655, new_n1662);
not_8  g1387(new_n1662, n770);
not_8  g1388(new_n1381_1, new_n1664);
xnor_4 g1389(new_n1402, new_n1664, n790);
xnor_4 g1390(new_n1100, new_n800, new_n1666);
nand_5 g1391(new_n1347_1, new_n807, new_n1667);
nand_5 g1392(new_n1428, new_n1411, new_n1668);
nand_5 g1393(new_n1668, new_n1667, new_n1669);
xnor_4 g1394(new_n1669, new_n1666, n792);
xnor_4 g1395(new_n1053, new_n1052, n813);
xnor_4 g1396(new_n1252, new_n1237_1, n823);
not_8  g1397(new_n472_1, new_n1673);
xnor_4 g1398(new_n475, new_n1673, n836);
xnor_4 g1399(new_n1619, new_n1612, n846);
xnor_4 g1400(new_n1258, new_n1220, n858);
xnor_4 g1401(new_n1268, new_n1066, n865);
xnor_4 g1402(new_n1407_1, new_n1377, n867);
not_8  g1403(new_n1344, new_n1679);
nand_5 g1404(new_n1679, new_n886, new_n1680);
xnor_4 g1405(new_n1680, new_n904, new_n1681);
not_8  g1406(new_n1345, new_n1682);
nand_5 g1407(new_n1682, new_n1100, new_n1683_1);
nand_5 g1408(new_n1373, new_n1346, new_n1684);
nand_5 g1409(new_n1684, new_n1683_1, new_n1685);
xnor_4 g1410(new_n1685, new_n1681, n883);
xnor_4 g1411(new_n745, new_n744, n888);
not_8  g1412(new_n1311, new_n1688_1);
nand_5 g1413(new_n1688_1, n1757, new_n1689);
not_8  g1414(new_n1689, new_n1690_1);
nand_5 g1415(new_n1690_1, n839, new_n1691);
nand_5 g1416(new_n1691, new_n1682, new_n1692);
xnor_4 g1417(new_n1691, new_n1345, new_n1693);
xnor_4 g1418(new_n1689, n839, new_n1694);
not_8  g1419(new_n1694, new_n1695);
nand_5 g1420(new_n1695, new_n1349_1, new_n1696);
xnor_4 g1421(new_n1695, new_n1348_1, new_n1697);
nand_5 g1422(new_n1313, new_n1353, new_n1698);
nand_5 g1423(new_n1317, new_n1314, new_n1699);
nand_5 g1424(new_n1699, new_n1698, new_n1700);
nand_5 g1425(new_n1700, new_n1697, new_n1701);
nand_5 g1426(new_n1701, new_n1696, new_n1702);
nand_5 g1427(new_n1702, new_n1693, new_n1703);
nand_5 g1428(new_n1703, new_n1692, new_n1704);
xnor_4 g1429(new_n1704, new_n1681, n891);
not_8  g1430(new_n1680, new_n1706);
nand_5 g1431(new_n1706, new_n904, new_n1707_1);
not_8  g1432(new_n1704, new_n1708);
nand_5 g1433(new_n1708, new_n1681, new_n1709);
nand_5 g1434(new_n1709, new_n1707_1, new_n1710);
not_8  g1435(new_n1710, new_n1711);
nand_5 g1436(new_n1711, new_n1600_1, new_n1712);
not_8  g1437(new_n1712, n892);
xnor_4 g1438(new_n1035, new_n1032, n902);
xnor_4 g1439(new_n706, new_n401_1, new_n1715);
xnor_4 g1440(new_n1715, new_n1148, n905);
xnor_4 g1441(new_n1127, new_n1122, n912);
xnor_4 g1442(n1149, new_n587, n935);
xnor_4 g1443(new_n1299, n1119, n942);
xnor_4 g1444(new_n1090, new_n1086, n944);
nand_5 g1445(n770, n547, new_n1721_1);
not_8  g1446(new_n1721_1, n974);
not_8  g1447(new_n395, new_n1723);
xnor_4 g1448(new_n434, new_n1723, n979);
not_8  g1449(new_n817, new_n1725);
nand_5 g1450(new_n1725, new_n795, new_n1726);
not_8  g1451(new_n779, new_n1727_1);
nand_5 g1452(new_n794, new_n1727_1, new_n1728);
not_8  g1453(new_n781, new_n1729_1);
nand_5 g1454(new_n792_1, new_n1729_1, new_n1730);
nand_5 g1455(new_n1730, new_n787, new_n1731_1);
nand_5 g1456(new_n1731_1, new_n1728, new_n1732);
not_8  g1457(new_n1732, new_n1733);
nand_5 g1458(new_n1733, new_n1726, new_n1734);
not_8  g1459(new_n1734, n980);
xnor_4 g1460(new_n1405, new_n1379, n989);
xnor_4 g1461(new_n1623, new_n1608, n991);
xnor_4 g1462(new_n1700, new_n1697, n1005);
xnor_4 g1463(new_n1371, new_n1351_1, n1012);
xnor_4 g1464(new_n1431, new_n960, n1015);
not_8  g1465(new_n1726, new_n1741);
not_8  g1466(new_n1731_1, new_n1742);
nand_5 g1467(new_n1742, new_n1741, new_n1743_1);
xnor_4 g1468(new_n1731_1, new_n1728, new_n1744);
nand_5 g1469(new_n1744, new_n1726, new_n1745);
nand_5 g1470(new_n1745, new_n1743_1, n1025);
xnor_4 g1471(new_n1702, new_n1693, n1030);
xnor_4 g1472(new_n813_1, new_n809, n1067);
not_8  g1473(new_n1600_1, new_n1749);
xnor_4 g1474(new_n1710, new_n1749, n1068);
xnor_4 g1475(new_n576, new_n575, n1103);
xnor_4 g1476(new_n468, new_n407, n1113);
not_8  g1477(new_n1659, new_n1753);
nand_5 g1478(new_n1753, n1422, new_n1754);
not_8  g1479(new_n1754, new_n1755);
nand_5 g1480(new_n1755, new_n1654_1, new_n1756);
nand_5 g1481(new_n1756, new_n1662, n1135);
not_8  g1482(new_n1571, new_n1758);
nand_5 g1483(new_n1630, new_n1758, new_n1759);
nand_5 g1484(new_n1632, new_n1571, new_n1760);
nand_5 g1485(new_n1760, new_n1759, n1142);
xnor_4 g1486(new_n1631, new_n1635_1, new_n1762);
xnor_4 g1487(new_n1762, new_n1625, n1161);
xnor_4 g1488(new_n1433, new_n1125, n1162);
not_8  g1489(n865, new_n1765);
nand_5 g1490(new_n1765, new_n1301, new_n1766);
nand_5 g1491(new_n1766, new_n1303, new_n1767);
not_8  g1492(new_n1767, n1175);
nand_5 g1493(new_n1100, new_n801_1, new_n1769);
nand_5 g1494(new_n1669, new_n1666, new_n1770);
nand_5 g1495(new_n1770, new_n1769, new_n1771);
not_8  g1496(new_n795, new_n1772);
nand_5 g1497(new_n1635_1, new_n1772, new_n1773);
nand_5 g1498(new_n1773, new_n1771, new_n1774);
nand_5 g1499(new_n1100, new_n795, new_n1775);
nand_5 g1500(new_n1775, new_n1770, new_n1776);
nand_5 g1501(new_n1776, new_n1774, new_n1777);
xnor_4 g1502(new_n1777, new_n1744, n1191);
xnor_4 g1503(new_n1435_1, new_n1122, n1194);
xnor_4 g1504(new_n432_1, new_n429_1, n1199);
xnor_4 g1505(new_n1394, new_n1386, n1201);
not_8  g1506(new_n929, new_n1782);
not_8  g1507(new_n661, new_n1783);
nand_5 g1508(new_n1783, new_n847, new_n1784);
nand_5 g1509(new_n1784, new_n1782, new_n1785);
nand_5 g1510(new_n1785, new_n1285, n1202);
xnor_4 g1511(n569, new_n1291, n1234);
xnor_4 g1512(new_n1653, new_n1120, n1235);
not_8  g1513(new_n1172_1, new_n1789);
nand_5 g1514(new_n1789, new_n791, new_n1790);
not_8  g1515(new_n1169, new_n1791);
nand_5 g1516(new_n1591, new_n1791, new_n1792);
nand_5 g1517(new_n1792, new_n1790, new_n1793);
nand_5 g1518(new_n1793, new_n787, new_n1794);
nand_5 g1519(new_n1794, new_n1175_1, n1260);
xnor_4 g1520(new_n1303, n1249, n1277);
not_8  g1521(new_n1685, new_n1797);
nand_5 g1522(new_n1797, new_n1681, new_n1798);
nand_5 g1523(new_n1798, new_n1707_1, new_n1799);
not_8  g1524(new_n1799, new_n1800);
nand_5 g1525(new_n1800, new_n1600_1, new_n1801);
not_8  g1526(new_n1801, n1278);
not_8  g1527(new_n414_1, new_n1803);
nand_5 g1528(new_n418, new_n1803, new_n1804);
not_8  g1529(new_n416_1, new_n1805);
nand_5 g1530(new_n1641, new_n1805, new_n1806);
nand_5 g1531(new_n1806, new_n422, new_n1807);
nand_5 g1532(new_n1807, new_n1804, new_n1808);
not_8  g1533(new_n1808, n1283);
nand_5 g1534(new_n1131, new_n1120, new_n1810);
nand_5 g1535(new_n1755, new_n1810, new_n1811);
nand_5 g1536(new_n1811, new_n1721_1, n1305);
xnor_4 g1537(new_n578, n1727, n1315);
xnor_4 g1538(new_n1565, new_n1540, n1330);
not_8  g1539(new_n1416, new_n1815);
xnor_4 g1540(new_n1420, new_n1815, n1338);
xnor_4 g1541(new_n732, new_n728, n1340);
xnor_4 g1542(new_n1569, new_n1520, n1347);
xnor_4 g1543(new_n1749, new_n1594, new_n1819);
not_8  g1544(new_n1819, n1348);
xnor_4 g1545(new_n1256, new_n1226, n1349);
xnor_4 g1546(new_n1659, n1422, new_n1822);
xnor_4 g1547(new_n1822, new_n1654_1, n1369);
xnor_4 g1548(new_n1822, new_n1810, n1383);
not_8  g1549(new_n1550, new_n1825);
xnor_4 g1550(new_n1560, new_n1825, n1393);
xnor_4 g1551(new_n1391, new_n1040, n1399);
xnor_4 g1552(new_n712_1, new_n406, new_n1828);
xnor_4 g1553(new_n1828, new_n1145_1, n1407);
nand_5 g1554(n643, new_n912_1, new_n1830);
not_8  g1555(new_n1830, n1440);
xnor_4 g1556(n1601, new_n961_1, n1453);
xnor_4 g1557(new_n1142_1, new_n728, n1460);
xnor_4 g1558(new_n1100, new_n795, new_n1834);
xnor_4 g1559(new_n1834, new_n1771, n1463);
xnor_4 g1560(new_n1129, new_n1121, n1470);
xnor_4 g1561(new_n1035, new_n407, n1481);
xnor_4 g1562(new_n736, new_n735, n1495);
xnor_4 g1563(new_n1050, new_n1023, n1498);
xnor_4 g1564(new_n1563, new_n1546, n1502);
xnor_4 g1565(new_n1254, new_n1232, n1507);
not_8  g1566(new_n1289, new_n1842);
xnor_4 g1567(n1683, new_n1842, n1525);
xnor_4 g1568(new_n738_1, new_n711, n1535);
xnor_4 g1569(n1601, n547, n1556);
not_8  g1570(new_n912_1, new_n1846);
xnor_4 g1571(new_n1819, new_n1846, n1595);
xnor_4 g1572(new_n1396, new_n1384, n1600);
not_8  g1573(new_n526, new_n1849);
nand_5 g1574(new_n459, new_n847, new_n1850);
nand_5 g1575(new_n1850, new_n1849, new_n1851);
nand_5 g1576(new_n1851, new_n567, n1613);
xnor_4 g1577(new_n1249_1, new_n1673, n1629);
nand_5 g1578(new_n1777, new_n1732, new_n1854);
not_8  g1579(new_n1728, new_n1855);
nand_5 g1580(new_n1742, new_n1855, new_n1856);
not_8  g1581(new_n1771, new_n1857);
not_8  g1582(new_n1775, new_n1858);
nand_5 g1583(new_n1858, new_n1857, new_n1859);
nand_5 g1584(new_n1859, new_n1856, new_n1860);
not_8  g1585(new_n1860, new_n1861);
nand_5 g1586(new_n1861, new_n1854, new_n1862);
not_8  g1587(new_n1862, n1633);
xnor_4 g1588(new_n966, new_n961_1, n1635);
xnor_4 g1589(new_n1366, new_n1364, n1654);
xnor_4 g1590(new_n582, n1138, n1657);
xnor_4 g1591(new_n1799, new_n1749, n1660);
xnor_4 g1592(new_n1044, new_n1040, n1675);
xnor_4 g1593(new_n1591, new_n1581, n1686);
xnor_4 g1594(new_n723, new_n407, n1688);
xnor_4 g1595(new_n1567, new_n1534, n1690);
xnor_4 g1596(new_n1621, new_n1610, n1729);
not_8  g1597(new_n1581, new_n1873);
nand_5 g1598(new_n1591, new_n1873, new_n1874);
nand_5 g1599(new_n1874, new_n1790, new_n1875);
nand_5 g1600(new_n1875, new_n787, new_n1876);
nand_5 g1601(new_n1876, new_n1582, n1737);
xnor_4 g1602(new_n1362, new_n1359, n1746);
xnor_4 g1603(new_n407, n347, n488);
xnor_4 g1604(new_n950, new_n949, n1677);
endmodule


