// Benchmark "top_809698493_843330999_809698999_896665269_4392119" written by ABC on Fri Jun 14 22:43:13 2024

module top_809698493_843330999_809698999_896665269_4392119 ( 
    n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753, n783,
    n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333, n1353,
    n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835, n1906,
    n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433, n2464,
    n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551, n2558,
    n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172, n3342,
    n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986, n3992,
    n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312, n4370,
    n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828, n4903,
    n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212, n5240,
    n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694, n5760,
    n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126, n6254,
    n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611, n6687,
    n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159, n7160,
    n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456, n7500,
    n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862, n7891,
    n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433, n8476,
    n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195, n9241,
    n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956, n10022,
    n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451, n10510,
    n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928, n10965,
    n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407, n11423,
    n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876, n11877,
    n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044, n12069,
    n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591, n12648,
    n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826, n12925,
    n12947,
    n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807  );
  input  n45, n137, n159, n217, n405, n447, n503, n521, n533, n615, n753,
    n783, n806, n996, n1067, n1094, n1097, n1198, n1199, n1209, n1333,
    n1353, n1357, n1471, n1478, n1510, n1512, n1564, n1576, n1798, n1835,
    n1906, n1980, n2024, n2087, n2226, n2253, n2278, n2347, n2393, n2433,
    n2464, n2498, n2507, n2508, n2509, n2512, n2515, n2522, n2530, n2551,
    n2558, n2564, n2577, n2585, n2749, n2802, n2879, n3022, n3146, n3172,
    n3342, n3602, n3616, n3627, n3719, n3754, n3842, n3865, n3932, n3986,
    n3992, n4005, n4086, n4094, n4141, n4187, n4189, n4190, n4203, n4312,
    n4370, n4436, n4499, n4516, n4634, n4722, n4805, n4817, n4826, n4828,
    n4903, n4921, n4928, n4938, n4970, n5069, n5105, n5153, n5198, n5212,
    n5240, n5283, n5305, n5314, n5319, n5320, n5331, n5579, n5645, n5694,
    n5760, n5767, n5798, n5814, n5857, n5860, n5964, n6016, n6038, n6126,
    n6254, n6294, n6358, n6359, n6429, n6431, n6441, n6578, n6604, n6611,
    n6687, n6703, n6770, n6776, n6797, n6806, n6826, n6877, n6986, n7159,
    n7160, n7236, n7265, n7270, n7294, n7320, n7354, n7388, n7436, n7456,
    n7500, n7523, n7546, n7610, n7646, n7690, n7730, n7733, n7823, n7862,
    n7891, n7946, n7965, n8028, n8065, n8236, n8276, n8336, n8384, n8433,
    n8476, n8595, n8665, n8717, n8759, n8819, n9080, n9111, n9189, n9195,
    n9241, n9400, n9457, n9583, n9637, n9640, n9725, n9763, n9920, n9956,
    n10022, n10174, n10217, n10223, n10278, n10327, n10391, n10439, n10451,
    n10510, n10545, n10547, n10644, n10678, n10685, n10848, n10898, n10928,
    n10965, n10990, n11023, n11153, n11222, n11257, n11296, n11311, n11407,
    n11423, n11478, n11536, n11662, n11728, n11757, n11791, n11821, n11876,
    n11877, n11892, n11917, n11922, n11967, n11999, n12000, n12025, n12044,
    n12069, n12145, n12221, n12247, n12299, n12391, n12489, n12511, n12591,
    n12648, n12704, n12705, n12706, n12709, n12720, n12753, n12777, n12826,
    n12925, n12947;
  output n112, n226, n381, n397, n658, n671, n837, n844, n911, n992, n1020,
    n1136, n1138, n1269, n1523, n1658, n1847, n2096, n2131, n2301, n2316,
    n2383, n2425, n2431, n2434, n2581, n2624, n2679, n2708, n2818, n2902,
    n3071, n3124, n3214, n3230, n3272, n3287, n3339, n3456, n3654, n3661,
    n3677, n3849, n4088, n4155, n4159, n4226, n4230, n4300, n4326, n4333,
    n4378, n4397, n4553, n4686, n4689, n4733, n4757, n4971, n5030, n5034,
    n5094, n5132, n5191, n5257, n5411, n5435, n5641, n5670, n5693, n5934,
    n6089, n6192, n6273, n6445, n6645, n6689, n6742, n6809, n6822, n6860,
    n7193, n7568, n7676, n7966, n7981, n8100, n8138, n8202, n8303, n8398,
    n9137, n9387, n9571, n9578, n9706, n9756, n9767, n9820, n9938, n10476,
    n10589, n10695, n10789, n10851, n10913, n10949, n11216, n11326, n11707,
    n11755, n11780, n11919, n12005, n12014, n12020, n12076, n12111, n12444,
    n12807;
  wire new_n377, new_n378, new_n379, new_n380, new_n381_1, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397_1,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405_1, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447_1, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503_1, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521_1, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533_1, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615_1, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658_1, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753_1, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783_1, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806_1, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837_1, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844_1, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911_1, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992_1,
    new_n993, new_n994, new_n995, new_n996_1, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020_1, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067_1, new_n1068, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094_1, new_n1095, new_n1096,
    new_n1097_1, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136_1, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198_1,
    new_n1199_1, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269_1, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333_1, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345, new_n1346, new_n1347, new_n1348, new_n1349, new_n1350,
    new_n1351, new_n1352, new_n1353_1, new_n1354, new_n1355, new_n1356,
    new_n1357_1, new_n1358, new_n1359, new_n1360, new_n1361, new_n1362,
    new_n1363, new_n1364, new_n1365, new_n1366, new_n1367, new_n1368,
    new_n1369, new_n1370, new_n1371, new_n1372, new_n1373, new_n1374,
    new_n1375, new_n1376, new_n1377, new_n1378, new_n1379, new_n1380,
    new_n1381, new_n1382, new_n1383, new_n1384, new_n1385, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1398,
    new_n1399, new_n1400, new_n1401, new_n1402, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1416,
    new_n1417, new_n1418, new_n1419, new_n1420, new_n1421, new_n1422,
    new_n1423, new_n1424, new_n1425, new_n1426, new_n1427, new_n1428,
    new_n1429, new_n1430, new_n1431, new_n1432, new_n1433, new_n1434,
    new_n1435, new_n1436, new_n1437, new_n1438, new_n1439, new_n1440,
    new_n1441, new_n1442, new_n1443, new_n1444, new_n1445, new_n1446,
    new_n1447, new_n1448, new_n1449, new_n1450, new_n1451, new_n1452,
    new_n1453, new_n1454, new_n1455, new_n1456, new_n1457, new_n1458,
    new_n1459, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1470,
    new_n1471_1, new_n1472, new_n1473, new_n1474, new_n1475, new_n1476,
    new_n1477, new_n1478_1, new_n1479, new_n1480, new_n1481, new_n1482,
    new_n1483, new_n1484, new_n1485, new_n1486, new_n1487, new_n1488,
    new_n1489, new_n1490, new_n1491, new_n1492, new_n1493, new_n1494,
    new_n1495, new_n1496, new_n1497, new_n1498, new_n1499, new_n1500,
    new_n1501, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507,
    new_n1508, new_n1509, new_n1510_1, new_n1511, new_n1512_1, new_n1513,
    new_n1514, new_n1515, new_n1516, new_n1517, new_n1518, new_n1519,
    new_n1520, new_n1521, new_n1522, new_n1523_1, new_n1524, new_n1525,
    new_n1526, new_n1527, new_n1528, new_n1529, new_n1530, new_n1531,
    new_n1532, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1540, new_n1541, new_n1542, new_n1543,
    new_n1544, new_n1545, new_n1546, new_n1547, new_n1548, new_n1549,
    new_n1550, new_n1551, new_n1552, new_n1553, new_n1554, new_n1555,
    new_n1556, new_n1557, new_n1558, new_n1559, new_n1560, new_n1561,
    new_n1562, new_n1563, new_n1564_1, new_n1565, new_n1566, new_n1567,
    new_n1568, new_n1569, new_n1570, new_n1571, new_n1572, new_n1573,
    new_n1574, new_n1575, new_n1576_1, new_n1577, new_n1578, new_n1579,
    new_n1580, new_n1581, new_n1582, new_n1583, new_n1584, new_n1585,
    new_n1586, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1600, new_n1601, new_n1602, new_n1603,
    new_n1604, new_n1605, new_n1606, new_n1607, new_n1608, new_n1609,
    new_n1610, new_n1611, new_n1612, new_n1613, new_n1614, new_n1615,
    new_n1616, new_n1617, new_n1618, new_n1619, new_n1620, new_n1621,
    new_n1622, new_n1623, new_n1624, new_n1625, new_n1626, new_n1627,
    new_n1628, new_n1629, new_n1630, new_n1631, new_n1632, new_n1633,
    new_n1634, new_n1635, new_n1636, new_n1637, new_n1638, new_n1639,
    new_n1640, new_n1641, new_n1642, new_n1643, new_n1644, new_n1645,
    new_n1646, new_n1647, new_n1648, new_n1649, new_n1650, new_n1651,
    new_n1652, new_n1653, new_n1654, new_n1655, new_n1656, new_n1657,
    new_n1658_1, new_n1659, new_n1660, new_n1661, new_n1662, new_n1663,
    new_n1664, new_n1665, new_n1666, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1678, new_n1679, new_n1680, new_n1681,
    new_n1682, new_n1683, new_n1684, new_n1685, new_n1686, new_n1687,
    new_n1688, new_n1689, new_n1690, new_n1691, new_n1692, new_n1693,
    new_n1694, new_n1695, new_n1696, new_n1697, new_n1698, new_n1699,
    new_n1700, new_n1701, new_n1702, new_n1703, new_n1704, new_n1705,
    new_n1706, new_n1707, new_n1708, new_n1709, new_n1710, new_n1711,
    new_n1712, new_n1713, new_n1714, new_n1715, new_n1716, new_n1717,
    new_n1718, new_n1719, new_n1720, new_n1721, new_n1722, new_n1723,
    new_n1724, new_n1725, new_n1726, new_n1727, new_n1728, new_n1729,
    new_n1730, new_n1731, new_n1732, new_n1733, new_n1734, new_n1735,
    new_n1736, new_n1737, new_n1738, new_n1739, new_n1740, new_n1741,
    new_n1742, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1753,
    new_n1754, new_n1755, new_n1756, new_n1757, new_n1758, new_n1759,
    new_n1760, new_n1761, new_n1762, new_n1763, new_n1764, new_n1765,
    new_n1766, new_n1767, new_n1768, new_n1769, new_n1770, new_n1771,
    new_n1772, new_n1773, new_n1774, new_n1775, new_n1776, new_n1777,
    new_n1778, new_n1779, new_n1780, new_n1781, new_n1782, new_n1783,
    new_n1784, new_n1785, new_n1786, new_n1787, new_n1788, new_n1789,
    new_n1790, new_n1791, new_n1792, new_n1793, new_n1794, new_n1795,
    new_n1796, new_n1797, new_n1798_1, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1806, new_n1807,
    new_n1808, new_n1809, new_n1810, new_n1811, new_n1812, new_n1813,
    new_n1814, new_n1815, new_n1816, new_n1817, new_n1818, new_n1819,
    new_n1820, new_n1821, new_n1822, new_n1823, new_n1824, new_n1825,
    new_n1826, new_n1827, new_n1828, new_n1829, new_n1830, new_n1831,
    new_n1832, new_n1833, new_n1834, new_n1835_1, new_n1836, new_n1837,
    new_n1838, new_n1839, new_n1840, new_n1841, new_n1842, new_n1843,
    new_n1844, new_n1845, new_n1846, new_n1847_1, new_n1848, new_n1849,
    new_n1850, new_n1851, new_n1852, new_n1853, new_n1854, new_n1855,
    new_n1856, new_n1857, new_n1858, new_n1859, new_n1860, new_n1861,
    new_n1862, new_n1863, new_n1864, new_n1865, new_n1866, new_n1867,
    new_n1868, new_n1869, new_n1870, new_n1871, new_n1872, new_n1873,
    new_n1874, new_n1875, new_n1876, new_n1877, new_n1878, new_n1879,
    new_n1880, new_n1881, new_n1882, new_n1883, new_n1884, new_n1885,
    new_n1886, new_n1887, new_n1888, new_n1889, new_n1890, new_n1891,
    new_n1892, new_n1893, new_n1894, new_n1895, new_n1896, new_n1897,
    new_n1898, new_n1899, new_n1900, new_n1901, new_n1902, new_n1903,
    new_n1904, new_n1905, new_n1906_1, new_n1907, new_n1908, new_n1909,
    new_n1910, new_n1911, new_n1912, new_n1913, new_n1914, new_n1915,
    new_n1916, new_n1917, new_n1918, new_n1919, new_n1920, new_n1921,
    new_n1922, new_n1923, new_n1924, new_n1925, new_n1926, new_n1927,
    new_n1928, new_n1929, new_n1930, new_n1931, new_n1932, new_n1933,
    new_n1934, new_n1935, new_n1936, new_n1937, new_n1938, new_n1939,
    new_n1940, new_n1941, new_n1942, new_n1943, new_n1944, new_n1945,
    new_n1946, new_n1947, new_n1948, new_n1949, new_n1950, new_n1951,
    new_n1952, new_n1953, new_n1954, new_n1955, new_n1956, new_n1957,
    new_n1958, new_n1959, new_n1960, new_n1961, new_n1962, new_n1963,
    new_n1964, new_n1965, new_n1966, new_n1967, new_n1968, new_n1969,
    new_n1970, new_n1971, new_n1972, new_n1973, new_n1974, new_n1975,
    new_n1976, new_n1977, new_n1978, new_n1979, new_n1980_1, new_n1981,
    new_n1982, new_n1983, new_n1984, new_n1985, new_n1986, new_n1987,
    new_n1988, new_n1989, new_n1990, new_n1991, new_n1992, new_n1993,
    new_n1994, new_n1995, new_n1996, new_n1997, new_n1998, new_n1999,
    new_n2000, new_n2001, new_n2002, new_n2003, new_n2004, new_n2005,
    new_n2006, new_n2007, new_n2008, new_n2009, new_n2010, new_n2011,
    new_n2012, new_n2013, new_n2014, new_n2015, new_n2016, new_n2017,
    new_n2018, new_n2019, new_n2020, new_n2021, new_n2022, new_n2023,
    new_n2024_1, new_n2025, new_n2026, new_n2027, new_n2028, new_n2029,
    new_n2030, new_n2031, new_n2032, new_n2033, new_n2034, new_n2035,
    new_n2036, new_n2037, new_n2038, new_n2039, new_n2040, new_n2041,
    new_n2042, new_n2043, new_n2044, new_n2045, new_n2046, new_n2047,
    new_n2048, new_n2049, new_n2050, new_n2051, new_n2052, new_n2053,
    new_n2054, new_n2055, new_n2056, new_n2057, new_n2058, new_n2059,
    new_n2060, new_n2061, new_n2062, new_n2063, new_n2064, new_n2065,
    new_n2066, new_n2067, new_n2068, new_n2069, new_n2070, new_n2071,
    new_n2072, new_n2073, new_n2074, new_n2075, new_n2076, new_n2077,
    new_n2078, new_n2079, new_n2080, new_n2081, new_n2082, new_n2083,
    new_n2084, new_n2085, new_n2086, new_n2087_1, new_n2088, new_n2089,
    new_n2090, new_n2091, new_n2092, new_n2093, new_n2094, new_n2095,
    new_n2096_1, new_n2097, new_n2098, new_n2099, new_n2100, new_n2101,
    new_n2102, new_n2103, new_n2104, new_n2105, new_n2106, new_n2107,
    new_n2108, new_n2109, new_n2110, new_n2111, new_n2112, new_n2113,
    new_n2114, new_n2115, new_n2116, new_n2117, new_n2118, new_n2119,
    new_n2120, new_n2121, new_n2122, new_n2123, new_n2124, new_n2125,
    new_n2126, new_n2127, new_n2128, new_n2129, new_n2130, new_n2131_1,
    new_n2132, new_n2133, new_n2134, new_n2135, new_n2136, new_n2137,
    new_n2138, new_n2139, new_n2140, new_n2141, new_n2142, new_n2143,
    new_n2144, new_n2145, new_n2146, new_n2147, new_n2148, new_n2149,
    new_n2150, new_n2151, new_n2152, new_n2153, new_n2154, new_n2155,
    new_n2156, new_n2157, new_n2158, new_n2159, new_n2160, new_n2161,
    new_n2162, new_n2163, new_n2164, new_n2165, new_n2166, new_n2167,
    new_n2168, new_n2169, new_n2170, new_n2171, new_n2172, new_n2173,
    new_n2174, new_n2175, new_n2176, new_n2177, new_n2178, new_n2179,
    new_n2180, new_n2181, new_n2182, new_n2183, new_n2184, new_n2185,
    new_n2186, new_n2187, new_n2188, new_n2189, new_n2190, new_n2191,
    new_n2192, new_n2193, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2213, new_n2214, new_n2215,
    new_n2216, new_n2217, new_n2218, new_n2219, new_n2220, new_n2221,
    new_n2222, new_n2223, new_n2224, new_n2225, new_n2226_1, new_n2227,
    new_n2228, new_n2229, new_n2230, new_n2231, new_n2232, new_n2233,
    new_n2234, new_n2235, new_n2236, new_n2237, new_n2238, new_n2239,
    new_n2240, new_n2241, new_n2242, new_n2243, new_n2244, new_n2245,
    new_n2246, new_n2247, new_n2248, new_n2249, new_n2250, new_n2251,
    new_n2252, new_n2253_1, new_n2254, new_n2255, new_n2256, new_n2257,
    new_n2258, new_n2259, new_n2260, new_n2261, new_n2262, new_n2263,
    new_n2264, new_n2265, new_n2266, new_n2267, new_n2268, new_n2269,
    new_n2270, new_n2271, new_n2272, new_n2273, new_n2274, new_n2275,
    new_n2276, new_n2277, new_n2278_1, new_n2279, new_n2280, new_n2281,
    new_n2282, new_n2283, new_n2284, new_n2285, new_n2286, new_n2287,
    new_n2288, new_n2289, new_n2290, new_n2291, new_n2292, new_n2293,
    new_n2294, new_n2295, new_n2296, new_n2297, new_n2298, new_n2299,
    new_n2300, new_n2301_1, new_n2302, new_n2303, new_n2304, new_n2305,
    new_n2306, new_n2307, new_n2308, new_n2309, new_n2310, new_n2311,
    new_n2312, new_n2313, new_n2314, new_n2315, new_n2316_1, new_n2317,
    new_n2318, new_n2319, new_n2320, new_n2321, new_n2322, new_n2323,
    new_n2324, new_n2325, new_n2326, new_n2327, new_n2328, new_n2329,
    new_n2330, new_n2331, new_n2332, new_n2333, new_n2334, new_n2335,
    new_n2336, new_n2337, new_n2338, new_n2339, new_n2340, new_n2341,
    new_n2342, new_n2343, new_n2344, new_n2345, new_n2346, new_n2347_1,
    new_n2348, new_n2349, new_n2350, new_n2351, new_n2352, new_n2353,
    new_n2354, new_n2355, new_n2356, new_n2357, new_n2358, new_n2359,
    new_n2360, new_n2361, new_n2362, new_n2363, new_n2364, new_n2365,
    new_n2366, new_n2367, new_n2368, new_n2369, new_n2370, new_n2371,
    new_n2372, new_n2373, new_n2374, new_n2375, new_n2376, new_n2377,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383_1, new_n2384,
    new_n2385, new_n2386, new_n2387, new_n2388, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393_1, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416, new_n2417, new_n2418, new_n2419, new_n2420,
    new_n2421, new_n2422, new_n2423, new_n2424, new_n2425_1, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431_1, new_n2432,
    new_n2433_1, new_n2434_1, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440, new_n2441, new_n2442, new_n2443, new_n2444,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464_1, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498_1,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507_1, new_n2508_1, new_n2509_1, new_n2510,
    new_n2511, new_n2512_1, new_n2513, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522_1,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530_1, new_n2531, new_n2532, new_n2533, new_n2534,
    new_n2535, new_n2536, new_n2537, new_n2538, new_n2539, new_n2540,
    new_n2541, new_n2542, new_n2543, new_n2544, new_n2545, new_n2546,
    new_n2547, new_n2548, new_n2549, new_n2550, new_n2551_1, new_n2552,
    new_n2553, new_n2554, new_n2555, new_n2556, new_n2557, new_n2558_1,
    new_n2559, new_n2560, new_n2561, new_n2562, new_n2563, new_n2564_1,
    new_n2565, new_n2566, new_n2567, new_n2568, new_n2569, new_n2570,
    new_n2571, new_n2572, new_n2573, new_n2574, new_n2575, new_n2576,
    new_n2577_1, new_n2578, new_n2579, new_n2580, new_n2581_1, new_n2582,
    new_n2583, new_n2584, new_n2585_1, new_n2586, new_n2587, new_n2588,
    new_n2589, new_n2590, new_n2591, new_n2592, new_n2593, new_n2594,
    new_n2595, new_n2596, new_n2597, new_n2598, new_n2599, new_n2600,
    new_n2601, new_n2602, new_n2603, new_n2604, new_n2605, new_n2606,
    new_n2607, new_n2608, new_n2609, new_n2610, new_n2611, new_n2612,
    new_n2613, new_n2614, new_n2615, new_n2616, new_n2617, new_n2618,
    new_n2619, new_n2620, new_n2621, new_n2622, new_n2623, new_n2624_1,
    new_n2625, new_n2626, new_n2627, new_n2628, new_n2629, new_n2630,
    new_n2631, new_n2632, new_n2633, new_n2634, new_n2635, new_n2636,
    new_n2637, new_n2638, new_n2639, new_n2640, new_n2641, new_n2642,
    new_n2643, new_n2644, new_n2645, new_n2646, new_n2647, new_n2648,
    new_n2649, new_n2650, new_n2651, new_n2652, new_n2653, new_n2654,
    new_n2655, new_n2656, new_n2657, new_n2658, new_n2659, new_n2660,
    new_n2661, new_n2662, new_n2663, new_n2664, new_n2665, new_n2666,
    new_n2667, new_n2668, new_n2669, new_n2670, new_n2671, new_n2672,
    new_n2673, new_n2674, new_n2675, new_n2676, new_n2677, new_n2678,
    new_n2679_1, new_n2680, new_n2681, new_n2682, new_n2683, new_n2684,
    new_n2685, new_n2686, new_n2687, new_n2688, new_n2689, new_n2690,
    new_n2691, new_n2692, new_n2693, new_n2694, new_n2695, new_n2696,
    new_n2697, new_n2698, new_n2699, new_n2700, new_n2701, new_n2702,
    new_n2703, new_n2704, new_n2705, new_n2706, new_n2707, new_n2708_1,
    new_n2709, new_n2710, new_n2711, new_n2712, new_n2713, new_n2714,
    new_n2715, new_n2716, new_n2717, new_n2718, new_n2719, new_n2720,
    new_n2721, new_n2722, new_n2723, new_n2724, new_n2725, new_n2726,
    new_n2727, new_n2728, new_n2729, new_n2730, new_n2731, new_n2732,
    new_n2733, new_n2734, new_n2735, new_n2736, new_n2737, new_n2738,
    new_n2739, new_n2740, new_n2741, new_n2742, new_n2743, new_n2744,
    new_n2745, new_n2746, new_n2747, new_n2748, new_n2749_1, new_n2750,
    new_n2751, new_n2752, new_n2753, new_n2754, new_n2755, new_n2756,
    new_n2757, new_n2758, new_n2759, new_n2760, new_n2761, new_n2762,
    new_n2763, new_n2764, new_n2765, new_n2766, new_n2767, new_n2768,
    new_n2769, new_n2770, new_n2771, new_n2772, new_n2773, new_n2774,
    new_n2775, new_n2776, new_n2777, new_n2778, new_n2779, new_n2780,
    new_n2781, new_n2782, new_n2783, new_n2784, new_n2785, new_n2786,
    new_n2787, new_n2788, new_n2789, new_n2790, new_n2791, new_n2792,
    new_n2793, new_n2794, new_n2795, new_n2796, new_n2797, new_n2798,
    new_n2799, new_n2800, new_n2801, new_n2802_1, new_n2803, new_n2804,
    new_n2805, new_n2806, new_n2807, new_n2808, new_n2809, new_n2810,
    new_n2811, new_n2812, new_n2813, new_n2814, new_n2815, new_n2816,
    new_n2817, new_n2818_1, new_n2819, new_n2820, new_n2821, new_n2822,
    new_n2823, new_n2824, new_n2825, new_n2826, new_n2827, new_n2828,
    new_n2829, new_n2830, new_n2831, new_n2832, new_n2833, new_n2834,
    new_n2835, new_n2836, new_n2837, new_n2838, new_n2839, new_n2840,
    new_n2841, new_n2842, new_n2843, new_n2844, new_n2845, new_n2846,
    new_n2847, new_n2848, new_n2849, new_n2850, new_n2851, new_n2852,
    new_n2853, new_n2854, new_n2855, new_n2856, new_n2857, new_n2858,
    new_n2859, new_n2860, new_n2861, new_n2862, new_n2863, new_n2864,
    new_n2865, new_n2866, new_n2867, new_n2868, new_n2869, new_n2870,
    new_n2871, new_n2872, new_n2873, new_n2874, new_n2875, new_n2876,
    new_n2877, new_n2878, new_n2879_1, new_n2880, new_n2881, new_n2882,
    new_n2883, new_n2884, new_n2885, new_n2886, new_n2887, new_n2888,
    new_n2889, new_n2890, new_n2891, new_n2892, new_n2893, new_n2894,
    new_n2895, new_n2896, new_n2897, new_n2898, new_n2899, new_n2900,
    new_n2901, new_n2902_1, new_n2903, new_n2904, new_n2905, new_n2906,
    new_n2907, new_n2908, new_n2909, new_n2910, new_n2911, new_n2912,
    new_n2913, new_n2914, new_n2915, new_n2916, new_n2917, new_n2918,
    new_n2919, new_n2920, new_n2921, new_n2922, new_n2923, new_n2924,
    new_n2925, new_n2926, new_n2927, new_n2928, new_n2929, new_n2930,
    new_n2931, new_n2932, new_n2933, new_n2934, new_n2935, new_n2936,
    new_n2937, new_n2938, new_n2939, new_n2940, new_n2941, new_n2942,
    new_n2943, new_n2944, new_n2945, new_n2946, new_n2947, new_n2948,
    new_n2949, new_n2950, new_n2951, new_n2952, new_n2953, new_n2954,
    new_n2955, new_n2956, new_n2957, new_n2958, new_n2959, new_n2960,
    new_n2961, new_n2962, new_n2963, new_n2964, new_n2965, new_n2966,
    new_n2967, new_n2968, new_n2969, new_n2970, new_n2971, new_n2972,
    new_n2973, new_n2974, new_n2975, new_n2976, new_n2977, new_n2978,
    new_n2979, new_n2980, new_n2981, new_n2982, new_n2983, new_n2984,
    new_n2985, new_n2986, new_n2987, new_n2988, new_n2989, new_n2990,
    new_n2991, new_n2992, new_n2993, new_n2994, new_n2995, new_n2996,
    new_n2997, new_n2998, new_n2999, new_n3000, new_n3001, new_n3002,
    new_n3003, new_n3004, new_n3005, new_n3006, new_n3007, new_n3008,
    new_n3009, new_n3010, new_n3011, new_n3012, new_n3013, new_n3014,
    new_n3015, new_n3016, new_n3017, new_n3018, new_n3019, new_n3020,
    new_n3021, new_n3022_1, new_n3023, new_n3024, new_n3025, new_n3026,
    new_n3027, new_n3028, new_n3029, new_n3030, new_n3031, new_n3032,
    new_n3033, new_n3034, new_n3035, new_n3036, new_n3037, new_n3038,
    new_n3039, new_n3040, new_n3041, new_n3042, new_n3043, new_n3044,
    new_n3045, new_n3046, new_n3047, new_n3048, new_n3049, new_n3050,
    new_n3051, new_n3052, new_n3053, new_n3054, new_n3055, new_n3056,
    new_n3057, new_n3058, new_n3059, new_n3060, new_n3061, new_n3062,
    new_n3063, new_n3064, new_n3065, new_n3066, new_n3067, new_n3068,
    new_n3069, new_n3070, new_n3071_1, new_n3072, new_n3073, new_n3074,
    new_n3075, new_n3076, new_n3077, new_n3078, new_n3079, new_n3080,
    new_n3081, new_n3082, new_n3083, new_n3084, new_n3085, new_n3086,
    new_n3087, new_n3088, new_n3089, new_n3090, new_n3091, new_n3092,
    new_n3093, new_n3094, new_n3095, new_n3096, new_n3097, new_n3098,
    new_n3099, new_n3100, new_n3101, new_n3102, new_n3103, new_n3104,
    new_n3105, new_n3106, new_n3107, new_n3108, new_n3109, new_n3110,
    new_n3111, new_n3112, new_n3113, new_n3114, new_n3115, new_n3116,
    new_n3117, new_n3118, new_n3119, new_n3120, new_n3121, new_n3122,
    new_n3123, new_n3124_1, new_n3125, new_n3126, new_n3127, new_n3128,
    new_n3129, new_n3130, new_n3131, new_n3132, new_n3133, new_n3134,
    new_n3135, new_n3136, new_n3137, new_n3138, new_n3139, new_n3140,
    new_n3141, new_n3142, new_n3143, new_n3144, new_n3145, new_n3146_1,
    new_n3147, new_n3148, new_n3149, new_n3150, new_n3151, new_n3152,
    new_n3153, new_n3154, new_n3155, new_n3156, new_n3157, new_n3158,
    new_n3159, new_n3160, new_n3161, new_n3162, new_n3163, new_n3164,
    new_n3165, new_n3166, new_n3167, new_n3168, new_n3169, new_n3170,
    new_n3171, new_n3172_1, new_n3173, new_n3174, new_n3175, new_n3176,
    new_n3177, new_n3178, new_n3179, new_n3180, new_n3181, new_n3182,
    new_n3183, new_n3184, new_n3185, new_n3186, new_n3187, new_n3188,
    new_n3189, new_n3190, new_n3191, new_n3192, new_n3193, new_n3194,
    new_n3195, new_n3196, new_n3197, new_n3198, new_n3199, new_n3200,
    new_n3201, new_n3202, new_n3203, new_n3204, new_n3205, new_n3206,
    new_n3207, new_n3208, new_n3209, new_n3210, new_n3211, new_n3212,
    new_n3213, new_n3214_1, new_n3215, new_n3216, new_n3217, new_n3218,
    new_n3219, new_n3220, new_n3221, new_n3222, new_n3223, new_n3224,
    new_n3225, new_n3226, new_n3227, new_n3228, new_n3229, new_n3230_1,
    new_n3231, new_n3232, new_n3233, new_n3234, new_n3235, new_n3236,
    new_n3237, new_n3238, new_n3239, new_n3240, new_n3241, new_n3242,
    new_n3243, new_n3244, new_n3245, new_n3246, new_n3247, new_n3248,
    new_n3249, new_n3250, new_n3251, new_n3252, new_n3253, new_n3254,
    new_n3255, new_n3256, new_n3257, new_n3258, new_n3259, new_n3260,
    new_n3261, new_n3262, new_n3263, new_n3264, new_n3265, new_n3266,
    new_n3267, new_n3268, new_n3269, new_n3270, new_n3271, new_n3272_1,
    new_n3273, new_n3274, new_n3275, new_n3276, new_n3277, new_n3278,
    new_n3279, new_n3280, new_n3282, new_n3283, new_n3284, new_n3285,
    new_n3286, new_n3287_1, new_n3288, new_n3289, new_n3290, new_n3291,
    new_n3292, new_n3293, new_n3294, new_n3295, new_n3296, new_n3297,
    new_n3298, new_n3299, new_n3300, new_n3301, new_n3302, new_n3303,
    new_n3304, new_n3305, new_n3306, new_n3307, new_n3308, new_n3309,
    new_n3310, new_n3311, new_n3312, new_n3313, new_n3314, new_n3315,
    new_n3316, new_n3317, new_n3318, new_n3319, new_n3320, new_n3321,
    new_n3322, new_n3323, new_n3324, new_n3325, new_n3326, new_n3327,
    new_n3328, new_n3329, new_n3330, new_n3331, new_n3332, new_n3333,
    new_n3334, new_n3335, new_n3336, new_n3337, new_n3338, new_n3339_1,
    new_n3340, new_n3341, new_n3342_1, new_n3343, new_n3344, new_n3345,
    new_n3346, new_n3347, new_n3348, new_n3349, new_n3350, new_n3351,
    new_n3352, new_n3353, new_n3354, new_n3355, new_n3356, new_n3357,
    new_n3358, new_n3359, new_n3360, new_n3361, new_n3362, new_n3363,
    new_n3364, new_n3365, new_n3366, new_n3367, new_n3368, new_n3369,
    new_n3370, new_n3371, new_n3372, new_n3373, new_n3374, new_n3375,
    new_n3376, new_n3377, new_n3378, new_n3379, new_n3380, new_n3381,
    new_n3382, new_n3383, new_n3384, new_n3385, new_n3386, new_n3387,
    new_n3388, new_n3389, new_n3390, new_n3391, new_n3392, new_n3393,
    new_n3394, new_n3395, new_n3396, new_n3397, new_n3398, new_n3399,
    new_n3400, new_n3401, new_n3402, new_n3403, new_n3404, new_n3405,
    new_n3406, new_n3407, new_n3408, new_n3409, new_n3410, new_n3411,
    new_n3412, new_n3413, new_n3414, new_n3415, new_n3416, new_n3417,
    new_n3418, new_n3419, new_n3420, new_n3421, new_n3422, new_n3423,
    new_n3424, new_n3425, new_n3426, new_n3427, new_n3428, new_n3429,
    new_n3430, new_n3431, new_n3432, new_n3433, new_n3434, new_n3435,
    new_n3436, new_n3437, new_n3438, new_n3439, new_n3440, new_n3441,
    new_n3442, new_n3443, new_n3444, new_n3445, new_n3446, new_n3447,
    new_n3448, new_n3449, new_n3450, new_n3451, new_n3452, new_n3453,
    new_n3454, new_n3455, new_n3456_1, new_n3457, new_n3458, new_n3459,
    new_n3460, new_n3461, new_n3462, new_n3463, new_n3464, new_n3465,
    new_n3466, new_n3467, new_n3468, new_n3469, new_n3470, new_n3471,
    new_n3472, new_n3473, new_n3474, new_n3475, new_n3476, new_n3477,
    new_n3478, new_n3479, new_n3480, new_n3481, new_n3482, new_n3483,
    new_n3484, new_n3485, new_n3486, new_n3487, new_n3488, new_n3489,
    new_n3490, new_n3491, new_n3492, new_n3493, new_n3494, new_n3495,
    new_n3496, new_n3497, new_n3498, new_n3499, new_n3500, new_n3501,
    new_n3502, new_n3503, new_n3504, new_n3505, new_n3506, new_n3507,
    new_n3508, new_n3509, new_n3510, new_n3511, new_n3512, new_n3513,
    new_n3514, new_n3515, new_n3516, new_n3517, new_n3518, new_n3519,
    new_n3520, new_n3521, new_n3522, new_n3523, new_n3524, new_n3525,
    new_n3526, new_n3527, new_n3528, new_n3529, new_n3530, new_n3531,
    new_n3532, new_n3533, new_n3534, new_n3535, new_n3536, new_n3537,
    new_n3538, new_n3539, new_n3540, new_n3541, new_n3542, new_n3543,
    new_n3544, new_n3545, new_n3546, new_n3547, new_n3548, new_n3549,
    new_n3550, new_n3551, new_n3552, new_n3553, new_n3554, new_n3555,
    new_n3556, new_n3557, new_n3558, new_n3559, new_n3560, new_n3561,
    new_n3562, new_n3563, new_n3564, new_n3565, new_n3566, new_n3567,
    new_n3568, new_n3569, new_n3570, new_n3571, new_n3572, new_n3573,
    new_n3574, new_n3575, new_n3576, new_n3577, new_n3578, new_n3579,
    new_n3580, new_n3581, new_n3582, new_n3583, new_n3584, new_n3585,
    new_n3586, new_n3587, new_n3588, new_n3589, new_n3590, new_n3591,
    new_n3592, new_n3593, new_n3594, new_n3595, new_n3596, new_n3597,
    new_n3598, new_n3599, new_n3600, new_n3601, new_n3602_1, new_n3603,
    new_n3604, new_n3605, new_n3606, new_n3607, new_n3608, new_n3609,
    new_n3610, new_n3611, new_n3612, new_n3613, new_n3614, new_n3615,
    new_n3616_1, new_n3617, new_n3618, new_n3619, new_n3620, new_n3621,
    new_n3622, new_n3623, new_n3624, new_n3625, new_n3626, new_n3627_1,
    new_n3628, new_n3629, new_n3630, new_n3631, new_n3632, new_n3633,
    new_n3634, new_n3635, new_n3636, new_n3637, new_n3638, new_n3639,
    new_n3640, new_n3641, new_n3642, new_n3643, new_n3644, new_n3645,
    new_n3646, new_n3647, new_n3648, new_n3649, new_n3650, new_n3651,
    new_n3652, new_n3653, new_n3654_1, new_n3655, new_n3656, new_n3657,
    new_n3658, new_n3659, new_n3660, new_n3661_1, new_n3662, new_n3663,
    new_n3664, new_n3665, new_n3666, new_n3667, new_n3668, new_n3669,
    new_n3670, new_n3671, new_n3672, new_n3673, new_n3674, new_n3675,
    new_n3676, new_n3677_1, new_n3678, new_n3679, new_n3680, new_n3681,
    new_n3682, new_n3683, new_n3684, new_n3685, new_n3686, new_n3687,
    new_n3688, new_n3689, new_n3690, new_n3691, new_n3692, new_n3693,
    new_n3694, new_n3695, new_n3696, new_n3697, new_n3698, new_n3699,
    new_n3700, new_n3701, new_n3702, new_n3703, new_n3704, new_n3705,
    new_n3706, new_n3707, new_n3708, new_n3709, new_n3710, new_n3711,
    new_n3712, new_n3713, new_n3714, new_n3715, new_n3716, new_n3717,
    new_n3718, new_n3719_1, new_n3720, new_n3721, new_n3722, new_n3723,
    new_n3724, new_n3725, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754_1, new_n3755, new_n3756, new_n3757, new_n3758, new_n3759,
    new_n3760, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781, new_n3782, new_n3783,
    new_n3784, new_n3785, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794, new_n3795,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849_1,
    new_n3850, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865_1, new_n3866, new_n3867,
    new_n3868, new_n3869, new_n3870, new_n3871, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925, new_n3926, new_n3927,
    new_n3928, new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933,
    new_n3934, new_n3935, new_n3936, new_n3937, new_n3938, new_n3939,
    new_n3940, new_n3941, new_n3942, new_n3943, new_n3944, new_n3945,
    new_n3946, new_n3947, new_n3948, new_n3949, new_n3950, new_n3951,
    new_n3952, new_n3953, new_n3954, new_n3955, new_n3956, new_n3957,
    new_n3958, new_n3959, new_n3960, new_n3961, new_n3962, new_n3963,
    new_n3964, new_n3965, new_n3966, new_n3967, new_n3968, new_n3969,
    new_n3970, new_n3971, new_n3972, new_n3973, new_n3974, new_n3975,
    new_n3976, new_n3977, new_n3978, new_n3979, new_n3980, new_n3981,
    new_n3982, new_n3983, new_n3984, new_n3985, new_n3986_1, new_n3987,
    new_n3988, new_n3989, new_n3990, new_n3991, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005_1, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010, new_n4011, new_n4012,
    new_n4013, new_n4014, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085, new_n4086_1, new_n4087, new_n4088_1, new_n4089, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094_1, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100, new_n4101, new_n4102,
    new_n4103, new_n4104, new_n4105, new_n4106, new_n4107, new_n4108,
    new_n4109, new_n4110, new_n4111, new_n4112, new_n4113, new_n4114,
    new_n4115, new_n4116, new_n4117, new_n4118, new_n4119, new_n4120,
    new_n4121, new_n4122, new_n4123, new_n4124, new_n4125, new_n4126,
    new_n4127, new_n4128, new_n4129, new_n4130, new_n4131, new_n4132,
    new_n4133, new_n4134, new_n4135, new_n4136, new_n4137, new_n4138,
    new_n4139, new_n4140, new_n4141_1, new_n4142, new_n4143, new_n4144,
    new_n4145, new_n4146, new_n4147, new_n4148, new_n4149, new_n4150,
    new_n4151, new_n4152, new_n4153, new_n4154, new_n4155_1, new_n4156,
    new_n4157, new_n4158, new_n4159_1, new_n4160, new_n4161, new_n4162,
    new_n4163, new_n4164, new_n4165, new_n4166, new_n4167, new_n4168,
    new_n4169, new_n4170, new_n4171, new_n4172, new_n4173, new_n4174,
    new_n4175, new_n4176, new_n4177, new_n4178, new_n4179, new_n4180,
    new_n4181, new_n4182, new_n4183, new_n4184, new_n4185, new_n4186,
    new_n4187_1, new_n4188, new_n4189_1, new_n4190_1, new_n4191, new_n4192,
    new_n4193, new_n4194, new_n4195, new_n4196, new_n4197, new_n4198,
    new_n4199, new_n4200, new_n4201, new_n4202, new_n4203_1, new_n4204,
    new_n4205, new_n4206, new_n4207, new_n4208, new_n4209, new_n4210,
    new_n4211, new_n4212, new_n4213, new_n4214, new_n4215, new_n4216,
    new_n4218, new_n4219, new_n4220, new_n4221, new_n4222, new_n4223,
    new_n4224, new_n4225, new_n4226_1, new_n4227, new_n4228, new_n4229,
    new_n4230_1, new_n4231, new_n4232, new_n4233, new_n4234, new_n4235,
    new_n4236, new_n4237, new_n4238, new_n4239, new_n4240, new_n4241,
    new_n4242, new_n4243, new_n4244, new_n4245, new_n4246, new_n4247,
    new_n4248, new_n4249, new_n4250, new_n4251, new_n4252, new_n4253,
    new_n4254, new_n4255, new_n4256, new_n4257, new_n4258, new_n4259,
    new_n4260, new_n4261, new_n4262, new_n4263, new_n4264, new_n4265,
    new_n4266, new_n4267, new_n4268, new_n4269, new_n4270, new_n4271,
    new_n4272, new_n4273, new_n4274, new_n4275, new_n4276, new_n4277,
    new_n4278, new_n4279, new_n4280, new_n4281, new_n4282, new_n4283,
    new_n4284, new_n4285, new_n4286, new_n4287, new_n4288, new_n4289,
    new_n4290, new_n4291, new_n4292, new_n4293, new_n4294, new_n4295,
    new_n4296, new_n4297, new_n4298, new_n4299, new_n4300_1, new_n4301,
    new_n4302, new_n4303, new_n4304, new_n4305, new_n4306, new_n4307,
    new_n4308, new_n4309, new_n4310, new_n4311, new_n4312_1, new_n4313,
    new_n4314, new_n4315, new_n4316, new_n4317, new_n4318, new_n4319,
    new_n4320, new_n4321, new_n4322, new_n4323, new_n4324, new_n4325,
    new_n4326_1, new_n4327, new_n4328, new_n4329, new_n4330, new_n4331,
    new_n4332, new_n4333_1, new_n4334, new_n4335, new_n4336, new_n4337,
    new_n4338, new_n4339, new_n4340, new_n4341, new_n4342, new_n4343,
    new_n4344, new_n4345, new_n4346, new_n4347, new_n4348, new_n4349,
    new_n4350, new_n4351, new_n4352, new_n4353, new_n4354, new_n4355,
    new_n4356, new_n4357, new_n4358, new_n4359, new_n4360, new_n4361,
    new_n4362, new_n4363, new_n4364, new_n4365, new_n4366, new_n4367,
    new_n4368, new_n4369, new_n4370_1, new_n4371, new_n4372, new_n4373,
    new_n4374, new_n4375, new_n4376, new_n4377, new_n4378_1, new_n4379,
    new_n4380, new_n4381, new_n4382, new_n4383, new_n4384, new_n4385,
    new_n4386, new_n4387, new_n4388, new_n4389, new_n4390, new_n4391,
    new_n4392, new_n4393, new_n4394, new_n4395, new_n4396, new_n4397_1,
    new_n4398, new_n4399, new_n4400, new_n4401, new_n4402, new_n4403,
    new_n4404, new_n4405, new_n4406, new_n4407, new_n4408, new_n4409,
    new_n4410, new_n4411, new_n4412, new_n4413, new_n4414, new_n4415,
    new_n4416, new_n4417, new_n4418, new_n4419, new_n4420, new_n4421,
    new_n4422, new_n4423, new_n4424, new_n4425, new_n4426, new_n4427,
    new_n4428, new_n4429, new_n4430, new_n4431, new_n4432, new_n4433,
    new_n4434, new_n4435, new_n4436_1, new_n4437, new_n4438, new_n4439,
    new_n4440, new_n4441, new_n4442, new_n4443, new_n4444, new_n4445,
    new_n4446, new_n4447, new_n4448, new_n4449, new_n4450, new_n4451,
    new_n4452, new_n4453, new_n4454, new_n4455, new_n4456, new_n4457,
    new_n4458, new_n4459, new_n4460, new_n4461, new_n4462, new_n4463,
    new_n4464, new_n4465, new_n4466, new_n4467, new_n4468, new_n4469,
    new_n4470, new_n4471, new_n4472, new_n4473, new_n4474, new_n4475,
    new_n4476, new_n4477, new_n4478, new_n4479, new_n4480, new_n4481,
    new_n4482, new_n4483, new_n4484, new_n4485, new_n4486, new_n4487,
    new_n4488, new_n4489, new_n4490, new_n4491, new_n4492, new_n4493,
    new_n4494, new_n4495, new_n4496, new_n4497, new_n4498, new_n4499_1,
    new_n4500, new_n4501, new_n4502, new_n4503, new_n4504, new_n4505,
    new_n4506, new_n4507, new_n4508, new_n4509, new_n4510, new_n4511,
    new_n4512, new_n4513, new_n4514, new_n4515, new_n4516_1, new_n4517,
    new_n4518, new_n4519, new_n4520, new_n4521, new_n4522, new_n4523,
    new_n4524, new_n4525, new_n4526, new_n4527, new_n4528, new_n4529,
    new_n4530, new_n4531, new_n4532, new_n4533, new_n4534, new_n4535,
    new_n4536, new_n4537, new_n4538, new_n4539, new_n4540, new_n4541,
    new_n4542, new_n4543, new_n4544, new_n4545, new_n4546, new_n4547,
    new_n4548, new_n4549, new_n4550, new_n4551, new_n4552, new_n4553_1,
    new_n4554, new_n4555, new_n4556, new_n4557, new_n4558, new_n4559,
    new_n4560, new_n4561, new_n4562, new_n4563, new_n4564, new_n4566,
    new_n4567, new_n4568, new_n4569, new_n4570, new_n4571, new_n4572,
    new_n4573, new_n4575, new_n4577, new_n4579, new_n4580, new_n4581,
    new_n4582, new_n4583, new_n4584, new_n4585, new_n4586, new_n4587,
    new_n4588, new_n4589, new_n4590, new_n4591, new_n4592, new_n4593,
    new_n4594, new_n4595, new_n4596, new_n4597, new_n4598, new_n4599,
    new_n4600, new_n4601, new_n4602, new_n4603, new_n4604, new_n4605,
    new_n4606, new_n4607, new_n4608, new_n4609, new_n4610, new_n4611,
    new_n4612, new_n4613, new_n4614, new_n4615, new_n4616, new_n4617,
    new_n4618, new_n4619, new_n4620, new_n4621, new_n4622, new_n4623,
    new_n4624, new_n4625, new_n4626, new_n4627, new_n4628, new_n4629,
    new_n4630, new_n4631, new_n4632, new_n4633, new_n4634_1, new_n4635,
    new_n4636, new_n4637, new_n4638, new_n4639, new_n4640, new_n4641,
    new_n4642, new_n4643, new_n4644, new_n4645, new_n4646, new_n4647,
    new_n4648, new_n4649, new_n4650, new_n4651, new_n4652, new_n4653,
    new_n4654, new_n4655, new_n4656, new_n4657, new_n4658, new_n4659,
    new_n4660, new_n4661, new_n4662, new_n4663, new_n4664, new_n4665,
    new_n4666, new_n4667, new_n4668, new_n4669, new_n4670, new_n4671,
    new_n4672, new_n4673, new_n4674, new_n4675, new_n4676, new_n4677,
    new_n4678, new_n4679, new_n4680, new_n4681, new_n4682, new_n4683,
    new_n4684, new_n4685, new_n4686_1, new_n4687, new_n4688, new_n4689_1,
    new_n4690, new_n4691, new_n4692, new_n4693, new_n4694, new_n4695,
    new_n4696, new_n4697, new_n4698, new_n4699, new_n4700, new_n4701,
    new_n4702, new_n4703, new_n4704, new_n4705, new_n4706, new_n4707,
    new_n4708, new_n4709, new_n4710, new_n4711, new_n4712, new_n4713,
    new_n4714, new_n4715, new_n4716, new_n4717, new_n4718, new_n4719,
    new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724, new_n4725,
    new_n4726, new_n4727, new_n4728, new_n4729, new_n4730, new_n4731,
    new_n4732, new_n4733_1, new_n4734, new_n4735, new_n4736, new_n4737,
    new_n4738, new_n4739, new_n4740, new_n4741, new_n4742, new_n4743,
    new_n4744, new_n4745, new_n4746, new_n4747, new_n4748, new_n4749,
    new_n4750, new_n4751, new_n4752, new_n4753, new_n4754, new_n4755,
    new_n4756, new_n4757_1, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766, new_n4767,
    new_n4768, new_n4769, new_n4770, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804, new_n4805_1, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810, new_n4811, new_n4812, new_n4813, new_n4814, new_n4815,
    new_n4816, new_n4817_1, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826_1, new_n4827,
    new_n4828_1, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903_1, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921_1, new_n4922, new_n4923,
    new_n4924, new_n4925, new_n4926, new_n4927, new_n4928_1, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938_1, new_n4939, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964, new_n4965,
    new_n4966, new_n4967, new_n4968, new_n4969, new_n4970_1, new_n4971_1,
    new_n4972, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020, new_n5021, new_n5022, new_n5023, new_n5024, new_n5025,
    new_n5026, new_n5027, new_n5028, new_n5029, new_n5030_1, new_n5031,
    new_n5032, new_n5033, new_n5034_1, new_n5035, new_n5036, new_n5037,
    new_n5038, new_n5039, new_n5040, new_n5041, new_n5042, new_n5043,
    new_n5044, new_n5045, new_n5046, new_n5047, new_n5048, new_n5049,
    new_n5050, new_n5051, new_n5052, new_n5053, new_n5054, new_n5055,
    new_n5056, new_n5057, new_n5058, new_n5059, new_n5060, new_n5061,
    new_n5062, new_n5063, new_n5064, new_n5065, new_n5066, new_n5067,
    new_n5068, new_n5069_1, new_n5070, new_n5071, new_n5072, new_n5073,
    new_n5074, new_n5075, new_n5076, new_n5077, new_n5078, new_n5079,
    new_n5080, new_n5081, new_n5082, new_n5083, new_n5084, new_n5085,
    new_n5086, new_n5087, new_n5088, new_n5089, new_n5090, new_n5091,
    new_n5092, new_n5093, new_n5094_1, new_n5095, new_n5096, new_n5097,
    new_n5098, new_n5099, new_n5100, new_n5101, new_n5102, new_n5103,
    new_n5104, new_n5105_1, new_n5106, new_n5107, new_n5108, new_n5109,
    new_n5110, new_n5111, new_n5112, new_n5113, new_n5114, new_n5115,
    new_n5116, new_n5117, new_n5118, new_n5119, new_n5120, new_n5121,
    new_n5122, new_n5123, new_n5124, new_n5125, new_n5126, new_n5127,
    new_n5128, new_n5129, new_n5130, new_n5131, new_n5132_1, new_n5133,
    new_n5134, new_n5135, new_n5136, new_n5137, new_n5138, new_n5139,
    new_n5140, new_n5141, new_n5142, new_n5143, new_n5144, new_n5145,
    new_n5146, new_n5147, new_n5148, new_n5149, new_n5150, new_n5151,
    new_n5152, new_n5153_1, new_n5154, new_n5155, new_n5156, new_n5157,
    new_n5158, new_n5159, new_n5160, new_n5161, new_n5162, new_n5163,
    new_n5164, new_n5165, new_n5166, new_n5167, new_n5168, new_n5169,
    new_n5170, new_n5171, new_n5172, new_n5173, new_n5174, new_n5175,
    new_n5176, new_n5177, new_n5178, new_n5179, new_n5180, new_n5181,
    new_n5182, new_n5183, new_n5184, new_n5185, new_n5186, new_n5187,
    new_n5188, new_n5189, new_n5190, new_n5191_1, new_n5192, new_n5193,
    new_n5194, new_n5195, new_n5196, new_n5197, new_n5198_1, new_n5199,
    new_n5200, new_n5201, new_n5202, new_n5203, new_n5204, new_n5205,
    new_n5206, new_n5207, new_n5208, new_n5209, new_n5210, new_n5211,
    new_n5212_1, new_n5213, new_n5214, new_n5215, new_n5216, new_n5217,
    new_n5218, new_n5219, new_n5220, new_n5221, new_n5222, new_n5223,
    new_n5224, new_n5225, new_n5226, new_n5227, new_n5228, new_n5229,
    new_n5230, new_n5231, new_n5232, new_n5233, new_n5234, new_n5235,
    new_n5236, new_n5237, new_n5238, new_n5239, new_n5240_1, new_n5241,
    new_n5242, new_n5243, new_n5244, new_n5245, new_n5246, new_n5247,
    new_n5248, new_n5249, new_n5250, new_n5251, new_n5252, new_n5253,
    new_n5254, new_n5255, new_n5256, new_n5257_1, new_n5258, new_n5259,
    new_n5260, new_n5261, new_n5262, new_n5263, new_n5264, new_n5265,
    new_n5266, new_n5267, new_n5268, new_n5269, new_n5270, new_n5271,
    new_n5272, new_n5273, new_n5274, new_n5275, new_n5276, new_n5277,
    new_n5278, new_n5279, new_n5280, new_n5281, new_n5282, new_n5283_1,
    new_n5284, new_n5285, new_n5286, new_n5287, new_n5288, new_n5289,
    new_n5290, new_n5291, new_n5292, new_n5293, new_n5294, new_n5295,
    new_n5296, new_n5297, new_n5298, new_n5299, new_n5300, new_n5301,
    new_n5302, new_n5303, new_n5304, new_n5305_1, new_n5306, new_n5307,
    new_n5308, new_n5309, new_n5310, new_n5311, new_n5312, new_n5313,
    new_n5314_1, new_n5315, new_n5316, new_n5317, new_n5318, new_n5319_1,
    new_n5320_1, new_n5321, new_n5322, new_n5323, new_n5324, new_n5325,
    new_n5326, new_n5327, new_n5328, new_n5329, new_n5330, new_n5331_1,
    new_n5332, new_n5333, new_n5334, new_n5335, new_n5336, new_n5337,
    new_n5338, new_n5339, new_n5340, new_n5341, new_n5342, new_n5343,
    new_n5344, new_n5345, new_n5346, new_n5347, new_n5348, new_n5349,
    new_n5350, new_n5351, new_n5352, new_n5353, new_n5354, new_n5355,
    new_n5356, new_n5357, new_n5358, new_n5359, new_n5360, new_n5361,
    new_n5362, new_n5363, new_n5364, new_n5365, new_n5366, new_n5367,
    new_n5368, new_n5369, new_n5370, new_n5371, new_n5372, new_n5373,
    new_n5374, new_n5375, new_n5376, new_n5377, new_n5378, new_n5379,
    new_n5380, new_n5381, new_n5382, new_n5383, new_n5384, new_n5385,
    new_n5386, new_n5387, new_n5388, new_n5389, new_n5390, new_n5391,
    new_n5392, new_n5393, new_n5394, new_n5395, new_n5396, new_n5397,
    new_n5398, new_n5399, new_n5400, new_n5401, new_n5402, new_n5403,
    new_n5404, new_n5405, new_n5406, new_n5407, new_n5408, new_n5409,
    new_n5410, new_n5411_1, new_n5412, new_n5413, new_n5414, new_n5415,
    new_n5416, new_n5417, new_n5418, new_n5419, new_n5420, new_n5421,
    new_n5422, new_n5423, new_n5424, new_n5425, new_n5426, new_n5427,
    new_n5428, new_n5429, new_n5430, new_n5431, new_n5432, new_n5433,
    new_n5434, new_n5435_1, new_n5436, new_n5437, new_n5438, new_n5439,
    new_n5440, new_n5441, new_n5442, new_n5443, new_n5444, new_n5445,
    new_n5446, new_n5447, new_n5448, new_n5449, new_n5450, new_n5451,
    new_n5452, new_n5453, new_n5454, new_n5455, new_n5456, new_n5457,
    new_n5458, new_n5459, new_n5460, new_n5461, new_n5462, new_n5463,
    new_n5464, new_n5465, new_n5466, new_n5467, new_n5468, new_n5469,
    new_n5470, new_n5471, new_n5472, new_n5473, new_n5474, new_n5475,
    new_n5476, new_n5477, new_n5478, new_n5479, new_n5481, new_n5482,
    new_n5483, new_n5484, new_n5485, new_n5486, new_n5487, new_n5488,
    new_n5489, new_n5490, new_n5491, new_n5492, new_n5493, new_n5494,
    new_n5495, new_n5496, new_n5497, new_n5498, new_n5499, new_n5500,
    new_n5501, new_n5502, new_n5503, new_n5504, new_n5505, new_n5506,
    new_n5507, new_n5508, new_n5509, new_n5510, new_n5511, new_n5512,
    new_n5513, new_n5514, new_n5515, new_n5516, new_n5517, new_n5518,
    new_n5519, new_n5520, new_n5521, new_n5522, new_n5523, new_n5524,
    new_n5525, new_n5526, new_n5527, new_n5528, new_n5529, new_n5530,
    new_n5531, new_n5532, new_n5533, new_n5534, new_n5535, new_n5536,
    new_n5537, new_n5538, new_n5539, new_n5540, new_n5541, new_n5542,
    new_n5543, new_n5544, new_n5545, new_n5546, new_n5547, new_n5548,
    new_n5549, new_n5550, new_n5551, new_n5552, new_n5553, new_n5554,
    new_n5555, new_n5556, new_n5557, new_n5558, new_n5559, new_n5560,
    new_n5561, new_n5562, new_n5563, new_n5564, new_n5565, new_n5566,
    new_n5567, new_n5568, new_n5569, new_n5570, new_n5571, new_n5572,
    new_n5573, new_n5574, new_n5575, new_n5576, new_n5577, new_n5578,
    new_n5579_1, new_n5580, new_n5581, new_n5582, new_n5583, new_n5584,
    new_n5585, new_n5586, new_n5587, new_n5588, new_n5589, new_n5590,
    new_n5591, new_n5592, new_n5593, new_n5594, new_n5595, new_n5596,
    new_n5597, new_n5598, new_n5599, new_n5600, new_n5601, new_n5602,
    new_n5603, new_n5604, new_n5605, new_n5606, new_n5607, new_n5608,
    new_n5609, new_n5610, new_n5611, new_n5612, new_n5613, new_n5614,
    new_n5615, new_n5616, new_n5617, new_n5618, new_n5619, new_n5620,
    new_n5621, new_n5622, new_n5623, new_n5624, new_n5625, new_n5626,
    new_n5627, new_n5628, new_n5629, new_n5630, new_n5631, new_n5632,
    new_n5633, new_n5634, new_n5635, new_n5636, new_n5637, new_n5638,
    new_n5639, new_n5640, new_n5641_1, new_n5642, new_n5643, new_n5644,
    new_n5645_1, new_n5646, new_n5647, new_n5648, new_n5649, new_n5650,
    new_n5651, new_n5652, new_n5653, new_n5654, new_n5655, new_n5656,
    new_n5657, new_n5658, new_n5659, new_n5660, new_n5661, new_n5662,
    new_n5663, new_n5664, new_n5665, new_n5666, new_n5667, new_n5668,
    new_n5669, new_n5670_1, new_n5671, new_n5672, new_n5673, new_n5674,
    new_n5675, new_n5676, new_n5677, new_n5678, new_n5679, new_n5680,
    new_n5681, new_n5682, new_n5683, new_n5684, new_n5685, new_n5686,
    new_n5687, new_n5688, new_n5689, new_n5690, new_n5691, new_n5692,
    new_n5693_1, new_n5694_1, new_n5695, new_n5696, new_n5697, new_n5698,
    new_n5699, new_n5700, new_n5701, new_n5702, new_n5703, new_n5704,
    new_n5705, new_n5706, new_n5707, new_n5708, new_n5709, new_n5710,
    new_n5711, new_n5712, new_n5713, new_n5714, new_n5715, new_n5716,
    new_n5717, new_n5718, new_n5719, new_n5720, new_n5721, new_n5722,
    new_n5723, new_n5724, new_n5725, new_n5726, new_n5727, new_n5728,
    new_n5729, new_n5730, new_n5731, new_n5732, new_n5733, new_n5734,
    new_n5735, new_n5736, new_n5737, new_n5738, new_n5739, new_n5740,
    new_n5741, new_n5742, new_n5743, new_n5744, new_n5745, new_n5746,
    new_n5747, new_n5748, new_n5749, new_n5750, new_n5751, new_n5752,
    new_n5753, new_n5754, new_n5755, new_n5756, new_n5757, new_n5758,
    new_n5759, new_n5760_1, new_n5761, new_n5762, new_n5763, new_n5764,
    new_n5765, new_n5766, new_n5767_1, new_n5768, new_n5769, new_n5770,
    new_n5771, new_n5772, new_n5773, new_n5774, new_n5775, new_n5776,
    new_n5777, new_n5778, new_n5779, new_n5780, new_n5781, new_n5782,
    new_n5783, new_n5784, new_n5785, new_n5786, new_n5787, new_n5788,
    new_n5789, new_n5790, new_n5791, new_n5792, new_n5793, new_n5794,
    new_n5795, new_n5796, new_n5797, new_n5798_1, new_n5799, new_n5800,
    new_n5801, new_n5802, new_n5803, new_n5804, new_n5805, new_n5806,
    new_n5807, new_n5808, new_n5809, new_n5810, new_n5811, new_n5812,
    new_n5813, new_n5814_1, new_n5815, new_n5816, new_n5817, new_n5818,
    new_n5819, new_n5820, new_n5821, new_n5822, new_n5823, new_n5824,
    new_n5825, new_n5826, new_n5827, new_n5828, new_n5829, new_n5830,
    new_n5831, new_n5832, new_n5833, new_n5834, new_n5835, new_n5836,
    new_n5837, new_n5838, new_n5839, new_n5840, new_n5841, new_n5842,
    new_n5843, new_n5844, new_n5845, new_n5846, new_n5847, new_n5848,
    new_n5849, new_n5850, new_n5851, new_n5852, new_n5853, new_n5854,
    new_n5855, new_n5856, new_n5857_1, new_n5858, new_n5859, new_n5860_1,
    new_n5861, new_n5862, new_n5863, new_n5864, new_n5865, new_n5866,
    new_n5867, new_n5868, new_n5869, new_n5870, new_n5871, new_n5872,
    new_n5873, new_n5874, new_n5875, new_n5876, new_n5877, new_n5878,
    new_n5879, new_n5880, new_n5881, new_n5882, new_n5883, new_n5884,
    new_n5885, new_n5886, new_n5887, new_n5888, new_n5889, new_n5890,
    new_n5891, new_n5892, new_n5893, new_n5894, new_n5895, new_n5896,
    new_n5897, new_n5898, new_n5899, new_n5900, new_n5901, new_n5902,
    new_n5903, new_n5904, new_n5905, new_n5906, new_n5907, new_n5908,
    new_n5909, new_n5910, new_n5911, new_n5912, new_n5913, new_n5914,
    new_n5915, new_n5916, new_n5917, new_n5918, new_n5919, new_n5920,
    new_n5921, new_n5922, new_n5923, new_n5924, new_n5925, new_n5926,
    new_n5927, new_n5928, new_n5929, new_n5930, new_n5931, new_n5932,
    new_n5933, new_n5934_1, new_n5935, new_n5936, new_n5937, new_n5938,
    new_n5939, new_n5940, new_n5941, new_n5942, new_n5944, new_n5945,
    new_n5946, new_n5947, new_n5948, new_n5949, new_n5950, new_n5951,
    new_n5952, new_n5953, new_n5954, new_n5955, new_n5956, new_n5957,
    new_n5958, new_n5959, new_n5960, new_n5961, new_n5962, new_n5963,
    new_n5964_1, new_n5965, new_n5966, new_n5967, new_n5968, new_n5969,
    new_n5970, new_n5971, new_n5972, new_n5973, new_n5974, new_n5975,
    new_n5976, new_n5977, new_n5978, new_n5979, new_n5980, new_n5981,
    new_n5982, new_n5983, new_n5984, new_n5985, new_n5986, new_n5987,
    new_n5988, new_n5989, new_n5990, new_n5991, new_n5992, new_n5993,
    new_n5994, new_n5995, new_n5996, new_n5997, new_n5998, new_n5999,
    new_n6000, new_n6001, new_n6002, new_n6003, new_n6004, new_n6005,
    new_n6006, new_n6007, new_n6008, new_n6009, new_n6010, new_n6011,
    new_n6012, new_n6013, new_n6014, new_n6015, new_n6016_1, new_n6017,
    new_n6018, new_n6019, new_n6020, new_n6021, new_n6022, new_n6023,
    new_n6024, new_n6025, new_n6026, new_n6027, new_n6028, new_n6029,
    new_n6030, new_n6031, new_n6032, new_n6033, new_n6034, new_n6035,
    new_n6036, new_n6037, new_n6038_1, new_n6039, new_n6040, new_n6041,
    new_n6042, new_n6043, new_n6044, new_n6045, new_n6046, new_n6047,
    new_n6048, new_n6049, new_n6050, new_n6051, new_n6052, new_n6053,
    new_n6054, new_n6055, new_n6056, new_n6057, new_n6058, new_n6059,
    new_n6060, new_n6061, new_n6062, new_n6063, new_n6064, new_n6065,
    new_n6066, new_n6067, new_n6068, new_n6069, new_n6070, new_n6071,
    new_n6072, new_n6073, new_n6074, new_n6075, new_n6076, new_n6077,
    new_n6078, new_n6079, new_n6080, new_n6081, new_n6082, new_n6083,
    new_n6084, new_n6085, new_n6086, new_n6087, new_n6088, new_n6089_1,
    new_n6090, new_n6091, new_n6092, new_n6093, new_n6094, new_n6095,
    new_n6096, new_n6097, new_n6098, new_n6099, new_n6100, new_n6101,
    new_n6102, new_n6103, new_n6104, new_n6105, new_n6106, new_n6107,
    new_n6108, new_n6109, new_n6110, new_n6111, new_n6112, new_n6113,
    new_n6114, new_n6115, new_n6116, new_n6117, new_n6118, new_n6119,
    new_n6120, new_n6121, new_n6122, new_n6123, new_n6124, new_n6125,
    new_n6126_1, new_n6127, new_n6128, new_n6129, new_n6130, new_n6131,
    new_n6132, new_n6133, new_n6134, new_n6135, new_n6136, new_n6137,
    new_n6138, new_n6139, new_n6140, new_n6141, new_n6142, new_n6143,
    new_n6144, new_n6145, new_n6146, new_n6147, new_n6148, new_n6149,
    new_n6150, new_n6151, new_n6152, new_n6153, new_n6154, new_n6155,
    new_n6156, new_n6157, new_n6158, new_n6159, new_n6160, new_n6161,
    new_n6162, new_n6163, new_n6164, new_n6165, new_n6166, new_n6167,
    new_n6168, new_n6169, new_n6170, new_n6171, new_n6172, new_n6173,
    new_n6174, new_n6175, new_n6176, new_n6177, new_n6178, new_n6179,
    new_n6180, new_n6181, new_n6182, new_n6183, new_n6184, new_n6185,
    new_n6186, new_n6187, new_n6188, new_n6189, new_n6190, new_n6191,
    new_n6192_1, new_n6193, new_n6194, new_n6195, new_n6196, new_n6197,
    new_n6198, new_n6199, new_n6200, new_n6201, new_n6202, new_n6203,
    new_n6204, new_n6205, new_n6206, new_n6207, new_n6208, new_n6209,
    new_n6210, new_n6211, new_n6212, new_n6213, new_n6214, new_n6215,
    new_n6216, new_n6217, new_n6218, new_n6219, new_n6220, new_n6221,
    new_n6222, new_n6223, new_n6224, new_n6225, new_n6226, new_n6227,
    new_n6228, new_n6229, new_n6230, new_n6231, new_n6232, new_n6233,
    new_n6234, new_n6235, new_n6236, new_n6237, new_n6238, new_n6239,
    new_n6240, new_n6241, new_n6242, new_n6243, new_n6244, new_n6245,
    new_n6246, new_n6247, new_n6248, new_n6249, new_n6250, new_n6251,
    new_n6252, new_n6253, new_n6254_1, new_n6255, new_n6256, new_n6257,
    new_n6258, new_n6259, new_n6260, new_n6261, new_n6262, new_n6263,
    new_n6264, new_n6265, new_n6266, new_n6267, new_n6268, new_n6269,
    new_n6270, new_n6271, new_n6272, new_n6273_1, new_n6274, new_n6275,
    new_n6276, new_n6277, new_n6278, new_n6279, new_n6280, new_n6281,
    new_n6282, new_n6283, new_n6284, new_n6285, new_n6286, new_n6287,
    new_n6289, new_n6290, new_n6291, new_n6292, new_n6293, new_n6294_1,
    new_n6295, new_n6296, new_n6297, new_n6298, new_n6299, new_n6300,
    new_n6301, new_n6302, new_n6303, new_n6304, new_n6305, new_n6306,
    new_n6307, new_n6308, new_n6309, new_n6310, new_n6311, new_n6312,
    new_n6313, new_n6314, new_n6315, new_n6316, new_n6317, new_n6318,
    new_n6319, new_n6320, new_n6321, new_n6322, new_n6323, new_n6324,
    new_n6325, new_n6326, new_n6327, new_n6328, new_n6329, new_n6330,
    new_n6331, new_n6332, new_n6333, new_n6334, new_n6335, new_n6336,
    new_n6337, new_n6338, new_n6339, new_n6340, new_n6341, new_n6342,
    new_n6343, new_n6344, new_n6345, new_n6346, new_n6347, new_n6348,
    new_n6349, new_n6350, new_n6351, new_n6352, new_n6353, new_n6354,
    new_n6355, new_n6356, new_n6357, new_n6358_1, new_n6359_1, new_n6360,
    new_n6361, new_n6362, new_n6363, new_n6364, new_n6365, new_n6366,
    new_n6367, new_n6368, new_n6369, new_n6370, new_n6371, new_n6372,
    new_n6373, new_n6374, new_n6375, new_n6376, new_n6377, new_n6378,
    new_n6379, new_n6380, new_n6381, new_n6382, new_n6383, new_n6384,
    new_n6385, new_n6386, new_n6387, new_n6388, new_n6389, new_n6390,
    new_n6391, new_n6392, new_n6393, new_n6394, new_n6395, new_n6396,
    new_n6397, new_n6398, new_n6399, new_n6400, new_n6401, new_n6402,
    new_n6403, new_n6404, new_n6405, new_n6406, new_n6407, new_n6408,
    new_n6409, new_n6410, new_n6411, new_n6412, new_n6413, new_n6414,
    new_n6415, new_n6416, new_n6417, new_n6418, new_n6419, new_n6420,
    new_n6421, new_n6422, new_n6423, new_n6424, new_n6425, new_n6426,
    new_n6427, new_n6428, new_n6429_1, new_n6430, new_n6431_1, new_n6432,
    new_n6433, new_n6434, new_n6435, new_n6436, new_n6437, new_n6438,
    new_n6439, new_n6440, new_n6441_1, new_n6442, new_n6443, new_n6444,
    new_n6445_1, new_n6446, new_n6447, new_n6448, new_n6449, new_n6450,
    new_n6451, new_n6452, new_n6453, new_n6454, new_n6455, new_n6456,
    new_n6457, new_n6458, new_n6459, new_n6460, new_n6461, new_n6462,
    new_n6463, new_n6464, new_n6465, new_n6466, new_n6467, new_n6468,
    new_n6469, new_n6470, new_n6471, new_n6472, new_n6473, new_n6474,
    new_n6475, new_n6476, new_n6477, new_n6478, new_n6479, new_n6480,
    new_n6481, new_n6482, new_n6483, new_n6484, new_n6485, new_n6486,
    new_n6487, new_n6488, new_n6489, new_n6490, new_n6491, new_n6492,
    new_n6493, new_n6494, new_n6495, new_n6496, new_n6497, new_n6498,
    new_n6499, new_n6500, new_n6501, new_n6502, new_n6503, new_n6504,
    new_n6505, new_n6506, new_n6507, new_n6508, new_n6509, new_n6510,
    new_n6511, new_n6512, new_n6513, new_n6514, new_n6515, new_n6516,
    new_n6517, new_n6518, new_n6519, new_n6520, new_n6521, new_n6522,
    new_n6523, new_n6524, new_n6525, new_n6526, new_n6528, new_n6529,
    new_n6530, new_n6531, new_n6532, new_n6533, new_n6534, new_n6535,
    new_n6536, new_n6537, new_n6538, new_n6539, new_n6540, new_n6541,
    new_n6542, new_n6543, new_n6544, new_n6545, new_n6546, new_n6547,
    new_n6548, new_n6549, new_n6550, new_n6551, new_n6552, new_n6553,
    new_n6554, new_n6555, new_n6556, new_n6557, new_n6558, new_n6559,
    new_n6560, new_n6561, new_n6564, new_n6565, new_n6566, new_n6567,
    new_n6568, new_n6569, new_n6570, new_n6571, new_n6572, new_n6573,
    new_n6574, new_n6575, new_n6576, new_n6577, new_n6578_1, new_n6579,
    new_n6580, new_n6581, new_n6582, new_n6583, new_n6584, new_n6585,
    new_n6586, new_n6587, new_n6588, new_n6589, new_n6590, new_n6591,
    new_n6592, new_n6593, new_n6594, new_n6595, new_n6596, new_n6597,
    new_n6598, new_n6599, new_n6600, new_n6601, new_n6602, new_n6603,
    new_n6604_1, new_n6605, new_n6606, new_n6607, new_n6608, new_n6609,
    new_n6610, new_n6611_1, new_n6612, new_n6613, new_n6614, new_n6615,
    new_n6616, new_n6617, new_n6618, new_n6619, new_n6620, new_n6621,
    new_n6622, new_n6623, new_n6624, new_n6625, new_n6626, new_n6627,
    new_n6628, new_n6629, new_n6630, new_n6631, new_n6632, new_n6633,
    new_n6634, new_n6635, new_n6636, new_n6637, new_n6638, new_n6639,
    new_n6640, new_n6641, new_n6642, new_n6643, new_n6644, new_n6645_1,
    new_n6646, new_n6647, new_n6648, new_n6649, new_n6650, new_n6651,
    new_n6652, new_n6653, new_n6654, new_n6655, new_n6656, new_n6657,
    new_n6658, new_n6659, new_n6660, new_n6661, new_n6662, new_n6663,
    new_n6664, new_n6665, new_n6666, new_n6667, new_n6668, new_n6669,
    new_n6670, new_n6671, new_n6672, new_n6673, new_n6674, new_n6675,
    new_n6676, new_n6677, new_n6678, new_n6679, new_n6680, new_n6681,
    new_n6682, new_n6683, new_n6684, new_n6685, new_n6686, new_n6687_1,
    new_n6688, new_n6689_1, new_n6690, new_n6691, new_n6692, new_n6693,
    new_n6694, new_n6695, new_n6696, new_n6697, new_n6698, new_n6699,
    new_n6700, new_n6701, new_n6702, new_n6703_1, new_n6704, new_n6705,
    new_n6706, new_n6707, new_n6708, new_n6709, new_n6710, new_n6711,
    new_n6712, new_n6713, new_n6714, new_n6715, new_n6716, new_n6717,
    new_n6718, new_n6719, new_n6720, new_n6721, new_n6722, new_n6723,
    new_n6724, new_n6725, new_n6726, new_n6727, new_n6728, new_n6729,
    new_n6730, new_n6731, new_n6732, new_n6733, new_n6734, new_n6735,
    new_n6736, new_n6737, new_n6738, new_n6739, new_n6740, new_n6741,
    new_n6742_1, new_n6743, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770_1, new_n6771,
    new_n6772, new_n6773, new_n6774, new_n6775, new_n6776_1, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790, new_n6791, new_n6792, new_n6793, new_n6794, new_n6795,
    new_n6796, new_n6797_1, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802, new_n6803, new_n6804, new_n6805, new_n6806_1, new_n6807,
    new_n6808, new_n6809_1, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822_1, new_n6823, new_n6824, new_n6825,
    new_n6826_1, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860_1, new_n6861,
    new_n6862, new_n6863, new_n6864, new_n6865, new_n6866, new_n6867,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877_1, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6965, new_n6966, new_n6967, new_n6968, new_n6969,
    new_n6970, new_n6971, new_n6972, new_n6973, new_n6974, new_n6975,
    new_n6976, new_n6977, new_n6978, new_n6979, new_n6980, new_n6981,
    new_n6982, new_n6983, new_n6984, new_n6985, new_n6986_1, new_n6987,
    new_n6988, new_n6989, new_n6990, new_n6991, new_n6992, new_n6993,
    new_n6994, new_n6995, new_n6996, new_n6997, new_n6998, new_n6999,
    new_n7000, new_n7001, new_n7002, new_n7003, new_n7004, new_n7005,
    new_n7006, new_n7007, new_n7008, new_n7009, new_n7010, new_n7011,
    new_n7012, new_n7013, new_n7014, new_n7015, new_n7016, new_n7017,
    new_n7018, new_n7019, new_n7020, new_n7021, new_n7022, new_n7023,
    new_n7024, new_n7025, new_n7026, new_n7027, new_n7028, new_n7029,
    new_n7030, new_n7031, new_n7032, new_n7033, new_n7034, new_n7035,
    new_n7036, new_n7037, new_n7038, new_n7039, new_n7042, new_n7043,
    new_n7044, new_n7045, new_n7046, new_n7047, new_n7048, new_n7049,
    new_n7050, new_n7051, new_n7052, new_n7053, new_n7054, new_n7055,
    new_n7056, new_n7057, new_n7058, new_n7059, new_n7060, new_n7061,
    new_n7062, new_n7063, new_n7064, new_n7065, new_n7066, new_n7067,
    new_n7068, new_n7069, new_n7070, new_n7071, new_n7072, new_n7073,
    new_n7074, new_n7075, new_n7076, new_n7077, new_n7078, new_n7079,
    new_n7080, new_n7081, new_n7082, new_n7083, new_n7084, new_n7085,
    new_n7086, new_n7087, new_n7088, new_n7089, new_n7090, new_n7091,
    new_n7092, new_n7093, new_n7094, new_n7095, new_n7096, new_n7097,
    new_n7098, new_n7099, new_n7100, new_n7101, new_n7102, new_n7103,
    new_n7104, new_n7105, new_n7106, new_n7107, new_n7108, new_n7109,
    new_n7110, new_n7111, new_n7112, new_n7113, new_n7114, new_n7115,
    new_n7116, new_n7117, new_n7118, new_n7119, new_n7120, new_n7121,
    new_n7122, new_n7123, new_n7124, new_n7125, new_n7126, new_n7127,
    new_n7128, new_n7129, new_n7130, new_n7131, new_n7132, new_n7133,
    new_n7134, new_n7135, new_n7136, new_n7137, new_n7138, new_n7139,
    new_n7140, new_n7141, new_n7142, new_n7143, new_n7144, new_n7145,
    new_n7146, new_n7147, new_n7148, new_n7149, new_n7150, new_n7151,
    new_n7152, new_n7153, new_n7154, new_n7155, new_n7156, new_n7157,
    new_n7158, new_n7159_1, new_n7160_1, new_n7161, new_n7162, new_n7163,
    new_n7164, new_n7165, new_n7166, new_n7167, new_n7168, new_n7169,
    new_n7170, new_n7171, new_n7172, new_n7173, new_n7174, new_n7175,
    new_n7176, new_n7177, new_n7178, new_n7179, new_n7180, new_n7181,
    new_n7182, new_n7183, new_n7184, new_n7185, new_n7186, new_n7187,
    new_n7188, new_n7189, new_n7190, new_n7191, new_n7192, new_n7193_1,
    new_n7194, new_n7195, new_n7196, new_n7197, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7202, new_n7203, new_n7204, new_n7205,
    new_n7206, new_n7207, new_n7208, new_n7209, new_n7210, new_n7211,
    new_n7212, new_n7213, new_n7214, new_n7215, new_n7216, new_n7217,
    new_n7218, new_n7219, new_n7220, new_n7221, new_n7222, new_n7223,
    new_n7224, new_n7225, new_n7226, new_n7227, new_n7228, new_n7229,
    new_n7230, new_n7231, new_n7232, new_n7233, new_n7234, new_n7235,
    new_n7236_1, new_n7237, new_n7238, new_n7239, new_n7240, new_n7241,
    new_n7242, new_n7243, new_n7244, new_n7245, new_n7246, new_n7247,
    new_n7248, new_n7249, new_n7250, new_n7251, new_n7252, new_n7253,
    new_n7254, new_n7255, new_n7256, new_n7257, new_n7258, new_n7259,
    new_n7260, new_n7261, new_n7262, new_n7263, new_n7264, new_n7265_1,
    new_n7266, new_n7267, new_n7268, new_n7269, new_n7270_1, new_n7271,
    new_n7272, new_n7273, new_n7274, new_n7275, new_n7276, new_n7277,
    new_n7278, new_n7279, new_n7280, new_n7281, new_n7282, new_n7283,
    new_n7284, new_n7285, new_n7286, new_n7287, new_n7288, new_n7289,
    new_n7290, new_n7291, new_n7292, new_n7293, new_n7294_1, new_n7295,
    new_n7296, new_n7297, new_n7298, new_n7299, new_n7300, new_n7301,
    new_n7302, new_n7303, new_n7304, new_n7305, new_n7306, new_n7307,
    new_n7308, new_n7309, new_n7310, new_n7311, new_n7312, new_n7313,
    new_n7314, new_n7315, new_n7316, new_n7317, new_n7318, new_n7319,
    new_n7320_1, new_n7321, new_n7322, new_n7323, new_n7324, new_n7325,
    new_n7326, new_n7327, new_n7328, new_n7329, new_n7330, new_n7331,
    new_n7332, new_n7333, new_n7334, new_n7335, new_n7336, new_n7337,
    new_n7338, new_n7339, new_n7340, new_n7341, new_n7342, new_n7343,
    new_n7344, new_n7345, new_n7346, new_n7347, new_n7348, new_n7349,
    new_n7350, new_n7351, new_n7352, new_n7353, new_n7354_1, new_n7355,
    new_n7356, new_n7357, new_n7358, new_n7359, new_n7360, new_n7361,
    new_n7362, new_n7363, new_n7364, new_n7365, new_n7366, new_n7367,
    new_n7368, new_n7369, new_n7370, new_n7371, new_n7372, new_n7373,
    new_n7374, new_n7375, new_n7376, new_n7377, new_n7378, new_n7379,
    new_n7380, new_n7381, new_n7382, new_n7383, new_n7384, new_n7385,
    new_n7386, new_n7387, new_n7388_1, new_n7389, new_n7390, new_n7391,
    new_n7392, new_n7393, new_n7394, new_n7395, new_n7396, new_n7397,
    new_n7398, new_n7399, new_n7400, new_n7401, new_n7402, new_n7403,
    new_n7404, new_n7405, new_n7406, new_n7407, new_n7408, new_n7409,
    new_n7410, new_n7411, new_n7412, new_n7413, new_n7414, new_n7415,
    new_n7416, new_n7417, new_n7418, new_n7419, new_n7420, new_n7421,
    new_n7422, new_n7423, new_n7424, new_n7425, new_n7426, new_n7427,
    new_n7428, new_n7429, new_n7430, new_n7431, new_n7432, new_n7433,
    new_n7434, new_n7435, new_n7436_1, new_n7437, new_n7438, new_n7439,
    new_n7440, new_n7441, new_n7442, new_n7443, new_n7444, new_n7445,
    new_n7446, new_n7447, new_n7448, new_n7449, new_n7450, new_n7451,
    new_n7452, new_n7453, new_n7454, new_n7455, new_n7456_1, new_n7457,
    new_n7458, new_n7459, new_n7460, new_n7461, new_n7462, new_n7463,
    new_n7464, new_n7465, new_n7466, new_n7467, new_n7468, new_n7469,
    new_n7470, new_n7471, new_n7472, new_n7473, new_n7474, new_n7475,
    new_n7476, new_n7477, new_n7478, new_n7479, new_n7480, new_n7481,
    new_n7482, new_n7483, new_n7484, new_n7485, new_n7486, new_n7487,
    new_n7488, new_n7489, new_n7490, new_n7491, new_n7492, new_n7493,
    new_n7494, new_n7495, new_n7496, new_n7497, new_n7498, new_n7499,
    new_n7500_1, new_n7501, new_n7502, new_n7503, new_n7504, new_n7505,
    new_n7506, new_n7507, new_n7508, new_n7509, new_n7510, new_n7511,
    new_n7512, new_n7513, new_n7514, new_n7515, new_n7516, new_n7517,
    new_n7518, new_n7519, new_n7520, new_n7521, new_n7522, new_n7523_1,
    new_n7524, new_n7525, new_n7526, new_n7527, new_n7528, new_n7529,
    new_n7530, new_n7531, new_n7532, new_n7533, new_n7534, new_n7535,
    new_n7536, new_n7537, new_n7538, new_n7539, new_n7540, new_n7541,
    new_n7542, new_n7543, new_n7544, new_n7545, new_n7546_1, new_n7547,
    new_n7548, new_n7549, new_n7550, new_n7551, new_n7552, new_n7553,
    new_n7554, new_n7555, new_n7556, new_n7557, new_n7558, new_n7559,
    new_n7560, new_n7561, new_n7562, new_n7563, new_n7564, new_n7565,
    new_n7566, new_n7567, new_n7568_1, new_n7569, new_n7570, new_n7571,
    new_n7572, new_n7573, new_n7574, new_n7575, new_n7576, new_n7577,
    new_n7578, new_n7579, new_n7580, new_n7581, new_n7582, new_n7583,
    new_n7584, new_n7585, new_n7586, new_n7587, new_n7588, new_n7589,
    new_n7590, new_n7591, new_n7592, new_n7593, new_n7594, new_n7595,
    new_n7596, new_n7597, new_n7598, new_n7599, new_n7600, new_n7601,
    new_n7602, new_n7603, new_n7604, new_n7605, new_n7606, new_n7607,
    new_n7608, new_n7609, new_n7610_1, new_n7611, new_n7612, new_n7613,
    new_n7614, new_n7615, new_n7616, new_n7617, new_n7618, new_n7619,
    new_n7620, new_n7621, new_n7622, new_n7623, new_n7624, new_n7625,
    new_n7626, new_n7627, new_n7628, new_n7629, new_n7630, new_n7631,
    new_n7632, new_n7633, new_n7634, new_n7635, new_n7636, new_n7637,
    new_n7638, new_n7639, new_n7640, new_n7641, new_n7642, new_n7643,
    new_n7644, new_n7645, new_n7646_1, new_n7647, new_n7648, new_n7649,
    new_n7650, new_n7651, new_n7652, new_n7653, new_n7654, new_n7655,
    new_n7656, new_n7657, new_n7658, new_n7659, new_n7660, new_n7661,
    new_n7662, new_n7663, new_n7664, new_n7665, new_n7666, new_n7667,
    new_n7668, new_n7669, new_n7670, new_n7671, new_n7672, new_n7673,
    new_n7674, new_n7675, new_n7676_1, new_n7677, new_n7678, new_n7679,
    new_n7680, new_n7681, new_n7682, new_n7683, new_n7684, new_n7685,
    new_n7686, new_n7687, new_n7688, new_n7689, new_n7690_1, new_n7691,
    new_n7692, new_n7693, new_n7694, new_n7695, new_n7696, new_n7697,
    new_n7698, new_n7699, new_n7700, new_n7701, new_n7702, new_n7703,
    new_n7704, new_n7705, new_n7706, new_n7707, new_n7708, new_n7709,
    new_n7710, new_n7712, new_n7714, new_n7715, new_n7718, new_n7720,
    new_n7722, new_n7723, new_n7724, new_n7725, new_n7726, new_n7727,
    new_n7728, new_n7729, new_n7730_1, new_n7731, new_n7732, new_n7733_1,
    new_n7734, new_n7735, new_n7736, new_n7737, new_n7738, new_n7739,
    new_n7740, new_n7741, new_n7742, new_n7743, new_n7744, new_n7745,
    new_n7746, new_n7747, new_n7748, new_n7749, new_n7750, new_n7751,
    new_n7752, new_n7753, new_n7754, new_n7755, new_n7756, new_n7757,
    new_n7758, new_n7759, new_n7760, new_n7761, new_n7762, new_n7763,
    new_n7764, new_n7765, new_n7766, new_n7767, new_n7768, new_n7769,
    new_n7770, new_n7771, new_n7772, new_n7773, new_n7774, new_n7775,
    new_n7776, new_n7777, new_n7778, new_n7779, new_n7780, new_n7781,
    new_n7782, new_n7783, new_n7784, new_n7785, new_n7786, new_n7787,
    new_n7788, new_n7789, new_n7790, new_n7791, new_n7792, new_n7793,
    new_n7794, new_n7795, new_n7796, new_n7797, new_n7798, new_n7799,
    new_n7800, new_n7801, new_n7802, new_n7803, new_n7804, new_n7805,
    new_n7806, new_n7807, new_n7808, new_n7809, new_n7810, new_n7811,
    new_n7812, new_n7813, new_n7814, new_n7815, new_n7816, new_n7817,
    new_n7818, new_n7819, new_n7820, new_n7821, new_n7822, new_n7823_1,
    new_n7824, new_n7825, new_n7826, new_n7827, new_n7828, new_n7829,
    new_n7830, new_n7831, new_n7832, new_n7833, new_n7834, new_n7835,
    new_n7836, new_n7837, new_n7838, new_n7839, new_n7840, new_n7841,
    new_n7842, new_n7843, new_n7844, new_n7845, new_n7846, new_n7847,
    new_n7848, new_n7849, new_n7850, new_n7851, new_n7852, new_n7853,
    new_n7854, new_n7855, new_n7856, new_n7857, new_n7858, new_n7859,
    new_n7860, new_n7861, new_n7862_1, new_n7863, new_n7864, new_n7865,
    new_n7866, new_n7867, new_n7868, new_n7869, new_n7870, new_n7871,
    new_n7872, new_n7873, new_n7874, new_n7875, new_n7876, new_n7877,
    new_n7878, new_n7879, new_n7880, new_n7881, new_n7882, new_n7883,
    new_n7884, new_n7885, new_n7886, new_n7887, new_n7888, new_n7889,
    new_n7890, new_n7891_1, new_n7892, new_n7893, new_n7894, new_n7895,
    new_n7896, new_n7897, new_n7898, new_n7899, new_n7900, new_n7901,
    new_n7902, new_n7903, new_n7904, new_n7905, new_n7906, new_n7907,
    new_n7908, new_n7909, new_n7910, new_n7911, new_n7912, new_n7913,
    new_n7914, new_n7915, new_n7916, new_n7917, new_n7918, new_n7919,
    new_n7920, new_n7921, new_n7922, new_n7923, new_n7924, new_n7925,
    new_n7926, new_n7927, new_n7928, new_n7929, new_n7930, new_n7931,
    new_n7932, new_n7933, new_n7934, new_n7935, new_n7936, new_n7937,
    new_n7938, new_n7939, new_n7940, new_n7941, new_n7942, new_n7943,
    new_n7944, new_n7945, new_n7946_1, new_n7947, new_n7948, new_n7949,
    new_n7950, new_n7951, new_n7952, new_n7953, new_n7954, new_n7955,
    new_n7956, new_n7957, new_n7958, new_n7959, new_n7960, new_n7961,
    new_n7962, new_n7963, new_n7964, new_n7965_1, new_n7966_1, new_n7967,
    new_n7968, new_n7969, new_n7970, new_n7971, new_n7972, new_n7973,
    new_n7974, new_n7975, new_n7976, new_n7977, new_n7978, new_n7979,
    new_n7980, new_n7981_1, new_n7982, new_n7983, new_n7984, new_n7985,
    new_n7986, new_n7987, new_n7988, new_n7989, new_n7990, new_n7991,
    new_n7992, new_n7993, new_n7994, new_n7995, new_n7996, new_n7997,
    new_n7998, new_n7999, new_n8000, new_n8001, new_n8002, new_n8003,
    new_n8004, new_n8005, new_n8006, new_n8007, new_n8008, new_n8009,
    new_n8010, new_n8011, new_n8012, new_n8013, new_n8014, new_n8015,
    new_n8016, new_n8017, new_n8018, new_n8019, new_n8020, new_n8021,
    new_n8022, new_n8023, new_n8024, new_n8025, new_n8026, new_n8027,
    new_n8028_1, new_n8029, new_n8030, new_n8031, new_n8032, new_n8033,
    new_n8034, new_n8035, new_n8036, new_n8037, new_n8038, new_n8039,
    new_n8040, new_n8041, new_n8042, new_n8043, new_n8044, new_n8045,
    new_n8046, new_n8047, new_n8048, new_n8049, new_n8050, new_n8051,
    new_n8052, new_n8053, new_n8054, new_n8055, new_n8056, new_n8057,
    new_n8058, new_n8059, new_n8060, new_n8061, new_n8062, new_n8063,
    new_n8064, new_n8065_1, new_n8066, new_n8067, new_n8068, new_n8069,
    new_n8070, new_n8071, new_n8072, new_n8073, new_n8074, new_n8075,
    new_n8076, new_n8077, new_n8078, new_n8079, new_n8080, new_n8081,
    new_n8082, new_n8083, new_n8084, new_n8085, new_n8086, new_n8087,
    new_n8088, new_n8089, new_n8090, new_n8091, new_n8092, new_n8093,
    new_n8094, new_n8095, new_n8096, new_n8097, new_n8098, new_n8099,
    new_n8100_1, new_n8101, new_n8102, new_n8103, new_n8104, new_n8105,
    new_n8106, new_n8107, new_n8108, new_n8109, new_n8110, new_n8111,
    new_n8112, new_n8113, new_n8114, new_n8115, new_n8116, new_n8117,
    new_n8118, new_n8119, new_n8120, new_n8121, new_n8122, new_n8123,
    new_n8124, new_n8125, new_n8126, new_n8127, new_n8128, new_n8129,
    new_n8130, new_n8131, new_n8132, new_n8133, new_n8134, new_n8135,
    new_n8136, new_n8137, new_n8138_1, new_n8139, new_n8140, new_n8141,
    new_n8142, new_n8143, new_n8144, new_n8145, new_n8146, new_n8147,
    new_n8148, new_n8149, new_n8150, new_n8151, new_n8152, new_n8153,
    new_n8154, new_n8155, new_n8156, new_n8157, new_n8158, new_n8159,
    new_n8160, new_n8161, new_n8162, new_n8163, new_n8164, new_n8165,
    new_n8166, new_n8167, new_n8168, new_n8169, new_n8170, new_n8171,
    new_n8172, new_n8173, new_n8174, new_n8175, new_n8176, new_n8177,
    new_n8178, new_n8179, new_n8180, new_n8181, new_n8182, new_n8183,
    new_n8184, new_n8185, new_n8186, new_n8187, new_n8188, new_n8189,
    new_n8190, new_n8191, new_n8192, new_n8193, new_n8194, new_n8195,
    new_n8196, new_n8197, new_n8198, new_n8199, new_n8200, new_n8201,
    new_n8202_1, new_n8203, new_n8204, new_n8205, new_n8206, new_n8207,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236_1, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255,
    new_n8256, new_n8257, new_n8258, new_n8259, new_n8260, new_n8261,
    new_n8263, new_n8264, new_n8265, new_n8266, new_n8267, new_n8268,
    new_n8269, new_n8270, new_n8271, new_n8272, new_n8273, new_n8274,
    new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279, new_n8280,
    new_n8281, new_n8282, new_n8283, new_n8284, new_n8285, new_n8286,
    new_n8287, new_n8288, new_n8289, new_n8290, new_n8291, new_n8292,
    new_n8293, new_n8294, new_n8295, new_n8296, new_n8297, new_n8298,
    new_n8299, new_n8300, new_n8301, new_n8302, new_n8303_1, new_n8304,
    new_n8305, new_n8306, new_n8307, new_n8308, new_n8309, new_n8310,
    new_n8311, new_n8312, new_n8313, new_n8314, new_n8315, new_n8316,
    new_n8317, new_n8318, new_n8319, new_n8320, new_n8321, new_n8322,
    new_n8323, new_n8324, new_n8325, new_n8326, new_n8327, new_n8328,
    new_n8329, new_n8330, new_n8331, new_n8332, new_n8333, new_n8334,
    new_n8335, new_n8336_1, new_n8337, new_n8338, new_n8339, new_n8340,
    new_n8341, new_n8342, new_n8343, new_n8344, new_n8345, new_n8346,
    new_n8347, new_n8348, new_n8349, new_n8350, new_n8351, new_n8352,
    new_n8353, new_n8354, new_n8355, new_n8356, new_n8357, new_n8358,
    new_n8359, new_n8360, new_n8361, new_n8362, new_n8363, new_n8364,
    new_n8365, new_n8366, new_n8367, new_n8368, new_n8369, new_n8370,
    new_n8371, new_n8372, new_n8373, new_n8374, new_n8375, new_n8376,
    new_n8377, new_n8378, new_n8379, new_n8380, new_n8381, new_n8382,
    new_n8383, new_n8384_1, new_n8385, new_n8386, new_n8387, new_n8388,
    new_n8389, new_n8390, new_n8391, new_n8392, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398_1, new_n8399, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405, new_n8406,
    new_n8407, new_n8408, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8427,
    new_n8428, new_n8429, new_n8430, new_n8431, new_n8432, new_n8433_1,
    new_n8434, new_n8435, new_n8436, new_n8438, new_n8440, new_n8441,
    new_n8442, new_n8443, new_n8444, new_n8445, new_n8446, new_n8447,
    new_n8448, new_n8449, new_n8450, new_n8451, new_n8452, new_n8453,
    new_n8454, new_n8455, new_n8456, new_n8457, new_n8458, new_n8459,
    new_n8460, new_n8461, new_n8462, new_n8463, new_n8464, new_n8465,
    new_n8466, new_n8467, new_n8468, new_n8469, new_n8470, new_n8471,
    new_n8472, new_n8473, new_n8474, new_n8475, new_n8476_1, new_n8477,
    new_n8478, new_n8479, new_n8480, new_n8481, new_n8482, new_n8483,
    new_n8484, new_n8485, new_n8486, new_n8487, new_n8488, new_n8489,
    new_n8490, new_n8491, new_n8492, new_n8493, new_n8494, new_n8495,
    new_n8496, new_n8497, new_n8498, new_n8499, new_n8500, new_n8501,
    new_n8502, new_n8503, new_n8504, new_n8505, new_n8506, new_n8507,
    new_n8508, new_n8509, new_n8510, new_n8511, new_n8512, new_n8513,
    new_n8514, new_n8515, new_n8516, new_n8517, new_n8518, new_n8519,
    new_n8520, new_n8521, new_n8522, new_n8523, new_n8524, new_n8525,
    new_n8526, new_n8527, new_n8528, new_n8529, new_n8530, new_n8531,
    new_n8532, new_n8533, new_n8534, new_n8535, new_n8536, new_n8537,
    new_n8538, new_n8539, new_n8540, new_n8541, new_n8542, new_n8543,
    new_n8544, new_n8545, new_n8546, new_n8547, new_n8548, new_n8549,
    new_n8550, new_n8551, new_n8552, new_n8554, new_n8555, new_n8557,
    new_n8558, new_n8560, new_n8561, new_n8562, new_n8563, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8571, new_n8572, new_n8573, new_n8574, new_n8575, new_n8576,
    new_n8577, new_n8578, new_n8579, new_n8580, new_n8581, new_n8582,
    new_n8583, new_n8584, new_n8585, new_n8586, new_n8587, new_n8588,
    new_n8589, new_n8590, new_n8591, new_n8592, new_n8593, new_n8594,
    new_n8595_1, new_n8596, new_n8597, new_n8598, new_n8599, new_n8600,
    new_n8601, new_n8602, new_n8603, new_n8604, new_n8605, new_n8606,
    new_n8607, new_n8608, new_n8609, new_n8610, new_n8611, new_n8612,
    new_n8613, new_n8614, new_n8615, new_n8616, new_n8617, new_n8618,
    new_n8619, new_n8620, new_n8621, new_n8622, new_n8623, new_n8624,
    new_n8625, new_n8626, new_n8627, new_n8628, new_n8629, new_n8630,
    new_n8631, new_n8632, new_n8633, new_n8634, new_n8635, new_n8636,
    new_n8637, new_n8638, new_n8639, new_n8640, new_n8641, new_n8642,
    new_n8643, new_n8644, new_n8645, new_n8646, new_n8647, new_n8648,
    new_n8649, new_n8650, new_n8651, new_n8652, new_n8653, new_n8654,
    new_n8655, new_n8656, new_n8657, new_n8658, new_n8659, new_n8660,
    new_n8661, new_n8662, new_n8663, new_n8664, new_n8665_1, new_n8666,
    new_n8667, new_n8668, new_n8669, new_n8670, new_n8671, new_n8672,
    new_n8673, new_n8674, new_n8675, new_n8676, new_n8677, new_n8678,
    new_n8679, new_n8680, new_n8681, new_n8682, new_n8683, new_n8684,
    new_n8685, new_n8686, new_n8687, new_n8688, new_n8689, new_n8690,
    new_n8691, new_n8692, new_n8693, new_n8694, new_n8695, new_n8696,
    new_n8697, new_n8698, new_n8699, new_n8700, new_n8701, new_n8702,
    new_n8703, new_n8704, new_n8705, new_n8706, new_n8707, new_n8708,
    new_n8709, new_n8710, new_n8711, new_n8712, new_n8713, new_n8714,
    new_n8715, new_n8716, new_n8717_1, new_n8718, new_n8719, new_n8720,
    new_n8721, new_n8722, new_n8723, new_n8724, new_n8725, new_n8726,
    new_n8727, new_n8728, new_n8729, new_n8730, new_n8731, new_n8732,
    new_n8733, new_n8734, new_n8735, new_n8736, new_n8737, new_n8738,
    new_n8739, new_n8740, new_n8741, new_n8742, new_n8743, new_n8744,
    new_n8745, new_n8746, new_n8747, new_n8748, new_n8749, new_n8750,
    new_n8751, new_n8752, new_n8753, new_n8754, new_n8755, new_n8756,
    new_n8757, new_n8758, new_n8759_1, new_n8760, new_n8761, new_n8762,
    new_n8763, new_n8764, new_n8765, new_n8766, new_n8767, new_n8768,
    new_n8769, new_n8770, new_n8771, new_n8772, new_n8773, new_n8774,
    new_n8775, new_n8776, new_n8777, new_n8778, new_n8779, new_n8780,
    new_n8781, new_n8782, new_n8783, new_n8784, new_n8785, new_n8786,
    new_n8787, new_n8788, new_n8789, new_n8790, new_n8791, new_n8792,
    new_n8793, new_n8794, new_n8795, new_n8796, new_n8797, new_n8798,
    new_n8799, new_n8800, new_n8801, new_n8802, new_n8803, new_n8804,
    new_n8805, new_n8806, new_n8807, new_n8808, new_n8809, new_n8810,
    new_n8811, new_n8812, new_n8813, new_n8814, new_n8815, new_n8816,
    new_n8817, new_n8818, new_n8819_1, new_n8820, new_n8821, new_n8822,
    new_n8823, new_n8824, new_n8825, new_n8826, new_n8827, new_n8828,
    new_n8829, new_n8830, new_n8831, new_n8832, new_n8833, new_n8834,
    new_n8835, new_n8836, new_n8837, new_n8838, new_n8839, new_n8840,
    new_n8841, new_n8842, new_n8843, new_n8844, new_n8845, new_n8846,
    new_n8847, new_n8848, new_n8849, new_n8850, new_n8851, new_n8852,
    new_n8853, new_n8854, new_n8855, new_n8856, new_n8857, new_n8858,
    new_n8859, new_n8860, new_n8861, new_n8862, new_n8863, new_n8864,
    new_n8865, new_n8866, new_n8867, new_n8868, new_n8869, new_n8870,
    new_n8871, new_n8872, new_n8873, new_n8874, new_n8875, new_n8876,
    new_n8877, new_n8878, new_n8879, new_n8880, new_n8881, new_n8882,
    new_n8883, new_n8884, new_n8885, new_n8886, new_n8887, new_n8888,
    new_n8889, new_n8890, new_n8891, new_n8892, new_n8893, new_n8894,
    new_n8895, new_n8896, new_n8897, new_n8898, new_n8899, new_n8900,
    new_n8901, new_n8902, new_n8903, new_n8904, new_n8905, new_n8906,
    new_n8907, new_n8908, new_n8909, new_n8910, new_n8911, new_n8912,
    new_n8913, new_n8914, new_n8915, new_n8916, new_n8917, new_n8918,
    new_n8919, new_n8920, new_n8921, new_n8922, new_n8923, new_n8924,
    new_n8925, new_n8926, new_n8927, new_n8928, new_n8929, new_n8930,
    new_n8931, new_n8932, new_n8933, new_n8934, new_n8935, new_n8936,
    new_n8937, new_n8938, new_n8939, new_n8940, new_n8941, new_n8942,
    new_n8943, new_n8944, new_n8945, new_n8946, new_n8947, new_n8948,
    new_n8949, new_n8950, new_n8951, new_n8952, new_n8953, new_n8954,
    new_n8955, new_n8956, new_n8957, new_n8958, new_n8959, new_n8960,
    new_n8961, new_n8962, new_n8963, new_n8964, new_n8965, new_n8966,
    new_n8967, new_n8968, new_n8969, new_n8970, new_n8971, new_n8972,
    new_n8973, new_n8974, new_n8975, new_n8976, new_n8977, new_n8978,
    new_n8979, new_n8980, new_n8981, new_n8982, new_n8983, new_n8984,
    new_n8985, new_n8986, new_n8987, new_n8988, new_n8989, new_n8990,
    new_n8991, new_n8992, new_n8993, new_n8994, new_n8995, new_n8996,
    new_n8997, new_n8998, new_n8999, new_n9000, new_n9001, new_n9002,
    new_n9003, new_n9004, new_n9005, new_n9006, new_n9007, new_n9008,
    new_n9009, new_n9010, new_n9011, new_n9012, new_n9013, new_n9014,
    new_n9015, new_n9016, new_n9017, new_n9018, new_n9019, new_n9020,
    new_n9021, new_n9022, new_n9023, new_n9024, new_n9025, new_n9026,
    new_n9027, new_n9028, new_n9029, new_n9030, new_n9031, new_n9032,
    new_n9033, new_n9034, new_n9035, new_n9036, new_n9037, new_n9038,
    new_n9039, new_n9040, new_n9041, new_n9042, new_n9043, new_n9044,
    new_n9045, new_n9046, new_n9047, new_n9048, new_n9049, new_n9050,
    new_n9051, new_n9052, new_n9053, new_n9054, new_n9055, new_n9056,
    new_n9057, new_n9058, new_n9059, new_n9060, new_n9061, new_n9062,
    new_n9063, new_n9064, new_n9065, new_n9066, new_n9067, new_n9068,
    new_n9069, new_n9070, new_n9071, new_n9072, new_n9073, new_n9074,
    new_n9075, new_n9076, new_n9077, new_n9078, new_n9079, new_n9080_1,
    new_n9081, new_n9082, new_n9083, new_n9084, new_n9085, new_n9086,
    new_n9087, new_n9088, new_n9089, new_n9090, new_n9091, new_n9092,
    new_n9093, new_n9094, new_n9095, new_n9096, new_n9097, new_n9098,
    new_n9099, new_n9100, new_n9101, new_n9102, new_n9103, new_n9104,
    new_n9105, new_n9106, new_n9107, new_n9108, new_n9109, new_n9110,
    new_n9111_1, new_n9112, new_n9113, new_n9114, new_n9115, new_n9116,
    new_n9117, new_n9118, new_n9119, new_n9120, new_n9121, new_n9122,
    new_n9123, new_n9124, new_n9125, new_n9126, new_n9127, new_n9128,
    new_n9129, new_n9130, new_n9131, new_n9132, new_n9133, new_n9134,
    new_n9135, new_n9136, new_n9137_1, new_n9138, new_n9139, new_n9140,
    new_n9141, new_n9142, new_n9143, new_n9144, new_n9145, new_n9146,
    new_n9147, new_n9148, new_n9149, new_n9150, new_n9151, new_n9152,
    new_n9153, new_n9154, new_n9155, new_n9156, new_n9157, new_n9158,
    new_n9159, new_n9160, new_n9161, new_n9162, new_n9163, new_n9164,
    new_n9165, new_n9166, new_n9167, new_n9168, new_n9169, new_n9170,
    new_n9171, new_n9172, new_n9173, new_n9174, new_n9175, new_n9176,
    new_n9177, new_n9178, new_n9179, new_n9180, new_n9181, new_n9182,
    new_n9183, new_n9184, new_n9185, new_n9186, new_n9187, new_n9188,
    new_n9189_1, new_n9190, new_n9191, new_n9192, new_n9193, new_n9194,
    new_n9195_1, new_n9196, new_n9197, new_n9198, new_n9199, new_n9200,
    new_n9201, new_n9202, new_n9203, new_n9204, new_n9205, new_n9206,
    new_n9207, new_n9208, new_n9209, new_n9210, new_n9211, new_n9212,
    new_n9213, new_n9214, new_n9215, new_n9216, new_n9217, new_n9218,
    new_n9219, new_n9220, new_n9221, new_n9222, new_n9223, new_n9224,
    new_n9225, new_n9226, new_n9227, new_n9228, new_n9229, new_n9230,
    new_n9231, new_n9232, new_n9233, new_n9234, new_n9235, new_n9236,
    new_n9237, new_n9238, new_n9239, new_n9240, new_n9241_1, new_n9242,
    new_n9243, new_n9244, new_n9245, new_n9246, new_n9247, new_n9248,
    new_n9249, new_n9250, new_n9251, new_n9252, new_n9253, new_n9254,
    new_n9255, new_n9256, new_n9257, new_n9258, new_n9259, new_n9260,
    new_n9261, new_n9262, new_n9263, new_n9264, new_n9265, new_n9266,
    new_n9267, new_n9268, new_n9269, new_n9270, new_n9271, new_n9272,
    new_n9273, new_n9274, new_n9275, new_n9276, new_n9277, new_n9278,
    new_n9279, new_n9280, new_n9281, new_n9282, new_n9283, new_n9284,
    new_n9285, new_n9286, new_n9287, new_n9288, new_n9289, new_n9290,
    new_n9291, new_n9292, new_n9293, new_n9294, new_n9295, new_n9296,
    new_n9297, new_n9298, new_n9299, new_n9300, new_n9301, new_n9302,
    new_n9303, new_n9304, new_n9305, new_n9306, new_n9307, new_n9308,
    new_n9309, new_n9310, new_n9311, new_n9312, new_n9313, new_n9314,
    new_n9315, new_n9316, new_n9317, new_n9318, new_n9319, new_n9320,
    new_n9321, new_n9322, new_n9323, new_n9324, new_n9325, new_n9326,
    new_n9327, new_n9328, new_n9329, new_n9330, new_n9331, new_n9332,
    new_n9333, new_n9334, new_n9335, new_n9336, new_n9337, new_n9338,
    new_n9339, new_n9340, new_n9341, new_n9342, new_n9343, new_n9346,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371,
    new_n9372, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380, new_n9381, new_n9382, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387_1, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9392, new_n9393, new_n9394, new_n9395,
    new_n9396, new_n9397, new_n9398, new_n9399, new_n9400_1, new_n9401,
    new_n9402, new_n9403, new_n9404, new_n9405, new_n9406, new_n9407,
    new_n9408, new_n9409, new_n9410, new_n9411, new_n9412, new_n9413,
    new_n9414, new_n9415, new_n9416, new_n9417, new_n9418, new_n9419,
    new_n9420, new_n9421, new_n9422, new_n9423, new_n9424, new_n9425,
    new_n9426, new_n9427, new_n9428, new_n9429, new_n9430, new_n9431,
    new_n9432, new_n9433, new_n9434, new_n9435, new_n9436, new_n9437,
    new_n9438, new_n9439, new_n9440, new_n9441, new_n9442, new_n9443,
    new_n9444, new_n9445, new_n9446, new_n9447, new_n9448, new_n9449,
    new_n9450, new_n9451, new_n9452, new_n9453, new_n9454, new_n9455,
    new_n9456, new_n9457_1, new_n9458, new_n9459, new_n9460, new_n9461,
    new_n9462, new_n9463, new_n9464, new_n9465, new_n9466, new_n9467,
    new_n9468, new_n9469, new_n9470, new_n9471, new_n9472, new_n9473,
    new_n9474, new_n9475, new_n9476, new_n9477, new_n9478, new_n9479,
    new_n9480, new_n9481, new_n9482, new_n9483, new_n9484, new_n9485,
    new_n9486, new_n9487, new_n9488, new_n9489, new_n9490, new_n9491,
    new_n9492, new_n9493, new_n9494, new_n9495, new_n9496, new_n9497,
    new_n9498, new_n9499, new_n9500, new_n9501, new_n9502, new_n9503,
    new_n9504, new_n9505, new_n9506, new_n9507, new_n9508, new_n9509,
    new_n9510, new_n9511, new_n9512, new_n9513, new_n9514, new_n9515,
    new_n9516, new_n9517, new_n9518, new_n9519, new_n9520, new_n9521,
    new_n9522, new_n9523, new_n9524, new_n9525, new_n9526, new_n9527,
    new_n9528, new_n9529, new_n9530, new_n9531, new_n9532, new_n9533,
    new_n9534, new_n9535, new_n9536, new_n9537, new_n9538, new_n9539,
    new_n9540, new_n9541, new_n9542, new_n9543, new_n9544, new_n9545,
    new_n9546, new_n9547, new_n9548, new_n9549, new_n9550, new_n9551,
    new_n9552, new_n9553, new_n9554, new_n9555, new_n9556, new_n9557,
    new_n9558, new_n9559, new_n9560, new_n9561, new_n9562, new_n9563,
    new_n9564, new_n9565, new_n9566, new_n9567, new_n9568, new_n9569,
    new_n9570, new_n9571_1, new_n9572, new_n9573, new_n9574, new_n9575,
    new_n9576, new_n9577, new_n9578_1, new_n9579, new_n9580, new_n9581,
    new_n9582, new_n9583_1, new_n9584, new_n9585, new_n9586, new_n9587,
    new_n9588, new_n9589, new_n9590, new_n9591, new_n9592, new_n9593,
    new_n9594, new_n9595, new_n9596, new_n9597, new_n9598, new_n9599,
    new_n9600, new_n9601, new_n9602, new_n9603, new_n9604, new_n9605,
    new_n9606, new_n9607, new_n9608, new_n9609, new_n9610, new_n9611,
    new_n9612, new_n9613, new_n9614, new_n9615, new_n9616, new_n9617,
    new_n9618, new_n9619, new_n9620, new_n9621, new_n9622, new_n9623,
    new_n9624, new_n9625, new_n9626, new_n9627, new_n9628, new_n9629,
    new_n9630, new_n9631, new_n9632, new_n9633, new_n9634, new_n9635,
    new_n9636, new_n9637_1, new_n9638, new_n9639, new_n9640_1, new_n9641,
    new_n9642, new_n9643, new_n9644, new_n9645, new_n9646, new_n9647,
    new_n9648, new_n9649, new_n9650, new_n9651, new_n9652, new_n9653,
    new_n9654, new_n9655, new_n9656, new_n9657, new_n9658, new_n9659,
    new_n9660, new_n9661, new_n9662, new_n9663, new_n9664, new_n9665,
    new_n9666, new_n9667, new_n9668, new_n9669, new_n9670, new_n9671,
    new_n9672, new_n9673, new_n9674, new_n9675, new_n9676, new_n9677,
    new_n9678, new_n9679, new_n9680, new_n9681, new_n9682, new_n9683,
    new_n9684, new_n9685, new_n9686, new_n9687, new_n9688, new_n9689,
    new_n9690, new_n9691, new_n9692, new_n9693, new_n9694, new_n9695,
    new_n9696, new_n9697, new_n9698, new_n9699, new_n9700, new_n9701,
    new_n9702, new_n9703, new_n9704, new_n9705, new_n9706_1, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9711, new_n9712, new_n9713,
    new_n9714, new_n9715, new_n9716, new_n9717, new_n9718, new_n9719,
    new_n9720, new_n9721, new_n9722, new_n9723, new_n9724, new_n9725_1,
    new_n9726, new_n9727, new_n9728, new_n9729, new_n9730, new_n9731,
    new_n9732, new_n9733, new_n9734, new_n9735, new_n9736, new_n9737,
    new_n9738, new_n9739, new_n9740, new_n9741, new_n9742, new_n9743,
    new_n9744, new_n9745, new_n9746, new_n9747, new_n9748, new_n9749,
    new_n9750, new_n9751, new_n9752, new_n9753, new_n9754, new_n9755,
    new_n9756_1, new_n9757, new_n9758, new_n9759, new_n9760, new_n9761,
    new_n9762, new_n9763_1, new_n9764, new_n9765, new_n9766, new_n9767_1,
    new_n9768, new_n9769, new_n9770, new_n9771, new_n9772, new_n9773,
    new_n9774, new_n9775, new_n9776, new_n9777, new_n9778, new_n9779,
    new_n9780, new_n9781, new_n9782, new_n9783, new_n9784, new_n9785,
    new_n9786, new_n9787, new_n9788, new_n9789, new_n9790, new_n9791,
    new_n9792, new_n9793, new_n9794, new_n9795, new_n9796, new_n9797,
    new_n9798, new_n9799, new_n9800, new_n9801, new_n9802, new_n9803,
    new_n9804, new_n9805, new_n9806, new_n9807, new_n9808, new_n9809,
    new_n9810, new_n9811, new_n9812, new_n9813, new_n9814, new_n9815,
    new_n9816, new_n9817, new_n9818, new_n9819, new_n9820_1, new_n9821,
    new_n9822, new_n9823, new_n9824, new_n9825, new_n9826, new_n9827,
    new_n9828, new_n9829, new_n9830, new_n9831, new_n9832, new_n9833,
    new_n9834, new_n9835, new_n9836, new_n9837, new_n9838, new_n9839,
    new_n9840, new_n9841, new_n9842, new_n9843, new_n9844, new_n9845,
    new_n9846, new_n9847, new_n9848, new_n9849, new_n9850, new_n9851,
    new_n9852, new_n9853, new_n9854, new_n9855, new_n9856, new_n9857,
    new_n9858, new_n9859, new_n9860, new_n9861, new_n9862, new_n9863,
    new_n9864, new_n9865, new_n9866, new_n9867, new_n9868, new_n9869,
    new_n9870, new_n9871, new_n9872, new_n9873, new_n9874, new_n9875,
    new_n9876, new_n9877, new_n9878, new_n9879, new_n9880, new_n9881,
    new_n9882, new_n9883, new_n9884, new_n9885, new_n9886, new_n9887,
    new_n9888, new_n9889, new_n9890, new_n9891, new_n9892, new_n9893,
    new_n9894, new_n9895, new_n9896, new_n9897, new_n9898, new_n9899,
    new_n9900, new_n9901, new_n9902, new_n9903, new_n9904, new_n9905,
    new_n9906, new_n9907, new_n9908, new_n9909, new_n9910, new_n9911,
    new_n9912, new_n9913, new_n9914, new_n9915, new_n9916, new_n9917,
    new_n9918, new_n9919, new_n9920_1, new_n9921, new_n9922, new_n9923,
    new_n9924, new_n9925, new_n9926, new_n9927, new_n9928, new_n9929,
    new_n9930, new_n9931, new_n9932, new_n9933, new_n9934, new_n9935,
    new_n9936, new_n9937, new_n9938_1, new_n9939, new_n9940, new_n9941,
    new_n9942, new_n9943, new_n9944, new_n9945, new_n9946, new_n9947,
    new_n9948, new_n9949, new_n9950, new_n9951, new_n9952, new_n9953,
    new_n9954, new_n9955, new_n9956_1, new_n9957, new_n9958, new_n9959,
    new_n9960, new_n9961, new_n9962, new_n9963, new_n9964, new_n9965,
    new_n9966, new_n9967, new_n9968, new_n9969, new_n9970, new_n9971,
    new_n9972, new_n9973, new_n9974, new_n9975, new_n9976, new_n9977,
    new_n9978, new_n9979, new_n9980, new_n9981, new_n9982, new_n9983,
    new_n9984, new_n9985, new_n9986, new_n9987, new_n9988, new_n9989,
    new_n9990, new_n9991, new_n9992, new_n9993, new_n9994, new_n9995,
    new_n9996, new_n9997, new_n9998, new_n9999, new_n10000, new_n10001,
    new_n10002, new_n10003, new_n10004, new_n10005, new_n10006, new_n10007,
    new_n10008, new_n10009, new_n10010, new_n10011, new_n10012, new_n10013,
    new_n10014, new_n10015, new_n10016, new_n10017, new_n10018, new_n10019,
    new_n10020, new_n10021, new_n10022_1, new_n10023, new_n10024,
    new_n10025, new_n10026, new_n10027, new_n10028, new_n10029, new_n10030,
    new_n10031, new_n10032, new_n10033, new_n10034, new_n10035, new_n10036,
    new_n10037, new_n10038, new_n10039, new_n10040, new_n10041, new_n10042,
    new_n10043, new_n10044, new_n10045, new_n10046, new_n10047, new_n10048,
    new_n10049, new_n10050, new_n10051, new_n10052, new_n10053, new_n10054,
    new_n10055, new_n10056, new_n10057, new_n10058, new_n10059, new_n10060,
    new_n10061, new_n10062, new_n10063, new_n10064, new_n10065, new_n10066,
    new_n10067, new_n10068, new_n10069, new_n10070, new_n10071, new_n10072,
    new_n10073, new_n10074, new_n10075, new_n10076, new_n10077, new_n10078,
    new_n10079, new_n10080, new_n10081, new_n10082, new_n10083, new_n10084,
    new_n10085, new_n10086, new_n10087, new_n10088, new_n10089, new_n10090,
    new_n10091, new_n10092, new_n10093, new_n10094, new_n10095, new_n10096,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101, new_n10102,
    new_n10103, new_n10104, new_n10105, new_n10106, new_n10107, new_n10108,
    new_n10109, new_n10110, new_n10111, new_n10112, new_n10113, new_n10114,
    new_n10115, new_n10116, new_n10117, new_n10118, new_n10119, new_n10120,
    new_n10121, new_n10122, new_n10123, new_n10124, new_n10125, new_n10126,
    new_n10127, new_n10128, new_n10129, new_n10130, new_n10131, new_n10132,
    new_n10133, new_n10134, new_n10135, new_n10136, new_n10137, new_n10138,
    new_n10139, new_n10140, new_n10141, new_n10142, new_n10143, new_n10144,
    new_n10145, new_n10146, new_n10147, new_n10148, new_n10149, new_n10150,
    new_n10151, new_n10152, new_n10153, new_n10154, new_n10155, new_n10156,
    new_n10157, new_n10158, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10164, new_n10165, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173,
    new_n10174_1, new_n10175, new_n10176, new_n10177, new_n10178,
    new_n10179, new_n10180, new_n10181, new_n10182, new_n10183, new_n10184,
    new_n10185, new_n10186, new_n10187, new_n10188, new_n10189, new_n10190,
    new_n10191, new_n10192, new_n10193, new_n10194, new_n10195, new_n10196,
    new_n10197, new_n10198, new_n10199, new_n10200, new_n10201, new_n10202,
    new_n10203, new_n10204, new_n10205, new_n10206, new_n10207, new_n10208,
    new_n10209, new_n10210, new_n10211, new_n10212, new_n10213, new_n10214,
    new_n10215, new_n10216, new_n10217_1, new_n10218, new_n10219,
    new_n10220, new_n10221, new_n10222, new_n10223_1, new_n10226,
    new_n10227, new_n10228, new_n10229, new_n10230, new_n10231, new_n10232,
    new_n10233, new_n10234, new_n10235, new_n10236, new_n10237, new_n10238,
    new_n10239, new_n10240, new_n10241, new_n10242, new_n10243, new_n10244,
    new_n10245, new_n10246, new_n10247, new_n10248, new_n10249, new_n10250,
    new_n10251, new_n10252, new_n10253, new_n10254, new_n10255, new_n10256,
    new_n10257, new_n10258, new_n10259, new_n10260, new_n10261, new_n10262,
    new_n10263, new_n10264, new_n10265, new_n10266, new_n10267, new_n10268,
    new_n10269, new_n10270, new_n10271, new_n10272, new_n10273, new_n10274,
    new_n10275, new_n10276, new_n10277, new_n10278_1, new_n10279,
    new_n10280, new_n10281, new_n10282, new_n10283, new_n10284, new_n10285,
    new_n10286, new_n10287, new_n10288, new_n10289, new_n10290, new_n10291,
    new_n10292, new_n10293, new_n10294, new_n10295, new_n10296, new_n10297,
    new_n10298, new_n10299, new_n10300, new_n10301, new_n10302, new_n10303,
    new_n10304, new_n10305, new_n10306, new_n10307, new_n10308, new_n10309,
    new_n10310, new_n10311, new_n10312, new_n10313, new_n10314, new_n10315,
    new_n10316, new_n10317, new_n10318, new_n10319, new_n10320, new_n10321,
    new_n10322, new_n10323, new_n10324, new_n10325, new_n10326,
    new_n10327_1, new_n10328, new_n10329, new_n10330, new_n10331,
    new_n10332, new_n10333, new_n10334, new_n10335, new_n10336, new_n10337,
    new_n10338, new_n10339, new_n10340, new_n10341, new_n10342, new_n10343,
    new_n10344, new_n10345, new_n10346, new_n10347, new_n10348, new_n10349,
    new_n10350, new_n10351, new_n10352, new_n10353, new_n10354, new_n10355,
    new_n10356, new_n10357, new_n10358, new_n10359, new_n10360, new_n10361,
    new_n10362, new_n10363, new_n10364, new_n10365, new_n10366, new_n10367,
    new_n10368, new_n10369, new_n10370, new_n10371, new_n10372, new_n10373,
    new_n10374, new_n10375, new_n10376, new_n10377, new_n10378, new_n10379,
    new_n10380, new_n10381, new_n10382, new_n10383, new_n10384, new_n10385,
    new_n10386, new_n10387, new_n10388, new_n10389, new_n10390,
    new_n10391_1, new_n10392, new_n10393, new_n10394, new_n10395,
    new_n10396, new_n10397, new_n10398, new_n10399, new_n10400, new_n10401,
    new_n10402, new_n10403, new_n10404, new_n10405, new_n10406, new_n10407,
    new_n10408, new_n10409, new_n10410, new_n10411, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420, new_n10421, new_n10422, new_n10423, new_n10424, new_n10425,
    new_n10426, new_n10427, new_n10428, new_n10429, new_n10430, new_n10431,
    new_n10432, new_n10433, new_n10434, new_n10435, new_n10436, new_n10437,
    new_n10438, new_n10439_1, new_n10440, new_n10441, new_n10442,
    new_n10443, new_n10444, new_n10445, new_n10446, new_n10447, new_n10448,
    new_n10449, new_n10450, new_n10451_1, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476_1,
    new_n10477, new_n10478, new_n10479, new_n10480, new_n10481, new_n10482,
    new_n10483, new_n10484, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489, new_n10490, new_n10491, new_n10492, new_n10493, new_n10494,
    new_n10495, new_n10496, new_n10497, new_n10498, new_n10499, new_n10500,
    new_n10501, new_n10502, new_n10503, new_n10504, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510_1, new_n10511,
    new_n10512, new_n10513, new_n10514, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525, new_n10526, new_n10527, new_n10528, new_n10529,
    new_n10530, new_n10531, new_n10532, new_n10533, new_n10534, new_n10535,
    new_n10536, new_n10537, new_n10538, new_n10539, new_n10540, new_n10541,
    new_n10542, new_n10543, new_n10544, new_n10545_1, new_n10546,
    new_n10547_1, new_n10548, new_n10549, new_n10550, new_n10551,
    new_n10552, new_n10553, new_n10554, new_n10555, new_n10556, new_n10557,
    new_n10558, new_n10559, new_n10560, new_n10562, new_n10566, new_n10567,
    new_n10570, new_n10571, new_n10572, new_n10573, new_n10574, new_n10575,
    new_n10576, new_n10577, new_n10578, new_n10579, new_n10580, new_n10581,
    new_n10582, new_n10583, new_n10584, new_n10585, new_n10586, new_n10587,
    new_n10588, new_n10589_1, new_n10590, new_n10591, new_n10592,
    new_n10593, new_n10594, new_n10595, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10606, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611, new_n10612, new_n10613, new_n10614, new_n10615, new_n10616,
    new_n10617, new_n10618, new_n10619, new_n10620, new_n10621, new_n10622,
    new_n10623, new_n10624, new_n10625, new_n10626, new_n10627, new_n10628,
    new_n10629, new_n10630, new_n10631, new_n10632, new_n10633, new_n10634,
    new_n10635, new_n10636, new_n10637, new_n10638, new_n10639, new_n10640,
    new_n10641, new_n10642, new_n10643, new_n10644_1, new_n10645,
    new_n10646, new_n10647, new_n10648, new_n10649, new_n10650, new_n10651,
    new_n10652, new_n10653, new_n10654, new_n10655, new_n10656, new_n10657,
    new_n10658, new_n10659, new_n10660, new_n10661, new_n10662, new_n10663,
    new_n10664, new_n10665, new_n10666, new_n10667, new_n10668, new_n10669,
    new_n10670, new_n10671, new_n10672, new_n10673, new_n10674, new_n10675,
    new_n10676, new_n10677, new_n10678_1, new_n10679, new_n10680,
    new_n10681, new_n10682, new_n10683, new_n10684, new_n10685_1,
    new_n10686, new_n10687, new_n10688, new_n10689, new_n10690, new_n10691,
    new_n10692, new_n10693, new_n10694, new_n10695_1, new_n10696,
    new_n10697, new_n10698, new_n10699, new_n10700, new_n10701, new_n10702,
    new_n10703, new_n10704, new_n10705, new_n10706, new_n10707, new_n10708,
    new_n10709, new_n10710, new_n10711, new_n10712, new_n10713, new_n10714,
    new_n10715, new_n10716, new_n10717, new_n10718, new_n10719, new_n10720,
    new_n10721, new_n10722, new_n10723, new_n10724, new_n10725, new_n10726,
    new_n10727, new_n10728, new_n10729, new_n10730, new_n10731, new_n10732,
    new_n10733, new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739, new_n10740, new_n10741, new_n10742, new_n10743, new_n10744,
    new_n10745, new_n10746, new_n10747, new_n10748, new_n10749, new_n10750,
    new_n10751, new_n10752, new_n10753, new_n10754, new_n10755, new_n10756,
    new_n10757, new_n10758, new_n10759, new_n10760, new_n10761, new_n10762,
    new_n10763, new_n10764, new_n10765, new_n10766, new_n10767, new_n10768,
    new_n10769, new_n10770, new_n10771, new_n10772, new_n10773, new_n10774,
    new_n10775, new_n10776, new_n10777, new_n10778, new_n10779, new_n10780,
    new_n10781, new_n10782, new_n10783, new_n10784, new_n10785, new_n10786,
    new_n10787, new_n10788, new_n10789_1, new_n10790, new_n10791,
    new_n10792, new_n10793, new_n10794, new_n10795, new_n10796, new_n10797,
    new_n10798, new_n10799, new_n10800, new_n10801, new_n10802, new_n10803,
    new_n10804, new_n10805, new_n10806, new_n10807, new_n10808, new_n10809,
    new_n10810, new_n10811, new_n10812, new_n10813, new_n10814, new_n10815,
    new_n10816, new_n10817, new_n10818, new_n10819, new_n10820, new_n10821,
    new_n10822, new_n10823, new_n10824, new_n10825, new_n10826, new_n10827,
    new_n10828, new_n10829, new_n10830, new_n10831, new_n10832, new_n10833,
    new_n10834, new_n10835, new_n10836, new_n10837, new_n10838, new_n10839,
    new_n10840, new_n10841, new_n10842, new_n10843, new_n10844, new_n10845,
    new_n10846, new_n10847, new_n10848_1, new_n10849, new_n10850,
    new_n10851_1, new_n10852, new_n10853, new_n10854, new_n10855,
    new_n10856, new_n10857, new_n10858, new_n10859, new_n10860, new_n10861,
    new_n10862, new_n10863, new_n10864, new_n10865, new_n10866, new_n10867,
    new_n10868, new_n10869, new_n10870, new_n10871, new_n10872, new_n10873,
    new_n10874, new_n10875, new_n10876, new_n10877, new_n10878, new_n10879,
    new_n10880, new_n10881, new_n10882, new_n10883, new_n10884, new_n10885,
    new_n10886, new_n10887, new_n10888, new_n10889, new_n10890, new_n10891,
    new_n10892, new_n10893, new_n10894, new_n10895, new_n10896, new_n10897,
    new_n10898_1, new_n10899, new_n10900, new_n10901, new_n10902,
    new_n10903, new_n10904, new_n10905, new_n10906, new_n10907, new_n10908,
    new_n10909, new_n10910, new_n10911, new_n10912, new_n10913_1,
    new_n10914, new_n10915, new_n10916, new_n10917, new_n10918, new_n10919,
    new_n10920, new_n10921, new_n10922, new_n10923, new_n10924, new_n10925,
    new_n10926, new_n10927, new_n10928_1, new_n10929, new_n10930,
    new_n10931, new_n10932, new_n10933, new_n10934, new_n10935, new_n10936,
    new_n10937, new_n10938, new_n10939, new_n10940, new_n10941, new_n10942,
    new_n10943, new_n10944, new_n10945, new_n10946, new_n10947, new_n10948,
    new_n10949_1, new_n10950, new_n10951, new_n10952, new_n10953,
    new_n10954, new_n10955, new_n10956, new_n10957, new_n10958, new_n10959,
    new_n10960, new_n10961, new_n10962, new_n10963, new_n10964,
    new_n10965_1, new_n10966, new_n10967, new_n10968, new_n10969,
    new_n10970, new_n10971, new_n10972, new_n10973, new_n10974, new_n10975,
    new_n10976, new_n10977, new_n10978, new_n10979, new_n10980, new_n10981,
    new_n10982, new_n10983, new_n10984, new_n10985, new_n10986, new_n10987,
    new_n10988, new_n10989, new_n10990_1, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005, new_n11006, new_n11007, new_n11008, new_n11009, new_n11010,
    new_n11011, new_n11012, new_n11013, new_n11014, new_n11015, new_n11016,
    new_n11017, new_n11018, new_n11019, new_n11020, new_n11021, new_n11022,
    new_n11023_1, new_n11024, new_n11025, new_n11026, new_n11027,
    new_n11028, new_n11029, new_n11030, new_n11031, new_n11032, new_n11033,
    new_n11034, new_n11035, new_n11036, new_n11037, new_n11038, new_n11039,
    new_n11040, new_n11041, new_n11042, new_n11043, new_n11044, new_n11045,
    new_n11046, new_n11047, new_n11048, new_n11049, new_n11050, new_n11051,
    new_n11052, new_n11053, new_n11054, new_n11055, new_n11056, new_n11057,
    new_n11058, new_n11059, new_n11060, new_n11061, new_n11062, new_n11063,
    new_n11064, new_n11065, new_n11066, new_n11067, new_n11068, new_n11069,
    new_n11070, new_n11071, new_n11072, new_n11073, new_n11074, new_n11075,
    new_n11076, new_n11077, new_n11078, new_n11079, new_n11080, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11091, new_n11092, new_n11093,
    new_n11094, new_n11096, new_n11098, new_n11100, new_n11101, new_n11102,
    new_n11103, new_n11104, new_n11105, new_n11106, new_n11107, new_n11108,
    new_n11109, new_n11110, new_n11111, new_n11112, new_n11113, new_n11114,
    new_n11115, new_n11116, new_n11117, new_n11118, new_n11119, new_n11120,
    new_n11121, new_n11122, new_n11123, new_n11124, new_n11125, new_n11126,
    new_n11127, new_n11128, new_n11129, new_n11130, new_n11131, new_n11132,
    new_n11133, new_n11134, new_n11135, new_n11136, new_n11137, new_n11138,
    new_n11139, new_n11140, new_n11141, new_n11142, new_n11143, new_n11144,
    new_n11145, new_n11146, new_n11147, new_n11148, new_n11149, new_n11150,
    new_n11151, new_n11152, new_n11153_1, new_n11154, new_n11155,
    new_n11156, new_n11157, new_n11158, new_n11159, new_n11160, new_n11161,
    new_n11162, new_n11163, new_n11164, new_n11165, new_n11166, new_n11167,
    new_n11168, new_n11169, new_n11170, new_n11171, new_n11172, new_n11173,
    new_n11174, new_n11175, new_n11176, new_n11177, new_n11178, new_n11179,
    new_n11180, new_n11181, new_n11182, new_n11183, new_n11184, new_n11185,
    new_n11186, new_n11187, new_n11188, new_n11189, new_n11190, new_n11191,
    new_n11192, new_n11193, new_n11194, new_n11195, new_n11196, new_n11197,
    new_n11198, new_n11199, new_n11200, new_n11201, new_n11202, new_n11203,
    new_n11204, new_n11205, new_n11206, new_n11207, new_n11208, new_n11209,
    new_n11210, new_n11211, new_n11212, new_n11213, new_n11214, new_n11215,
    new_n11216_1, new_n11217, new_n11218, new_n11219, new_n11220,
    new_n11221, new_n11222_1, new_n11223, new_n11224, new_n11225,
    new_n11226, new_n11227, new_n11228, new_n11229, new_n11230, new_n11231,
    new_n11232, new_n11233, new_n11234, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245, new_n11246, new_n11247, new_n11248, new_n11249,
    new_n11250, new_n11251, new_n11252, new_n11253, new_n11254, new_n11256,
    new_n11257_1, new_n11258, new_n11259, new_n11260, new_n11261,
    new_n11262, new_n11263, new_n11264, new_n11265, new_n11266, new_n11267,
    new_n11268, new_n11269, new_n11270, new_n11271, new_n11272, new_n11273,
    new_n11274, new_n11275, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290, new_n11291,
    new_n11292, new_n11293, new_n11294, new_n11295, new_n11296_1,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301, new_n11302,
    new_n11303, new_n11304, new_n11305, new_n11306, new_n11307, new_n11308,
    new_n11309, new_n11310, new_n11311_1, new_n11312, new_n11313,
    new_n11314, new_n11315, new_n11316, new_n11317, new_n11318, new_n11319,
    new_n11320, new_n11321, new_n11322, new_n11323, new_n11324, new_n11325,
    new_n11326_1, new_n11327, new_n11328, new_n11329, new_n11330,
    new_n11331, new_n11332, new_n11333, new_n11334, new_n11335, new_n11336,
    new_n11337, new_n11338, new_n11339, new_n11340, new_n11341, new_n11342,
    new_n11343, new_n11344, new_n11345, new_n11346, new_n11347, new_n11348,
    new_n11349, new_n11350, new_n11351, new_n11352, new_n11353, new_n11354,
    new_n11355, new_n11356, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375, new_n11376, new_n11377, new_n11378,
    new_n11379, new_n11380, new_n11381, new_n11382, new_n11383, new_n11384,
    new_n11385, new_n11386, new_n11387, new_n11388, new_n11389, new_n11390,
    new_n11391, new_n11392, new_n11393, new_n11394, new_n11395, new_n11396,
    new_n11397, new_n11398, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403, new_n11404, new_n11405, new_n11406, new_n11407_1,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11414, new_n11415, new_n11416, new_n11417, new_n11418, new_n11419,
    new_n11420, new_n11421, new_n11422, new_n11423_1, new_n11424,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439, new_n11440, new_n11441, new_n11442,
    new_n11443, new_n11444, new_n11445, new_n11446, new_n11447, new_n11448,
    new_n11449, new_n11450, new_n11451, new_n11452, new_n11453, new_n11454,
    new_n11455, new_n11456, new_n11457, new_n11458, new_n11459, new_n11460,
    new_n11461, new_n11462, new_n11463, new_n11464, new_n11465, new_n11466,
    new_n11467, new_n11468, new_n11469, new_n11470, new_n11471, new_n11472,
    new_n11473, new_n11474, new_n11475, new_n11476, new_n11477,
    new_n11478_1, new_n11479, new_n11480, new_n11481, new_n11482,
    new_n11483, new_n11484, new_n11485, new_n11486, new_n11487, new_n11488,
    new_n11489, new_n11490, new_n11491, new_n11492, new_n11493, new_n11494,
    new_n11495, new_n11496, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503, new_n11504, new_n11505, new_n11506,
    new_n11507, new_n11508, new_n11509, new_n11510, new_n11511, new_n11512,
    new_n11513, new_n11514, new_n11515, new_n11516, new_n11517, new_n11518,
    new_n11519, new_n11520, new_n11521, new_n11522, new_n11523, new_n11524,
    new_n11525, new_n11526, new_n11527, new_n11528, new_n11529, new_n11530,
    new_n11531, new_n11532, new_n11533, new_n11534, new_n11535,
    new_n11536_1, new_n11537, new_n11538, new_n11539, new_n11540,
    new_n11541, new_n11542, new_n11543, new_n11544, new_n11545, new_n11546,
    new_n11547, new_n11548, new_n11549, new_n11550, new_n11551, new_n11552,
    new_n11553, new_n11554, new_n11555, new_n11556, new_n11557, new_n11558,
    new_n11559, new_n11560, new_n11561, new_n11562, new_n11563, new_n11564,
    new_n11565, new_n11566, new_n11567, new_n11568, new_n11569, new_n11570,
    new_n11571, new_n11572, new_n11573, new_n11574, new_n11575, new_n11576,
    new_n11577, new_n11578, new_n11579, new_n11580, new_n11581, new_n11582,
    new_n11583, new_n11584, new_n11585, new_n11586, new_n11587, new_n11588,
    new_n11589, new_n11590, new_n11591, new_n11592, new_n11593, new_n11594,
    new_n11595, new_n11596, new_n11597, new_n11598, new_n11599, new_n11600,
    new_n11601, new_n11602, new_n11603, new_n11604, new_n11605, new_n11606,
    new_n11607, new_n11608, new_n11609, new_n11610, new_n11611, new_n11612,
    new_n11613, new_n11614, new_n11615, new_n11616, new_n11617, new_n11618,
    new_n11619, new_n11620, new_n11621, new_n11622, new_n11623, new_n11624,
    new_n11625, new_n11626, new_n11627, new_n11628, new_n11629, new_n11630,
    new_n11631, new_n11632, new_n11633, new_n11634, new_n11635, new_n11636,
    new_n11637, new_n11638, new_n11639, new_n11640, new_n11641, new_n11642,
    new_n11643, new_n11644, new_n11645, new_n11646, new_n11647, new_n11648,
    new_n11649, new_n11650, new_n11651, new_n11652, new_n11653, new_n11654,
    new_n11655, new_n11656, new_n11657, new_n11658, new_n11659, new_n11660,
    new_n11661, new_n11662_1, new_n11663, new_n11664, new_n11665,
    new_n11666, new_n11667, new_n11668, new_n11669, new_n11670, new_n11671,
    new_n11672, new_n11673, new_n11674, new_n11675, new_n11676, new_n11677,
    new_n11678, new_n11679, new_n11680, new_n11681, new_n11682, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706,
    new_n11707_1, new_n11708, new_n11709, new_n11710, new_n11711,
    new_n11712, new_n11713, new_n11714, new_n11715, new_n11716, new_n11717,
    new_n11718, new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724, new_n11725, new_n11726, new_n11727, new_n11728_1,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736, new_n11737, new_n11738, new_n11739, new_n11740,
    new_n11741, new_n11742, new_n11743, new_n11744, new_n11745, new_n11746,
    new_n11747, new_n11748, new_n11749, new_n11750, new_n11751, new_n11752,
    new_n11753, new_n11754, new_n11755_1, new_n11756, new_n11757_1,
    new_n11758, new_n11759, new_n11760, new_n11761, new_n11762, new_n11763,
    new_n11764, new_n11765, new_n11766, new_n11767, new_n11768, new_n11769,
    new_n11770, new_n11771, new_n11772, new_n11773, new_n11774, new_n11775,
    new_n11776, new_n11777, new_n11778, new_n11779, new_n11780_1,
    new_n11781, new_n11782, new_n11783, new_n11784, new_n11785, new_n11786,
    new_n11787, new_n11788, new_n11789, new_n11790, new_n11791_1,
    new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818, new_n11819, new_n11820,
    new_n11821_1, new_n11822, new_n11823, new_n11824, new_n11825,
    new_n11826, new_n11827, new_n11828, new_n11829, new_n11830, new_n11831,
    new_n11832, new_n11833, new_n11834, new_n11835, new_n11836, new_n11837,
    new_n11838, new_n11839, new_n11840, new_n11841, new_n11842, new_n11843,
    new_n11844, new_n11845, new_n11846, new_n11847, new_n11848, new_n11849,
    new_n11850, new_n11851, new_n11852, new_n11853, new_n11854, new_n11855,
    new_n11856, new_n11857, new_n11858, new_n11859, new_n11860, new_n11861,
    new_n11862, new_n11863, new_n11864, new_n11865, new_n11866, new_n11867,
    new_n11868, new_n11869, new_n11870, new_n11871, new_n11872, new_n11873,
    new_n11874, new_n11875, new_n11876_1, new_n11877_1, new_n11878,
    new_n11879, new_n11880, new_n11881, new_n11882, new_n11883, new_n11884,
    new_n11885, new_n11886, new_n11887, new_n11888, new_n11889, new_n11890,
    new_n11891, new_n11892_1, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898, new_n11899, new_n11900, new_n11901,
    new_n11902, new_n11903, new_n11904, new_n11905, new_n11906, new_n11907,
    new_n11908, new_n11909, new_n11910, new_n11911, new_n11912, new_n11913,
    new_n11914, new_n11915, new_n11916, new_n11917_1, new_n11918,
    new_n11919_1, new_n11920, new_n11921, new_n11922_1, new_n11923,
    new_n11924, new_n11925, new_n11926, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964, new_n11965,
    new_n11966, new_n11967_1, new_n11968, new_n11969, new_n11970,
    new_n11971, new_n11972, new_n11973, new_n11974, new_n11975, new_n11976,
    new_n11977, new_n11978, new_n11979, new_n11980, new_n11981, new_n11982,
    new_n11983, new_n11984, new_n11985, new_n11986, new_n11987, new_n11988,
    new_n11989, new_n11990, new_n11991, new_n11992, new_n11993, new_n11994,
    new_n11995, new_n11996, new_n11997, new_n11998, new_n11999_1,
    new_n12000_1, new_n12001, new_n12002, new_n12003, new_n12004,
    new_n12005_1, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011, new_n12012, new_n12013, new_n12014_1,
    new_n12015, new_n12016, new_n12017, new_n12018, new_n12019,
    new_n12020_1, new_n12021, new_n12022, new_n12023, new_n12024,
    new_n12025_1, new_n12026, new_n12027, new_n12028, new_n12029,
    new_n12030, new_n12031, new_n12032, new_n12033, new_n12034, new_n12035,
    new_n12036, new_n12037, new_n12038, new_n12039, new_n12040, new_n12041,
    new_n12042, new_n12043, new_n12044_1, new_n12045, new_n12046,
    new_n12047, new_n12048, new_n12049, new_n12050, new_n12051, new_n12052,
    new_n12053, new_n12054, new_n12055, new_n12056, new_n12057, new_n12058,
    new_n12059, new_n12060, new_n12061, new_n12062, new_n12063, new_n12064,
    new_n12065, new_n12066, new_n12067, new_n12068, new_n12069_1,
    new_n12070, new_n12071, new_n12072, new_n12073, new_n12074, new_n12075,
    new_n12076_1, new_n12077, new_n12078, new_n12079, new_n12080,
    new_n12081, new_n12082, new_n12083, new_n12084, new_n12085, new_n12086,
    new_n12087, new_n12088, new_n12089, new_n12090, new_n12091, new_n12092,
    new_n12093, new_n12094, new_n12095, new_n12096, new_n12097, new_n12098,
    new_n12099, new_n12100, new_n12101, new_n12102, new_n12103, new_n12104,
    new_n12105, new_n12106, new_n12107, new_n12108, new_n12109, new_n12110,
    new_n12111_1, new_n12112, new_n12113, new_n12114, new_n12115,
    new_n12116, new_n12117, new_n12118, new_n12119, new_n12120, new_n12121,
    new_n12122, new_n12123, new_n12124, new_n12125, new_n12126, new_n12127,
    new_n12128, new_n12129, new_n12130, new_n12131, new_n12132, new_n12133,
    new_n12134, new_n12135, new_n12136, new_n12137, new_n12138, new_n12139,
    new_n12140, new_n12141, new_n12142, new_n12143, new_n12144,
    new_n12145_1, new_n12146, new_n12147, new_n12148, new_n12149,
    new_n12150, new_n12151, new_n12152, new_n12153, new_n12154, new_n12155,
    new_n12156, new_n12157, new_n12158, new_n12159, new_n12160, new_n12161,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12177, new_n12178,
    new_n12181, new_n12184, new_n12186, new_n12188, new_n12189, new_n12190,
    new_n12191, new_n12192, new_n12193, new_n12194, new_n12195, new_n12196,
    new_n12197, new_n12198, new_n12199, new_n12200, new_n12201, new_n12202,
    new_n12203, new_n12204, new_n12205, new_n12206, new_n12207, new_n12208,
    new_n12209, new_n12210, new_n12211, new_n12212, new_n12213, new_n12214,
    new_n12215, new_n12216, new_n12217, new_n12218, new_n12219, new_n12220,
    new_n12221_1, new_n12222, new_n12223, new_n12224, new_n12225,
    new_n12226, new_n12227, new_n12228, new_n12229, new_n12230, new_n12231,
    new_n12232, new_n12233, new_n12234, new_n12235, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247_1, new_n12248,
    new_n12249, new_n12250, new_n12251, new_n12252, new_n12253, new_n12254,
    new_n12255, new_n12256, new_n12257, new_n12258, new_n12259, new_n12260,
    new_n12261, new_n12262, new_n12263, new_n12264, new_n12265, new_n12266,
    new_n12267, new_n12268, new_n12269, new_n12270, new_n12271, new_n12272,
    new_n12273, new_n12274, new_n12275, new_n12276, new_n12277, new_n12278,
    new_n12279, new_n12280, new_n12281, new_n12282, new_n12283, new_n12284,
    new_n12285, new_n12286, new_n12287, new_n12288, new_n12289, new_n12290,
    new_n12291, new_n12292, new_n12293, new_n12294, new_n12295, new_n12296,
    new_n12297, new_n12298, new_n12299_1, new_n12300, new_n12301,
    new_n12302, new_n12303, new_n12304, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315, new_n12316, new_n12317, new_n12318, new_n12319,
    new_n12320, new_n12321, new_n12322, new_n12323, new_n12324, new_n12325,
    new_n12326, new_n12327, new_n12328, new_n12329, new_n12330, new_n12331,
    new_n12332, new_n12333, new_n12334, new_n12335, new_n12336, new_n12337,
    new_n12338, new_n12339, new_n12340, new_n12341, new_n12342, new_n12343,
    new_n12344, new_n12345, new_n12346, new_n12347, new_n12348, new_n12349,
    new_n12350, new_n12351, new_n12352, new_n12353, new_n12354, new_n12355,
    new_n12356, new_n12357, new_n12358, new_n12359, new_n12360, new_n12361,
    new_n12362, new_n12363, new_n12364, new_n12365, new_n12366, new_n12367,
    new_n12368, new_n12369, new_n12370, new_n12371, new_n12372, new_n12373,
    new_n12374, new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380, new_n12381, new_n12382, new_n12383, new_n12384, new_n12385,
    new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391_1, new_n12392, new_n12393, new_n12394, new_n12395,
    new_n12396, new_n12397, new_n12398, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408, new_n12409, new_n12410, new_n12411, new_n12412, new_n12413,
    new_n12414, new_n12415, new_n12416, new_n12417, new_n12418, new_n12419,
    new_n12420, new_n12421, new_n12422, new_n12423, new_n12424, new_n12425,
    new_n12426, new_n12427, new_n12428, new_n12429, new_n12430, new_n12431,
    new_n12432, new_n12433, new_n12434, new_n12435, new_n12436, new_n12437,
    new_n12438, new_n12439, new_n12440, new_n12441, new_n12442, new_n12443,
    new_n12444_1, new_n12445, new_n12446, new_n12447, new_n12448,
    new_n12449, new_n12450, new_n12451, new_n12452, new_n12453, new_n12454,
    new_n12455, new_n12456, new_n12457, new_n12458, new_n12459, new_n12460,
    new_n12461, new_n12462, new_n12463, new_n12464, new_n12465, new_n12466,
    new_n12467, new_n12468, new_n12469, new_n12470, new_n12471, new_n12472,
    new_n12473, new_n12474, new_n12475, new_n12476, new_n12477, new_n12478,
    new_n12479, new_n12480, new_n12481, new_n12482, new_n12483, new_n12484,
    new_n12485, new_n12486, new_n12487, new_n12488, new_n12489_1,
    new_n12490, new_n12491, new_n12492, new_n12493, new_n12494, new_n12495,
    new_n12496, new_n12497, new_n12498, new_n12499, new_n12500, new_n12501,
    new_n12502, new_n12503, new_n12504, new_n12505, new_n12506, new_n12507,
    new_n12508, new_n12509, new_n12510, new_n12511_1, new_n12512,
    new_n12513, new_n12514, new_n12515, new_n12516, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12533, new_n12534, new_n12535, new_n12536, new_n12537, new_n12538,
    new_n12539, new_n12540, new_n12541, new_n12542, new_n12543, new_n12544,
    new_n12545, new_n12546, new_n12547, new_n12548, new_n12549, new_n12550,
    new_n12551, new_n12552, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561, new_n12562,
    new_n12563, new_n12564, new_n12565, new_n12566, new_n12567, new_n12568,
    new_n12569, new_n12570, new_n12571, new_n12572, new_n12573, new_n12574,
    new_n12575, new_n12576, new_n12577, new_n12578, new_n12579, new_n12580,
    new_n12581, new_n12582, new_n12583, new_n12584, new_n12585, new_n12586,
    new_n12587, new_n12588, new_n12589, new_n12590, new_n12591_1,
    new_n12592, new_n12593, new_n12594, new_n12595, new_n12596, new_n12597,
    new_n12598, new_n12599, new_n12600, new_n12601, new_n12602, new_n12603,
    new_n12604, new_n12605, new_n12606, new_n12607, new_n12608, new_n12609,
    new_n12610, new_n12611, new_n12612, new_n12613, new_n12614, new_n12615,
    new_n12616, new_n12617, new_n12618, new_n12619, new_n12620, new_n12621,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626, new_n12627,
    new_n12628, new_n12629, new_n12630, new_n12631, new_n12632, new_n12633,
    new_n12634, new_n12635, new_n12636, new_n12637, new_n12638, new_n12639,
    new_n12640, new_n12641, new_n12642, new_n12643, new_n12644, new_n12645,
    new_n12646, new_n12647, new_n12648_1, new_n12649, new_n12650,
    new_n12651, new_n12652, new_n12653, new_n12654, new_n12655, new_n12656,
    new_n12657, new_n12658, new_n12659, new_n12660, new_n12661, new_n12662,
    new_n12663, new_n12664, new_n12665, new_n12666, new_n12667, new_n12668,
    new_n12669, new_n12670, new_n12671, new_n12672, new_n12673, new_n12674,
    new_n12675, new_n12676, new_n12677, new_n12678, new_n12679, new_n12680,
    new_n12681, new_n12682, new_n12683, new_n12684, new_n12685, new_n12686,
    new_n12687, new_n12688, new_n12689, new_n12690, new_n12691, new_n12692,
    new_n12693, new_n12694, new_n12695, new_n12696, new_n12697, new_n12698,
    new_n12699, new_n12700, new_n12701, new_n12702, new_n12703,
    new_n12704_1, new_n12705_1, new_n12706_1, new_n12707, new_n12708,
    new_n12709_1, new_n12710, new_n12711, new_n12712, new_n12713,
    new_n12714, new_n12715, new_n12716, new_n12717, new_n12718, new_n12719,
    new_n12720_1, new_n12721, new_n12722, new_n12723, new_n12724,
    new_n12725, new_n12726, new_n12727, new_n12728, new_n12729, new_n12730,
    new_n12731, new_n12732, new_n12733, new_n12734, new_n12735, new_n12736,
    new_n12737, new_n12738, new_n12739, new_n12741, new_n12745, new_n12747,
    new_n12749, new_n12751, new_n12753_1, new_n12754, new_n12755,
    new_n12756, new_n12757, new_n12758, new_n12759, new_n12760, new_n12761,
    new_n12762, new_n12763, new_n12764, new_n12765, new_n12766, new_n12767,
    new_n12768, new_n12769, new_n12770, new_n12771, new_n12772, new_n12773,
    new_n12774, new_n12775, new_n12776, new_n12777_1, new_n12778,
    new_n12779, new_n12780, new_n12781, new_n12782, new_n12783, new_n12784,
    new_n12785, new_n12786, new_n12787, new_n12788, new_n12789, new_n12790,
    new_n12791, new_n12792, new_n12793, new_n12794, new_n12795, new_n12796,
    new_n12797, new_n12798, new_n12799, new_n12800, new_n12801, new_n12802,
    new_n12803, new_n12804, new_n12805, new_n12806, new_n12807_1,
    new_n12808, new_n12809, new_n12810, new_n12811, new_n12812, new_n12813,
    new_n12814, new_n12815, new_n12816, new_n12817, new_n12818, new_n12819,
    new_n12820, new_n12821, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826_1, new_n12827, new_n12828, new_n12829, new_n12830,
    new_n12831, new_n12832, new_n12833, new_n12834, new_n12835, new_n12836,
    new_n12837, new_n12838, new_n12839, new_n12840, new_n12841, new_n12842,
    new_n12843, new_n12844, new_n12845, new_n12846, new_n12847, new_n12848,
    new_n12849, new_n12850, new_n12851, new_n12852, new_n12853, new_n12854,
    new_n12855, new_n12856, new_n12857, new_n12858, new_n12859, new_n12860,
    new_n12861, new_n12862, new_n12863, new_n12864, new_n12865, new_n12866,
    new_n12867, new_n12868, new_n12869, new_n12870, new_n12871, new_n12872,
    new_n12873, new_n12874, new_n12875, new_n12876, new_n12877, new_n12878,
    new_n12879, new_n12880, new_n12881, new_n12882, new_n12883, new_n12884,
    new_n12885, new_n12886, new_n12887, new_n12888, new_n12889, new_n12890,
    new_n12891, new_n12892, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900, new_n12901, new_n12902,
    new_n12903, new_n12904, new_n12905, new_n12906, new_n12907, new_n12908,
    new_n12909, new_n12910, new_n12911, new_n12912, new_n12913, new_n12914,
    new_n12915, new_n12916, new_n12917, new_n12918, new_n12919, new_n12920,
    new_n12921, new_n12922, new_n12923, new_n12924, new_n12925_1,
    new_n12926, new_n12927, new_n12928, new_n12929, new_n12930, new_n12931,
    new_n12932, new_n12933, new_n12934, new_n12935, new_n12936, new_n12937,
    new_n12938, new_n12939, new_n12940, new_n12941, new_n12942, new_n12943,
    new_n12944, new_n12945, new_n12946, new_n12947_1, new_n12948,
    new_n12949, new_n12950, new_n12951, new_n12952, new_n12953, new_n12954,
    new_n12955, new_n12956, new_n12957, new_n12958, new_n12959, new_n12960,
    new_n12961, new_n12962, new_n12963, new_n12964, new_n12965, new_n12966,
    new_n12967, new_n12968, new_n12969, new_n12970, new_n12971, new_n12972,
    new_n12973, new_n12974, new_n12975, new_n12976, new_n12977, new_n12978,
    new_n12979, new_n12980, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985, new_n12986, new_n12987, new_n12988, new_n12989, new_n12990,
    new_n12991, new_n12992, new_n12993, new_n12994, new_n12995, new_n12996,
    new_n12997, new_n12998, new_n12999, new_n13000, new_n13001, new_n13002,
    new_n13003, new_n13004, new_n13005, new_n13006, new_n13007, new_n13008,
    new_n13009, new_n13010, new_n13011, new_n13012, new_n13013, new_n13014,
    new_n13015, new_n13016, new_n13017, new_n13018, new_n13019, new_n13020,
    new_n13021, new_n13022, new_n13023, new_n13024, new_n13025, new_n13026,
    new_n13027, new_n13028, new_n13029, new_n13030, new_n13031, new_n13032,
    new_n13033, new_n13034, new_n13035, new_n13036, new_n13037, new_n13038,
    new_n13039, new_n13040, new_n13041, new_n13042, new_n13043, new_n13044,
    new_n13045, new_n13046, new_n13047, new_n13048, new_n13049, new_n13050,
    new_n13051, new_n13052, new_n13053, new_n13054, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073, new_n13074,
    new_n13075, new_n13076, new_n13077, new_n13078, new_n13079, new_n13080,
    new_n13081, new_n13082, new_n13083, new_n13084, new_n13085, new_n13086,
    new_n13087, new_n13088, new_n13089, new_n13090, new_n13091, new_n13092,
    new_n13093, new_n13094, new_n13095, new_n13096, new_n13097, new_n13098,
    new_n13099, new_n13100, new_n13101, new_n13102, new_n13103, new_n13104,
    new_n13105, new_n13106, new_n13107, new_n13108, new_n13109, new_n13110,
    new_n13111, new_n13112, new_n13113, new_n13114, new_n13115, new_n13116,
    new_n13117, new_n13118, new_n13119, new_n13120, new_n13121, new_n13122,
    new_n13123, new_n13124, new_n13125, new_n13129, new_n13131, new_n13134,
    new_n13136, new_n13138, new_n13140, new_n13142, new_n13144, new_n13146,
    new_n13147, new_n13148, new_n13149, new_n13150, new_n13151, new_n13152,
    new_n13153, new_n13154, new_n13155, new_n13156, new_n13157, new_n13158,
    new_n13159, new_n13160, new_n13161, new_n13162, new_n13163, new_n13164,
    new_n13165, new_n13166, new_n13167, new_n13168, new_n13169, new_n13170,
    new_n13171, new_n13172, new_n13173, new_n13174, new_n13175, new_n13176,
    new_n13177, new_n13178, new_n13179, new_n13180, new_n13181, new_n13182,
    new_n13183, new_n13184, new_n13185, new_n13186, new_n13187, new_n13188,
    new_n13189, new_n13190, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198, new_n13199, new_n13200,
    new_n13201, new_n13202, new_n13203, new_n13204, new_n13205, new_n13206,
    new_n13207, new_n13208, new_n13209, new_n13210, new_n13211, new_n13212,
    new_n13213, new_n13214, new_n13215, new_n13216, new_n13217, new_n13218,
    new_n13219, new_n13220, new_n13221, new_n13222, new_n13223, new_n13224,
    new_n13225, new_n13226, new_n13227, new_n13228, new_n13229, new_n13230,
    new_n13231, new_n13232, new_n13233, new_n13234, new_n13235, new_n13236,
    new_n13237, new_n13238, new_n13239, new_n13240, new_n13241, new_n13242,
    new_n13243, new_n13244, new_n13245, new_n13246, new_n13247, new_n13248,
    new_n13249, new_n13250, new_n13251, new_n13252, new_n13253, new_n13254,
    new_n13255, new_n13256, new_n13257, new_n13258, new_n13259, new_n13260,
    new_n13261, new_n13262, new_n13263, new_n13264, new_n13265, new_n13266,
    new_n13267, new_n13268, new_n13269, new_n13270, new_n13271, new_n13272,
    new_n13273, new_n13274, new_n13275, new_n13276, new_n13277, new_n13278,
    new_n13279, new_n13280, new_n13281, new_n13282, new_n13283, new_n13284,
    new_n13285, new_n13286, new_n13287, new_n13288, new_n13289, new_n13290,
    new_n13291, new_n13292, new_n13293, new_n13294, new_n13295, new_n13296,
    new_n13297, new_n13298, new_n13299, new_n13300, new_n13301, new_n13302,
    new_n13303, new_n13304, new_n13305, new_n13306, new_n13307, new_n13308,
    new_n13309, new_n13310, new_n13311, new_n13312, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319, new_n13320,
    new_n13321, new_n13322, new_n13323, new_n13324, new_n13325, new_n13326,
    new_n13327, new_n13328, new_n13329, new_n13330, new_n13331, new_n13332,
    new_n13333, new_n13334, new_n13335, new_n13336, new_n13337, new_n13338,
    new_n13339, new_n13340, new_n13341, new_n13342, new_n13343, new_n13344,
    new_n13345, new_n13347, new_n13348, new_n13350, new_n13351, new_n13352,
    new_n13353, new_n13354, new_n13355, new_n13356, new_n13357, new_n13358,
    new_n13359, new_n13360, new_n13361, new_n13362, new_n13363, new_n13364,
    new_n13365, new_n13366, new_n13367, new_n13368, new_n13369, new_n13370,
    new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13376,
    new_n13377, new_n13378, new_n13379, new_n13380, new_n13381, new_n13382,
    new_n13383, new_n13384, new_n13385, new_n13386, new_n13387, new_n13388,
    new_n13389, new_n13390, new_n13391, new_n13392, new_n13393, new_n13394,
    new_n13395, new_n13396, new_n13397, new_n13398, new_n13399, new_n13400,
    new_n13401, new_n13402, new_n13403, new_n13404, new_n13405, new_n13406,
    new_n13407, new_n13408, new_n13409, new_n13410, new_n13411, new_n13412,
    new_n13413, new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419, new_n13420, new_n13421, new_n13422, new_n13423, new_n13424,
    new_n13425, new_n13426, new_n13427, new_n13428, new_n13429, new_n13430,
    new_n13431, new_n13432, new_n13433, new_n13434, new_n13435, new_n13436,
    new_n13437, new_n13438, new_n13439, new_n13440, new_n13441, new_n13442,
    new_n13443, new_n13444, new_n13445, new_n13446, new_n13447, new_n13448,
    new_n13449, new_n13450, new_n13451, new_n13452, new_n13453, new_n13454,
    new_n13455, new_n13456, new_n13457, new_n13458, new_n13459, new_n13460,
    new_n13461, new_n13462, new_n13463, new_n13464, new_n13465, new_n13466,
    new_n13467, new_n13468, new_n13469, new_n13470, new_n13471, new_n13472,
    new_n13473, new_n13474, new_n13475, new_n13476, new_n13477, new_n13478,
    new_n13479, new_n13480, new_n13481, new_n13482, new_n13483, new_n13484,
    new_n13485, new_n13486, new_n13487, new_n13488, new_n13489, new_n13490,
    new_n13491, new_n13492, new_n13493, new_n13494, new_n13495, new_n13496,
    new_n13497, new_n13498, new_n13499, new_n13500, new_n13501, new_n13502,
    new_n13503, new_n13504, new_n13505, new_n13506, new_n13507, new_n13508,
    new_n13509, new_n13510, new_n13511, new_n13512, new_n13513, new_n13514,
    new_n13515, new_n13516, new_n13517, new_n13518, new_n13519, new_n13520,
    new_n13521, new_n13522, new_n13523, new_n13524, new_n13525, new_n13526,
    new_n13527, new_n13528, new_n13529, new_n13530, new_n13531, new_n13532,
    new_n13533, new_n13534, new_n13535, new_n13536, new_n13537, new_n13538,
    new_n13539, new_n13540, new_n13541, new_n13542, new_n13543, new_n13544,
    new_n13545, new_n13547, new_n13549, new_n13552, new_n13554, new_n13556,
    new_n13558, new_n13560, new_n13563, new_n13565, new_n13566, new_n13567,
    new_n13568, new_n13569, new_n13570, new_n13571, new_n13572, new_n13573,
    new_n13574, new_n13575, new_n13576, new_n13577, new_n13578, new_n13579,
    new_n13580, new_n13581, new_n13582, new_n13583, new_n13584, new_n13585,
    new_n13586, new_n13587, new_n13588, new_n13589, new_n13590, new_n13591,
    new_n13592, new_n13593, new_n13594, new_n13595, new_n13596, new_n13597,
    new_n13598, new_n13599, new_n13600, new_n13601, new_n13602, new_n13603,
    new_n13604, new_n13605, new_n13606, new_n13607, new_n13608, new_n13609,
    new_n13610, new_n13611, new_n13612, new_n13613, new_n13614, new_n13615,
    new_n13616, new_n13617, new_n13618, new_n13619, new_n13620, new_n13621,
    new_n13622, new_n13623, new_n13624, new_n13625, new_n13626, new_n13627,
    new_n13628, new_n13629, new_n13630, new_n13631, new_n13632, new_n13633,
    new_n13634, new_n13635, new_n13636, new_n13637, new_n13638, new_n13639,
    new_n13640, new_n13641, new_n13642, new_n13643, new_n13644, new_n13645,
    new_n13646, new_n13647, new_n13648, new_n13649, new_n13650, new_n13651,
    new_n13652, new_n13653, new_n13654, new_n13655, new_n13656, new_n13657,
    new_n13658, new_n13659, new_n13660, new_n13661, new_n13662, new_n13663,
    new_n13664, new_n13665, new_n13666, new_n13667, new_n13668, new_n13669,
    new_n13670, new_n13671, new_n13672, new_n13673, new_n13674, new_n13675,
    new_n13676, new_n13677, new_n13678, new_n13679, new_n13680, new_n13681,
    new_n13682, new_n13683, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708, new_n13709, new_n13710, new_n13711,
    new_n13712, new_n13713, new_n13714, new_n13715, new_n13716, new_n13717,
    new_n13718, new_n13719, new_n13720, new_n13721, new_n13722, new_n13723,
    new_n13724, new_n13725, new_n13726, new_n13727, new_n13728, new_n13729,
    new_n13730, new_n13731, new_n13732, new_n13733, new_n13734, new_n13735,
    new_n13736, new_n13737, new_n13738, new_n13739, new_n13740, new_n13741,
    new_n13742, new_n13743, new_n13744, new_n13745, new_n13746, new_n13747,
    new_n13748, new_n13749, new_n13750, new_n13751, new_n13752, new_n13753,
    new_n13754, new_n13755, new_n13756, new_n13757, new_n13758, new_n13759,
    new_n13760, new_n13761, new_n13762, new_n13764, new_n13766, new_n13770,
    new_n13772, new_n13773, new_n13776, new_n13781, new_n13782, new_n13783,
    new_n13784, new_n13785, new_n13786, new_n13787, new_n13788, new_n13789,
    new_n13790, new_n13791, new_n13792, new_n13793, new_n13794, new_n13795,
    new_n13796, new_n13797, new_n13798, new_n13799, new_n13800, new_n13801,
    new_n13802, new_n13803, new_n13804, new_n13805, new_n13806, new_n13807,
    new_n13808, new_n13809, new_n13810, new_n13811, new_n13812, new_n13813,
    new_n13814, new_n13815, new_n13816, new_n13817, new_n13818, new_n13819,
    new_n13820, new_n13821, new_n13822, new_n13823, new_n13824, new_n13825,
    new_n13826, new_n13827, new_n13828, new_n13829, new_n13830, new_n13831,
    new_n13832, new_n13833, new_n13834, new_n13835, new_n13836, new_n13837,
    new_n13838, new_n13839, new_n13840, new_n13841, new_n13842, new_n13843,
    new_n13844, new_n13845, new_n13846, new_n13847, new_n13848, new_n13849,
    new_n13850, new_n13851, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912, new_n13913, new_n13914, new_n13915,
    new_n13916, new_n13917, new_n13918, new_n13919, new_n13920, new_n13921,
    new_n13922, new_n13923, new_n13924, new_n13925, new_n13926, new_n13927,
    new_n13928, new_n13929, new_n13930, new_n13931, new_n13932, new_n13933,
    new_n13934, new_n13935, new_n13936, new_n13937, new_n13938, new_n13939,
    new_n13940, new_n13941, new_n13942, new_n13943, new_n13944, new_n13945,
    new_n13946, new_n13947, new_n13948, new_n13949, new_n13950, new_n13951,
    new_n13952, new_n13953, new_n13954, new_n13955, new_n13956, new_n13957,
    new_n13958, new_n13959, new_n13960, new_n13961, new_n13962, new_n13963,
    new_n13964, new_n13965, new_n13966, new_n13967, new_n13968, new_n13969,
    new_n13970, new_n13971, new_n13972, new_n13973, new_n13974, new_n13975,
    new_n13976, new_n13977, new_n13978, new_n13979, new_n13981, new_n13984,
    new_n13988, new_n13990, new_n13994;
nand_4 g00000(new_n377, n6687, n6038);
not_3  g00001(new_n378, new_n377);
nand_4 g00002(new_n379, n8336, n7354);
not_3  g00003(new_n380, new_n379);
nand_4 g00004(new_n381_1, n11222, n8028);
nand_4 g00005(new_n382, n12069, n1564);
not_3  g00006(new_n383, new_n382);
xor_3  g00007(new_n384, new_n383, new_n381_1);
not_3  g00008(new_n385, new_n384);
xor_3  g00009(new_n386, new_n385, new_n380);
xor_3  g00010(n112, new_n386, new_n378);
nand_4 g00011(new_n388, n7436, n1209);
nand_4 g00012(new_n389, n8276, n7500);
nand_4 g00013(new_n390, n9241, n7354);
xnor_3 g00014(new_n391, new_n390, new_n389);
nor_4  g00015(new_n392, new_n391, new_n388);
not_3  g00016(new_n393, new_n388);
not_3  g00017(new_n394, new_n391);
nor_4  g00018(new_n395, new_n394, new_n393);
nor_4  g00019(new_n396, new_n395, new_n392);
nand_4 g00020(new_n397_1, n8276, n7354);
not_3  g00021(new_n398, new_n397_1);
nand_4 g00022(new_n399, n12299, n1209);
not_3  g00023(new_n400, new_n399);
nor_4  g00024(new_n401, new_n400, new_n398);
nand_4 g00025(new_n402, n7500, n7436);
not_3  g00026(new_n403, new_n402);
xnor_3 g00027(new_n404, new_n399, new_n397_1);
nor_4  g00028(new_n405_1, new_n404, new_n403);
nor_4  g00029(new_n406, new_n405_1, new_n401);
xnor_3 g00030(new_n407, new_n406, new_n396);
nand_4 g00031(new_n408, n6776, n4141);
nand_4 g00032(new_n409, n12299, n5105);
xor_3  g00033(new_n410, new_n409, new_n408);
xnor_3 g00034(new_n411, new_n410, new_n407);
nand_4 g00035(new_n412, n6776, n5105);
not_3  g00036(new_n413, new_n412);
nand_4 g00037(new_n414, n7436, n7354);
not_3  g00038(new_n415, new_n414);
nand_4 g00039(new_n416, n6776, n1209);
not_3  g00040(new_n417, new_n416);
nor_4  g00041(new_n418, new_n417, new_n415);
nand_4 g00042(new_n419, n12299, n7500);
not_3  g00043(new_n420, new_n419);
xnor_3 g00044(new_n421, new_n416, new_n414);
nor_4  g00045(new_n422, new_n421, new_n420);
nor_4  g00046(new_n423, new_n422, new_n418);
nand_4 g00047(new_n424, new_n423, new_n413);
xnor_3 g00048(new_n425, new_n423, new_n413);
not_3  g00049(new_n426, new_n425);
xnor_3 g00050(new_n427, new_n404, new_n402);
not_3  g00051(new_n428, new_n427);
nand_4 g00052(new_n429, new_n428, new_n426);
nand_4 g00053(new_n430, new_n429, new_n424);
xnor_3 g00054(new_n431, new_n430, new_n411);
not_3  g00055(new_n432, new_n431);
nand_4 g00056(new_n433, n8759, n4141);
not_3  g00057(new_n434, new_n433);
xnor_3 g00058(new_n435, new_n427, new_n425);
not_3  g00059(new_n436, new_n435);
nand_4 g00060(new_n437, new_n436, new_n434);
not_3  g00061(new_n438, new_n437);
nor_4  g00062(new_n439, new_n436, new_n434);
nor_4  g00063(new_n440, new_n439, new_n438);
nand_4 g00064(new_n441, n8759, n5105);
not_3  g00065(new_n442, new_n441);
nand_4 g00066(new_n443, n12299, n7354);
nand_4 g00067(new_n444, n8759, n1209);
nand_4 g00068(new_n445, new_n444, new_n443);
not_3  g00069(new_n446, new_n445);
nor_4  g00070(new_n447_1, new_n444, new_n443);
nand_4 g00071(new_n448, n7500, n6776);
not_3  g00072(new_n449, new_n448);
nor_4  g00073(new_n450, new_n449, new_n447_1);
nor_4  g00074(new_n451, new_n450, new_n446);
nand_4 g00075(new_n452, new_n451, new_n442);
not_3  g00076(new_n453, new_n452);
xnor_3 g00077(new_n454, new_n451, new_n442);
xnor_3 g00078(new_n455, new_n421, new_n419);
nor_4  g00079(new_n456, new_n455, new_n454);
nor_4  g00080(new_n457, new_n456, new_n453);
not_3  g00081(new_n458, new_n457);
nand_4 g00082(new_n459, new_n458, new_n440);
nand_4 g00083(new_n460, new_n459, new_n437);
nand_4 g00084(new_n461, new_n460, new_n432);
nand_4 g00085(new_n462, new_n406, new_n396);
not_3  g00086(new_n463, new_n462);
nor_4  g00087(new_n464, new_n463, new_n392);
not_3  g00088(new_n465, new_n464);
nand_4 g00089(new_n466, n6776, n4928);
nand_4 g00090(new_n467, n12299, n4141);
nand_4 g00091(new_n468, n8759, n8236);
not_3  g00092(new_n469, new_n468);
xor_3  g00093(new_n470, new_n469, new_n467);
xnor_3 g00094(new_n471, new_n470, new_n466);
xnor_3 g00095(new_n472, new_n471, new_n465);
nor_4  g00096(new_n473, new_n390, new_n389);
not_3  g00097(new_n474, new_n473);
nand_4 g00098(new_n475, n7436, n5105);
xor_3  g00099(new_n476, new_n475, new_n474);
nand_4 g00100(new_n477, n9241, n7500);
not_3  g00101(new_n478, new_n477);
nand_4 g00102(new_n479, n8276, n1209);
nand_4 g00103(new_n480, n10510, n7354);
xor_3  g00104(new_n481, new_n480, new_n479);
xnor_3 g00105(new_n482, new_n481, new_n478);
xnor_3 g00106(new_n483, new_n482, new_n476);
xnor_3 g00107(new_n484, new_n483, new_n472);
not_3  g00108(new_n485, new_n407);
nand_4 g00109(new_n486, new_n410, new_n485);
nor_4  g00110(new_n487, new_n409, new_n408);
not_3  g00111(new_n488, new_n487);
nand_4 g00112(new_n489, new_n430, new_n411);
xnor_3 g00113(new_n490, new_n489, new_n488);
nand_4 g00114(new_n491, new_n490, new_n486);
xnor_3 g00115(new_n492, new_n491, new_n484);
xnor_3 g00116(new_n493, new_n492, new_n461);
nand_4 g00117(new_n494, n8759, n4928);
not_3  g00118(new_n495, new_n494);
xnor_3 g00119(new_n496, new_n460, new_n431);
nand_4 g00120(new_n497, new_n496, new_n495);
xnor_3 g00121(new_n498, new_n455, new_n454);
nand_4 g00122(new_n499, n8759, n7354);
not_3  g00123(new_n500, new_n499);
nor_4  g00124(new_n501, new_n500, new_n448);
nor_4  g00125(new_n502, new_n501, new_n445);
nor_4  g00126(new_n503_1, new_n502, new_n447_1);
nor_4  g00127(new_n504, new_n503_1, new_n448);
not_3  g00128(new_n505, new_n504);
nor_4  g00129(new_n506, new_n505, new_n498);
not_3  g00130(new_n507, new_n506);
xnor_3 g00131(new_n508, new_n458, new_n440);
nor_4  g00132(new_n509, new_n508, new_n507);
xnor_3 g00133(new_n510, new_n496, new_n494);
nand_4 g00134(new_n511, new_n510, new_n509);
nand_4 g00135(new_n512, new_n511, new_n497);
xnor_3 g00136(new_n513, new_n512, new_n493);
nand_4 g00137(new_n514, n12648, n533);
nand_4 g00138(new_n515, n10545, n1512);
nand_4 g00139(new_n516, n7690, n1564);
xnor_3 g00140(new_n517, new_n516, new_n515);
nor_4  g00141(new_n518, new_n517, new_n514);
not_3  g00142(new_n519, new_n514);
not_3  g00143(new_n520, new_n517);
nor_4  g00144(new_n521_1, new_n520, new_n519);
nor_4  g00145(new_n522, new_n521_1, new_n518);
nand_4 g00146(new_n523, n10545, n1564);
not_3  g00147(new_n524, new_n523);
nand_4 g00148(new_n525, n2530, n533);
not_3  g00149(new_n526, new_n525);
nor_4  g00150(new_n527, new_n526, new_n524);
nand_4 g00151(new_n528, n12648, n1512);
not_3  g00152(new_n529, new_n528);
xnor_3 g00153(new_n530, new_n525, new_n523);
nor_4  g00154(new_n531, new_n530, new_n529);
nor_4  g00155(new_n532, new_n531, new_n527);
xnor_3 g00156(new_n533_1, new_n532, new_n522);
nand_4 g00157(new_n534, n8476, n6806);
nand_4 g00158(new_n535, n2802, n2530);
xor_3  g00159(new_n536, new_n535, new_n534);
xnor_3 g00160(new_n537, new_n536, new_n533_1);
nand_4 g00161(new_n538, n8476, n2802);
not_3  g00162(new_n539, new_n538);
nand_4 g00163(new_n540, n12648, n1564);
not_3  g00164(new_n541, new_n540);
nand_4 g00165(new_n542, n8476, n533);
not_3  g00166(new_n543, new_n542);
nor_4  g00167(new_n544, new_n543, new_n541);
nand_4 g00168(new_n545, n2530, n1512);
not_3  g00169(new_n546, new_n545);
xnor_3 g00170(new_n547, new_n542, new_n540);
nor_4  g00171(new_n548, new_n547, new_n546);
nor_4  g00172(new_n549, new_n548, new_n544);
nand_4 g00173(new_n550, new_n549, new_n539);
not_3  g00174(new_n551, new_n550);
nor_4  g00175(new_n552, new_n549, new_n539);
nor_4  g00176(new_n553, new_n552, new_n551);
xnor_3 g00177(new_n554, new_n530, new_n528);
not_3  g00178(new_n555, new_n554);
nand_4 g00179(new_n556, new_n555, new_n553);
nand_4 g00180(new_n557, new_n556, new_n550);
xnor_3 g00181(new_n558, new_n557, new_n537);
nand_4 g00182(new_n559, n6806, n5331);
not_3  g00183(new_n560, new_n559);
xnor_3 g00184(new_n561, new_n555, new_n553);
not_3  g00185(new_n562, new_n561);
nand_4 g00186(new_n563, new_n562, new_n560);
xnor_3 g00187(new_n564, new_n561, new_n560);
nand_4 g00188(new_n565, n5331, n2802);
not_3  g00189(new_n566, new_n565);
nand_4 g00190(new_n567, n2530, n1564);
nand_4 g00191(new_n568, n5331, n533);
nand_4 g00192(new_n569, new_n568, new_n567);
not_3  g00193(new_n570, new_n569);
nor_4  g00194(new_n571, new_n568, new_n567);
nand_4 g00195(new_n572, n8476, n1512);
not_3  g00196(new_n573, new_n572);
nor_4  g00197(new_n574, new_n573, new_n571);
nor_4  g00198(new_n575, new_n574, new_n570);
nand_4 g00199(new_n576, new_n575, new_n566);
not_3  g00200(new_n577, new_n576);
xnor_3 g00201(new_n578, new_n575, new_n566);
xnor_3 g00202(new_n579, new_n547, new_n545);
nor_4  g00203(new_n580, new_n579, new_n578);
nor_4  g00204(new_n581, new_n580, new_n577);
not_3  g00205(new_n582, new_n581);
nand_4 g00206(new_n583, new_n582, new_n564);
nand_4 g00207(new_n584, new_n583, new_n563);
not_3  g00208(new_n585, new_n584);
nor_4  g00209(new_n586, new_n585, new_n558);
not_3  g00210(new_n587, new_n586);
nand_4 g00211(new_n588, new_n532, new_n522);
not_3  g00212(new_n589, new_n588);
nor_4  g00213(new_n590, new_n589, new_n518);
not_3  g00214(new_n591, new_n590);
nand_4 g00215(new_n592, n8476, n5069);
nand_4 g00216(new_n593, n6806, n2530);
nand_4 g00217(new_n594, n12044, n5331);
not_3  g00218(new_n595, new_n594);
xor_3  g00219(new_n596, new_n595, new_n593);
xnor_3 g00220(new_n597, new_n596, new_n592);
xnor_3 g00221(new_n598, new_n597, new_n591);
nor_4  g00222(new_n599, new_n516, new_n515);
nand_4 g00223(new_n600, n12648, n2802);
not_3  g00224(new_n601, new_n600);
xor_3  g00225(new_n602, new_n601, new_n599);
not_3  g00226(new_n603, new_n602);
nand_4 g00227(new_n604, n7690, n1512);
not_3  g00228(new_n605, new_n604);
nand_4 g00229(new_n606, n10545, n533);
nand_4 g00230(new_n607, n3616, n1564);
not_3  g00231(new_n608, new_n607);
xor_3  g00232(new_n609, new_n608, new_n606);
xnor_3 g00233(new_n610, new_n609, new_n605);
xnor_3 g00234(new_n611, new_n610, new_n603);
xnor_3 g00235(new_n612, new_n611, new_n598);
not_3  g00236(new_n613, new_n533_1);
nand_4 g00237(new_n614, new_n536, new_n613);
nor_4  g00238(new_n615_1, new_n535, new_n534);
nand_4 g00239(new_n616, new_n557, new_n537);
not_3  g00240(new_n617, new_n616);
xnor_3 g00241(new_n618, new_n617, new_n615_1);
nand_4 g00242(new_n619, new_n618, new_n614);
xnor_3 g00243(new_n620, new_n619, new_n612);
xnor_3 g00244(new_n621, new_n620, new_n587);
nand_4 g00245(new_n622, n5331, n5069);
xnor_3 g00246(new_n623, new_n585, new_n558);
nand_4 g00247(new_n624, new_n623, new_n622);
xnor_3 g00248(new_n625, new_n579, new_n578);
nand_4 g00249(new_n626, n5331, n1564);
not_3  g00250(new_n627, new_n626);
nor_4  g00251(new_n628, new_n627, new_n572);
not_3  g00252(new_n629, new_n628);
xnor_3 g00253(new_n630, new_n568, new_n567);
nand_4 g00254(new_n631, new_n630, new_n629);
nor_4  g00255(new_n632, new_n631, new_n572);
not_3  g00256(new_n633, new_n632);
nor_4  g00257(new_n634, new_n633, new_n625);
not_3  g00258(new_n635, new_n634);
xnor_3 g00259(new_n636, new_n582, new_n564);
nor_4  g00260(new_n637, new_n636, new_n635);
not_3  g00261(new_n638, new_n637);
xnor_3 g00262(new_n639, new_n623, new_n622);
not_3  g00263(new_n640, new_n639);
nand_4 g00264(new_n641, new_n640, new_n638);
nand_4 g00265(new_n642, new_n641, new_n624);
xnor_3 g00266(new_n643, new_n642, new_n621);
nand_4 g00267(new_n644, n2393, n1980);
nand_4 g00268(new_n645, n8028, n3986);
nand_4 g00269(new_n646, n10848, n5860);
xnor_3 g00270(new_n647, new_n646, new_n645);
nor_4  g00271(new_n648, new_n647, new_n644);
not_3  g00272(new_n649, new_n644);
not_3  g00273(new_n650, new_n647);
nor_4  g00274(new_n651, new_n650, new_n649);
nor_4  g00275(new_n652, new_n651, new_n648);
nand_4 g00276(new_n653, n8028, n5860);
not_3  g00277(new_n654, new_n653);
nand_4 g00278(new_n655, n11892, n1980);
not_3  g00279(new_n656, new_n655);
nor_4  g00280(new_n657, new_n656, new_n654);
nor_4  g00281(new_n658_1, new_n655, new_n653);
nand_4 g00282(new_n659, n10848, n2393);
not_3  g00283(new_n660, new_n659);
nor_4  g00284(new_n661, new_n660, new_n658_1);
nor_4  g00285(new_n662, new_n661, new_n657);
xnor_3 g00286(new_n663, new_n662, new_n652);
nand_4 g00287(new_n664, n12704, n7388);
nand_4 g00288(new_n665, n11892, n7294);
not_3  g00289(new_n666, new_n665);
xor_3  g00290(new_n667, new_n666, new_n664);
xnor_3 g00291(new_n668, new_n667, new_n663);
nand_4 g00292(new_n669, n7388, n7294);
not_3  g00293(new_n670, new_n669);
nand_4 g00294(new_n671_1, n7388, n1980);
not_3  g00295(new_n672, new_n671_1);
nand_4 g00296(new_n673, n8028, n2393);
not_3  g00297(new_n674, new_n673);
nor_4  g00298(new_n675, new_n674, new_n672);
nor_4  g00299(new_n676, new_n673, new_n671_1);
nand_4 g00300(new_n677, n11892, n10848);
not_3  g00301(new_n678, new_n677);
nor_4  g00302(new_n679, new_n678, new_n676);
nor_4  g00303(new_n680, new_n679, new_n675);
and_4  g00304(new_n681, new_n680, new_n670);
xnor_3 g00305(new_n682, new_n680, new_n670);
nor_4  g00306(new_n683, new_n658_1, new_n657);
xnor_3 g00307(new_n684, new_n683, new_n660);
nor_4  g00308(new_n685, new_n684, new_n682);
nor_4  g00309(new_n686, new_n685, new_n681);
xnor_3 g00310(new_n687, new_n686, new_n668);
nand_4 g00311(new_n688, n12704, n7965);
xnor_3 g00312(new_n689, new_n684, new_n682);
nor_4  g00313(new_n690, new_n689, new_n688);
not_3  g00314(new_n691, new_n690);
not_3  g00315(new_n692, new_n688);
not_3  g00316(new_n693, new_n689);
nor_4  g00317(new_n694, new_n693, new_n692);
nor_4  g00318(new_n695, new_n694, new_n690);
nand_4 g00319(new_n696, n7965, n7294);
not_3  g00320(new_n697, new_n696);
nand_4 g00321(new_n698, n11892, n8028);
not_3  g00322(new_n699, new_n698);
nand_4 g00323(new_n700, n7965, n1980);
not_3  g00324(new_n701, new_n700);
nor_4  g00325(new_n702, new_n701, new_n699);
nor_4  g00326(new_n703, new_n700, new_n698);
nand_4 g00327(new_n704, n10848, n7388);
not_3  g00328(new_n705, new_n704);
nor_4  g00329(new_n706, new_n705, new_n703);
nor_4  g00330(new_n707, new_n706, new_n702);
nand_4 g00331(new_n708, new_n707, new_n697);
xnor_3 g00332(new_n709, new_n707, new_n697);
not_3  g00333(new_n710, new_n709);
xnor_3 g00334(new_n711, new_n673, new_n671_1);
xnor_3 g00335(new_n712, new_n711, new_n677);
not_3  g00336(new_n713, new_n712);
nand_4 g00337(new_n714, new_n713, new_n710);
nand_4 g00338(new_n715, new_n714, new_n708);
nand_4 g00339(new_n716, new_n715, new_n695);
nand_4 g00340(new_n717, new_n716, new_n691);
not_3  g00341(new_n718, new_n717);
nor_4  g00342(new_n719, new_n718, new_n687);
not_3  g00343(new_n720, new_n648);
nand_4 g00344(new_n721, new_n662, new_n652);
nand_4 g00345(new_n722, new_n721, new_n720);
nand_4 g00346(new_n723, n7388, n5814);
nand_4 g00347(new_n724, n12704, n11892);
nand_4 g00348(new_n725, n7965, n4903);
not_3  g00349(new_n726, new_n725);
xor_3  g00350(new_n727, new_n726, new_n724);
xnor_3 g00351(new_n728, new_n727, new_n723);
not_3  g00352(new_n729, new_n728);
and_4  g00353(new_n730, new_n729, new_n722);
nor_4  g00354(new_n731, new_n729, new_n722);
nor_4  g00355(new_n732, new_n731, new_n730);
nor_4  g00356(new_n733, new_n646, new_n645);
not_3  g00357(new_n734, new_n733);
nand_4 g00358(new_n735, n7294, n2393);
xor_3  g00359(new_n736, new_n735, new_n734);
nand_4 g00360(new_n737, n10848, n3986);
nand_4 g00361(new_n738, n5860, n1980);
nand_4 g00362(new_n739, n8028, n5857);
not_3  g00363(new_n740, new_n739);
xor_3  g00364(new_n741, new_n740, new_n738);
xnor_3 g00365(new_n742, new_n741, new_n737);
xnor_3 g00366(new_n743, new_n742, new_n736);
xnor_3 g00367(new_n744, new_n743, new_n732);
nor_4  g00368(new_n745, new_n667, new_n663);
not_3  g00369(new_n746, new_n745);
nor_4  g00370(new_n747, new_n665, new_n664);
nor_4  g00371(new_n748, new_n686, new_n668);
xnor_3 g00372(new_n749, new_n748, new_n747);
nand_4 g00373(new_n750, new_n749, new_n746);
xnor_3 g00374(new_n751, new_n750, new_n744);
xnor_3 g00375(new_n752, new_n751, new_n719);
nand_4 g00376(new_n753_1, n7965, n5814);
not_3  g00377(new_n754, new_n753_1);
xnor_3 g00378(new_n755, new_n717, new_n687);
nand_4 g00379(new_n756, new_n755, new_n754);
not_3  g00380(new_n757, new_n755);
nand_4 g00381(new_n758, new_n757, new_n753_1);
xnor_3 g00382(new_n759, new_n712, new_n709);
not_3  g00383(new_n760, new_n703);
nand_4 g00384(new_n761, n8028, n7965);
nand_4 g00385(new_n762, new_n761, new_n705);
nand_4 g00386(new_n763, new_n762, new_n702);
nand_4 g00387(new_n764, new_n763, new_n760);
not_3  g00388(new_n765, new_n764);
nor_4  g00389(new_n766, new_n765, new_n704);
not_3  g00390(new_n767, new_n766);
nor_4  g00391(new_n768, new_n767, new_n759);
not_3  g00392(new_n769, new_n768);
xnor_3 g00393(new_n770, new_n715, new_n695);
nor_4  g00394(new_n771, new_n770, new_n769);
nand_4 g00395(new_n772, new_n771, new_n758);
nand_4 g00396(new_n773, new_n772, new_n756);
xnor_3 g00397(new_n774, new_n773, new_n752);
xnor_3 g00398(new_n775, new_n774, new_n643);
xnor_3 g00399(new_n776, new_n636, new_n635);
not_3  g00400(new_n777, new_n625);
nor_4  g00401(new_n778, new_n632, new_n777);
nor_4  g00402(new_n779, new_n778, new_n634);
not_3  g00403(new_n780, new_n759);
nor_4  g00404(new_n781, new_n766, new_n780);
nor_4  g00405(new_n782, new_n781, new_n768);
nor_4  g00406(new_n783_1, new_n782, new_n779);
not_3  g00407(new_n784, new_n783_1);
not_3  g00408(new_n785, new_n782);
xnor_3 g00409(new_n786, new_n785, new_n779);
nor_4  g00410(new_n787, new_n762, new_n702);
nor_4  g00411(new_n788, new_n787, new_n764);
nand_4 g00412(new_n789, new_n628, new_n569);
nand_4 g00413(new_n790, new_n789, new_n631);
not_3  g00414(new_n791, new_n790);
nand_4 g00415(new_n792, new_n791, new_n788);
not_3  g00416(new_n793, new_n792);
xnor_3 g00417(new_n794, new_n791, new_n788);
not_3  g00418(new_n795, new_n761);
nand_4 g00419(new_n796, new_n795, new_n627);
nand_4 g00420(new_n797, n5331, n1512);
nand_4 g00421(new_n798, n8476, n1564);
xnor_3 g00422(new_n799, new_n798, new_n797);
nor_4  g00423(new_n800, new_n799, new_n796);
xnor_3 g00424(new_n801, new_n799, new_n796);
nand_4 g00425(new_n802, n8028, n7388);
nand_4 g00426(new_n803, n10848, n7965);
xnor_3 g00427(new_n804, new_n803, new_n802);
nor_4  g00428(new_n805, new_n804, new_n801);
nor_4  g00429(new_n806_1, new_n805, new_n800);
nor_4  g00430(new_n807, new_n806_1, new_n794);
nor_4  g00431(new_n808, new_n807, new_n793);
nand_4 g00432(new_n809, new_n808, new_n786);
nand_4 g00433(new_n810, new_n809, new_n784);
nand_4 g00434(new_n811, new_n810, new_n776);
not_3  g00435(new_n812, new_n811);
not_3  g00436(new_n813, new_n770);
nor_4  g00437(new_n814, new_n813, new_n768);
nor_4  g00438(new_n815, new_n814, new_n771);
xnor_3 g00439(new_n816, new_n810, new_n776);
nor_4  g00440(new_n817, new_n816, new_n815);
nor_4  g00441(new_n818, new_n817, new_n812);
xnor_3 g00442(new_n819, new_n639, new_n638);
not_3  g00443(new_n820, new_n819);
nand_4 g00444(new_n821, new_n820, new_n818);
xnor_3 g00445(new_n822, new_n819, new_n818);
nand_4 g00446(new_n823, new_n758, new_n756);
xnor_3 g00447(new_n824, new_n823, new_n771);
nand_4 g00448(new_n825, new_n824, new_n822);
nand_4 g00449(new_n826, new_n825, new_n821);
xnor_3 g00450(new_n827, new_n826, new_n775);
xnor_3 g00451(new_n828, new_n827, new_n513);
not_3  g00452(new_n829, new_n510);
xnor_3 g00453(new_n830, new_n829, new_n509);
xnor_3 g00454(new_n831, new_n508, new_n507);
not_3  g00455(new_n832, new_n498);
nor_4  g00456(new_n833, new_n504, new_n832);
nor_4  g00457(new_n834, new_n833, new_n506);
not_3  g00458(new_n835, new_n834);
xnor_3 g00459(new_n836, new_n761, new_n626);
nor_4  g00460(new_n837_1, new_n836, new_n499);
not_3  g00461(new_n838, new_n837_1);
nand_4 g00462(new_n839, n7354, n6776);
nand_4 g00463(new_n840, n8759, n7500);
xnor_3 g00464(new_n841, new_n840, new_n839);
nand_4 g00465(new_n842, new_n841, new_n838);
xnor_3 g00466(new_n843, new_n804, new_n801);
xnor_3 g00467(new_n844_1, new_n841, new_n837_1);
nand_4 g00468(new_n845, new_n844_1, new_n843);
nand_4 g00469(new_n846, new_n845, new_n842);
not_3  g00470(new_n847, new_n503_1);
not_3  g00471(new_n848, new_n501);
nor_4  g00472(new_n849, new_n848, new_n446);
nor_4  g00473(new_n850, new_n849, new_n847);
not_3  g00474(new_n851, new_n850);
nand_4 g00475(new_n852, new_n851, new_n846);
xnor_3 g00476(new_n853, new_n806_1, new_n794);
xnor_3 g00477(new_n854, new_n850, new_n846);
nand_4 g00478(new_n855, new_n854, new_n853);
nand_4 g00479(new_n856, new_n855, new_n852);
nand_4 g00480(new_n857, new_n856, new_n835);
not_3  g00481(new_n858, new_n808);
xnor_3 g00482(new_n859, new_n858, new_n786);
xnor_3 g00483(new_n860, new_n856, new_n834);
nand_4 g00484(new_n861, new_n860, new_n859);
nand_4 g00485(new_n862, new_n861, new_n857);
nand_4 g00486(new_n863, new_n862, new_n831);
not_3  g00487(new_n864, new_n815);
xnor_3 g00488(new_n865, new_n816, new_n864);
not_3  g00489(new_n866, new_n863);
nor_4  g00490(new_n867, new_n862, new_n831);
nor_4  g00491(new_n868, new_n867, new_n866);
nand_4 g00492(new_n869, new_n868, new_n865);
nand_4 g00493(new_n870, new_n869, new_n863);
not_3  g00494(new_n871, new_n870);
nor_4  g00495(new_n872, new_n871, new_n830);
xnor_3 g00496(new_n873, new_n870, new_n830);
not_3  g00497(new_n874, new_n873);
xnor_3 g00498(new_n875, new_n820, new_n818);
xnor_3 g00499(new_n876, new_n824, new_n875);
nor_4  g00500(new_n877, new_n876, new_n874);
nor_4  g00501(new_n878, new_n877, new_n872);
xnor_3 g00502(new_n879, new_n878, new_n828);
nand_4 g00503(new_n880, n12720, n4312);
not_3  g00504(new_n881, new_n880);
nand_4 g00505(new_n882, n12025, n6038);
nand_4 g00506(new_n883, n12705, n2509);
not_3  g00507(new_n884, new_n883);
xor_3  g00508(new_n885, new_n884, new_n882);
not_3  g00509(new_n886, new_n885);
xor_3  g00510(new_n887, new_n886, new_n881);
nand_4 g00511(new_n888, n12705, n6038);
not_3  g00512(new_n889, new_n888);
nand_4 g00513(new_n890, n12720, n1097);
not_3  g00514(new_n891, new_n890);
nor_4  g00515(new_n892, new_n891, new_n889);
nand_4 g00516(new_n893, n4312, n2509);
not_3  g00517(new_n894, new_n893);
xor_3  g00518(new_n895, new_n891, new_n888);
nor_4  g00519(new_n896, new_n895, new_n894);
nor_4  g00520(new_n897, new_n896, new_n892);
xnor_3 g00521(new_n898, new_n897, new_n887);
nand_4 g00522(new_n899, n2508, n1097);
nand_4 g00523(new_n900, n5964, n2585);
xor_3  g00524(new_n901, new_n900, new_n899);
not_3  g00525(new_n902, new_n901);
nor_4  g00526(new_n903, new_n902, new_n898);
not_3  g00527(new_n904, new_n898);
nor_4  g00528(new_n905, new_n901, new_n904);
nor_4  g00529(new_n906, new_n905, new_n903);
nand_4 g00530(new_n907, n5964, n2508);
not_3  g00531(new_n908, new_n907);
xnor_3 g00532(new_n909, new_n895, new_n893);
not_3  g00533(new_n910, new_n909);
nor_4  g00534(new_n911_1, new_n910, new_n908);
xor_3  g00535(new_n912, new_n910, new_n907);
nand_4 g00536(new_n913, n6038, n4312);
not_3  g00537(new_n914, new_n913);
nand_4 g00538(new_n915, n12720, n5964);
not_3  g00539(new_n916, new_n915);
nor_4  g00540(new_n917, new_n916, new_n914);
nor_4  g00541(new_n918, new_n915, new_n913);
nand_4 g00542(new_n919, n2509, n1097);
not_3  g00543(new_n920, new_n919);
nor_4  g00544(new_n921, new_n920, new_n918);
nor_4  g00545(new_n922, new_n921, new_n917);
nor_4  g00546(new_n923, new_n922, new_n912);
nor_4  g00547(new_n924, new_n923, new_n911_1);
not_3  g00548(new_n925, new_n924);
xnor_3 g00549(new_n926, new_n925, new_n906);
nand_4 g00550(new_n927, n5305, n2585);
not_3  g00551(new_n928, new_n922);
xnor_3 g00552(new_n929, new_n928, new_n912);
nand_4 g00553(new_n930, new_n929, new_n927);
not_3  g00554(new_n931, new_n930);
nor_4  g00555(new_n932, new_n929, new_n927);
nor_4  g00556(new_n933, new_n932, new_n931);
nand_4 g00557(new_n934, n5305, n2508);
nand_4 g00558(new_n935, n6038, n1097);
not_3  g00559(new_n936, new_n935);
nand_4 g00560(new_n937, n12720, n5305);
not_3  g00561(new_n938, new_n937);
nand_4 g00562(new_n939, new_n938, new_n936);
nand_4 g00563(new_n940, new_n937, new_n935);
nand_4 g00564(new_n941, n5964, n2509);
not_3  g00565(new_n942, new_n941);
nand_4 g00566(new_n943, new_n942, new_n940);
nand_4 g00567(new_n944, new_n943, new_n939);
not_3  g00568(new_n945, new_n944);
nor_4  g00569(new_n946, new_n945, new_n934);
xor_3  g00570(new_n947, new_n944, new_n934);
nor_4  g00571(new_n948, new_n918, new_n917);
xor_3  g00572(new_n949, new_n948, new_n919);
nor_4  g00573(new_n950, new_n949, new_n947);
nor_4  g00574(new_n951, new_n950, new_n946);
nand_4 g00575(new_n952, new_n951, new_n933);
nand_4 g00576(new_n953, new_n952, new_n930);
not_3  g00577(new_n954, new_n953);
nand_4 g00578(new_n955, new_n954, new_n926);
nor_4  g00579(new_n956, new_n885, new_n880);
nand_4 g00580(new_n957, new_n897, new_n887);
not_3  g00581(new_n958, new_n957);
nor_4  g00582(new_n959, new_n958, new_n956);
not_3  g00583(new_n960, new_n959);
nand_4 g00584(new_n961, n5964, n4005);
nand_4 g00585(new_n962, n2585, n1097);
nand_4 g00586(new_n963, n12706, n5305);
nand_4 g00587(new_n964, new_n963, new_n962);
not_3  g00588(new_n965, new_n962);
not_3  g00589(new_n966, new_n963);
nand_4 g00590(new_n967, new_n966, new_n965);
and_4  g00591(new_n968, new_n967, new_n964);
xor_3  g00592(new_n969, new_n968, new_n961);
xnor_3 g00593(new_n970, new_n969, new_n960);
nor_4  g00594(new_n971, new_n883, new_n882);
nand_4 g00595(new_n972, n4312, n2508);
not_3  g00596(new_n973, new_n972);
xor_3  g00597(new_n974, new_n973, new_n971);
nand_4 g00598(new_n975, n12025, n2509);
not_3  g00599(new_n976, new_n975);
nand_4 g00600(new_n977, n12720, n12705);
nand_4 g00601(new_n978, n11257, n6038);
not_3  g00602(new_n979, new_n978);
xor_3  g00603(new_n980, new_n979, new_n977);
xnor_3 g00604(new_n981, new_n980, new_n976);
xnor_3 g00605(new_n982, new_n981, new_n974);
not_3  g00606(new_n983, new_n982);
xnor_3 g00607(new_n984, new_n983, new_n970);
nor_4  g00608(new_n985, new_n900, new_n899);
nand_4 g00609(new_n986, new_n924, new_n906);
xnor_3 g00610(new_n987, new_n986, new_n985);
nor_4  g00611(new_n988, new_n987, new_n903);
xnor_3 g00612(new_n989, new_n988, new_n984);
xnor_3 g00613(new_n990, new_n989, new_n955);
nand_4 g00614(new_n991, n5305, n4005);
not_3  g00615(new_n992_1, new_n926);
xnor_3 g00616(new_n993, new_n953, new_n992_1);
nor_4  g00617(new_n994, new_n993, new_n991);
not_3  g00618(new_n995, new_n994);
nand_4 g00619(new_n996_1, new_n993, new_n991);
and_4  g00620(new_n997, new_n940, new_n939);
nand_4 g00621(new_n998, n6038, n5964);
nand_4 g00622(new_n999, n5305, n2509);
nor_4  g00623(new_n1000, new_n999, new_n998);
not_3  g00624(new_n1001, new_n1000);
nor_4  g00625(new_n1002, new_n1001, new_n997);
not_3  g00626(new_n1003, new_n1002);
xnor_3 g00627(new_n1004, new_n949, new_n947);
nor_4  g00628(new_n1005, new_n1004, new_n1003);
xnor_3 g00629(new_n1006, new_n951, new_n933);
nand_4 g00630(new_n1007, new_n1006, new_n1005);
not_3  g00631(new_n1008, new_n1007);
nand_4 g00632(new_n1009, new_n1008, new_n996_1);
nand_4 g00633(new_n1010, new_n1009, new_n995);
xnor_3 g00634(new_n1011, new_n1010, new_n990);
xnor_3 g00635(new_n1012, new_n876, new_n874);
xnor_3 g00636(new_n1013, new_n993, new_n991);
xnor_3 g00637(new_n1014, new_n1013, new_n1008);
nor_4  g00638(new_n1015, new_n1014, new_n1012);
xnor_3 g00639(new_n1016, new_n876, new_n873);
xnor_3 g00640(new_n1017, new_n1013, new_n1007);
nor_4  g00641(new_n1018, new_n1017, new_n1016);
xnor_3 g00642(new_n1019, new_n1006, new_n1005);
xnor_3 g00643(new_n1020_1, new_n868, new_n865);
not_3  g00644(new_n1021, new_n1020_1);
nor_4  g00645(new_n1022, new_n1021, new_n1019);
not_3  g00646(new_n1023, new_n1022);
xnor_3 g00647(new_n1024, new_n1020_1, new_n1019);
not_3  g00648(new_n1025, new_n1004);
xor_3  g00649(new_n1026, new_n1025, new_n1003);
xnor_3 g00650(new_n1027, new_n860, new_n859);
not_3  g00651(new_n1028, new_n1027);
nor_4  g00652(new_n1029, new_n1028, new_n1026);
not_3  g00653(new_n1030, new_n1029);
not_3  g00654(new_n1031, new_n853);
xor_3  g00655(new_n1032, new_n854, new_n1031);
nand_4 g00656(new_n1033, n6038, n5305);
not_3  g00657(new_n1034, new_n1033);
nor_4  g00658(new_n1035, new_n1034, new_n941);
nor_4  g00659(new_n1036, new_n1035, new_n997);
nor_4  g00660(new_n1037, new_n1034, new_n943);
nor_4  g00661(new_n1038, new_n1037, new_n1036);
nor_4  g00662(new_n1039, new_n1038, new_n1032);
not_3  g00663(new_n1040, new_n1032);
xor_3  g00664(new_n1041, new_n1038, new_n1040);
xor_3  g00665(new_n1042, new_n836, new_n499);
not_3  g00666(new_n1043, new_n1042);
nor_4  g00667(new_n1044, new_n1043, new_n1033);
not_3  g00668(new_n1045, new_n1044);
xor_3  g00669(new_n1046, new_n999, new_n998);
not_3  g00670(new_n1047, new_n1046);
nor_4  g00671(new_n1048, new_n1047, new_n1045);
xor_3  g00672(new_n1049, new_n844_1, new_n843);
xor_3  g00673(new_n1050, new_n1047, new_n1044);
nor_4  g00674(new_n1051, new_n1050, new_n1049);
nor_4  g00675(new_n1052, new_n1051, new_n1048);
not_3  g00676(new_n1053, new_n1052);
nor_4  g00677(new_n1054, new_n1053, new_n1041);
nor_4  g00678(new_n1055, new_n1054, new_n1039);
not_3  g00679(new_n1056, new_n1026);
nor_4  g00680(new_n1057, new_n1027, new_n1056);
nor_4  g00681(new_n1058, new_n1057, new_n1029);
nand_4 g00682(new_n1059, new_n1058, new_n1055);
nand_4 g00683(new_n1060, new_n1059, new_n1030);
nand_4 g00684(new_n1061, new_n1060, new_n1024);
nand_4 g00685(new_n1062, new_n1061, new_n1023);
nor_4  g00686(new_n1063, new_n1062, new_n1018);
nor_4  g00687(new_n1064, new_n1063, new_n1015);
nor_4  g00688(new_n1065, new_n1064, new_n1011);
nand_4 g00689(new_n1066, new_n1064, new_n1011);
not_3  g00690(new_n1067_1, new_n1066);
nor_4  g00691(new_n1068, new_n1067_1, new_n1065);
xnor_3 g00692(n226, new_n1068, new_n879);
nand_4 g00693(new_n1070, n5305, n4634);
not_3  g00694(new_n1071, new_n1070);
nand_4 g00695(new_n1072, n10223, n5305);
not_3  g00696(new_n1073, new_n1072);
nand_4 g00697(new_n1074, n7265, n1097);
not_3  g00698(new_n1075, new_n1074);
nor_4  g00699(new_n1076, new_n1075, new_n1073);
nor_4  g00700(new_n1077, new_n1074, new_n1072);
nand_4 g00701(new_n1078, n5964, n2879);
not_3  g00702(new_n1079, new_n1078);
nor_4  g00703(new_n1080, new_n1079, new_n1077);
nor_4  g00704(new_n1081, new_n1080, new_n1076);
nand_4 g00705(new_n1082, new_n1081, new_n1071);
not_3  g00706(new_n1083, new_n1082);
nor_4  g00707(new_n1084, new_n1081, new_n1071);
nor_4  g00708(new_n1085, new_n1084, new_n1083);
nand_4 g00709(new_n1086, n2879, n1097);
not_3  g00710(new_n1087, new_n1086);
nand_4 g00711(new_n1088, n10223, n5964);
nand_4 g00712(new_n1089, n7265, n4312);
xnor_3 g00713(new_n1090, new_n1089, new_n1088);
xnor_3 g00714(new_n1091, new_n1090, new_n1087);
xor_3  g00715(new_n1092, new_n1091, new_n1085);
not_3  g00716(new_n1093, new_n1092);
nand_4 g00717(new_n1094_1, n7265, n5305);
not_3  g00718(new_n1095, new_n1094_1);
nor_4  g00719(new_n1096, new_n1095, new_n1078);
nor_4  g00720(new_n1097_1, new_n1077, new_n1076);
nor_4  g00721(new_n1098, new_n1097_1, new_n1096);
not_3  g00722(new_n1099, new_n1098);
nor_4  g00723(new_n1100, new_n1099, new_n1078);
not_3  g00724(new_n1101, new_n1100);
xor_3  g00725(new_n1102, new_n1101, new_n1093);
nand_4 g00726(new_n1103, n8759, n7946);
nand_4 g00727(new_n1104, n5331, n2558);
nand_4 g00728(new_n1105, n9763, n7965);
xnor_3 g00729(new_n1106, new_n1105, new_n1104);
nor_4  g00730(new_n1107, new_n1106, new_n1103);
not_3  g00731(new_n1108, new_n1107);
nand_4 g00732(new_n1109, n7946, n6776);
nand_4 g00733(new_n1110, n8759, n2024);
xnor_3 g00734(new_n1111, new_n1110, new_n1109);
nor_4  g00735(new_n1112, new_n1111, new_n1108);
not_3  g00736(new_n1113, new_n1112);
nor_4  g00737(new_n1114, new_n1105, new_n1104);
nand_4 g00738(new_n1115, n9111, n7965);
nand_4 g00739(new_n1116, n9763, n7388);
xnor_3 g00740(new_n1117, new_n1116, new_n1115);
not_3  g00741(new_n1118, new_n1117);
xnor_3 g00742(new_n1119, new_n1118, new_n1114);
nand_4 g00743(new_n1120, n5331, n2498);
nand_4 g00744(new_n1121, n8476, n2558);
and_4  g00745(new_n1122, new_n1121, new_n1120);
nor_4  g00746(new_n1123, new_n1121, new_n1120);
nor_4  g00747(new_n1124, new_n1123, new_n1122);
xnor_3 g00748(new_n1125, new_n1124, new_n1119);
not_3  g00749(new_n1126, new_n1111);
nor_4  g00750(new_n1127, new_n1126, new_n1107);
nor_4  g00751(new_n1128, new_n1127, new_n1112);
nand_4 g00752(new_n1129, new_n1128, new_n1125);
nand_4 g00753(new_n1130, new_n1129, new_n1113);
not_3  g00754(new_n1131, new_n1130);
not_3  g00755(new_n1132, new_n1103);
nand_4 g00756(new_n1133, n6776, n2024);
nor_4  g00757(new_n1134, new_n1133, new_n1132);
nand_4 g00758(new_n1135, n12299, n7946);
not_3  g00759(new_n1136_1, new_n1135);
nand_4 g00760(new_n1137, n9189, n8759);
not_3  g00761(new_n1138_1, new_n1137);
nand_4 g00762(new_n1139, new_n1138_1, new_n1136_1);
nand_4 g00763(new_n1140, new_n1137, new_n1135);
nand_4 g00764(new_n1141, new_n1140, new_n1139);
not_3  g00765(new_n1142, new_n1141);
nor_4  g00766(new_n1143, new_n1142, new_n1134);
not_3  g00767(new_n1144, new_n1133);
nand_4 g00768(new_n1145, new_n1140, new_n1144);
nor_4  g00769(new_n1146, new_n1145, new_n1132);
nor_4  g00770(new_n1147, new_n1146, new_n1143);
not_3  g00771(new_n1148, new_n1147);
nor_4  g00772(new_n1149, new_n1148, new_n1131);
nor_4  g00773(new_n1150, new_n1147, new_n1130);
nor_4  g00774(new_n1151, new_n1150, new_n1149);
nor_4  g00775(new_n1152, new_n1118, new_n1114);
nor_4  g00776(new_n1153, new_n1124, new_n1119);
nor_4  g00777(new_n1154, new_n1153, new_n1152);
not_3  g00778(new_n1155, new_n1105);
nand_4 g00779(new_n1156, n9111, n7388);
nor_4  g00780(new_n1157, new_n1156, new_n1155);
nand_4 g00781(new_n1158, n11892, n9763);
nand_4 g00782(new_n1159, n7965, n3342);
nand_4 g00783(new_n1160, new_n1159, new_n1158);
nor_4  g00784(new_n1161, new_n1159, new_n1158);
not_3  g00785(new_n1162, new_n1161);
nand_4 g00786(new_n1163, new_n1162, new_n1160);
not_3  g00787(new_n1164, new_n1163);
nor_4  g00788(new_n1165, new_n1164, new_n1157);
not_3  g00789(new_n1166, new_n1156);
nand_4 g00790(new_n1167, new_n1160, new_n1166);
nor_4  g00791(new_n1168, new_n1167, new_n1155);
nor_4  g00792(new_n1169, new_n1168, new_n1165);
xnor_3 g00793(new_n1170, new_n1169, new_n1154);
not_3  g00794(new_n1171, new_n1104);
nand_4 g00795(new_n1172, n8476, n2498);
nor_4  g00796(new_n1173, new_n1172, new_n1171);
not_3  g00797(new_n1174, new_n1173);
nand_4 g00798(new_n1175, n2558, n2530);
nand_4 g00799(new_n1176, n5579, n5331);
nand_4 g00800(new_n1177, new_n1176, new_n1175);
nor_4  g00801(new_n1178, new_n1177, new_n1174);
not_3  g00802(new_n1179, new_n1177);
nor_4  g00803(new_n1180, new_n1176, new_n1175);
nor_4  g00804(new_n1181, new_n1180, new_n1179);
not_3  g00805(new_n1182, new_n1181);
nor_4  g00806(new_n1183, new_n1182, new_n1173);
nor_4  g00807(new_n1184, new_n1183, new_n1178);
not_3  g00808(new_n1185, new_n1184);
nor_4  g00809(new_n1186, new_n1185, new_n1170);
not_3  g00810(new_n1187, new_n1170);
nor_4  g00811(new_n1188, new_n1184, new_n1187);
nor_4  g00812(new_n1189, new_n1188, new_n1186);
xnor_3 g00813(new_n1190, new_n1189, new_n1151);
not_3  g00814(new_n1191, new_n1190);
not_3  g00815(new_n1192, new_n1076);
nand_4 g00816(new_n1193, new_n1096, new_n1192);
nand_4 g00817(new_n1194, new_n1193, new_n1099);
nor_4  g00818(new_n1195, new_n1194, new_n1191);
not_3  g00819(new_n1196, new_n1195);
xor_3  g00820(new_n1197, new_n1106, new_n1103);
nand_4 g00821(new_n1198_1, new_n1197, new_n1095);
nand_4 g00822(new_n1199_1, n7265, n5964);
nand_4 g00823(new_n1200, n5305, n2879);
not_3  g00824(new_n1201, new_n1200);
xor_3  g00825(new_n1202, new_n1201, new_n1199_1);
nand_4 g00826(new_n1203, new_n1202, new_n1198_1);
not_3  g00827(new_n1204, new_n1203);
xor_3  g00828(new_n1205, new_n1128, new_n1125);
not_3  g00829(new_n1206, new_n1198_1);
xor_3  g00830(new_n1207, new_n1202, new_n1206);
nor_4  g00831(new_n1208, new_n1207, new_n1205);
nor_4  g00832(new_n1209_1, new_n1208, new_n1204);
not_3  g00833(new_n1210, new_n1194);
nor_4  g00834(new_n1211, new_n1210, new_n1190);
nor_4  g00835(new_n1212, new_n1211, new_n1195);
nand_4 g00836(new_n1213, new_n1212, new_n1209_1);
nand_4 g00837(new_n1214, new_n1213, new_n1196);
xnor_3 g00838(new_n1215, new_n1214, new_n1102);
nand_4 g00839(new_n1216, n8759, n2522);
nand_4 g00840(new_n1217, new_n1145, new_n1139);
xnor_3 g00841(new_n1218, new_n1217, new_n1216);
not_3  g00842(new_n1219, new_n1218);
nand_4 g00843(new_n1220, n12299, n2024);
not_3  g00844(new_n1221, new_n1220);
nand_4 g00845(new_n1222, n7946, n7436);
nand_4 g00846(new_n1223, n9189, n6776);
xnor_3 g00847(new_n1224, new_n1223, new_n1222);
xnor_3 g00848(new_n1225, new_n1224, new_n1221);
xor_3  g00849(new_n1226, new_n1225, new_n1219);
not_3  g00850(new_n1227, new_n1143);
nor_4  g00851(new_n1228, new_n1227, new_n1133);
not_3  g00852(new_n1229, new_n1228);
xnor_3 g00853(new_n1230, new_n1229, new_n1226);
not_3  g00854(new_n1231, new_n1150);
nand_4 g00855(new_n1232, new_n1189, new_n1151);
nand_4 g00856(new_n1233, new_n1232, new_n1231);
xnor_3 g00857(new_n1234, new_n1233, new_n1230);
nand_4 g00858(new_n1235, n5331, n521);
not_3  g00859(new_n1236, new_n1172);
nand_4 g00860(new_n1237, new_n1177, new_n1236);
not_3  g00861(new_n1238, new_n1237);
nor_4  g00862(new_n1239, new_n1238, new_n1180);
xnor_3 g00863(new_n1240, new_n1239, new_n1235);
nand_4 g00864(new_n1241, n12648, n2558);
nand_4 g00865(new_n1242, n8476, n5579);
not_3  g00866(new_n1243, new_n1242);
nand_4 g00867(new_n1244, n2530, n2498);
not_3  g00868(new_n1245, new_n1244);
nor_4  g00869(new_n1246, new_n1245, new_n1243);
nor_4  g00870(new_n1247, new_n1244, new_n1242);
nor_4  g00871(new_n1248, new_n1247, new_n1246);
xnor_3 g00872(new_n1249, new_n1248, new_n1241);
not_3  g00873(new_n1250, new_n1249);
xnor_3 g00874(new_n1251, new_n1250, new_n1240);
not_3  g00875(new_n1252, new_n1123);
nor_4  g00876(new_n1253, new_n1181, new_n1252);
not_3  g00877(new_n1254, new_n1253);
nor_4  g00878(new_n1255, new_n1254, new_n1251);
not_3  g00879(new_n1256, new_n1251);
nor_4  g00880(new_n1257, new_n1253, new_n1256);
nor_4  g00881(new_n1258, new_n1257, new_n1255);
nand_4 g00882(new_n1259, n7965, n806);
not_3  g00883(new_n1260, new_n1167);
nor_4  g00884(new_n1261, new_n1260, new_n1161);
xnor_3 g00885(new_n1262, new_n1261, new_n1259);
nand_4 g00886(new_n1263, n9763, n2393);
nand_4 g00887(new_n1264, n7388, n3342);
not_3  g00888(new_n1265, new_n1264);
nand_4 g00889(new_n1266, n11892, n9111);
not_3  g00890(new_n1267, new_n1266);
nor_4  g00891(new_n1268, new_n1267, new_n1265);
nor_4  g00892(new_n1269_1, new_n1266, new_n1264);
nor_4  g00893(new_n1270, new_n1269_1, new_n1268);
xnor_3 g00894(new_n1271, new_n1270, new_n1263);
not_3  g00895(new_n1272, new_n1271);
xnor_3 g00896(new_n1273, new_n1272, new_n1262);
not_3  g00897(new_n1274, new_n1165);
nor_4  g00898(new_n1275, new_n1274, new_n1156);
not_3  g00899(new_n1276, new_n1275);
nor_4  g00900(new_n1277, new_n1276, new_n1273);
not_3  g00901(new_n1278, new_n1273);
nor_4  g00902(new_n1279, new_n1275, new_n1278);
nor_4  g00903(new_n1280, new_n1279, new_n1277);
xnor_3 g00904(new_n1281, new_n1280, new_n1258);
not_3  g00905(new_n1282, new_n1281);
nor_4  g00906(new_n1283, new_n1169, new_n1154);
nor_4  g00907(new_n1284, new_n1186, new_n1283);
not_3  g00908(new_n1285, new_n1284);
nor_4  g00909(new_n1286, new_n1285, new_n1282);
nor_4  g00910(new_n1287, new_n1284, new_n1281);
nor_4  g00911(new_n1288, new_n1287, new_n1286);
xnor_3 g00912(new_n1289, new_n1288, new_n1234);
xor_3  g00913(n381, new_n1289, new_n1215);
nand_4 g00914(new_n1291, n7862, n6038);
nand_4 g00915(new_n1292, n7354, n6877);
nand_4 g00916(new_n1293, n4805, n1564);
nand_4 g00917(new_n1294, n8028, n7236);
not_3  g00918(new_n1295, new_n1294);
xor_3  g00919(new_n1296, new_n1295, new_n1293);
xor_3  g00920(new_n1297, new_n1296, new_n1292);
not_3  g00921(new_n1298, new_n1297);
xor_3  g00922(n397, new_n1298, new_n1291);
nand_4 g00923(new_n1300, n6687, n4370);
nand_4 g00924(new_n1301, n11407, n4189);
nand_4 g00925(new_n1302, n11877, n6687);
nand_4 g00926(new_n1303, new_n1302, new_n1301);
not_3  g00927(new_n1304, new_n1303);
nor_4  g00928(new_n1305, new_n1302, new_n1301);
nand_4 g00929(new_n1306, n5212, n2564);
not_3  g00930(new_n1307, new_n1306);
nor_4  g00931(new_n1308, new_n1307, new_n1305);
nor_4  g00932(new_n1309, new_n1308, new_n1304);
xor_3  g00933(new_n1310, new_n1309, new_n1300);
nand_4 g00934(new_n1311, n5212, n4189);
not_3  g00935(new_n1312, new_n1311);
nand_4 g00936(new_n1313, n11407, n6770);
nand_4 g00937(new_n1314, n11877, n2564);
xnor_3 g00938(new_n1315, new_n1314, new_n1313);
xor_3  g00939(new_n1316, new_n1315, new_n1312);
xnor_3 g00940(new_n1317, new_n1316, new_n1310);
not_3  g00941(new_n1318, new_n1317);
nand_4 g00942(new_n1319, n11407, n6687);
not_3  g00943(new_n1320, new_n1319);
nor_4  g00944(new_n1321, new_n1320, new_n1306);
nor_4  g00945(new_n1322, new_n1321, new_n1303);
nor_4  g00946(new_n1323, new_n1322, new_n1305);
nor_4  g00947(new_n1324, new_n1323, new_n1306);
xor_3  g00948(new_n1325, new_n1324, new_n1318);
not_3  g00949(new_n1326, new_n1325);
nand_4 g00950(new_n1327, n12709, n8336);
nand_4 g00951(new_n1328, n11222, n10990);
nand_4 g00952(new_n1329, n12489, n12069);
xnor_3 g00953(new_n1330, new_n1329, new_n1328);
nor_4  g00954(new_n1331, new_n1330, new_n1327);
not_3  g00955(new_n1332, new_n1331);
nand_4 g00956(new_n1333_1, n11728, n8336);
nand_4 g00957(new_n1334, n12709, n10928);
not_3  g00958(new_n1335, new_n1334);
xor_3  g00959(new_n1336, new_n1335, new_n1333_1);
nand_4 g00960(new_n1337, new_n1336, new_n1332);
nor_4  g00961(new_n1338, new_n1329, new_n1328);
not_3  g00962(new_n1339, new_n1338);
nand_4 g00963(new_n1340, n11222, n5760);
nand_4 g00964(new_n1341, n11153, n10990);
xnor_3 g00965(new_n1342, new_n1341, new_n1340);
xnor_3 g00966(new_n1343, new_n1342, new_n1339);
nand_4 g00967(new_n1344, n12069, n7159);
nand_4 g00968(new_n1345, n12489, n12391);
xor_3  g00969(new_n1346, new_n1345, new_n1344);
not_3  g00970(new_n1347, new_n1346);
xnor_3 g00971(new_n1348, new_n1347, new_n1343);
not_3  g00972(new_n1349, new_n1337);
nor_4  g00973(new_n1350, new_n1336, new_n1332);
nor_4  g00974(new_n1351, new_n1350, new_n1349);
nand_4 g00975(new_n1352, new_n1351, new_n1348);
nand_4 g00976(new_n1353_1, new_n1352, new_n1337);
not_3  g00977(new_n1354, new_n1327);
nand_4 g00978(new_n1355, n11728, n10928);
nor_4  g00979(new_n1356, new_n1355, new_n1354);
nand_4 g00980(new_n1357_1, n12709, n6986);
not_3  g00981(new_n1358, new_n1357_1);
nand_4 g00982(new_n1359, n8336, n6429);
not_3  g00983(new_n1360, new_n1359);
nor_4  g00984(new_n1361, new_n1360, new_n1358);
nor_4  g00985(new_n1362, new_n1359, new_n1357_1);
nor_4  g00986(new_n1363, new_n1362, new_n1361);
nor_4  g00987(new_n1364, new_n1363, new_n1356);
not_3  g00988(new_n1365, new_n1364);
not_3  g00989(new_n1366, new_n1361);
nand_4 g00990(new_n1367, new_n1366, new_n1356);
nand_4 g00991(new_n1368, new_n1367, new_n1365);
xnor_3 g00992(new_n1369, new_n1368, new_n1353_1);
not_3  g00993(new_n1370, new_n1329);
nand_4 g00994(new_n1371, n12391, n7159);
nor_4  g00995(new_n1372, new_n1371, new_n1370);
nand_4 g00996(new_n1373, n12489, n7891);
nand_4 g00997(new_n1374, n12777, n12069);
nand_4 g00998(new_n1375, new_n1374, new_n1373);
nor_4  g00999(new_n1376, new_n1375, new_n1372);
nor_4  g01000(new_n1377, new_n1374, new_n1373);
nor_4  g01001(new_n1378, new_n1377, new_n1376);
nand_4 g01002(new_n1379, new_n1375, new_n1372);
nand_4 g01003(new_n1380, new_n1379, new_n1378);
nand_4 g01004(new_n1381, n11153, n5760);
not_3  g01005(new_n1382, new_n1381);
nand_4 g01006(new_n1383, new_n1382, new_n1328);
nand_4 g01007(new_n1384, n10990, n5314);
not_3  g01008(new_n1385, new_n1384);
nand_4 g01009(new_n1386, n11222, n1478);
not_3  g01010(new_n1387, new_n1386);
nand_4 g01011(new_n1388, new_n1387, new_n1385);
nand_4 g01012(new_n1389, new_n1386, new_n1384);
nand_4 g01013(new_n1390, new_n1389, new_n1388);
nand_4 g01014(new_n1391, new_n1390, new_n1383);
nand_4 g01015(new_n1392, new_n1389, new_n1382);
not_3  g01016(new_n1393, new_n1392);
nand_4 g01017(new_n1394, new_n1393, new_n1328);
nand_4 g01018(new_n1395, new_n1394, new_n1391);
xnor_3 g01019(new_n1396, new_n1395, new_n1380);
nor_4  g01020(new_n1397, new_n1342, new_n1339);
nor_4  g01021(new_n1398, new_n1347, new_n1343);
nor_4  g01022(new_n1399, new_n1398, new_n1397);
nor_4  g01023(new_n1400, new_n1399, new_n1396);
and_4  g01024(new_n1401, new_n1399, new_n1396);
nor_4  g01025(new_n1402, new_n1401, new_n1400);
xnor_3 g01026(new_n1403, new_n1402, new_n1369);
not_3  g01027(new_n1404, new_n1403);
not_3  g01028(new_n1405, new_n1323);
not_3  g01029(new_n1406, new_n1321);
nor_4  g01030(new_n1407, new_n1406, new_n1304);
nor_4  g01031(new_n1408, new_n1407, new_n1405);
not_3  g01032(new_n1409, new_n1408);
nand_4 g01033(new_n1410, new_n1409, new_n1404);
xnor_3 g01034(new_n1411, new_n1409, new_n1403);
xor_3  g01035(new_n1412, new_n1330, new_n1327);
nand_4 g01036(new_n1413, new_n1412, new_n1320);
not_3  g01037(new_n1414, new_n1413);
nand_4 g01038(new_n1415, n11407, n2564);
nand_4 g01039(new_n1416, n6687, n5212);
xor_3  g01040(new_n1417, new_n1416, new_n1415);
nor_4  g01041(new_n1418, new_n1417, new_n1414);
not_3  g01042(new_n1419, new_n1418);
not_3  g01043(new_n1420, new_n1348);
xnor_3 g01044(new_n1421, new_n1351, new_n1420);
xor_3  g01045(new_n1422, new_n1417, new_n1414);
nand_4 g01046(new_n1423, new_n1422, new_n1421);
nand_4 g01047(new_n1424, new_n1423, new_n1419);
nand_4 g01048(new_n1425, new_n1424, new_n1411);
nand_4 g01049(new_n1426, new_n1425, new_n1410);
nor_4  g01050(new_n1427, new_n1426, new_n1326);
not_3  g01051(new_n1428, new_n1426);
nor_4  g01052(new_n1429, new_n1428, new_n1325);
nor_4  g01053(new_n1430, new_n1429, new_n1427);
nand_4 g01054(new_n1431, n8819, n8336);
nand_4 g01055(new_n1432, n11728, n6986);
not_3  g01056(new_n1433, new_n1432);
nand_4 g01057(new_n1434, n10928, n6429);
nand_4 g01058(new_n1435, n12709, n2226);
xnor_3 g01059(new_n1436, new_n1435, new_n1434);
xnor_3 g01060(new_n1437, new_n1436, new_n1433);
not_3  g01061(new_n1438, new_n1437);
xor_3  g01062(new_n1439, new_n1438, new_n1431);
not_3  g01063(new_n1440, new_n1355);
nor_4  g01064(new_n1441, new_n1362, new_n1440);
nor_4  g01065(new_n1442, new_n1441, new_n1361);
xnor_3 g01066(new_n1443, new_n1442, new_n1439);
nor_4  g01067(new_n1444, new_n1365, new_n1355);
xnor_3 g01068(new_n1445, new_n1444, new_n1443);
nand_4 g01069(new_n1446, n12069, n6254);
not_3  g01070(new_n1447, new_n1446);
not_3  g01071(new_n1448, new_n1375);
not_3  g01072(new_n1449, new_n1371);
nor_4  g01073(new_n1450, new_n1377, new_n1449);
nor_4  g01074(new_n1451, new_n1450, new_n1448);
xnor_3 g01075(new_n1452, new_n1451, new_n1447);
nand_4 g01076(new_n1453, n12489, n7160);
nand_4 g01077(new_n1454, n12777, n12391);
not_3  g01078(new_n1455, new_n1454);
nand_4 g01079(new_n1456, n7891, n7159);
not_3  g01080(new_n1457, new_n1456);
nor_4  g01081(new_n1458, new_n1457, new_n1455);
nor_4  g01082(new_n1459, new_n1456, new_n1454);
nor_4  g01083(new_n1460, new_n1459, new_n1458);
xnor_3 g01084(new_n1461, new_n1460, new_n1453);
not_3  g01085(new_n1462, new_n1461);
xnor_3 g01086(new_n1463, new_n1462, new_n1452);
nor_4  g01087(new_n1464, new_n1378, new_n1371);
not_3  g01088(new_n1465, new_n1464);
nor_4  g01089(new_n1466, new_n1465, new_n1463);
not_3  g01090(new_n1467, new_n1463);
nor_4  g01091(new_n1468, new_n1464, new_n1467);
nor_4  g01092(new_n1469, new_n1468, new_n1466);
nand_4 g01093(new_n1470, n11791, n11222);
nand_4 g01094(new_n1471_1, new_n1392, new_n1388);
not_3  g01095(new_n1472, new_n1471_1);
xnor_3 g01096(new_n1473, new_n1472, new_n1470);
nand_4 g01097(new_n1474, n5760, n5314);
nand_4 g01098(new_n1475, n10990, n996);
nand_4 g01099(new_n1476, n11153, n1478);
xnor_3 g01100(new_n1477, new_n1476, new_n1475);
xnor_3 g01101(new_n1478_1, new_n1477, new_n1474);
xnor_3 g01102(new_n1479, new_n1478_1, new_n1473);
nor_4  g01103(new_n1480, new_n1391, new_n1381);
not_3  g01104(new_n1481, new_n1480);
nor_4  g01105(new_n1482, new_n1481, new_n1479);
not_3  g01106(new_n1483, new_n1479);
nor_4  g01107(new_n1484, new_n1480, new_n1483);
nor_4  g01108(new_n1485, new_n1484, new_n1482);
xnor_3 g01109(new_n1486, new_n1485, new_n1469);
nor_4  g01110(new_n1487, new_n1395, new_n1380);
not_3  g01111(new_n1488, new_n1487);
not_3  g01112(new_n1489, new_n1400);
nand_4 g01113(new_n1490, new_n1489, new_n1488);
xnor_3 g01114(new_n1491, new_n1490, new_n1486);
xnor_3 g01115(new_n1492, new_n1491, new_n1445);
nand_4 g01116(new_n1493, new_n1368, new_n1353_1);
not_3  g01117(new_n1494, new_n1493);
nor_4  g01118(new_n1495, new_n1402, new_n1369);
nor_4  g01119(new_n1496, new_n1495, new_n1494);
not_3  g01120(new_n1497, new_n1496);
nor_4  g01121(new_n1498, new_n1497, new_n1492);
not_3  g01122(new_n1499, new_n1492);
nor_4  g01123(new_n1500, new_n1496, new_n1499);
nor_4  g01124(new_n1501, new_n1500, new_n1498);
xor_3  g01125(n658, new_n1501, new_n1430);
nand_4 g01126(new_n1503, n7862, n2585);
not_3  g01127(new_n1504, new_n1503);
nand_4 g01128(new_n1505, n2508, n1333);
not_3  g01129(new_n1506, new_n1505);
nand_4 g01130(new_n1507, n11757, n6038);
not_3  g01131(new_n1508, new_n1507);
nand_4 g01132(new_n1509, n12720, n1333);
not_3  g01133(new_n1510_1, new_n1509);
nor_4  g01134(new_n1511, new_n1510_1, new_n1508);
nor_4  g01135(new_n1512_1, new_n1509, new_n1507);
nand_4 g01136(new_n1513, n3172, n2509);
not_3  g01137(new_n1514, new_n1513);
nor_4  g01138(new_n1515, new_n1514, new_n1512_1);
nor_4  g01139(new_n1516, new_n1515, new_n1511);
xnor_3 g01140(new_n1517, new_n1516, new_n1506);
nand_4 g01141(new_n1518, n11757, n2509);
nand_4 g01142(new_n1519, n6038, n5240);
nand_4 g01143(new_n1520, n12720, n3172);
xnor_3 g01144(new_n1521, new_n1520, new_n1519);
xnor_3 g01145(new_n1522, new_n1521, new_n1518);
xnor_3 g01146(new_n1523_1, new_n1522, new_n1517);
not_3  g01147(new_n1524, new_n1523_1);
nor_4  g01148(new_n1525, new_n1524, new_n1504);
not_3  g01149(new_n1526, new_n1525);
nor_4  g01150(new_n1527, new_n1523_1, new_n1503);
nor_4  g01151(new_n1528, new_n1527, new_n1525);
nand_4 g01152(new_n1529, n7862, n2508);
nand_4 g01153(new_n1530, n2509, n1333);
not_3  g01154(new_n1531, new_n1530);
nand_4 g01155(new_n1532, n6038, n3172);
nand_4 g01156(new_n1533, n12720, n7862);
nand_4 g01157(new_n1534, new_n1533, new_n1532);
nand_4 g01158(new_n1535, new_n1534, new_n1531);
not_3  g01159(new_n1536, new_n1532);
not_3  g01160(new_n1537, new_n1533);
nand_4 g01161(new_n1538, new_n1537, new_n1536);
nand_4 g01162(new_n1539, new_n1538, new_n1535);
not_3  g01163(new_n1540, new_n1539);
nor_4  g01164(new_n1541, new_n1540, new_n1529);
xor_3  g01165(new_n1542, new_n1539, new_n1529);
nor_4  g01166(new_n1543, new_n1512_1, new_n1511);
xor_3  g01167(new_n1544, new_n1543, new_n1513);
nor_4  g01168(new_n1545, new_n1544, new_n1542);
nor_4  g01169(new_n1546, new_n1545, new_n1541);
nand_4 g01170(new_n1547, new_n1546, new_n1528);
nand_4 g01171(new_n1548, new_n1547, new_n1526);
not_3  g01172(new_n1549, new_n1548);
nand_4 g01173(new_n1550, n12720, n11757);
nand_4 g01174(new_n1551, n5240, n2509);
nand_4 g01175(new_n1552, n11821, n6038);
xnor_3 g01176(new_n1553, new_n1552, new_n1551);
nor_4  g01177(new_n1554, new_n1553, new_n1550);
not_3  g01178(new_n1555, new_n1550);
not_3  g01179(new_n1556, new_n1553);
nor_4  g01180(new_n1557, new_n1556, new_n1555);
nor_4  g01181(new_n1558, new_n1557, new_n1554);
not_3  g01182(new_n1559, new_n1519);
not_3  g01183(new_n1560, new_n1520);
nor_4  g01184(new_n1561, new_n1560, new_n1559);
not_3  g01185(new_n1562, new_n1518);
nor_4  g01186(new_n1563, new_n1521, new_n1562);
nor_4  g01187(new_n1564_1, new_n1563, new_n1561);
xnor_3 g01188(new_n1565, new_n1564_1, new_n1558);
not_3  g01189(new_n1566, new_n1565);
nand_4 g01190(new_n1567, new_n1516, new_n1506);
not_3  g01191(new_n1568, new_n1567);
nor_4  g01192(new_n1569, new_n1522, new_n1517);
nor_4  g01193(new_n1570, new_n1569, new_n1568);
not_3  g01194(new_n1571, new_n1570);
nand_4 g01195(new_n1572, n2585, n1333);
nand_4 g01196(new_n1573, n3172, n2508);
xor_3  g01197(new_n1574, new_n1573, new_n1572);
nor_4  g01198(new_n1575, new_n1574, new_n1571);
not_3  g01199(new_n1576_1, new_n1574);
nor_4  g01200(new_n1577, new_n1576_1, new_n1570);
nor_4  g01201(new_n1578, new_n1577, new_n1575);
xnor_3 g01202(new_n1579, new_n1578, new_n1566);
not_3  g01203(new_n1580, new_n1579);
nand_4 g01204(new_n1581, new_n1580, new_n1549);
not_3  g01205(new_n1582, new_n1577);
nor_4  g01206(new_n1583, new_n1573, new_n1572);
nor_4  g01207(new_n1584, new_n1575, new_n1565);
xnor_3 g01208(new_n1585, new_n1584, new_n1583);
nand_4 g01209(new_n1586, new_n1585, new_n1582);
nor_4  g01210(new_n1587, new_n1552, new_n1551);
nand_4 g01211(new_n1588, n11757, n2508);
not_3  g01212(new_n1589, new_n1588);
xor_3  g01213(new_n1590, new_n1589, new_n1587);
nand_4 g01214(new_n1591, n11821, n2509);
not_3  g01215(new_n1592, new_n1591);
nand_4 g01216(new_n1593, n12720, n5240);
nand_4 g01217(new_n1594, n9080, n6038);
xnor_3 g01218(new_n1595, new_n1594, new_n1593);
xnor_3 g01219(new_n1596, new_n1595, new_n1592);
not_3  g01220(new_n1597, new_n1596);
xnor_3 g01221(new_n1598, new_n1597, new_n1590);
not_3  g01222(new_n1599, new_n1554);
nand_4 g01223(new_n1600, new_n1564_1, new_n1558);
nand_4 g01224(new_n1601, new_n1600, new_n1599);
nand_4 g01225(new_n1602, n4005, n1333);
nand_4 g01226(new_n1603, n3172, n2585);
nand_4 g01227(new_n1604, n12706, n7862);
nand_4 g01228(new_n1605, new_n1604, new_n1603);
not_3  g01229(new_n1606, new_n1603);
not_3  g01230(new_n1607, new_n1604);
nand_4 g01231(new_n1608, new_n1607, new_n1606);
nand_4 g01232(new_n1609, new_n1608, new_n1605);
xor_3  g01233(new_n1610, new_n1609, new_n1602);
xnor_3 g01234(new_n1611, new_n1610, new_n1601);
xnor_3 g01235(new_n1612, new_n1611, new_n1598);
not_3  g01236(new_n1613, new_n1612);
xnor_3 g01237(new_n1614, new_n1613, new_n1586);
xnor_3 g01238(new_n1615, new_n1614, new_n1581);
nand_4 g01239(new_n1616, n7862, n4005);
not_3  g01240(new_n1617, new_n1616);
xnor_3 g01241(new_n1618, new_n1579, new_n1548);
not_3  g01242(new_n1619, new_n1618);
nand_4 g01243(new_n1620, new_n1619, new_n1617);
and_4  g01244(new_n1621, new_n1538, new_n1534);
nand_4 g01245(new_n1622, n6038, n1333);
nand_4 g01246(new_n1623, n7862, n2509);
nor_4  g01247(new_n1624, new_n1623, new_n1622);
not_3  g01248(new_n1625, new_n1624);
nor_4  g01249(new_n1626, new_n1625, new_n1621);
not_3  g01250(new_n1627, new_n1542);
not_3  g01251(new_n1628, new_n1544);
xor_3  g01252(new_n1629, new_n1628, new_n1627);
nand_4 g01253(new_n1630, new_n1629, new_n1626);
not_3  g01254(new_n1631, new_n1547);
nor_4  g01255(new_n1632, new_n1546, new_n1528);
nor_4  g01256(new_n1633, new_n1632, new_n1631);
nor_4  g01257(new_n1634, new_n1633, new_n1630);
nor_4  g01258(new_n1635, new_n1618, new_n1616);
nor_4  g01259(new_n1636, new_n1619, new_n1617);
nor_4  g01260(new_n1637, new_n1636, new_n1635);
nand_4 g01261(new_n1638, new_n1637, new_n1634);
nand_4 g01262(new_n1639, new_n1638, new_n1620);
xnor_3 g01263(new_n1640, new_n1639, new_n1615);
not_3  g01264(new_n1641, new_n1640);
nand_4 g01265(new_n1642, n2464, n1209);
nor_4  g01266(new_n1643, new_n1642, new_n1292);
nand_4 g01267(new_n1644, n7354, n2464);
nand_4 g01268(new_n1645, n6877, n1209);
nand_4 g01269(new_n1646, new_n1645, new_n1644);
not_3  g01270(new_n1647, new_n1646);
nor_4  g01271(new_n1648, new_n1647, new_n1643);
nand_4 g01272(new_n1649, n9400, n7354);
nand_4 g01273(new_n1650, n7500, n6877);
nor_4  g01274(new_n1651, new_n1650, new_n1649);
not_3  g01275(new_n1652, new_n1651);
nor_4  g01276(new_n1653, new_n1652, new_n1648);
not_3  g01277(new_n1654, new_n1653);
nand_4 g01278(new_n1655, n6877, n5105);
not_3  g01279(new_n1656, new_n1655);
not_3  g01280(new_n1657, new_n1643);
nand_4 g01281(new_n1658_1, n9400, n7500);
not_3  g01282(new_n1659, new_n1658_1);
nand_4 g01283(new_n1660, new_n1659, new_n1646);
nand_4 g01284(new_n1661, new_n1660, new_n1657);
nand_4 g01285(new_n1662, new_n1661, new_n1656);
not_3  g01286(new_n1663, new_n1662);
nor_4  g01287(new_n1664, new_n1661, new_n1656);
nor_4  g01288(new_n1665, new_n1664, new_n1663);
nand_4 g01289(new_n1666, n7500, n2464);
nand_4 g01290(new_n1667, n9400, n1209);
not_3  g01291(new_n1668, new_n1667);
nand_4 g01292(new_n1669, n11311, n7354);
not_3  g01293(new_n1670, new_n1669);
nor_4  g01294(new_n1671, new_n1670, new_n1668);
nor_4  g01295(new_n1672, new_n1669, new_n1667);
nor_4  g01296(new_n1673, new_n1672, new_n1671);
xnor_3 g01297(new_n1674, new_n1673, new_n1666);
xor_3  g01298(new_n1675, new_n1674, new_n1665);
not_3  g01299(new_n1676, new_n1675);
nor_4  g01300(new_n1677, new_n1676, new_n1654);
not_3  g01301(new_n1678, new_n1677);
nand_4 g01302(new_n1679, n11311, n7500);
not_3  g01303(new_n1680, new_n1679);
nand_4 g01304(new_n1681, n7354, n4187);
xnor_3 g01305(new_n1682, new_n1681, new_n1642);
xnor_3 g01306(new_n1683, new_n1682, new_n1680);
not_3  g01307(new_n1684, new_n1683);
nand_4 g01308(new_n1685, n9400, n5105);
not_3  g01309(new_n1686, new_n1666);
nor_4  g01310(new_n1687, new_n1672, new_n1686);
nor_4  g01311(new_n1688, new_n1687, new_n1671);
xnor_3 g01312(new_n1689, new_n1688, new_n1685);
xnor_3 g01313(new_n1690, new_n1689, new_n1684);
nand_4 g01314(new_n1691, n6877, n4141);
not_3  g01315(new_n1692, new_n1691);
nand_4 g01316(new_n1693, new_n1674, new_n1665);
nand_4 g01317(new_n1694, new_n1693, new_n1662);
xnor_3 g01318(new_n1695, new_n1694, new_n1692);
xor_3  g01319(new_n1696, new_n1695, new_n1690);
nor_4  g01320(new_n1697, new_n1696, new_n1678);
not_3  g01321(new_n1698, new_n1697);
nand_4 g01322(new_n1699, n6877, n4928);
nor_4  g01323(new_n1700, new_n1694, new_n1692);
nor_4  g01324(new_n1701, new_n1695, new_n1690);
nor_4  g01325(new_n1702, new_n1701, new_n1700);
not_3  g01326(new_n1703, new_n1702);
nand_4 g01327(new_n1704, n11311, n1209);
nand_4 g01328(new_n1705, n7500, n4187);
nand_4 g01329(new_n1706, n7354, n4203);
xnor_3 g01330(new_n1707, new_n1706, new_n1705);
nor_4  g01331(new_n1708, new_n1707, new_n1704);
not_3  g01332(new_n1709, new_n1704);
not_3  g01333(new_n1710, new_n1707);
nor_4  g01334(new_n1711, new_n1710, new_n1709);
nor_4  g01335(new_n1712, new_n1711, new_n1708);
and_4  g01336(new_n1713, new_n1681, new_n1642);
nor_4  g01337(new_n1714, new_n1682, new_n1680);
nor_4  g01338(new_n1715, new_n1714, new_n1713);
xnor_3 g01339(new_n1716, new_n1715, new_n1712);
not_3  g01340(new_n1717, new_n1685);
nand_4 g01341(new_n1718, new_n1688, new_n1717);
nand_4 g01342(new_n1719, new_n1689, new_n1683);
nand_4 g01343(new_n1720, new_n1719, new_n1718);
nand_4 g01344(new_n1721, n9400, n4141);
nand_4 g01345(new_n1722, n5105, n2464);
xor_3  g01346(new_n1723, new_n1722, new_n1721);
xnor_3 g01347(new_n1724, new_n1723, new_n1720);
xnor_3 g01348(new_n1725, new_n1724, new_n1716);
nor_4  g01349(new_n1726, new_n1725, new_n1703);
not_3  g01350(new_n1727, new_n1725);
nor_4  g01351(new_n1728, new_n1727, new_n1702);
nor_4  g01352(new_n1729, new_n1728, new_n1726);
xnor_3 g01353(new_n1730, new_n1729, new_n1699);
xnor_3 g01354(new_n1731, new_n1730, new_n1698);
not_3  g01355(new_n1732, new_n1731);
nand_4 g01356(new_n1733, n7294, n7236);
not_3  g01357(new_n1734, new_n1733);
nand_4 g01358(new_n1735, n10848, n3992);
not_3  g01359(new_n1736, new_n1735);
nand_4 g01360(new_n1737, n8384, n8028);
nand_4 g01361(new_n1738, n7236, n1980);
nand_4 g01362(new_n1739, new_n1738, new_n1737);
nand_4 g01363(new_n1740, new_n1739, new_n1736);
not_3  g01364(new_n1741, new_n1737);
not_3  g01365(new_n1742, new_n1738);
nand_4 g01366(new_n1743, new_n1742, new_n1741);
nand_4 g01367(new_n1744, new_n1743, new_n1740);
nand_4 g01368(new_n1745, new_n1744, new_n1734);
not_3  g01369(new_n1746, new_n1745);
nor_4  g01370(new_n1747, new_n1744, new_n1734);
nor_4  g01371(new_n1748, new_n1747, new_n1746);
nand_4 g01372(new_n1749, n8028, n6358);
nand_4 g01373(new_n1750, n3992, n1980);
nand_4 g01374(new_n1751, n10848, n8384);
xnor_3 g01375(new_n1752, new_n1751, new_n1750);
xnor_3 g01376(new_n1753, new_n1752, new_n1749);
not_3  g01377(new_n1754, new_n1753);
xnor_3 g01378(new_n1755, new_n1754, new_n1748);
nand_4 g01379(new_n1756, new_n1743, new_n1739);
not_3  g01380(new_n1757, new_n1756);
nand_4 g01381(new_n1758, n10848, n7236);
nand_4 g01382(new_n1759, n8028, n3992);
nor_4  g01383(new_n1760, new_n1759, new_n1758);
not_3  g01384(new_n1761, new_n1760);
nor_4  g01385(new_n1762, new_n1761, new_n1757);
not_3  g01386(new_n1763, new_n1762);
nor_4  g01387(new_n1764, new_n1763, new_n1755);
nand_4 g01388(new_n1765, n10848, n6358);
not_3  g01389(new_n1766, new_n1765);
nand_4 g01390(new_n1767, n8384, n1980);
nand_4 g01391(new_n1768, n8028, n5198);
xnor_3 g01392(new_n1769, new_n1768, new_n1767);
nor_4  g01393(new_n1770, new_n1769, new_n1766);
not_3  g01394(new_n1771, new_n1769);
nor_4  g01395(new_n1772, new_n1771, new_n1765);
nor_4  g01396(new_n1773, new_n1772, new_n1770);
nand_4 g01397(new_n1774, n7294, n3992);
not_3  g01398(new_n1775, new_n1750);
not_3  g01399(new_n1776, new_n1751);
nor_4  g01400(new_n1777, new_n1776, new_n1775);
not_3  g01401(new_n1778, new_n1749);
nor_4  g01402(new_n1779, new_n1752, new_n1778);
nor_4  g01403(new_n1780, new_n1779, new_n1777);
xnor_3 g01404(new_n1781, new_n1780, new_n1774);
xnor_3 g01405(new_n1782, new_n1781, new_n1773);
nand_4 g01406(new_n1783, n12704, n7236);
not_3  g01407(new_n1784, new_n1783);
nand_4 g01408(new_n1785, new_n1754, new_n1748);
nand_4 g01409(new_n1786, new_n1785, new_n1745);
xnor_3 g01410(new_n1787, new_n1786, new_n1784);
xnor_3 g01411(new_n1788, new_n1787, new_n1782);
nand_4 g01412(new_n1789, new_n1788, new_n1764);
nand_4 g01413(new_n1790, n7236, n5814);
not_3  g01414(new_n1791, new_n1790);
not_3  g01415(new_n1792, new_n1774);
nand_4 g01416(new_n1793, new_n1780, new_n1792);
not_3  g01417(new_n1794, new_n1773);
nand_4 g01418(new_n1795, new_n1781, new_n1794);
nand_4 g01419(new_n1796, new_n1795, new_n1793);
nand_4 g01420(new_n1797, n8384, n7294);
nand_4 g01421(new_n1798_1, n12704, n3992);
xor_3  g01422(new_n1799, new_n1798_1, new_n1797);
xnor_3 g01423(new_n1800, new_n1799, new_n1796);
nand_4 g01424(new_n1801, n6358, n1980);
not_3  g01425(new_n1802, new_n1767);
not_3  g01426(new_n1803, new_n1768);
nor_4  g01427(new_n1804, new_n1803, new_n1802);
nor_4  g01428(new_n1805, new_n1770, new_n1804);
xnor_3 g01429(new_n1806, new_n1805, new_n1801);
nand_4 g01430(new_n1807, n10848, n5198);
nand_4 g01431(new_n1808, n8028, n1471);
xor_3  g01432(new_n1809, new_n1808, new_n1807);
xnor_3 g01433(new_n1810, new_n1809, new_n1806);
xnor_3 g01434(new_n1811, new_n1810, new_n1800);
nor_4  g01435(new_n1812, new_n1786, new_n1784);
nor_4  g01436(new_n1813, new_n1787, new_n1782);
nor_4  g01437(new_n1814, new_n1813, new_n1812);
xnor_3 g01438(new_n1815, new_n1814, new_n1811);
xnor_3 g01439(new_n1816, new_n1815, new_n1791);
nor_4  g01440(new_n1817, new_n1816, new_n1789);
not_3  g01441(new_n1818, new_n1789);
not_3  g01442(new_n1819, new_n1816);
nor_4  g01443(new_n1820, new_n1819, new_n1818);
nor_4  g01444(new_n1821, new_n1820, new_n1817);
nand_4 g01445(new_n1822, n4805, n533);
nand_4 g01446(new_n1823, n5283, n1564);
nand_4 g01447(new_n1824, new_n1823, new_n1822);
nor_4  g01448(new_n1825, new_n1823, new_n1822);
not_3  g01449(new_n1826, new_n1825);
nand_4 g01450(new_n1827, new_n1826, new_n1824);
not_3  g01451(new_n1828, new_n1827);
nand_4 g01452(new_n1829, n11478, n1564);
nand_4 g01453(new_n1830, n4805, n1512);
nor_4  g01454(new_n1831, new_n1830, new_n1829);
not_3  g01455(new_n1832, new_n1831);
nor_4  g01456(new_n1833, new_n1832, new_n1828);
not_3  g01457(new_n1834, new_n1833);
nand_4 g01458(new_n1835_1, n4805, n2802);
nand_4 g01459(new_n1836, n11478, n1512);
not_3  g01460(new_n1837, new_n1836);
nand_4 g01461(new_n1838, new_n1837, new_n1824);
nand_4 g01462(new_n1839, new_n1838, new_n1826);
not_3  g01463(new_n1840, new_n1839);
xnor_3 g01464(new_n1841, new_n1840, new_n1835_1);
nand_4 g01465(new_n1842, n1564, n137);
nand_4 g01466(new_n1843, n5283, n1512);
nand_4 g01467(new_n1844, n11478, n533);
xnor_3 g01468(new_n1845, new_n1844, new_n1843);
xnor_3 g01469(new_n1846, new_n1845, new_n1842);
xnor_3 g01470(new_n1847_1, new_n1846, new_n1841);
nor_4  g01471(new_n1848, new_n1847_1, new_n1834);
not_3  g01472(new_n1849, new_n1848);
nand_4 g01473(new_n1850, n6806, n4805);
nand_4 g01474(new_n1851, n11478, n2802);
not_3  g01475(new_n1852, new_n1851);
not_3  g01476(new_n1853, new_n1843);
not_3  g01477(new_n1854, new_n1844);
nor_4  g01478(new_n1855, new_n1854, new_n1853);
not_3  g01479(new_n1856, new_n1842);
nor_4  g01480(new_n1857, new_n1845, new_n1856);
nor_4  g01481(new_n1858, new_n1857, new_n1855);
xnor_3 g01482(new_n1859, new_n1858, new_n1852);
nand_4 g01483(new_n1860, n1512, n137);
nand_4 g01484(new_n1861, n5283, n533);
nand_4 g01485(new_n1862, n6294, n1564);
xnor_3 g01486(new_n1863, new_n1862, new_n1861);
xnor_3 g01487(new_n1864, new_n1863, new_n1860);
xnor_3 g01488(new_n1865, new_n1864, new_n1859);
nand_4 g01489(new_n1866, new_n1865, new_n1850);
not_3  g01490(new_n1867, new_n1866);
nor_4  g01491(new_n1868, new_n1865, new_n1850);
nor_4  g01492(new_n1869, new_n1868, new_n1867);
nor_4  g01493(new_n1870, new_n1840, new_n1835_1);
nor_4  g01494(new_n1871, new_n1846, new_n1841);
nor_4  g01495(new_n1872, new_n1871, new_n1870);
nand_4 g01496(new_n1873, new_n1872, new_n1869);
not_3  g01497(new_n1874, new_n1873);
nor_4  g01498(new_n1875, new_n1872, new_n1869);
nor_4  g01499(new_n1876, new_n1875, new_n1874);
nor_4  g01500(new_n1877, new_n1876, new_n1849);
nand_4 g01501(new_n1878, n5069, n4805);
nand_4 g01502(new_n1879, n533, n137);
nand_4 g01503(new_n1880, n6294, n1512);
nand_4 g01504(new_n1881, n6797, n1564);
xnor_3 g01505(new_n1882, new_n1881, new_n1880);
nor_4  g01506(new_n1883, new_n1882, new_n1879);
not_3  g01507(new_n1884, new_n1879);
not_3  g01508(new_n1885, new_n1882);
nor_4  g01509(new_n1886, new_n1885, new_n1884);
nor_4  g01510(new_n1887, new_n1886, new_n1883);
and_4  g01511(new_n1888, new_n1862, new_n1861);
not_3  g01512(new_n1889, new_n1860);
nor_4  g01513(new_n1890, new_n1863, new_n1889);
nor_4  g01514(new_n1891, new_n1890, new_n1888);
xnor_3 g01515(new_n1892, new_n1891, new_n1887);
not_3  g01516(new_n1893, new_n1892);
nand_4 g01517(new_n1894, n11478, n6806);
nand_4 g01518(new_n1895, n5283, n2802);
xor_3  g01519(new_n1896, new_n1895, new_n1894);
xnor_3 g01520(new_n1897, new_n1896, new_n1893);
nand_4 g01521(new_n1898, new_n1858, new_n1852);
not_3  g01522(new_n1899, new_n1898);
nor_4  g01523(new_n1900, new_n1864, new_n1859);
nor_4  g01524(new_n1901, new_n1900, new_n1899);
xnor_3 g01525(new_n1902, new_n1901, new_n1897);
nand_4 g01526(new_n1903, new_n1873, new_n1866);
xnor_3 g01527(new_n1904, new_n1903, new_n1902);
nor_4  g01528(new_n1905, new_n1904, new_n1878);
not_3  g01529(new_n1906_1, new_n1878);
not_3  g01530(new_n1907, new_n1904);
nor_4  g01531(new_n1908, new_n1907, new_n1906_1);
nor_4  g01532(new_n1909, new_n1908, new_n1905);
xnor_3 g01533(new_n1910, new_n1909, new_n1877);
xnor_3 g01534(new_n1911, new_n1910, new_n1821);
nor_4  g01535(new_n1912, new_n1788, new_n1764);
nor_4  g01536(new_n1913, new_n1912, new_n1818);
xnor_3 g01537(new_n1914, new_n1847_1, new_n1834);
not_3  g01538(new_n1915, new_n1914);
not_3  g01539(new_n1916, new_n1755);
nor_4  g01540(new_n1917, new_n1762, new_n1916);
nor_4  g01541(new_n1918, new_n1917, new_n1764);
nor_4  g01542(new_n1919, new_n1918, new_n1915);
nor_4  g01543(new_n1920, new_n1294, new_n1293);
xnor_3 g01544(new_n1921, new_n1830, new_n1829);
not_3  g01545(new_n1922, new_n1921);
nor_4  g01546(new_n1923, new_n1922, new_n1920);
not_3  g01547(new_n1924, new_n1923);
not_3  g01548(new_n1925, new_n1920);
nor_4  g01549(new_n1926, new_n1921, new_n1925);
nor_4  g01550(new_n1927, new_n1926, new_n1923);
not_3  g01551(new_n1928, new_n1759);
xor_3  g01552(new_n1929, new_n1928, new_n1758);
nand_4 g01553(new_n1930, new_n1929, new_n1927);
nand_4 g01554(new_n1931, new_n1930, new_n1924);
not_3  g01555(new_n1932, new_n1293);
nor_4  g01556(new_n1933, new_n1836, new_n1932);
nor_4  g01557(new_n1934, new_n1933, new_n1828);
nor_4  g01558(new_n1935, new_n1838, new_n1932);
nor_4  g01559(new_n1936, new_n1935, new_n1934);
not_3  g01560(new_n1937, new_n1936);
nand_4 g01561(new_n1938, new_n1937, new_n1931);
not_3  g01562(new_n1939, new_n1938);
xnor_3 g01563(new_n1940, new_n1937, new_n1931);
nor_4  g01564(new_n1941, new_n1735, new_n1295);
nor_4  g01565(new_n1942, new_n1941, new_n1757);
nor_4  g01566(new_n1943, new_n1740, new_n1295);
nor_4  g01567(new_n1944, new_n1943, new_n1942);
nor_4  g01568(new_n1945, new_n1944, new_n1940);
nor_4  g01569(new_n1946, new_n1945, new_n1939);
not_3  g01570(new_n1947, new_n1918);
nor_4  g01571(new_n1948, new_n1947, new_n1914);
nor_4  g01572(new_n1949, new_n1948, new_n1919);
not_3  g01573(new_n1950, new_n1949);
nor_4  g01574(new_n1951, new_n1950, new_n1946);
nor_4  g01575(new_n1952, new_n1951, new_n1919);
nor_4  g01576(new_n1953, new_n1952, new_n1913);
not_3  g01577(new_n1954, new_n1876);
nor_4  g01578(new_n1955, new_n1954, new_n1848);
nor_4  g01579(new_n1956, new_n1955, new_n1877);
not_3  g01580(new_n1957, new_n1913);
not_3  g01581(new_n1958, new_n1919);
nor_4  g01582(new_n1959, new_n1937, new_n1931);
nor_4  g01583(new_n1960, new_n1959, new_n1939);
not_3  g01584(new_n1961, new_n1944);
nand_4 g01585(new_n1962, new_n1961, new_n1960);
nand_4 g01586(new_n1963, new_n1962, new_n1938);
nand_4 g01587(new_n1964, new_n1949, new_n1963);
nand_4 g01588(new_n1965, new_n1964, new_n1958);
xnor_3 g01589(new_n1966, new_n1965, new_n1957);
nor_4  g01590(new_n1967, new_n1966, new_n1956);
nor_4  g01591(new_n1968, new_n1967, new_n1953);
xnor_3 g01592(new_n1969, new_n1968, new_n1911);
nand_4 g01593(new_n1970, new_n1969, new_n1732);
xnor_3 g01594(new_n1971, new_n1969, new_n1731);
not_3  g01595(new_n1972, new_n1696);
nor_4  g01596(new_n1973, new_n1972, new_n1677);
nor_4  g01597(new_n1974, new_n1973, new_n1697);
not_3  g01598(new_n1975, new_n1974);
not_3  g01599(new_n1976, new_n1956);
xnor_3 g01600(new_n1977, new_n1966, new_n1976);
nor_4  g01601(new_n1978, new_n1977, new_n1975);
xnor_3 g01602(new_n1979, new_n1966, new_n1956);
xnor_3 g01603(new_n1980_1, new_n1979, new_n1974);
xor_3  g01604(new_n1981, new_n1676, new_n1654);
not_3  g01605(new_n1982, new_n1981);
nor_4  g01606(new_n1983, new_n1949, new_n1963);
nor_4  g01607(new_n1984, new_n1983, new_n1951);
nor_4  g01608(new_n1985, new_n1984, new_n1982);
xnor_3 g01609(new_n1986, new_n1984, new_n1982);
xnor_3 g01610(new_n1987, new_n1944, new_n1940);
not_3  g01611(new_n1988, new_n1987);
not_3  g01612(new_n1989, new_n1292);
nor_4  g01613(new_n1990, new_n1658_1, new_n1989);
nor_4  g01614(new_n1991, new_n1990, new_n1648);
nor_4  g01615(new_n1992, new_n1660, new_n1989);
nor_4  g01616(new_n1993, new_n1992, new_n1991);
not_3  g01617(new_n1994, new_n1993);
nor_4  g01618(new_n1995, new_n1994, new_n1988);
xor_3  g01619(new_n1996, new_n1994, new_n1988);
not_3  g01620(new_n1997, new_n1996);
xnor_3 g01621(new_n1998, new_n1929, new_n1927);
not_3  g01622(new_n1999, new_n1998);
xor_3  g01623(new_n2000, new_n1650, new_n1649);
not_3  g01624(new_n2001, new_n2000);
nor_4  g01625(new_n2002, new_n2001, new_n1999);
nor_4  g01626(new_n2003, new_n1296, new_n1292);
not_3  g01627(new_n2004, new_n2003);
xor_3  g01628(new_n2005, new_n2000, new_n1999);
nor_4  g01629(new_n2006, new_n2005, new_n2004);
nor_4  g01630(new_n2007, new_n2006, new_n2002);
nor_4  g01631(new_n2008, new_n2007, new_n1997);
nor_4  g01632(new_n2009, new_n2008, new_n1995);
nor_4  g01633(new_n2010, new_n2009, new_n1986);
nor_4  g01634(new_n2011, new_n2010, new_n1985);
nor_4  g01635(new_n2012, new_n2011, new_n1980_1);
nor_4  g01636(new_n2013, new_n2012, new_n1978);
nand_4 g01637(new_n2014, new_n2013, new_n1971);
nand_4 g01638(new_n2015, new_n2014, new_n1970);
not_3  g01639(new_n2016, new_n1726);
nand_4 g01640(new_n2017, new_n1715, new_n1712);
not_3  g01641(new_n2018, new_n2017);
nor_4  g01642(new_n2019, new_n2018, new_n1708);
not_3  g01643(new_n2020, new_n2019);
nand_4 g01644(new_n2021, n9400, n4928);
not_3  g01645(new_n2022, new_n2021);
nand_4 g01646(new_n2023, n4141, n2464);
nand_4 g01647(new_n2024_1, n8236, n6877);
nand_4 g01648(new_n2025, new_n2024_1, new_n2023);
not_3  g01649(new_n2026, new_n2023);
not_3  g01650(new_n2027, new_n2024_1);
nand_4 g01651(new_n2028, new_n2027, new_n2026);
nand_4 g01652(new_n2029, new_n2028, new_n2025);
xor_3  g01653(new_n2030, new_n2029, new_n2022);
xnor_3 g01654(new_n2031, new_n2030, new_n2020);
nor_4  g01655(new_n2032, new_n1706, new_n1705);
nand_4 g01656(new_n2033, n11311, n5105);
xnor_3 g01657(new_n2034, new_n2033, new_n2032);
nand_4 g01658(new_n2035, n7500, n4203);
not_3  g01659(new_n2036, new_n2035);
nand_4 g01660(new_n2037, n4187, n1209);
nand_4 g01661(new_n2038, n12753, n7354);
xnor_3 g01662(new_n2039, new_n2038, new_n2037);
xnor_3 g01663(new_n2040, new_n2039, new_n2036);
not_3  g01664(new_n2041, new_n2040);
xor_3  g01665(new_n2042, new_n2041, new_n2034);
xnor_3 g01666(new_n2043, new_n2042, new_n2031);
not_3  g01667(new_n2044, new_n2043);
nand_4 g01668(new_n2045, new_n1723, new_n1720);
nor_4  g01669(new_n2046, new_n1722, new_n1721);
nor_4  g01670(new_n2047, new_n1723, new_n1720);
nor_4  g01671(new_n2048, new_n2047, new_n1716);
xnor_3 g01672(new_n2049, new_n2048, new_n2046);
nand_4 g01673(new_n2050, new_n2049, new_n2045);
xnor_3 g01674(new_n2051, new_n2050, new_n2044);
xnor_3 g01675(new_n2052, new_n2051, new_n2016);
not_3  g01676(new_n2053, new_n1699);
nand_4 g01677(new_n2054, new_n1729, new_n2053);
nand_4 g01678(new_n2055, new_n1730, new_n1697);
nand_4 g01679(new_n2056, new_n2055, new_n2054);
xnor_3 g01680(new_n2057, new_n2056, new_n2052);
not_3  g01681(new_n2058, new_n2057);
not_3  g01682(new_n2059, new_n1811);
nand_4 g01683(new_n2060, new_n1814, new_n2059);
not_3  g01684(new_n2061, new_n1805);
nand_4 g01685(new_n2062, new_n2061, new_n1801);
not_3  g01686(new_n2063, new_n1809);
nand_4 g01687(new_n2064, new_n2063, new_n1806);
nand_4 g01688(new_n2065, new_n2064, new_n2062);
nand_4 g01689(new_n2066, n5814, n3992);
not_3  g01690(new_n2067, new_n2066);
nand_4 g01691(new_n2068, n12704, n8384);
nand_4 g01692(new_n2069, n7236, n4903);
xnor_3 g01693(new_n2070, new_n2069, new_n2068);
xor_3  g01694(new_n2071, new_n2070, new_n2067);
not_3  g01695(new_n2072, new_n2071);
xnor_3 g01696(new_n2073, new_n2072, new_n2065);
nor_4  g01697(new_n2074, new_n1808, new_n1807);
nand_4 g01698(new_n2075, n7294, n6358);
not_3  g01699(new_n2076, new_n2075);
xor_3  g01700(new_n2077, new_n2076, new_n2074);
nand_4 g01701(new_n2078, n10848, n1471);
nand_4 g01702(new_n2079, n5198, n1980);
nand_4 g01703(new_n2080, n8028, n7646);
not_3  g01704(new_n2081, new_n2080);
xor_3  g01705(new_n2082, new_n2081, new_n2079);
xnor_3 g01706(new_n2083, new_n2082, new_n2078);
not_3  g01707(new_n2084, new_n2083);
xnor_3 g01708(new_n2085, new_n2084, new_n2077);
xnor_3 g01709(new_n2086, new_n2085, new_n2073);
nand_4 g01710(new_n2087_1, new_n1799, new_n1796);
nor_4  g01711(new_n2088, new_n1798_1, new_n1797);
nor_4  g01712(new_n2089, new_n1810, new_n1800);
xnor_3 g01713(new_n2090, new_n2089, new_n2088);
nand_4 g01714(new_n2091, new_n2090, new_n2087_1);
xnor_3 g01715(new_n2092, new_n2091, new_n2086);
xnor_3 g01716(new_n2093, new_n2092, new_n2060);
nand_4 g01717(new_n2094, new_n1815, new_n1791);
not_3  g01718(new_n2095, new_n2094);
nor_4  g01719(new_n2096_1, new_n1817, new_n2095);
xnor_3 g01720(new_n2097, new_n2096_1, new_n2093);
not_3  g01721(new_n2098, new_n1905);
nand_4 g01722(new_n2099, new_n1909, new_n1877);
nand_4 g01723(new_n2100, new_n2099, new_n2098);
nor_4  g01724(new_n2101, new_n1903, new_n1902);
not_3  g01725(new_n2102, new_n2101);
not_3  g01726(new_n2103, new_n1883);
nand_4 g01727(new_n2104, new_n1891, new_n1887);
nand_4 g01728(new_n2105, new_n2104, new_n2103);
nand_4 g01729(new_n2106, n11478, n5069);
not_3  g01730(new_n2107, new_n2106);
nand_4 g01731(new_n2108, n6806, n5283);
nand_4 g01732(new_n2109, n12044, n4805);
nand_4 g01733(new_n2110, new_n2109, new_n2108);
not_3  g01734(new_n2111, new_n2108);
not_3  g01735(new_n2112, new_n2109);
nand_4 g01736(new_n2113, new_n2112, new_n2111);
nand_4 g01737(new_n2114, new_n2113, new_n2110);
xor_3  g01738(new_n2115, new_n2114, new_n2107);
xnor_3 g01739(new_n2116, new_n2115, new_n2105);
nor_4  g01740(new_n2117, new_n1881, new_n1880);
nand_4 g01741(new_n2118, n2802, n137);
not_3  g01742(new_n2119, new_n2118);
xor_3  g01743(new_n2120, new_n2119, new_n2117);
nand_4 g01744(new_n2121, n6797, n1512);
not_3  g01745(new_n2122, new_n2121);
nand_4 g01746(new_n2123, n6294, n533);
nand_4 g01747(new_n2124, n3146, n1564);
xnor_3 g01748(new_n2125, new_n2124, new_n2123);
xor_3  g01749(new_n2126, new_n2125, new_n2122);
not_3  g01750(new_n2127, new_n2126);
nor_4  g01751(new_n2128, new_n2127, new_n2120);
not_3  g01752(new_n2129, new_n2120);
nor_4  g01753(new_n2130, new_n2126, new_n2129);
nor_4  g01754(new_n2131_1, new_n2130, new_n2128);
xnor_3 g01755(new_n2132, new_n2131_1, new_n2116);
nand_4 g01756(new_n2133, new_n1896, new_n1893);
nor_4  g01757(new_n2134, new_n1895, new_n1894);
xnor_3 g01758(new_n2135, new_n1896, new_n1892);
not_3  g01759(new_n2136, new_n1901);
nand_4 g01760(new_n2137, new_n2136, new_n2135);
not_3  g01761(new_n2138, new_n2137);
xnor_3 g01762(new_n2139, new_n2138, new_n2134);
nand_4 g01763(new_n2140, new_n2139, new_n2133);
xnor_3 g01764(new_n2141, new_n2140, new_n2132);
xnor_3 g01765(new_n2142, new_n2141, new_n2102);
xnor_3 g01766(new_n2143, new_n2142, new_n2100);
xnor_3 g01767(new_n2144, new_n2143, new_n2097);
not_3  g01768(new_n2145, new_n1821);
nand_4 g01769(new_n2146, new_n1910, new_n2145);
not_3  g01770(new_n2147, new_n1968);
nand_4 g01771(new_n2148, new_n2147, new_n1911);
nand_4 g01772(new_n2149, new_n2148, new_n2146);
xnor_3 g01773(new_n2150, new_n2149, new_n2144);
xnor_3 g01774(new_n2151, new_n2150, new_n2058);
xnor_3 g01775(new_n2152, new_n2151, new_n2015);
nand_4 g01776(new_n2153, new_n2152, new_n1641);
xnor_3 g01777(new_n2154, new_n2152, new_n1640);
xor_3  g01778(new_n2155, new_n1637, new_n1634);
xnor_3 g01779(new_n2156, new_n2013, new_n1971);
nand_4 g01780(new_n2157, new_n2156, new_n2155);
not_3  g01781(new_n2158, new_n1630);
xor_3  g01782(new_n2159, new_n1633, new_n2158);
not_3  g01783(new_n2160, new_n2159);
not_3  g01784(new_n2161, new_n1980_1);
xnor_3 g01785(new_n2162, new_n2011, new_n2161);
nor_4  g01786(new_n2163, new_n2162, new_n2160);
xnor_3 g01787(new_n2164, new_n2162, new_n2160);
xor_3  g01788(new_n2165, new_n1629, new_n1626);
not_3  g01789(new_n2166, new_n1986);
xnor_3 g01790(new_n2167, new_n2009, new_n2166);
nor_4  g01791(new_n2168, new_n2167, new_n2165);
xnor_3 g01792(new_n2169, new_n2007, new_n1996);
not_3  g01793(new_n2170, new_n1291);
nor_4  g01794(new_n2171, new_n1530, new_n2170);
nor_4  g01795(new_n2172, new_n2171, new_n1621);
nor_4  g01796(new_n2173, new_n1535, new_n2170);
nor_4  g01797(new_n2174, new_n2173, new_n2172);
nor_4  g01798(new_n2175, new_n2174, new_n2169);
xnor_3 g01799(new_n2176, new_n2174, new_n2169);
nor_4  g01800(new_n2177, new_n1298, new_n1291);
xor_3  g01801(new_n2178, new_n1623, new_n1622);
nor_4  g01802(new_n2179, new_n2178, new_n2177);
xnor_3 g01803(new_n2180, new_n2005, new_n2003);
not_3  g01804(new_n2181, new_n2178);
xor_3  g01805(new_n2182, new_n2181, new_n2177);
nor_4  g01806(new_n2183, new_n2182, new_n2180);
nor_4  g01807(new_n2184, new_n2183, new_n2179);
nor_4  g01808(new_n2185, new_n2184, new_n2176);
nor_4  g01809(new_n2186, new_n2185, new_n2175);
xnor_3 g01810(new_n2187, new_n2167, new_n2165);
nor_4  g01811(new_n2188, new_n2187, new_n2186);
nor_4  g01812(new_n2189, new_n2188, new_n2168);
nor_4  g01813(new_n2190, new_n2189, new_n2164);
nor_4  g01814(new_n2191, new_n2190, new_n2163);
not_3  g01815(new_n2192, new_n2155);
xnor_3 g01816(new_n2193, new_n2156, new_n2192);
nand_4 g01817(new_n2194, new_n2193, new_n2191);
nand_4 g01818(new_n2195, new_n2194, new_n2157);
nand_4 g01819(new_n2196, new_n2195, new_n2154);
nand_4 g01820(new_n2197, new_n2196, new_n2153);
nand_4 g01821(new_n2198, new_n2076, new_n2074);
nand_4 g01822(new_n2199, new_n2084, new_n2077);
nand_4 g01823(new_n2200, new_n2199, new_n2198);
nand_4 g01824(new_n2201, new_n2025, new_n2022);
nand_4 g01825(new_n2202, new_n2201, new_n2028);
nand_4 g01826(new_n2203, n6294, n2802);
nand_4 g01827(new_n2204, n6797, n533);
xor_3  g01828(new_n2205, new_n2204, new_n2203);
xor_3  g01829(new_n2206, new_n2205, new_n2202);
xor_3  g01830(new_n2207, new_n2206, new_n2200);
nand_4 g01831(new_n2208, new_n2143, new_n2097);
not_3  g01832(new_n2209, new_n2097);
xnor_3 g01833(new_n2210, new_n2143, new_n2209);
nand_4 g01834(new_n2211, new_n2149, new_n2210);
nand_4 g01835(new_n2212, new_n2211, new_n2208);
not_3  g01836(new_n2213, new_n1581);
nand_4 g01837(new_n2214, new_n1614, new_n2213);
nand_4 g01838(new_n2215, new_n1639, new_n1615);
nand_4 g01839(new_n2216, new_n2215, new_n2214);
nand_4 g01840(new_n2217, new_n2051, new_n1726);
nand_4 g01841(new_n2218, new_n2056, new_n2052);
nand_4 g01842(new_n2219, new_n2218, new_n2217);
xnor_3 g01843(new_n2220, new_n2219, new_n2216);
xnor_3 g01844(new_n2221, new_n2220, new_n2212);
not_3  g01845(new_n2222, new_n2105);
nand_4 g01846(new_n2223, new_n2115, new_n2222);
not_3  g01847(new_n2224, new_n2131_1);
nand_4 g01848(new_n2225, new_n2224, new_n2116);
nand_4 g01849(new_n2226_1, new_n2225, new_n2223);
nand_4 g01850(new_n2227, new_n2119, new_n2117);
nand_4 g01851(new_n2228, new_n2127, new_n2120);
nand_4 g01852(new_n2229, new_n2228, new_n2227);
nand_4 g01853(new_n2230, n6826, n6038);
not_3  g01854(new_n2231, new_n2230);
nand_4 g01855(new_n2232, new_n2110, new_n2107);
nand_4 g01856(new_n2233, new_n2232, new_n2113);
xor_3  g01857(new_n2234, new_n2233, new_n2231);
xor_3  g01858(new_n2235, new_n2234, new_n2229);
xnor_3 g01859(new_n2236, new_n2235, new_n2226_1);
nand_4 g01860(new_n2237, new_n2030, new_n2019);
nand_4 g01861(new_n2238, new_n2042, new_n2031);
nand_4 g01862(new_n2239, new_n2238, new_n2237);
nand_4 g01863(new_n2240, n5283, n5069);
nand_4 g01864(new_n2241, n4928, n2464);
not_3  g01865(new_n2242, new_n2241);
xor_3  g01866(new_n2243, new_n2242, new_n2240);
xnor_3 g01867(new_n2244, new_n2243, new_n2239);
xnor_3 g01868(new_n2245, new_n2244, new_n2236);
nand_4 g01869(new_n2246, new_n2138, new_n2134);
not_3  g01870(new_n2247, new_n2132);
nand_4 g01871(new_n2248, new_n2140, new_n2247);
nand_4 g01872(new_n2249, new_n2248, new_n2246);
not_3  g01873(new_n2250, new_n2079);
nor_4  g01874(new_n2251, new_n2081, new_n2250);
not_3  g01875(new_n2252, new_n2078);
nor_4  g01876(new_n2253_1, new_n2082, new_n2252);
nor_4  g01877(new_n2254, new_n2253_1, new_n2251);
nand_4 g01878(new_n2255, n10848, n7646);
not_3  g01879(new_n2256, new_n2255);
nand_4 g01880(new_n2257, n6806, n137);
nand_4 g01881(new_n2258, n8384, n5814);
xor_3  g01882(new_n2259, new_n2258, new_n2257);
xor_3  g01883(new_n2260, new_n2259, new_n2256);
xnor_3 g01884(new_n2261, new_n2260, new_n2254);
xnor_3 g01885(new_n2262, new_n2261, new_n2249);
xnor_3 g01886(new_n2263, new_n2262, new_n2245);
nand_4 g01887(new_n2264, new_n2141, new_n2101);
nand_4 g01888(new_n2265, new_n2142, new_n2100);
nand_4 g01889(new_n2266, new_n2265, new_n2264);
nand_4 g01890(new_n2267, new_n1584, new_n1583);
nand_4 g01891(new_n2268, new_n1612, new_n1586);
nand_4 g01892(new_n2269, new_n2268, new_n2267);
nand_4 g01893(new_n2270, new_n2089, new_n2088);
nand_4 g01894(new_n2271, new_n2091, new_n2086);
nand_4 g01895(new_n2272, new_n2271, new_n2270);
xnor_3 g01896(new_n2273, new_n2272, new_n2269);
nand_4 g01897(new_n2274, new_n2048, new_n2046);
nand_4 g01898(new_n2275, new_n2050, new_n2043);
nand_4 g01899(new_n2276, new_n2275, new_n2274);
nor_4  g01900(new_n2277, new_n1610, new_n1601);
nor_4  g01901(new_n2278_1, new_n1611, new_n1598);
nor_4  g01902(new_n2279, new_n2278_1, new_n2277);
and_4  g01903(new_n2280, new_n1594, new_n1593);
nor_4  g01904(new_n2281, new_n1595, new_n1592);
nor_4  g01905(new_n2282, new_n2281, new_n2280);
nand_4 g01906(new_n2283, n12706, n1333);
nand_4 g01907(new_n2284, n5240, n2508);
nand_4 g01908(new_n2285, n4005, n3172);
xnor_3 g01909(new_n2286, new_n2285, new_n2284);
xnor_3 g01910(new_n2287, new_n2286, new_n2283);
xnor_3 g01911(new_n2288, new_n2287, new_n2282);
and_4  g01912(new_n2289, new_n2038, new_n2037);
nor_4  g01913(new_n2290, new_n2039, new_n2036);
nor_4  g01914(new_n2291, new_n2290, new_n2289);
nand_4 g01915(new_n2292, n4203, n1209);
nand_4 g01916(new_n2293, n9400, n8236);
nand_4 g01917(new_n2294, n5105, n4187);
xnor_3 g01918(new_n2295, new_n2294, new_n2293);
xnor_3 g01919(new_n2296, new_n2295, new_n2292);
xnor_3 g01920(new_n2297, new_n2296, new_n2291);
xnor_3 g01921(new_n2298, new_n2297, new_n2288);
nand_4 g01922(new_n2299, n12720, n11821);
nand_4 g01923(new_n2300, n6877, n783);
xnor_3 g01924(new_n2301_1, new_n2300, new_n2299);
nand_4 g01925(new_n2302, n9080, n2509);
nand_4 g01926(new_n2303, n11757, n2585);
xnor_3 g01927(new_n2304, new_n2303, new_n2302);
xnor_3 g01928(new_n2305, new_n2304, new_n2301_1);
not_3  g01929(new_n2306, new_n1602);
nand_4 g01930(new_n2307, new_n1605, new_n2306);
nand_4 g01931(new_n2308, new_n2307, new_n1608);
nand_4 g01932(new_n2309, n12753, n7500);
nand_4 g01933(new_n2310, n10174, n7354);
xnor_3 g01934(new_n2311, new_n2310, new_n2309);
xnor_3 g01935(new_n2312, new_n2311, new_n2308);
xnor_3 g01936(new_n2313, new_n2312, new_n2305);
xnor_3 g01937(new_n2314, new_n2313, new_n2298);
and_4  g01938(new_n2315, new_n2124, new_n2123);
nor_4  g01939(new_n2316_1, new_n2125, new_n2122);
nor_4  g01940(new_n2317, new_n2316_1, new_n2315);
nand_4 g01941(new_n2318, n11311, n4141);
nand_4 g01942(new_n2319, n12044, n11478);
nand_4 g01943(new_n2320, n7862, n615);
xnor_3 g01944(new_n2321, new_n2320, new_n2319);
xnor_3 g01945(new_n2322, new_n2321, new_n2318);
xnor_3 g01946(new_n2323, new_n2322, new_n2317);
nand_4 g01947(new_n2324, n1980, n1471);
not_3  g01948(new_n2325, new_n2033);
nand_4 g01949(new_n2326, new_n2325, new_n2032);
nand_4 g01950(new_n2327, new_n2040, new_n2034);
nand_4 g01951(new_n2328, new_n2327, new_n2326);
xnor_3 g01952(new_n2329, new_n2328, new_n2324);
xnor_3 g01953(new_n2330, new_n2329, new_n2323);
xnor_3 g01954(new_n2331, new_n2330, new_n2314);
xnor_3 g01955(new_n2332, new_n2331, new_n2279);
xnor_3 g01956(new_n2333, new_n2332, new_n2276);
nand_4 g01957(new_n2334, n8028, n4722);
not_3  g01958(new_n2335, new_n2334);
nand_4 g01959(new_n2336, new_n2071, new_n2065);
nand_4 g01960(new_n2337, new_n2085, new_n2073);
nand_4 g01961(new_n2338, new_n2337, new_n2336);
nand_4 g01962(new_n2339, n3146, n1512);
not_3  g01963(new_n2340, new_n2339);
nand_4 g01964(new_n2341, n5694, n4805);
nand_4 g01965(new_n2342, n4903, n3992);
xnor_3 g01966(new_n2343, new_n2342, new_n2341);
nand_4 g01967(new_n2344, n4938, n1564);
nand_4 g01968(new_n2345, n12704, n6358);
xnor_3 g01969(new_n2346, new_n2345, new_n2344);
xnor_3 g01970(new_n2347_1, new_n2346, new_n2343);
xnor_3 g01971(new_n2348, new_n2347_1, new_n2340);
nand_4 g01972(new_n2349, n7294, n5198);
not_3  g01973(new_n2350, new_n2349);
and_4  g01974(new_n2351, new_n2069, new_n2068);
nor_4  g01975(new_n2352, new_n2070, new_n2067);
nor_4  g01976(new_n2353, new_n2352, new_n2351);
xnor_3 g01977(new_n2354, new_n2353, new_n2350);
xnor_3 g01978(new_n2355, new_n2354, new_n2348);
nand_4 g01979(new_n2356, n7236, n1906);
nand_4 g01980(new_n2357, new_n1589, new_n1587);
nand_4 g01981(new_n2358, new_n1596, new_n1590);
nand_4 g01982(new_n2359, new_n2358, new_n2357);
xnor_3 g01983(new_n2360, new_n2359, new_n2356);
xnor_3 g01984(new_n2361, new_n2360, new_n2355);
xnor_3 g01985(new_n2362, new_n2361, new_n2338);
xnor_3 g01986(new_n2363, new_n2362, new_n2335);
xnor_3 g01987(new_n2364, new_n2363, new_n2333);
xnor_3 g01988(new_n2365, new_n2364, new_n2273);
xnor_3 g01989(new_n2366, new_n2365, new_n2266);
xnor_3 g01990(new_n2367, new_n2366, new_n2263);
xnor_3 g01991(new_n2368, new_n2367, new_n2221);
xnor_3 g01992(new_n2369, new_n2368, new_n2207);
nor_4  g01993(new_n2370, new_n2092, new_n2060);
nor_4  g01994(new_n2371, new_n2096_1, new_n2093);
nor_4  g01995(new_n2372, new_n2371, new_n2370);
nand_4 g01996(new_n2373, new_n2150, new_n2057);
nand_4 g01997(new_n2374, new_n2151, new_n2015);
nand_4 g01998(new_n2375, new_n2374, new_n2373);
xnor_3 g01999(new_n2376, new_n2375, new_n2372);
xnor_3 g02000(new_n2377, new_n2376, new_n2369);
xnor_3 g02001(n671, new_n2377, new_n2197);
nand_4 g02002(new_n2379, n5964, n2577);
nand_4 g02003(new_n2380, n3842, n1097);
nor_4  g02004(new_n2381, new_n2380, new_n2379);
nand_4 g02005(new_n2382, n11917, n4312);
nand_4 g02006(new_n2383_1, n12705, n4921);
nand_4 g02007(new_n2384, n12025, n9956);
xnor_3 g02008(new_n2385, new_n2384, new_n2383_1);
xnor_3 g02009(new_n2386, new_n2385, new_n2382);
nand_4 g02010(new_n2387, n12705, n9956);
not_3  g02011(new_n2388, new_n2387);
nand_4 g02012(new_n2389, n11917, n1097);
not_3  g02013(new_n2390, new_n2389);
nor_4  g02014(new_n2391, new_n2390, new_n2388);
nor_4  g02015(new_n2392, new_n2389, new_n2387);
nand_4 g02016(new_n2393_1, n4921, n4312);
not_3  g02017(new_n2394, new_n2393_1);
nor_4  g02018(new_n2395, new_n2394, new_n2392);
nor_4  g02019(new_n2396, new_n2395, new_n2391);
xnor_3 g02020(new_n2397, new_n2396, new_n2386);
xor_3  g02021(new_n2398, new_n2380, new_n2379);
xnor_3 g02022(new_n2399, new_n2398, new_n2397);
nand_4 g02023(new_n2400, n5964, n3842);
not_3  g02024(new_n2401, new_n2400);
nand_4 g02025(new_n2402, n9956, n4312);
not_3  g02026(new_n2403, new_n2402);
nand_4 g02027(new_n2404, n11917, n5964);
not_3  g02028(new_n2405, new_n2404);
nor_4  g02029(new_n2406, new_n2405, new_n2403);
nor_4  g02030(new_n2407, new_n2404, new_n2402);
nand_4 g02031(new_n2408, n4921, n1097);
not_3  g02032(new_n2409, new_n2408);
nor_4  g02033(new_n2410, new_n2409, new_n2407);
nor_4  g02034(new_n2411, new_n2410, new_n2406);
nand_4 g02035(new_n2412, new_n2411, new_n2401);
not_3  g02036(new_n2413, new_n2412);
nor_4  g02037(new_n2414, new_n2411, new_n2401);
nor_4  g02038(new_n2415, new_n2414, new_n2413);
not_3  g02039(new_n2416, new_n2391);
not_3  g02040(new_n2417, new_n2392);
nand_4 g02041(new_n2418, new_n2417, new_n2416);
xnor_3 g02042(new_n2419, new_n2418, new_n2393_1);
not_3  g02043(new_n2420, new_n2419);
nand_4 g02044(new_n2421, new_n2420, new_n2415);
nand_4 g02045(new_n2422, new_n2421, new_n2412);
not_3  g02046(new_n2423, new_n2422);
nor_4  g02047(new_n2424, new_n2423, new_n2399);
and_4  g02048(new_n2425_1, new_n2424, new_n2381);
nand_4 g02049(new_n2426, new_n2385, new_n2382);
not_3  g02050(new_n2427, new_n2386);
not_3  g02051(new_n2428, new_n2396);
nand_4 g02052(new_n2429, new_n2428, new_n2427);
and_4  g02053(new_n2430, new_n2429, new_n2426);
nand_4 g02054(new_n2431_1, n9637, n5964);
not_3  g02055(new_n2432, new_n2431_1);
nand_4 g02056(new_n2433_1, n2577, n1097);
nand_4 g02057(new_n2434_1, n5305, n1835);
xnor_3 g02058(new_n2435, new_n2434_1, new_n2433_1);
xor_3  g02059(new_n2436, new_n2435, new_n2432);
xnor_3 g02060(new_n2437, new_n2436, new_n2430);
not_3  g02061(new_n2438, new_n2437);
nor_4  g02062(new_n2439, new_n2384, new_n2383_1);
not_3  g02063(new_n2440, new_n2439);
nand_4 g02064(new_n2441, n4312, n3842);
xor_3  g02065(new_n2442, new_n2441, new_n2440);
not_3  g02066(new_n2443, new_n2442);
nand_4 g02067(new_n2444, n12025, n4921);
not_3  g02068(new_n2445, new_n2444);
nand_4 g02069(new_n2446, n12705, n11917);
nand_4 g02070(new_n2447, n11257, n9956);
xnor_3 g02071(new_n2448, new_n2447, new_n2446);
and_4  g02072(new_n2449, new_n2448, new_n2445);
nor_4  g02073(new_n2450, new_n2448, new_n2445);
nor_4  g02074(new_n2451, new_n2450, new_n2449);
xnor_3 g02075(new_n2452, new_n2451, new_n2443);
xnor_3 g02076(new_n2453, new_n2452, new_n2438);
not_3  g02077(new_n2454, new_n2453);
nand_4 g02078(new_n2455, new_n2398, new_n2397);
xnor_3 g02079(new_n2456, new_n2424, new_n2381);
nand_4 g02080(new_n2457, new_n2456, new_n2455);
and_4  g02081(new_n2458, new_n2457, new_n2454);
nor_4  g02082(new_n2459, new_n2458, new_n2425_1);
nand_4 g02083(new_n2460, n8759, n8065);
not_3  g02084(new_n2461, new_n2460);
nand_4 g02085(new_n2462, n7436, n6126);
nand_4 g02086(new_n2463, n8276, n3602);
nand_4 g02087(new_n2464_1, n9241, n3719);
xnor_3 g02088(new_n2465, new_n2464_1, new_n2463);
nor_4  g02089(new_n2466, new_n2465, new_n2462);
not_3  g02090(new_n2467, new_n2462);
not_3  g02091(new_n2468, new_n2465);
nor_4  g02092(new_n2469, new_n2468, new_n2467);
nor_4  g02093(new_n2470, new_n2469, new_n2466);
nand_4 g02094(new_n2471, n8276, n3719);
not_3  g02095(new_n2472, new_n2471);
nand_4 g02096(new_n2473, n12299, n6126);
not_3  g02097(new_n2474, new_n2473);
nor_4  g02098(new_n2475, new_n2474, new_n2472);
nor_4  g02099(new_n2476, new_n2473, new_n2471);
nand_4 g02100(new_n2477, n7436, n3602);
not_3  g02101(new_n2478, new_n2477);
nor_4  g02102(new_n2479, new_n2478, new_n2476);
nor_4  g02103(new_n2480, new_n2479, new_n2475);
xnor_3 g02104(new_n2481, new_n2480, new_n2470);
nand_4 g02105(new_n2482, n10439, n6776);
nand_4 g02106(new_n2483, n12299, n8595);
xor_3  g02107(new_n2484, new_n2483, new_n2482);
xnor_3 g02108(new_n2485, new_n2484, new_n2481);
nand_4 g02109(new_n2486, n8595, n6776);
not_3  g02110(new_n2487, new_n2486);
nand_4 g02111(new_n2488, n7436, n3719);
not_3  g02112(new_n2489, new_n2488);
nand_4 g02113(new_n2490, n6776, n6126);
not_3  g02114(new_n2491, new_n2490);
nor_4  g02115(new_n2492, new_n2491, new_n2489);
nor_4  g02116(new_n2493, new_n2490, new_n2488);
nand_4 g02117(new_n2494, n12299, n3602);
not_3  g02118(new_n2495, new_n2494);
nor_4  g02119(new_n2496, new_n2495, new_n2493);
nor_4  g02120(new_n2497, new_n2496, new_n2492);
nand_4 g02121(new_n2498_1, new_n2497, new_n2487);
not_3  g02122(new_n2499, new_n2498_1);
xnor_3 g02123(new_n2500, new_n2497, new_n2487);
nor_4  g02124(new_n2501, new_n2476, new_n2475);
xnor_3 g02125(new_n2502, new_n2501, new_n2478);
nor_4  g02126(new_n2503, new_n2502, new_n2500);
nor_4  g02127(new_n2504, new_n2503, new_n2499);
not_3  g02128(new_n2505, new_n2504);
nand_4 g02129(new_n2506, new_n2505, new_n2485);
not_3  g02130(new_n2507_1, new_n2506);
nor_4  g02131(new_n2508_1, new_n2505, new_n2485);
nor_4  g02132(new_n2509_1, new_n2508_1, new_n2507_1);
not_3  g02133(new_n2510, new_n2509_1);
nand_4 g02134(new_n2511, n10439, n8759);
not_3  g02135(new_n2512_1, new_n2511);
xnor_3 g02136(new_n2513, new_n2502, new_n2500);
not_3  g02137(new_n2514, new_n2513);
nor_4  g02138(new_n2515_1, new_n2514, new_n2512_1);
not_3  g02139(new_n2516, new_n2515_1);
nor_4  g02140(new_n2517, new_n2513, new_n2511);
nor_4  g02141(new_n2518, new_n2517, new_n2515_1);
nand_4 g02142(new_n2519, n8759, n8595);
nand_4 g02143(new_n2520, n12299, n3719);
not_3  g02144(new_n2521, new_n2520);
nand_4 g02145(new_n2522_1, n8759, n6126);
not_3  g02146(new_n2523, new_n2522_1);
nand_4 g02147(new_n2524, new_n2523, new_n2521);
nand_4 g02148(new_n2525, new_n2522_1, new_n2520);
nand_4 g02149(new_n2526, n6776, n3602);
not_3  g02150(new_n2527, new_n2526);
nand_4 g02151(new_n2528, new_n2527, new_n2525);
nand_4 g02152(new_n2529, new_n2528, new_n2524);
not_3  g02153(new_n2530_1, new_n2529);
nor_4  g02154(new_n2531, new_n2530_1, new_n2519);
xor_3  g02155(new_n2532, new_n2529, new_n2519);
nor_4  g02156(new_n2533, new_n2493, new_n2492);
xor_3  g02157(new_n2534, new_n2533, new_n2494);
nor_4  g02158(new_n2535, new_n2534, new_n2532);
nor_4  g02159(new_n2536, new_n2535, new_n2531);
nand_4 g02160(new_n2537, new_n2536, new_n2518);
nand_4 g02161(new_n2538, new_n2537, new_n2516);
nor_4  g02162(new_n2539, new_n2538, new_n2510);
not_3  g02163(new_n2540, new_n2538);
nor_4  g02164(new_n2541, new_n2540, new_n2509_1);
nor_4  g02165(new_n2542, new_n2541, new_n2539);
nand_4 g02166(new_n2543, new_n2542, new_n2461);
and_4  g02167(new_n2544, new_n2525, new_n2524);
nand_4 g02168(new_n2545, n6776, n3719);
nand_4 g02169(new_n2546, n8759, n3602);
nor_4  g02170(new_n2547, new_n2546, new_n2545);
not_3  g02171(new_n2548, new_n2547);
nor_4  g02172(new_n2549, new_n2548, new_n2544);
not_3  g02173(new_n2550, new_n2549);
xnor_3 g02174(new_n2551_1, new_n2534, new_n2532);
nor_4  g02175(new_n2552, new_n2551_1, new_n2550);
not_3  g02176(new_n2553, new_n2552);
xnor_3 g02177(new_n2554, new_n2536, new_n2518);
not_3  g02178(new_n2555, new_n2554);
nor_4  g02179(new_n2556, new_n2555, new_n2553);
xnor_3 g02180(new_n2557, new_n2542, new_n2460);
nand_4 g02181(new_n2558_1, new_n2557, new_n2556);
nand_4 g02182(new_n2559, new_n2558_1, new_n2543);
not_3  g02183(new_n2560, new_n2466);
nand_4 g02184(new_n2561, new_n2480, new_n2470);
nand_4 g02185(new_n2562, new_n2561, new_n2560);
nand_4 g02186(new_n2563, n8065, n6776);
nand_4 g02187(new_n2564_1, n12299, n10439);
nand_4 g02188(new_n2565, n10391, n8759);
not_3  g02189(new_n2566, new_n2565);
xor_3  g02190(new_n2567, new_n2566, new_n2564_1);
xnor_3 g02191(new_n2568, new_n2567, new_n2563);
not_3  g02192(new_n2569, new_n2568);
xor_3  g02193(new_n2570, new_n2569, new_n2562);
nor_4  g02194(new_n2571, new_n2464_1, new_n2463);
not_3  g02195(new_n2572, new_n2571);
nand_4 g02196(new_n2573, n8595, n7436);
xor_3  g02197(new_n2574, new_n2573, new_n2572);
nand_4 g02198(new_n2575, n9241, n3602);
not_3  g02199(new_n2576, new_n2575);
nand_4 g02200(new_n2577_1, n8276, n6126);
nand_4 g02201(new_n2578, n10510, n3719);
xor_3  g02202(new_n2579, new_n2578, new_n2577_1);
xnor_3 g02203(new_n2580, new_n2579, new_n2576);
xnor_3 g02204(new_n2581_1, new_n2580, new_n2574);
xnor_3 g02205(new_n2582, new_n2581_1, new_n2570);
not_3  g02206(new_n2583, new_n2481);
nand_4 g02207(new_n2584, new_n2484, new_n2583);
nor_4  g02208(new_n2585_1, new_n2483, new_n2482);
xnor_3 g02209(new_n2586, new_n2507_1, new_n2585_1);
nand_4 g02210(new_n2587, new_n2586, new_n2584);
xnor_3 g02211(new_n2588, new_n2587, new_n2582);
xnor_3 g02212(new_n2589, new_n2588, new_n2539);
xnor_3 g02213(new_n2590, new_n2589, new_n2559);
nand_4 g02214(new_n2591, n12648, n4826);
nand_4 g02215(new_n2592, n10545, n7733);
nand_4 g02216(new_n2593, n12925, n7690);
xnor_3 g02217(new_n2594, new_n2593, new_n2592);
nor_4  g02218(new_n2595, new_n2594, new_n2591);
not_3  g02219(new_n2596, new_n2591);
not_3  g02220(new_n2597, new_n2594);
nor_4  g02221(new_n2598, new_n2597, new_n2596);
nor_4  g02222(new_n2599, new_n2598, new_n2595);
nand_4 g02223(new_n2600, n12925, n10545);
not_3  g02224(new_n2601, new_n2600);
nand_4 g02225(new_n2602, n4826, n2530);
not_3  g02226(new_n2603, new_n2602);
nor_4  g02227(new_n2604, new_n2603, new_n2601);
nand_4 g02228(new_n2605, n12648, n7733);
not_3  g02229(new_n2606, new_n2605);
xnor_3 g02230(new_n2607, new_n2602, new_n2600);
nor_4  g02231(new_n2608, new_n2607, new_n2606);
nor_4  g02232(new_n2609, new_n2608, new_n2604);
xnor_3 g02233(new_n2610, new_n2609, new_n2599);
nand_4 g02234(new_n2611, n8476, n4970);
nand_4 g02235(new_n2612, n7610, n2530);
xor_3  g02236(new_n2613, new_n2612, new_n2611);
xnor_3 g02237(new_n2614, new_n2613, new_n2610);
nand_4 g02238(new_n2615, n8476, n7610);
not_3  g02239(new_n2616, new_n2615);
nand_4 g02240(new_n2617, n12925, n12648);
not_3  g02241(new_n2618, new_n2617);
nand_4 g02242(new_n2619, n8476, n4826);
not_3  g02243(new_n2620, new_n2619);
nor_4  g02244(new_n2621, new_n2620, new_n2618);
nand_4 g02245(new_n2622, n7733, n2530);
not_3  g02246(new_n2623, new_n2622);
xnor_3 g02247(new_n2624_1, new_n2619, new_n2617);
nor_4  g02248(new_n2625, new_n2624_1, new_n2623);
nor_4  g02249(new_n2626, new_n2625, new_n2621);
nand_4 g02250(new_n2627, new_n2626, new_n2616);
not_3  g02251(new_n2628, new_n2627);
nor_4  g02252(new_n2629, new_n2626, new_n2616);
nor_4  g02253(new_n2630, new_n2629, new_n2628);
xnor_3 g02254(new_n2631, new_n2607, new_n2605);
not_3  g02255(new_n2632, new_n2631);
nand_4 g02256(new_n2633, new_n2632, new_n2630);
nand_4 g02257(new_n2634, new_n2633, new_n2627);
xnor_3 g02258(new_n2635, new_n2634, new_n2614);
nand_4 g02259(new_n2636, n5331, n4970);
not_3  g02260(new_n2637, new_n2636);
nand_4 g02261(new_n2638, n7610, n5331);
not_3  g02262(new_n2639, new_n2638);
nand_4 g02263(new_n2640, n12925, n2530);
not_3  g02264(new_n2641, new_n2640);
nand_4 g02265(new_n2642, n5331, n4826);
not_3  g02266(new_n2643, new_n2642);
nor_4  g02267(new_n2644, new_n2643, new_n2641);
nor_4  g02268(new_n2645, new_n2642, new_n2640);
nand_4 g02269(new_n2646, n8476, n7733);
not_3  g02270(new_n2647, new_n2646);
nor_4  g02271(new_n2648, new_n2647, new_n2645);
nor_4  g02272(new_n2649, new_n2648, new_n2644);
nand_4 g02273(new_n2650, new_n2649, new_n2639);
not_3  g02274(new_n2651, new_n2650);
nor_4  g02275(new_n2652, new_n2649, new_n2639);
nor_4  g02276(new_n2653, new_n2652, new_n2651);
xnor_3 g02277(new_n2654, new_n2624_1, new_n2622);
not_3  g02278(new_n2655, new_n2654);
nand_4 g02279(new_n2656, new_n2655, new_n2653);
nand_4 g02280(new_n2657, new_n2656, new_n2650);
nor_4  g02281(new_n2658, new_n2657, new_n2637);
not_3  g02282(new_n2659, new_n2658);
xnor_3 g02283(new_n2660, new_n2632, new_n2630);
not_3  g02284(new_n2661, new_n2657);
nor_4  g02285(new_n2662, new_n2661, new_n2636);
nor_4  g02286(new_n2663, new_n2662, new_n2658);
nand_4 g02287(new_n2664, new_n2663, new_n2660);
nand_4 g02288(new_n2665, new_n2664, new_n2659);
nor_4  g02289(new_n2666, new_n2665, new_n2635);
not_3  g02290(new_n2667, new_n2610);
nand_4 g02291(new_n2668, new_n2613, new_n2667);
nor_4  g02292(new_n2669, new_n2612, new_n2611);
nand_4 g02293(new_n2670, new_n2634, new_n2614);
not_3  g02294(new_n2671, new_n2670);
xnor_3 g02295(new_n2672, new_n2671, new_n2669);
nand_4 g02296(new_n2673, new_n2672, new_n2668);
not_3  g02297(new_n2674, new_n2595);
nand_4 g02298(new_n2675, new_n2609, new_n2599);
nand_4 g02299(new_n2676, new_n2675, new_n2674);
nand_4 g02300(new_n2677, n8476, n503);
nand_4 g02301(new_n2678, n4970, n2530);
nand_4 g02302(new_n2679_1, n10965, n5331);
xnor_3 g02303(new_n2680, new_n2679_1, new_n2678);
xor_3  g02304(new_n2681, new_n2680, new_n2677);
xnor_3 g02305(new_n2682, new_n2681, new_n2676);
nor_4  g02306(new_n2683, new_n2593, new_n2592);
nand_4 g02307(new_n2684, n12648, n7610);
not_3  g02308(new_n2685, new_n2684);
xor_3  g02309(new_n2686, new_n2685, new_n2683);
not_3  g02310(new_n2687, new_n2686);
nand_4 g02311(new_n2688, n7733, n7690);
not_3  g02312(new_n2689, new_n2688);
nand_4 g02313(new_n2690, n10545, n4826);
nand_4 g02314(new_n2691, n12925, n3616);
xnor_3 g02315(new_n2692, new_n2691, new_n2690);
xnor_3 g02316(new_n2693, new_n2692, new_n2689);
not_3  g02317(new_n2694, new_n2693);
xor_3  g02318(new_n2695, new_n2694, new_n2687);
xnor_3 g02319(new_n2696, new_n2695, new_n2682);
xnor_3 g02320(new_n2697, new_n2696, new_n2673);
xnor_3 g02321(new_n2698, new_n2697, new_n2666);
nand_4 g02322(new_n2699, n5331, n503);
not_3  g02323(new_n2700, new_n2699);
not_3  g02324(new_n2701, new_n2665);
xnor_3 g02325(new_n2702, new_n2701, new_n2635);
nand_4 g02326(new_n2703, new_n2702, new_n2700);
xnor_3 g02327(new_n2704, new_n2649, new_n2639);
xnor_3 g02328(new_n2705, new_n2654, new_n2704);
not_3  g02329(new_n2706, new_n2644);
nand_4 g02330(new_n2707, n12925, n5331);
not_3  g02331(new_n2708_1, new_n2707);
nor_4  g02332(new_n2709, new_n2708_1, new_n2646);
nor_4  g02333(new_n2710, new_n2709, new_n2706);
nor_4  g02334(new_n2711, new_n2710, new_n2645);
nor_4  g02335(new_n2712, new_n2711, new_n2646);
not_3  g02336(new_n2713, new_n2712);
nor_4  g02337(new_n2714, new_n2713, new_n2705);
xnor_3 g02338(new_n2715, new_n2663, new_n2660);
nand_4 g02339(new_n2716, new_n2715, new_n2714);
not_3  g02340(new_n2717, new_n2716);
xnor_3 g02341(new_n2718, new_n2702, new_n2699);
nand_4 g02342(new_n2719, new_n2718, new_n2717);
nand_4 g02343(new_n2720, new_n2719, new_n2703);
xnor_3 g02344(new_n2721, new_n2720, new_n2698);
nand_4 g02345(new_n2722, n4086, n2393);
nand_4 g02346(new_n2723, n5860, n405);
nand_4 g02347(new_n2724, n8433, n3986);
xnor_3 g02348(new_n2725, new_n2724, new_n2723);
nor_4  g02349(new_n2726, new_n2725, new_n2722);
not_3  g02350(new_n2727, new_n2722);
not_3  g02351(new_n2728, new_n2725);
nor_4  g02352(new_n2729, new_n2728, new_n2727);
nor_4  g02353(new_n2730, new_n2729, new_n2726);
nand_4 g02354(new_n2731, n8433, n5860);
not_3  g02355(new_n2732, new_n2731);
nand_4 g02356(new_n2733, n11892, n4086);
not_3  g02357(new_n2734, new_n2733);
nor_4  g02358(new_n2735, new_n2734, new_n2732);
nand_4 g02359(new_n2736, n2393, n405);
not_3  g02360(new_n2737, new_n2736);
xnor_3 g02361(new_n2738, new_n2733, new_n2731);
nor_4  g02362(new_n2739, new_n2738, new_n2737);
nor_4  g02363(new_n2740, new_n2739, new_n2735);
xnor_3 g02364(new_n2741, new_n2740, new_n2730);
not_3  g02365(new_n2742, new_n2741);
nand_4 g02366(new_n2743, n7388, n6611);
nand_4 g02367(new_n2744, n11892, n217);
xor_3  g02368(new_n2745, new_n2744, new_n2743);
xnor_3 g02369(new_n2746, new_n2745, new_n2742);
nand_4 g02370(new_n2747, n7388, n217);
not_3  g02371(new_n2748, new_n2747);
nand_4 g02372(new_n2749_1, n8433, n2393);
not_3  g02373(new_n2750, new_n2749_1);
nand_4 g02374(new_n2751, n7388, n4086);
not_3  g02375(new_n2752, new_n2751);
nor_4  g02376(new_n2753, new_n2752, new_n2750);
nor_4  g02377(new_n2754, new_n2751, new_n2749_1);
nand_4 g02378(new_n2755, n11892, n405);
not_3  g02379(new_n2756, new_n2755);
nor_4  g02380(new_n2757, new_n2756, new_n2754);
nor_4  g02381(new_n2758, new_n2757, new_n2753);
nand_4 g02382(new_n2759, new_n2758, new_n2748);
not_3  g02383(new_n2760, new_n2759);
xnor_3 g02384(new_n2761, new_n2758, new_n2748);
xnor_3 g02385(new_n2762, new_n2738, new_n2736);
nor_4  g02386(new_n2763, new_n2762, new_n2761);
nor_4  g02387(new_n2764, new_n2763, new_n2760);
xnor_3 g02388(new_n2765, new_n2764, new_n2746);
nand_4 g02389(new_n2766, n7965, n6611);
xnor_3 g02390(new_n2767, new_n2762, new_n2761);
nor_4  g02391(new_n2768, new_n2767, new_n2766);
xnor_3 g02392(new_n2769, new_n2767, new_n2766);
nand_4 g02393(new_n2770, n7965, n217);
nand_4 g02394(new_n2771, n11892, n8433);
not_3  g02395(new_n2772, new_n2771);
nand_4 g02396(new_n2773, n7965, n4086);
not_3  g02397(new_n2774, new_n2773);
nand_4 g02398(new_n2775, new_n2774, new_n2772);
nand_4 g02399(new_n2776, new_n2773, new_n2771);
nand_4 g02400(new_n2777, n7388, n405);
not_3  g02401(new_n2778, new_n2777);
nand_4 g02402(new_n2779, new_n2778, new_n2776);
nand_4 g02403(new_n2780, new_n2779, new_n2775);
not_3  g02404(new_n2781, new_n2780);
nor_4  g02405(new_n2782, new_n2781, new_n2770);
xnor_3 g02406(new_n2783, new_n2781, new_n2770);
nor_4  g02407(new_n2784, new_n2754, new_n2753);
xnor_3 g02408(new_n2785, new_n2784, new_n2756);
nor_4  g02409(new_n2786, new_n2785, new_n2783);
nor_4  g02410(new_n2787, new_n2786, new_n2782);
nor_4  g02411(new_n2788, new_n2787, new_n2769);
nor_4  g02412(new_n2789, new_n2788, new_n2768);
nor_4  g02413(new_n2790, new_n2789, new_n2765);
not_3  g02414(new_n2791, new_n2790);
nand_4 g02415(new_n2792, new_n2745, new_n2742);
nor_4  g02416(new_n2793, new_n2744, new_n2743);
xnor_3 g02417(new_n2794, new_n2745, new_n2741);
not_3  g02418(new_n2795, new_n2764);
nand_4 g02419(new_n2796, new_n2795, new_n2794);
not_3  g02420(new_n2797, new_n2796);
xnor_3 g02421(new_n2798, new_n2797, new_n2793);
nand_4 g02422(new_n2799, new_n2798, new_n2792);
nor_4  g02423(new_n2800, new_n2724, new_n2723);
nand_4 g02424(new_n2801, n2393, n217);
xor_3  g02425(new_n2802_1, new_n2801, new_n2800);
nand_4 g02426(new_n2803, n3986, n405);
not_3  g02427(new_n2804, new_n2803);
nand_4 g02428(new_n2805, n5860, n4086);
nand_4 g02429(new_n2806, n8433, n5857);
xnor_3 g02430(new_n2807, new_n2806, new_n2805);
and_4  g02431(new_n2808, new_n2807, new_n2804);
nor_4  g02432(new_n2809, new_n2807, new_n2804);
nor_4  g02433(new_n2810, new_n2809, new_n2808);
xnor_3 g02434(new_n2811, new_n2810, new_n2802_1);
not_3  g02435(new_n2812, new_n2811);
nand_4 g02436(new_n2813, new_n2740, new_n2730);
not_3  g02437(new_n2814, new_n2813);
nor_4  g02438(new_n2815, new_n2814, new_n2726);
not_3  g02439(new_n2816, new_n2815);
nand_4 g02440(new_n2817, n11296, n7965);
not_3  g02441(new_n2818_1, new_n2817);
nand_4 g02442(new_n2819, n11892, n6611);
nand_4 g02443(new_n2820, n7388, n6359);
xnor_3 g02444(new_n2821, new_n2820, new_n2819);
xor_3  g02445(new_n2822, new_n2821, new_n2818_1);
xnor_3 g02446(new_n2823, new_n2822, new_n2816);
xnor_3 g02447(new_n2824, new_n2823, new_n2812);
xnor_3 g02448(new_n2825, new_n2824, new_n2799);
xnor_3 g02449(new_n2826, new_n2825, new_n2791);
nand_4 g02450(new_n2827, n7965, n6359);
not_3  g02451(new_n2828, new_n2827);
not_3  g02452(new_n2829, new_n2765);
xnor_3 g02453(new_n2830, new_n2789, new_n2829);
nand_4 g02454(new_n2831, new_n2830, new_n2828);
nand_4 g02455(new_n2832, new_n2776, new_n2775);
not_3  g02456(new_n2833, new_n2832);
nand_4 g02457(new_n2834, n8433, n7388);
nand_4 g02458(new_n2835, n7965, n405);
nor_4  g02459(new_n2836, new_n2835, new_n2834);
not_3  g02460(new_n2837, new_n2836);
nor_4  g02461(new_n2838, new_n2837, new_n2833);
not_3  g02462(new_n2839, new_n2838);
xnor_3 g02463(new_n2840, new_n2785, new_n2783);
nor_4  g02464(new_n2841, new_n2840, new_n2839);
not_3  g02465(new_n2842, new_n2841);
xnor_3 g02466(new_n2843, new_n2787, new_n2769);
nor_4  g02467(new_n2844, new_n2843, new_n2842);
xnor_3 g02468(new_n2845, new_n2830, new_n2827);
nand_4 g02469(new_n2846, new_n2845, new_n2844);
nand_4 g02470(new_n2847, new_n2846, new_n2831);
xnor_3 g02471(new_n2848, new_n2847, new_n2826);
xnor_3 g02472(new_n2849, new_n2848, new_n2721);
xnor_3 g02473(new_n2850, new_n2702, new_n2700);
nor_4  g02474(new_n2851, new_n2850, new_n2716);
nor_4  g02475(new_n2852, new_n2718, new_n2717);
nor_4  g02476(new_n2853, new_n2852, new_n2851);
not_3  g02477(new_n2854, new_n2853);
xnor_3 g02478(new_n2855, new_n2845, new_n2844);
nand_4 g02479(new_n2856, new_n2855, new_n2854);
xnor_3 g02480(new_n2857, new_n2843, new_n2842);
not_3  g02481(new_n2858, new_n2857);
not_3  g02482(new_n2859, new_n2705);
nor_4  g02483(new_n2860, new_n2712, new_n2859);
nor_4  g02484(new_n2861, new_n2860, new_n2714);
xnor_3 g02485(new_n2862, new_n2840, new_n2839);
not_3  g02486(new_n2863, new_n2862);
nor_4  g02487(new_n2864, new_n2863, new_n2861);
not_3  g02488(new_n2865, new_n2864);
nand_4 g02489(new_n2866, n8433, n7965);
nor_4  g02490(new_n2867, new_n2866, new_n2707);
xnor_3 g02491(new_n2868, new_n2835, new_n2834);
not_3  g02492(new_n2869, new_n2868);
nor_4  g02493(new_n2870, new_n2869, new_n2867);
not_3  g02494(new_n2871, new_n2870);
not_3  g02495(new_n2872, new_n2867);
nor_4  g02496(new_n2873, new_n2868, new_n2872);
nor_4  g02497(new_n2874, new_n2873, new_n2870);
nand_4 g02498(new_n2875, n12925, n8476);
nand_4 g02499(new_n2876, n7733, n5331);
xnor_3 g02500(new_n2877, new_n2876, new_n2875);
nand_4 g02501(new_n2878, new_n2877, new_n2874);
nand_4 g02502(new_n2879_1, new_n2878, new_n2871);
not_3  g02503(new_n2880, new_n2879_1);
not_3  g02504(new_n2881, new_n2711);
not_3  g02505(new_n2882, new_n2709);
nor_4  g02506(new_n2883, new_n2882, new_n2644);
nor_4  g02507(new_n2884, new_n2883, new_n2881);
nor_4  g02508(new_n2885, new_n2884, new_n2880);
not_3  g02509(new_n2886, new_n2885);
not_3  g02510(new_n2887, new_n2884);
nor_4  g02511(new_n2888, new_n2887, new_n2879_1);
nor_4  g02512(new_n2889, new_n2888, new_n2885);
not_3  g02513(new_n2890, new_n2866);
nor_4  g02514(new_n2891, new_n2890, new_n2777);
nor_4  g02515(new_n2892, new_n2891, new_n2833);
nor_4  g02516(new_n2893, new_n2890, new_n2779);
nor_4  g02517(new_n2894, new_n2893, new_n2892);
not_3  g02518(new_n2895, new_n2894);
nand_4 g02519(new_n2896, new_n2895, new_n2889);
nand_4 g02520(new_n2897, new_n2896, new_n2886);
not_3  g02521(new_n2898, new_n2861);
nor_4  g02522(new_n2899, new_n2862, new_n2898);
nor_4  g02523(new_n2900, new_n2899, new_n2864);
nand_4 g02524(new_n2901, new_n2900, new_n2897);
nand_4 g02525(new_n2902_1, new_n2901, new_n2865);
not_3  g02526(new_n2903, new_n2902_1);
nor_4  g02527(new_n2904, new_n2903, new_n2858);
nor_4  g02528(new_n2905, new_n2715, new_n2714);
nor_4  g02529(new_n2906, new_n2905, new_n2717);
xnor_3 g02530(new_n2907, new_n2902_1, new_n2857);
nor_4  g02531(new_n2908, new_n2907, new_n2906);
nor_4  g02532(new_n2909, new_n2908, new_n2904);
not_3  g02533(new_n2910, new_n2909);
xnor_3 g02534(new_n2911, new_n2855, new_n2853);
nand_4 g02535(new_n2912, new_n2911, new_n2910);
nand_4 g02536(new_n2913, new_n2912, new_n2856);
xnor_3 g02537(new_n2914, new_n2913, new_n2849);
not_3  g02538(new_n2915, new_n2914);
nand_4 g02539(new_n2916, new_n2915, new_n2590);
xnor_3 g02540(new_n2917, new_n2914, new_n2590);
not_3  g02541(new_n2918, new_n2556);
xnor_3 g02542(new_n2919, new_n2557, new_n2918);
xnor_3 g02543(new_n2920, new_n2911, new_n2910);
nor_4  g02544(new_n2921, new_n2920, new_n2919);
not_3  g02545(new_n2922, new_n2921);
not_3  g02546(new_n2923, new_n2919);
xnor_3 g02547(new_n2924, new_n2911, new_n2909);
nor_4  g02548(new_n2925, new_n2924, new_n2923);
nor_4  g02549(new_n2926, new_n2925, new_n2921);
xnor_3 g02550(new_n2927, new_n2554, new_n2552);
xnor_3 g02551(new_n2928, new_n2907, new_n2906);
not_3  g02552(new_n2929, new_n2928);
nor_4  g02553(new_n2930, new_n2929, new_n2927);
not_3  g02554(new_n2931, new_n2930);
xnor_3 g02555(new_n2932, new_n2928, new_n2927);
not_3  g02556(new_n2933, new_n2551_1);
xor_3  g02557(new_n2934, new_n2933, new_n2550);
not_3  g02558(new_n2935, new_n2901);
nor_4  g02559(new_n2936, new_n2900, new_n2897);
nor_4  g02560(new_n2937, new_n2936, new_n2935);
nor_4  g02561(new_n2938, new_n2937, new_n2934);
not_3  g02562(new_n2939, new_n2938);
xnor_3 g02563(new_n2940, new_n2937, new_n2934);
xnor_3 g02564(new_n2941, new_n2895, new_n2889);
not_3  g02565(new_n2942, new_n2941);
not_3  g02566(new_n2943, new_n2544);
nand_4 g02567(new_n2944, n8759, n3719);
not_3  g02568(new_n2945, new_n2944);
nor_4  g02569(new_n2946, new_n2945, new_n2526);
not_3  g02570(new_n2947, new_n2946);
nand_4 g02571(new_n2948, new_n2947, new_n2943);
nand_4 g02572(new_n2949, new_n2946, new_n2525);
nand_4 g02573(new_n2950, new_n2949, new_n2948);
nor_4  g02574(new_n2951, new_n2950, new_n2942);
not_3  g02575(new_n2952, new_n2950);
nor_4  g02576(new_n2953, new_n2952, new_n2941);
nor_4  g02577(new_n2954, new_n2953, new_n2951);
not_3  g02578(new_n2955, new_n2954);
xor_3  g02579(new_n2956, new_n2877, new_n2874);
xor_3  g02580(new_n2957, new_n2546, new_n2545);
not_3  g02581(new_n2958, new_n2957);
nor_4  g02582(new_n2959, new_n2958, new_n2956);
xor_3  g02583(new_n2960, new_n2890, new_n2707);
nor_4  g02584(new_n2961, new_n2960, new_n2944);
not_3  g02585(new_n2962, new_n2961);
not_3  g02586(new_n2963, new_n2956);
xor_3  g02587(new_n2964, new_n2958, new_n2963);
nor_4  g02588(new_n2965, new_n2964, new_n2962);
nor_4  g02589(new_n2966, new_n2965, new_n2959);
nor_4  g02590(new_n2967, new_n2966, new_n2955);
nor_4  g02591(new_n2968, new_n2967, new_n2951);
nor_4  g02592(new_n2969, new_n2968, new_n2940);
not_3  g02593(new_n2970, new_n2969);
nand_4 g02594(new_n2971, new_n2970, new_n2939);
nand_4 g02595(new_n2972, new_n2971, new_n2932);
nand_4 g02596(new_n2973, new_n2972, new_n2931);
not_3  g02597(new_n2974, new_n2973);
nand_4 g02598(new_n2975, new_n2974, new_n2926);
nand_4 g02599(new_n2976, new_n2975, new_n2922);
not_3  g02600(new_n2977, new_n2976);
nand_4 g02601(new_n2978, new_n2977, new_n2917);
nand_4 g02602(new_n2979, new_n2978, new_n2916);
xnor_3 g02603(new_n2980, new_n2979, new_n2459);
not_3  g02604(new_n2981, new_n2980);
xnor_3 g02605(new_n2982, new_n2422, new_n2399);
not_3  g02606(new_n2983, new_n2982);
nand_4 g02607(new_n2984, n5305, n2577);
not_3  g02608(new_n2985, new_n2984);
xnor_3 g02609(new_n2986, new_n2420, new_n2415);
not_3  g02610(new_n2987, new_n2986);
nor_4  g02611(new_n2988, new_n2987, new_n2985);
not_3  g02612(new_n2989, new_n2988);
nor_4  g02613(new_n2990, new_n2986, new_n2984);
nor_4  g02614(new_n2991, new_n2990, new_n2988);
nand_4 g02615(new_n2992, n5305, n3842);
nand_4 g02616(new_n2993, n9956, n1097);
not_3  g02617(new_n2994, new_n2993);
nand_4 g02618(new_n2995, n11917, n5305);
not_3  g02619(new_n2996, new_n2995);
nand_4 g02620(new_n2997, new_n2996, new_n2994);
nand_4 g02621(new_n2998, new_n2995, new_n2993);
nand_4 g02622(new_n2999, n5964, n4921);
not_3  g02623(new_n3000, new_n2999);
nand_4 g02624(new_n3001, new_n3000, new_n2998);
nand_4 g02625(new_n3002, new_n3001, new_n2997);
not_3  g02626(new_n3003, new_n3002);
nor_4  g02627(new_n3004, new_n3003, new_n2992);
not_3  g02628(new_n3005, new_n2992);
xnor_3 g02629(new_n3006, new_n3002, new_n3005);
nor_4  g02630(new_n3007, new_n2407, new_n2406);
xnor_3 g02631(new_n3008, new_n3007, new_n2409);
nor_4  g02632(new_n3009, new_n3008, new_n3006);
nor_4  g02633(new_n3010, new_n3009, new_n3004);
nand_4 g02634(new_n3011, new_n3010, new_n2991);
nand_4 g02635(new_n3012, new_n3011, new_n2989);
nor_4  g02636(new_n3013, new_n3012, new_n2983);
not_3  g02637(new_n3014, new_n3013);
xnor_3 g02638(new_n3015, new_n2457, new_n2453);
xnor_3 g02639(new_n3016, new_n3015, new_n3014);
nand_4 g02640(new_n3017, n9637, n5305);
not_3  g02641(new_n3018, new_n3017);
not_3  g02642(new_n3019, new_n3012);
nor_4  g02643(new_n3020, new_n3019, new_n2982);
nor_4  g02644(new_n3021, new_n3020, new_n3013);
nand_4 g02645(new_n3022_1, new_n3021, new_n3018);
and_4  g02646(new_n3023, new_n2998, new_n2997);
nand_4 g02647(new_n3024, n9956, n5964);
nand_4 g02648(new_n3025, n5305, n4921);
nor_4  g02649(new_n3026, new_n3025, new_n3024);
not_3  g02650(new_n3027, new_n3026);
nor_4  g02651(new_n3028, new_n3027, new_n3023);
xor_3  g02652(new_n3029, new_n3008, new_n3006);
nand_4 g02653(new_n3030, new_n3029, new_n3028);
not_3  g02654(new_n3031, new_n3011);
nor_4  g02655(new_n3032, new_n3010, new_n2991);
nor_4  g02656(new_n3033, new_n3032, new_n3031);
nor_4  g02657(new_n3034, new_n3033, new_n3030);
xnor_3 g02658(new_n3035, new_n3021, new_n3017);
nand_4 g02659(new_n3036, new_n3035, new_n3034);
nand_4 g02660(new_n3037, new_n3036, new_n3022_1);
xnor_3 g02661(new_n3038, new_n3037, new_n3016);
not_3  g02662(new_n3039, new_n3038);
xnor_3 g02663(new_n3040, new_n2976, new_n2917);
nor_4  g02664(new_n3041, new_n3040, new_n3039);
not_3  g02665(new_n3042, new_n3041);
nand_4 g02666(new_n3043, new_n3040, new_n3039);
xor_3  g02667(new_n3044, new_n3035, new_n3034);
not_3  g02668(new_n3045, new_n3044);
xnor_3 g02669(new_n3046, new_n2974, new_n2926);
not_3  g02670(new_n3047, new_n3046);
nand_4 g02671(new_n3048, new_n3047, new_n3045);
nand_4 g02672(new_n3049, new_n3046, new_n3044);
xor_3  g02673(new_n3050, new_n3033, new_n3030);
not_3  g02674(new_n3051, new_n3050);
xnor_3 g02675(new_n3052, new_n2971, new_n2932);
nand_4 g02676(new_n3053, new_n3052, new_n3051);
not_3  g02677(new_n3054, new_n3053);
nor_4  g02678(new_n3055, new_n3052, new_n3051);
nor_4  g02679(new_n3056, new_n3055, new_n3054);
not_3  g02680(new_n3057, new_n3029);
xor_3  g02681(new_n3058, new_n3057, new_n3028);
xnor_3 g02682(new_n3059, new_n2968, new_n2940);
nand_4 g02683(new_n3060, new_n3059, new_n3058);
xnor_3 g02684(new_n3061, new_n2966, new_n2955);
not_3  g02685(new_n3062, new_n3023);
nand_4 g02686(new_n3063, n9956, n5305);
not_3  g02687(new_n3064, new_n3063);
nor_4  g02688(new_n3065, new_n3064, new_n2999);
not_3  g02689(new_n3066, new_n3065);
nand_4 g02690(new_n3067, new_n3066, new_n3062);
nand_4 g02691(new_n3068, new_n3065, new_n2998);
nand_4 g02692(new_n3069, new_n3068, new_n3067);
nand_4 g02693(new_n3070, new_n3069, new_n3061);
not_3  g02694(new_n3071_1, new_n3070);
nor_4  g02695(new_n3072, new_n3069, new_n3061);
nor_4  g02696(new_n3073, new_n3072, new_n3071_1);
xor_3  g02697(new_n3074, new_n2960, new_n2944);
nand_4 g02698(new_n3075, new_n3074, new_n3064);
not_3  g02699(new_n3076, new_n3075);
xor_3  g02700(new_n3077, new_n3025, new_n3024);
or_4   g02701(new_n3078, new_n3077, new_n3076);
xnor_3 g02702(new_n3079, new_n2964, new_n2962);
xor_3  g02703(new_n3080, new_n3077, new_n3076);
nand_4 g02704(new_n3081, new_n3080, new_n3079);
nand_4 g02705(new_n3082, new_n3081, new_n3078);
nand_4 g02706(new_n3083, new_n3082, new_n3073);
nand_4 g02707(new_n3084, new_n3083, new_n3070);
not_3  g02708(new_n3085, new_n3060);
nor_4  g02709(new_n3086, new_n3059, new_n3058);
nor_4  g02710(new_n3087, new_n3086, new_n3085);
nand_4 g02711(new_n3088, new_n3087, new_n3084);
nand_4 g02712(new_n3089, new_n3088, new_n3060);
nand_4 g02713(new_n3090, new_n3089, new_n3056);
nand_4 g02714(new_n3091, new_n3090, new_n3053);
nand_4 g02715(new_n3092, new_n3091, new_n3049);
nand_4 g02716(new_n3093, new_n3092, new_n3048);
nand_4 g02717(new_n3094, new_n3093, new_n3043);
nand_4 g02718(new_n3095, new_n3094, new_n3042);
xnor_3 g02719(new_n3096, new_n3095, new_n2981);
nand_4 g02720(new_n3097, n11536, n5305);
not_3  g02721(new_n3098, new_n3097);
nand_4 g02722(new_n3099, n10545, n7610);
nand_4 g02723(new_n3100, n7690, n4826);
not_3  g02724(new_n3101, new_n3100);
xor_3  g02725(new_n3102, new_n3101, new_n3099);
nand_4 g02726(new_n3103, new_n2848, new_n2721);
not_3  g02727(new_n3104, new_n2849);
nand_4 g02728(new_n3105, new_n2913, new_n3104);
nand_4 g02729(new_n3106, new_n3105, new_n3103);
nand_4 g02730(new_n3107, n10510, n3602);
nand_4 g02731(new_n3108, new_n2507_1, new_n2585_1);
not_3  g02732(new_n3109, new_n2582);
nand_4 g02733(new_n3110, new_n2587, new_n3109);
nand_4 g02734(new_n3111, new_n3110, new_n3108);
xnor_3 g02735(new_n3112, new_n3111, new_n3107);
nor_4  g02736(new_n3113, new_n2569, new_n2562);
not_3  g02737(new_n3114, new_n2570);
nor_4  g02738(new_n3115, new_n2581_1, new_n3114);
nor_4  g02739(new_n3116, new_n3115, new_n3113);
nor_4  g02740(new_n3117, new_n2573, new_n2572);
not_3  g02741(new_n3118, new_n2574);
nor_4  g02742(new_n3119, new_n2580, new_n3118);
nor_4  g02743(new_n3120, new_n3119, new_n3117);
not_3  g02744(new_n3121, new_n2564_1);
nor_4  g02745(new_n3122, new_n2566, new_n3121);
not_3  g02746(new_n3123, new_n2563);
nor_4  g02747(new_n3124_1, new_n2567, new_n3123);
nor_4  g02748(new_n3125, new_n3124_1, new_n3122);
nand_4 g02749(new_n3126, n10439, n7436);
not_3  g02750(new_n3127, new_n3126);
nand_4 g02751(new_n3128, n10391, n6776);
nand_4 g02752(new_n3129, n8595, n8276);
xor_3  g02753(new_n3130, new_n3129, new_n3128);
xnor_3 g02754(new_n3131, new_n3130, new_n3127);
xnor_3 g02755(new_n3132, new_n3131, new_n3125);
xnor_3 g02756(new_n3133, new_n3132, new_n3120);
nor_4  g02757(new_n3134, new_n2578, new_n2577_1);
nand_4 g02758(new_n3135, new_n2578, new_n2577_1);
nand_4 g02759(new_n3136, new_n3135, new_n2576);
not_3  g02760(new_n3137, new_n3136);
or_4   g02761(new_n3138, new_n3137, new_n3134);
nand_4 g02762(new_n3139, n9241, n6126);
nand_4 g02763(new_n3140, n12299, n8065);
xor_3  g02764(new_n3141, new_n3140, new_n3139);
nand_4 g02765(new_n3142, n10644, n3719);
nand_4 g02766(new_n3143, n8759, n4190);
xor_3  g02767(new_n3144, new_n3143, new_n3142);
xnor_3 g02768(new_n3145, new_n3144, new_n3141);
xnor_3 g02769(new_n3146_1, new_n3145, new_n3138);
xnor_3 g02770(new_n3147, new_n3146_1, new_n3133);
xnor_3 g02771(new_n3148, new_n3147, new_n3116);
nand_4 g02772(new_n3149, new_n2797, new_n2793);
not_3  g02773(new_n3150, new_n2824);
nand_4 g02774(new_n3151, new_n3150, new_n2799);
nand_4 g02775(new_n3152, new_n3151, new_n3149);
not_3  g02776(new_n3153, new_n2430);
nand_4 g02777(new_n3154, new_n2436, new_n3153);
nand_4 g02778(new_n3155, new_n2452, new_n2437);
nand_4 g02779(new_n3156, new_n3155, new_n3154);
nand_4 g02780(new_n3157, n11257, n4921);
nand_4 g02781(new_n3158, n5964, n1835);
xor_3  g02782(new_n3159, new_n3158, new_n3157);
nand_4 g02783(new_n3160, n4312, n2577);
nand_4 g02784(new_n3161, n12025, n11917);
xor_3  g02785(new_n3162, new_n3161, new_n3160);
xnor_3 g02786(new_n3163, new_n3162, new_n3159);
and_4  g02787(new_n3164, new_n2447, new_n2446);
nor_4  g02788(new_n3165, new_n2450, new_n3164);
and_4  g02789(new_n3166, new_n2434_1, new_n2433_1);
nor_4  g02790(new_n3167, new_n2435, new_n2432);
nor_4  g02791(new_n3168, new_n3167, new_n3166);
xnor_3 g02792(new_n3169, new_n3168, new_n3165);
xnor_3 g02793(new_n3170, new_n3169, new_n3163);
nand_4 g02794(new_n3171, new_n2441, new_n2440);
nand_4 g02795(new_n3172_1, new_n2451, new_n2442);
nand_4 g02796(new_n3173, new_n3172_1, new_n3171);
nand_4 g02797(new_n3174, n9637, n1097);
xnor_3 g02798(new_n3175, new_n3174, new_n3173);
xnor_3 g02799(new_n3176, new_n3175, new_n3170);
xnor_3 g02800(new_n3177, new_n3176, new_n3156);
nand_4 g02801(new_n3178, n4086, n3986);
nand_4 g02802(new_n3179, n12705, n3842);
not_3  g02803(new_n3180, new_n3179);
xor_3  g02804(new_n3181, new_n3180, new_n3178);
xnor_3 g02805(new_n3182, new_n3181, new_n3177);
xnor_3 g02806(new_n3183, new_n3182, new_n3152);
xnor_3 g02807(new_n3184, new_n3183, new_n3148);
xnor_3 g02808(new_n3185, new_n3184, new_n3112);
xnor_3 g02809(new_n3186, new_n3185, new_n3106);
nand_4 g02810(new_n3187, new_n2588, new_n2539);
not_3  g02811(new_n3188, new_n2589);
nand_4 g02812(new_n3189, new_n3188, new_n2559);
nand_4 g02813(new_n3190, new_n3189, new_n3187);
not_3  g02814(new_n3191, new_n2697);
nand_4 g02815(new_n3192, new_n3191, new_n2666);
nand_4 g02816(new_n3193, new_n2720, new_n2698);
nand_4 g02817(new_n3194, new_n3193, new_n3192);
xnor_3 g02818(new_n3195, new_n3194, new_n3190);
nand_4 g02819(new_n3196, n8433, n45);
not_3  g02820(new_n3197, new_n3196);
nand_4 g02821(new_n3198, n5857, n405);
nand_4 g02822(new_n3199, n7965, n1357);
xor_3  g02823(new_n3200, new_n3199, new_n3198);
xor_3  g02824(new_n3201, new_n3200, new_n3197);
and_4  g02825(new_n3202, new_n2820, new_n2819);
nor_4  g02826(new_n3203, new_n2821, new_n2818_1);
nor_4  g02827(new_n3204, new_n3203, new_n3202);
and_4  g02828(new_n3205, new_n2806, new_n2805);
nor_4  g02829(new_n3206, new_n2809, new_n3205);
xnor_3 g02830(new_n3207, new_n3206, new_n3204);
nand_4 g02831(new_n3208, n10965, n8476);
and_4  g02832(new_n3209, new_n2691, new_n2690);
nor_4  g02833(new_n3210, new_n2692, new_n2689);
nor_4  g02834(new_n3211, new_n3210, new_n3209);
xnor_3 g02835(new_n3212, new_n3211, new_n3208);
xnor_3 g02836(new_n3213, new_n3212, new_n3207);
nand_4 g02837(new_n3214_1, new_n2685, new_n2683);
nand_4 g02838(new_n3215, new_n2693, new_n2686);
nand_4 g02839(new_n3216, new_n3215, new_n3214_1);
nand_4 g02840(new_n3217, n5860, n217);
nand_4 g02841(new_n3218, n6611, n2393);
not_3  g02842(new_n3219, new_n3218);
xor_3  g02843(new_n3220, new_n3219, new_n3217);
nand_4 g02844(new_n3221, n7546, n5331);
nand_4 g02845(new_n3222, n12925, n4499);
xnor_3 g02846(new_n3223, new_n3222, new_n3221);
nand_4 g02847(new_n3224, n11892, n6359);
nand_4 g02848(new_n3225, n11296, n7388);
xnor_3 g02849(new_n3226, new_n3225, new_n3224);
xnor_3 g02850(new_n3227, new_n3226, new_n3223);
xnor_3 g02851(new_n3228, new_n3227, new_n3220);
xnor_3 g02852(new_n3229, new_n3228, new_n3216);
xnor_3 g02853(new_n3230_1, new_n3229, new_n3213);
nand_4 g02854(new_n3231, n2530, n503);
not_3  g02855(new_n3232, new_n2800);
nor_4  g02856(new_n3233, new_n2801, new_n3232);
nor_4  g02857(new_n3234, new_n2810, new_n2802_1);
nor_4  g02858(new_n3235, new_n3234, new_n3233);
and_4  g02859(new_n3236, new_n2679_1, new_n2678);
not_3  g02860(new_n3237, new_n2677);
nor_4  g02861(new_n3238, new_n2680, new_n3237);
nor_4  g02862(new_n3239, new_n3238, new_n3236);
nand_4 g02863(new_n3240, n7733, n3616);
nand_4 g02864(new_n3241, n12648, n4970);
not_3  g02865(new_n3242, new_n3241);
xor_3  g02866(new_n3243, new_n3242, new_n3240);
xnor_3 g02867(new_n3244, new_n3243, new_n3239);
xnor_3 g02868(new_n3245, new_n3244, new_n3235);
xnor_3 g02869(new_n3246, new_n3245, new_n3231);
xnor_3 g02870(new_n3247, new_n3246, new_n3230_1);
nand_4 g02871(new_n3248, new_n2822, new_n2815);
nand_4 g02872(new_n3249, new_n2823, new_n2811);
nand_4 g02873(new_n3250, new_n3249, new_n3248);
nand_4 g02874(new_n3251, new_n2681, new_n2676);
not_3  g02875(new_n3252, new_n2682);
nand_4 g02876(new_n3253, new_n2695, new_n3252);
nand_4 g02877(new_n3254, new_n3253, new_n3251);
xnor_3 g02878(new_n3255, new_n3254, new_n3250);
xnor_3 g02879(new_n3256, new_n3255, new_n3247);
nand_4 g02880(new_n3257, new_n2671, new_n2669);
nand_4 g02881(new_n3258, new_n2696, new_n2673);
nand_4 g02882(new_n3259, new_n3258, new_n3257);
nand_4 g02883(new_n3260, n10547, n9956);
not_3  g02884(new_n3261, new_n3260);
xnor_3 g02885(new_n3262, new_n3261, new_n3259);
xnor_3 g02886(new_n3263, new_n3262, new_n3256);
xnor_3 g02887(new_n3264, new_n3263, new_n3201);
nand_4 g02888(new_n3265, new_n3015, new_n3013);
nand_4 g02889(new_n3266, new_n3037, new_n3016);
nand_4 g02890(new_n3267, new_n3266, new_n3265);
nand_4 g02891(new_n3268, new_n2825, new_n2790);
nand_4 g02892(new_n3269, new_n2847, new_n2826);
nand_4 g02893(new_n3270, new_n3269, new_n3268);
xnor_3 g02894(new_n3271, new_n3270, new_n3267);
xnor_3 g02895(new_n3272_1, new_n3271, new_n3264);
xnor_3 g02896(new_n3273, new_n3272_1, new_n3195);
xnor_3 g02897(new_n3274, new_n3273, new_n3186);
xnor_3 g02898(new_n3275, new_n3274, new_n3102);
xnor_3 g02899(new_n3276, new_n3275, new_n3098);
nand_4 g02900(new_n3277, new_n3276, new_n3096);
xnor_3 g02901(new_n3278, new_n3095, new_n2980);
xnor_3 g02902(new_n3279, new_n3275, new_n3097);
nand_4 g02903(new_n3280, new_n3279, new_n3278);
nand_4 g02904(n837, new_n3280, new_n3277);
nand_4 g02905(new_n3282, n11917, n11757);
not_3  g02906(new_n3283, new_n3282);
nand_4 g02907(new_n3284, n9956, n5240);
nand_4 g02908(new_n3285, n11757, n4921);
not_3  g02909(new_n3286, new_n3285);
nand_4 g02910(new_n3287_1, n11917, n3172);
xnor_3 g02911(new_n3288, new_n3287_1, new_n3284);
nor_4  g02912(new_n3289, new_n3288, new_n3286);
nor_4  g02913(new_n3290, new_n3289, new_n3284);
nor_4  g02914(new_n3291, new_n3290, new_n3283);
nand_4 g02915(new_n3292, n4921, n3172);
not_3  g02916(new_n3293, new_n3292);
nor_4  g02917(new_n3294, new_n3293, new_n3290);
nor_4  g02918(new_n3295, new_n3294, new_n3282);
nor_4  g02919(new_n3296, new_n3295, new_n3291);
nand_4 g02920(new_n3297, n5240, n4921);
nand_4 g02921(new_n3298, n11821, n9956);
xor_3  g02922(new_n3299, new_n3298, new_n3297);
xnor_3 g02923(new_n3300, new_n3299, new_n3296);
not_3  g02924(new_n3301, new_n3300);
nand_4 g02925(new_n3302, n2577, n1333);
nand_4 g02926(new_n3303, n3842, n3172);
xor_3  g02927(new_n3304, new_n3303, new_n3302);
xnor_3 g02928(new_n3305, new_n3304, new_n3301);
nand_4 g02929(new_n3306, n3842, n1333);
not_3  g02930(new_n3307, new_n3306);
nand_4 g02931(new_n3308, n11757, n9956);
not_3  g02932(new_n3309, new_n3308);
nand_4 g02933(new_n3310, n11917, n1333);
not_3  g02934(new_n3311, new_n3310);
nor_4  g02935(new_n3312, new_n3311, new_n3309);
nor_4  g02936(new_n3313, new_n3310, new_n3308);
nor_4  g02937(new_n3314, new_n3313, new_n3293);
nor_4  g02938(new_n3315, new_n3314, new_n3312);
and_4  g02939(new_n3316, new_n3315, new_n3307);
not_3  g02940(new_n3317, new_n3288);
nor_4  g02941(new_n3318, new_n3317, new_n3285);
nor_4  g02942(new_n3319, new_n3318, new_n3289);
xnor_3 g02943(new_n3320, new_n3315, new_n3307);
nor_4  g02944(new_n3321, new_n3320, new_n3319);
nor_4  g02945(new_n3322, new_n3321, new_n3316);
xnor_3 g02946(new_n3323, new_n3322, new_n3305);
not_3  g02947(new_n3324, new_n3323);
nand_4 g02948(new_n3325, n7862, n2577);
xnor_3 g02949(new_n3326, new_n3320, new_n3319);
nor_4  g02950(new_n3327, new_n3326, new_n3325);
not_3  g02951(new_n3328, new_n3327);
nand_4 g02952(new_n3329, n7862, n3842);
nand_4 g02953(new_n3330, n9956, n3172);
not_3  g02954(new_n3331, new_n3330);
nand_4 g02955(new_n3332, n11917, n7862);
not_3  g02956(new_n3333, new_n3332);
nand_4 g02957(new_n3334, new_n3333, new_n3331);
nand_4 g02958(new_n3335, new_n3332, new_n3330);
nand_4 g02959(new_n3336, n4921, n1333);
not_3  g02960(new_n3337, new_n3336);
nand_4 g02961(new_n3338, new_n3337, new_n3335);
nand_4 g02962(new_n3339_1, new_n3338, new_n3334);
not_3  g02963(new_n3340, new_n3339_1);
nor_4  g02964(new_n3341, new_n3340, new_n3329);
not_3  g02965(new_n3342_1, new_n3341);
xor_3  g02966(new_n3343, new_n3340, new_n3329);
nor_4  g02967(new_n3344, new_n3313, new_n3312);
xor_3  g02968(new_n3345, new_n3344, new_n3293);
nand_4 g02969(new_n3346, new_n3345, new_n3343);
nand_4 g02970(new_n3347, new_n3346, new_n3342_1);
xnor_3 g02971(new_n3348, new_n3326, new_n3325);
not_3  g02972(new_n3349, new_n3348);
nand_4 g02973(new_n3350, new_n3349, new_n3347);
nand_4 g02974(new_n3351, new_n3350, new_n3328);
nand_4 g02975(new_n3352, new_n3351, new_n3324);
not_3  g02976(new_n3353, new_n3295);
nand_4 g02977(new_n3354, new_n3299, new_n3296);
nand_4 g02978(new_n3355, new_n3354, new_n3353);
nand_4 g02979(new_n3356, n9637, n1333);
not_3  g02980(new_n3357, new_n3356);
nand_4 g02981(new_n3358, n3172, n2577);
nand_4 g02982(new_n3359, n7862, n1835);
xor_3  g02983(new_n3360, new_n3359, new_n3358);
xnor_3 g02984(new_n3361, new_n3360, new_n3357);
xnor_3 g02985(new_n3362, new_n3361, new_n3355);
nor_4  g02986(new_n3363, new_n3298, new_n3297);
not_3  g02987(new_n3364, new_n3363);
nand_4 g02988(new_n3365, n11757, n3842);
xor_3  g02989(new_n3366, new_n3365, new_n3364);
nand_4 g02990(new_n3367, n11821, n4921);
nand_4 g02991(new_n3368, n9956, n9080);
nand_4 g02992(new_n3369, n11917, n5240);
not_3  g02993(new_n3370, new_n3369);
xor_3  g02994(new_n3371, new_n3370, new_n3368);
xnor_3 g02995(new_n3372, new_n3371, new_n3367);
not_3  g02996(new_n3373, new_n3372);
nor_4  g02997(new_n3374, new_n3373, new_n3366);
not_3  g02998(new_n3375, new_n3366);
nor_4  g02999(new_n3376, new_n3372, new_n3375);
nor_4  g03000(new_n3377, new_n3376, new_n3374);
xnor_3 g03001(new_n3378, new_n3377, new_n3362);
nand_4 g03002(new_n3379, new_n3304, new_n3301);
nor_4  g03003(new_n3380, new_n3303, new_n3302);
nor_4  g03004(new_n3381, new_n3322, new_n3305);
xnor_3 g03005(new_n3382, new_n3381, new_n3380);
nand_4 g03006(new_n3383, new_n3382, new_n3379);
xnor_3 g03007(new_n3384, new_n3383, new_n3378);
xnor_3 g03008(new_n3385, new_n3384, new_n3352);
nand_4 g03009(new_n3386, n9637, n7862);
not_3  g03010(new_n3387, new_n3386);
xnor_3 g03011(new_n3388, new_n3351, new_n3324);
not_3  g03012(new_n3389, new_n3388);
nand_4 g03013(new_n3390, new_n3389, new_n3387);
and_4  g03014(new_n3391, new_n3335, new_n3334);
nand_4 g03015(new_n3392, n9956, n1333);
nand_4 g03016(new_n3393, n7862, n4921);
nor_4  g03017(new_n3394, new_n3393, new_n3392);
not_3  g03018(new_n3395, new_n3394);
nor_4  g03019(new_n3396, new_n3395, new_n3391);
xor_3  g03020(new_n3397, new_n3339_1, new_n3329);
xor_3  g03021(new_n3398, new_n3344, new_n3292);
nor_4  g03022(new_n3399, new_n3398, new_n3397);
nor_4  g03023(new_n3400, new_n3345, new_n3343);
nor_4  g03024(new_n3401, new_n3400, new_n3399);
nand_4 g03025(new_n3402, new_n3401, new_n3396);
xnor_3 g03026(new_n3403, new_n3349, new_n3347);
nor_4  g03027(new_n3404, new_n3403, new_n3402);
xnor_3 g03028(new_n3405, new_n3388, new_n3387);
nand_4 g03029(new_n3406, new_n3405, new_n3404);
nand_4 g03030(new_n3407, new_n3406, new_n3390);
xor_3  g03031(new_n3408, new_n3407, new_n3385);
not_3  g03032(new_n3409, new_n3405);
xor_3  g03033(new_n3410, new_n3409, new_n3404);
not_3  g03034(new_n3411, new_n3410);
nand_4 g03035(new_n3412, n8595, n6877);
nand_4 g03036(new_n3413, n6877, n6126);
not_3  g03037(new_n3414, new_n3413);
nand_4 g03038(new_n3415, n3719, n2464);
not_3  g03039(new_n3416, new_n3415);
nor_4  g03040(new_n3417, new_n3416, new_n3414);
nor_4  g03041(new_n3418, new_n3415, new_n3413);
nand_4 g03042(new_n3419, n9400, n3602);
not_3  g03043(new_n3420, new_n3419);
nor_4  g03044(new_n3421, new_n3420, new_n3418);
nor_4  g03045(new_n3422, new_n3421, new_n3417);
xor_3  g03046(new_n3423, new_n3422, new_n3412);
nand_4 g03047(new_n3424, n3602, n2464);
nand_4 g03048(new_n3425, n9400, n6126);
not_3  g03049(new_n3426, new_n3425);
nand_4 g03050(new_n3427, n11311, n3719);
not_3  g03051(new_n3428, new_n3427);
nor_4  g03052(new_n3429, new_n3428, new_n3426);
nor_4  g03053(new_n3430, new_n3427, new_n3425);
nor_4  g03054(new_n3431, new_n3430, new_n3429);
xor_3  g03055(new_n3432, new_n3431, new_n3424);
xnor_3 g03056(new_n3433, new_n3432, new_n3423);
nand_4 g03057(new_n3434, n6877, n3719);
not_3  g03058(new_n3435, new_n3434);
nor_4  g03059(new_n3436, new_n3435, new_n3419);
nor_4  g03060(new_n3437, new_n3418, new_n3417);
nor_4  g03061(new_n3438, new_n3437, new_n3436);
not_3  g03062(new_n3439, new_n3438);
nor_4  g03063(new_n3440, new_n3439, new_n3419);
not_3  g03064(new_n3441, new_n3440);
nor_4  g03065(new_n3442, new_n3441, new_n3433);
not_3  g03066(new_n3443, new_n3442);
nand_4 g03067(new_n3444, n10439, n6877);
nand_4 g03068(new_n3445, n9400, n8595);
not_3  g03069(new_n3446, new_n3445);
not_3  g03070(new_n3447, new_n3424);
nor_4  g03071(new_n3448, new_n3430, new_n3447);
nor_4  g03072(new_n3449, new_n3448, new_n3429);
xnor_3 g03073(new_n3450, new_n3449, new_n3446);
nand_4 g03074(new_n3451, n11311, n3602);
not_3  g03075(new_n3452, new_n3451);
nand_4 g03076(new_n3453, n6126, n2464);
nand_4 g03077(new_n3454, n4187, n3719);
xnor_3 g03078(new_n3455, new_n3454, new_n3453);
xor_3  g03079(new_n3456_1, new_n3455, new_n3452);
xnor_3 g03080(new_n3457, new_n3456_1, new_n3450);
xnor_3 g03081(new_n3458, new_n3457, new_n3444);
not_3  g03082(new_n3459, new_n3412);
and_4  g03083(new_n3460, new_n3422, new_n3459);
nor_4  g03084(new_n3461, new_n3432, new_n3423);
nor_4  g03085(new_n3462, new_n3461, new_n3460);
xnor_3 g03086(new_n3463, new_n3462, new_n3458);
nor_4  g03087(new_n3464, new_n3463, new_n3443);
not_3  g03088(new_n3465, new_n3464);
nand_4 g03089(new_n3466, n8065, n6877);
nand_4 g03090(new_n3467, n11311, n6126);
nand_4 g03091(new_n3468, n4203, n3719);
nand_4 g03092(new_n3469, n4187, n3602);
xnor_3 g03093(new_n3470, new_n3469, new_n3468);
nor_4  g03094(new_n3471, new_n3470, new_n3467);
not_3  g03095(new_n3472, new_n3467);
not_3  g03096(new_n3473, new_n3470);
nor_4  g03097(new_n3474, new_n3473, new_n3472);
nor_4  g03098(new_n3475, new_n3474, new_n3471);
and_4  g03099(new_n3476, new_n3454, new_n3453);
nor_4  g03100(new_n3477, new_n3455, new_n3452);
nor_4  g03101(new_n3478, new_n3477, new_n3476);
not_3  g03102(new_n3479, new_n3478);
xor_3  g03103(new_n3480, new_n3479, new_n3475);
nand_4 g03104(new_n3481, n10439, n9400);
nand_4 g03105(new_n3482, n8595, n2464);
xor_3  g03106(new_n3483, new_n3482, new_n3481);
not_3  g03107(new_n3484, new_n3483);
xnor_3 g03108(new_n3485, new_n3484, new_n3480);
and_4  g03109(new_n3486, new_n3449, new_n3446);
not_3  g03110(new_n3487, new_n3486);
not_3  g03111(new_n3488, new_n3450);
not_3  g03112(new_n3489, new_n3456_1);
nand_4 g03113(new_n3490, new_n3489, new_n3488);
and_4  g03114(new_n3491, new_n3490, new_n3487);
xnor_3 g03115(new_n3492, new_n3491, new_n3485);
not_3  g03116(new_n3493, new_n3444);
not_3  g03117(new_n3494, new_n3457);
nand_4 g03118(new_n3495, new_n3494, new_n3493);
xor_3  g03119(new_n3496, new_n3494, new_n3493);
not_3  g03120(new_n3497, new_n3462);
nand_4 g03121(new_n3498, new_n3497, new_n3496);
nand_4 g03122(new_n3499, new_n3498, new_n3495);
not_3  g03123(new_n3500, new_n3499);
xnor_3 g03124(new_n3501, new_n3500, new_n3492);
xnor_3 g03125(new_n3502, new_n3501, new_n3466);
xnor_3 g03126(new_n3503, new_n3502, new_n3465);
not_3  g03127(new_n3504, new_n3463);
xor_3  g03128(new_n3505, new_n3504, new_n3443);
not_3  g03129(new_n3506, new_n3505);
not_3  g03130(new_n3507, new_n3433);
xor_3  g03131(new_n3508, new_n3440, new_n3507);
not_3  g03132(new_n3509, new_n3508);
nand_4 g03133(new_n3510, n8433, n7236);
nand_4 g03134(new_n3511, n12925, n4805);
nor_4  g03135(new_n3512, new_n3511, new_n3510);
nand_4 g03136(new_n3513, n7733, n4805);
nand_4 g03137(new_n3514, n12925, n11478);
xnor_3 g03138(new_n3515, new_n3514, new_n3513);
not_3  g03139(new_n3516, new_n3515);
nor_4  g03140(new_n3517, new_n3516, new_n3512);
not_3  g03141(new_n3518, new_n3517);
not_3  g03142(new_n3519, new_n3512);
nor_4  g03143(new_n3520, new_n3515, new_n3519);
nor_4  g03144(new_n3521, new_n3520, new_n3517);
nand_4 g03145(new_n3522, n7236, n405);
nand_4 g03146(new_n3523, n8433, n3992);
xnor_3 g03147(new_n3524, new_n3523, new_n3522);
nand_4 g03148(new_n3525, new_n3524, new_n3521);
nand_4 g03149(new_n3526, new_n3525, new_n3518);
not_3  g03150(new_n3527, new_n3510);
nand_4 g03151(new_n3528, n3992, n405);
nor_4  g03152(new_n3529, new_n3528, new_n3527);
nand_4 g03153(new_n3530, n8433, n8384);
not_3  g03154(new_n3531, new_n3530);
nand_4 g03155(new_n3532, n7236, n4086);
not_3  g03156(new_n3533, new_n3532);
nor_4  g03157(new_n3534, new_n3533, new_n3531);
not_3  g03158(new_n3535, new_n3534);
nor_4  g03159(new_n3536, new_n3535, new_n3529);
nor_4  g03160(new_n3537, new_n3532, new_n3530);
nor_4  g03161(new_n3538, new_n3537, new_n3536);
not_3  g03162(new_n3539, new_n3529);
nor_4  g03163(new_n3540, new_n3534, new_n3539);
not_3  g03164(new_n3541, new_n3540);
nand_4 g03165(new_n3542, new_n3541, new_n3538);
xnor_3 g03166(new_n3543, new_n3542, new_n3526);
not_3  g03167(new_n3544, new_n3511);
nand_4 g03168(new_n3545, n11478, n7733);
nor_4  g03169(new_n3546, new_n3545, new_n3544);
not_3  g03170(new_n3547, new_n3546);
nand_4 g03171(new_n3548, n12925, n5283);
nand_4 g03172(new_n3549, n4826, n4805);
nand_4 g03173(new_n3550, new_n3549, new_n3548);
nor_4  g03174(new_n3551, new_n3550, new_n3547);
not_3  g03175(new_n3552, new_n3550);
not_3  g03176(new_n3553, new_n3548);
not_3  g03177(new_n3554, new_n3549);
nand_4 g03178(new_n3555, new_n3554, new_n3553);
not_3  g03179(new_n3556, new_n3555);
nor_4  g03180(new_n3557, new_n3556, new_n3552);
not_3  g03181(new_n3558, new_n3557);
nor_4  g03182(new_n3559, new_n3558, new_n3546);
nor_4  g03183(new_n3560, new_n3559, new_n3551);
not_3  g03184(new_n3561, new_n3560);
xnor_3 g03185(new_n3562, new_n3561, new_n3543);
not_3  g03186(new_n3563, new_n3562);
not_3  g03187(new_n3564, new_n3417);
nand_4 g03188(new_n3565, new_n3436, new_n3564);
nand_4 g03189(new_n3566, new_n3565, new_n3439);
nor_4  g03190(new_n3567, new_n3566, new_n3563);
not_3  g03191(new_n3568, new_n3566);
nor_4  g03192(new_n3569, new_n3568, new_n3562);
nor_4  g03193(new_n3570, new_n3569, new_n3567);
not_3  g03194(new_n3571, new_n3570);
xnor_3 g03195(new_n3572, new_n3524, new_n3521);
not_3  g03196(new_n3573, new_n3572);
nand_4 g03197(new_n3574, n9400, n3719);
nand_4 g03198(new_n3575, n6877, n3602);
not_3  g03199(new_n3576, new_n3575);
xor_3  g03200(new_n3577, new_n3576, new_n3574);
nor_4  g03201(new_n3578, new_n3577, new_n3573);
xor_3  g03202(new_n3579, new_n3511, new_n3510);
nand_4 g03203(new_n3580, new_n3579, new_n3435);
xnor_3 g03204(new_n3581, new_n3577, new_n3572);
not_3  g03205(new_n3582, new_n3581);
nor_4  g03206(new_n3583, new_n3582, new_n3580);
nor_4  g03207(new_n3584, new_n3583, new_n3578);
nor_4  g03208(new_n3585, new_n3584, new_n3571);
nor_4  g03209(new_n3586, new_n3585, new_n3567);
nor_4  g03210(new_n3587, new_n3586, new_n3509);
not_3  g03211(new_n3588, new_n3587);
nand_4 g03212(new_n3589, new_n3586, new_n3509);
nand_4 g03213(new_n3590, n7610, n4805);
not_3  g03214(new_n3591, new_n3545);
nand_4 g03215(new_n3592, new_n3550, new_n3591);
nand_4 g03216(new_n3593, new_n3592, new_n3555);
not_3  g03217(new_n3594, new_n3593);
xnor_3 g03218(new_n3595, new_n3594, new_n3590);
nand_4 g03219(new_n3596, n7733, n5283);
nand_4 g03220(new_n3597, n12925, n137);
nand_4 g03221(new_n3598, n11478, n4826);
xnor_3 g03222(new_n3599, new_n3598, new_n3597);
xnor_3 g03223(new_n3600, new_n3599, new_n3596);
xnor_3 g03224(new_n3601, new_n3600, new_n3595);
not_3  g03225(new_n3602_1, new_n3601);
nor_4  g03226(new_n3603, new_n3514, new_n3513);
not_3  g03227(new_n3604, new_n3603);
nor_4  g03228(new_n3605, new_n3557, new_n3604);
nor_4  g03229(new_n3606, new_n3605, new_n3602_1);
not_3  g03230(new_n3607, new_n3605);
nor_4  g03231(new_n3608, new_n3607, new_n3601);
nor_4  g03232(new_n3609, new_n3608, new_n3606);
nand_4 g03233(new_n3610, n7236, n217);
not_3  g03234(new_n3611, new_n3610);
not_3  g03235(new_n3612, new_n3528);
nor_4  g03236(new_n3613, new_n3537, new_n3612);
nor_4  g03237(new_n3614, new_n3613, new_n3534);
xnor_3 g03238(new_n3615, new_n3614, new_n3611);
nand_4 g03239(new_n3616_1, n8384, n405);
nand_4 g03240(new_n3617, n8433, n6358);
nand_4 g03241(new_n3618, n4086, n3992);
xnor_3 g03242(new_n3619, new_n3618, new_n3617);
xnor_3 g03243(new_n3620, new_n3619, new_n3616_1);
xnor_3 g03244(new_n3621, new_n3620, new_n3615);
not_3  g03245(new_n3622, new_n3621);
nor_4  g03246(new_n3623, new_n3538, new_n3528);
nor_4  g03247(new_n3624, new_n3623, new_n3622);
not_3  g03248(new_n3625, new_n3623);
nor_4  g03249(new_n3626, new_n3625, new_n3621);
nor_4  g03250(new_n3627_1, new_n3626, new_n3624);
xnor_3 g03251(new_n3628, new_n3627_1, new_n3609);
not_3  g03252(new_n3629, new_n3628);
and_4  g03253(new_n3630, new_n3542, new_n3526);
nor_4  g03254(new_n3631, new_n3561, new_n3543);
nor_4  g03255(new_n3632, new_n3631, new_n3630);
not_3  g03256(new_n3633, new_n3632);
nor_4  g03257(new_n3634, new_n3633, new_n3629);
nor_4  g03258(new_n3635, new_n3632, new_n3628);
nor_4  g03259(new_n3636, new_n3635, new_n3634);
not_3  g03260(new_n3637, new_n3636);
nand_4 g03261(new_n3638, new_n3637, new_n3589);
nand_4 g03262(new_n3639, new_n3638, new_n3588);
nand_4 g03263(new_n3640, new_n3639, new_n3506);
not_3  g03264(new_n3641, new_n3586);
nor_4  g03265(new_n3642, new_n3641, new_n3508);
nor_4  g03266(new_n3643, new_n3636, new_n3642);
nor_4  g03267(new_n3644, new_n3643, new_n3587);
nand_4 g03268(new_n3645, new_n3644, new_n3505);
nand_4 g03269(new_n3646, n7236, n6611);
nand_4 g03270(new_n3647, n3992, n217);
not_3  g03271(new_n3648, new_n3647);
not_3  g03272(new_n3649, new_n3617);
not_3  g03273(new_n3650, new_n3618);
nor_4  g03274(new_n3651, new_n3650, new_n3649);
not_3  g03275(new_n3652, new_n3616_1);
nor_4  g03276(new_n3653, new_n3619, new_n3652);
nor_4  g03277(new_n3654_1, new_n3653, new_n3651);
xnor_3 g03278(new_n3655, new_n3654_1, new_n3648);
nand_4 g03279(new_n3656, n6358, n405);
nand_4 g03280(new_n3657, n8384, n4086);
nand_4 g03281(new_n3658, n8433, n5198);
xnor_3 g03282(new_n3659, new_n3658, new_n3657);
xnor_3 g03283(new_n3660, new_n3659, new_n3656);
xnor_3 g03284(new_n3661_1, new_n3660, new_n3655);
nor_4  g03285(new_n3662, new_n3661_1, new_n3646);
not_3  g03286(new_n3663, new_n3646);
not_3  g03287(new_n3664, new_n3661_1);
nor_4  g03288(new_n3665, new_n3664, new_n3663);
nor_4  g03289(new_n3666, new_n3665, new_n3662);
nand_4 g03290(new_n3667, new_n3614, new_n3611);
not_3  g03291(new_n3668, new_n3667);
nor_4  g03292(new_n3669, new_n3620, new_n3615);
nor_4  g03293(new_n3670, new_n3669, new_n3668);
not_3  g03294(new_n3671, new_n3670);
nand_4 g03295(new_n3672, new_n3671, new_n3666);
not_3  g03296(new_n3673, new_n3672);
nor_4  g03297(new_n3674, new_n3671, new_n3666);
nor_4  g03298(new_n3675, new_n3674, new_n3673);
nor_4  g03299(new_n3676, new_n3675, new_n3626);
nand_4 g03300(new_n3677_1, new_n3675, new_n3626);
not_3  g03301(new_n3678, new_n3677_1);
nor_4  g03302(new_n3679, new_n3678, new_n3676);
nand_4 g03303(new_n3680, n4970, n4805);
nand_4 g03304(new_n3681, n11478, n7610);
not_3  g03305(new_n3682, new_n3681);
not_3  g03306(new_n3683, new_n3597);
not_3  g03307(new_n3684, new_n3598);
nor_4  g03308(new_n3685, new_n3684, new_n3683);
not_3  g03309(new_n3686, new_n3596);
nor_4  g03310(new_n3687, new_n3599, new_n3686);
nor_4  g03311(new_n3688, new_n3687, new_n3685);
xnor_3 g03312(new_n3689, new_n3688, new_n3682);
nand_4 g03313(new_n3690, n7733, n137);
nand_4 g03314(new_n3691, n5283, n4826);
nand_4 g03315(new_n3692, n12925, n6294);
xnor_3 g03316(new_n3693, new_n3692, new_n3691);
xnor_3 g03317(new_n3694, new_n3693, new_n3690);
xnor_3 g03318(new_n3695, new_n3694, new_n3689);
nor_4  g03319(new_n3696, new_n3695, new_n3680);
not_3  g03320(new_n3697, new_n3680);
not_3  g03321(new_n3698, new_n3695);
nor_4  g03322(new_n3699, new_n3698, new_n3697);
nor_4  g03323(new_n3700, new_n3699, new_n3696);
nor_4  g03324(new_n3701, new_n3594, new_n3590);
nor_4  g03325(new_n3702, new_n3600, new_n3595);
nor_4  g03326(new_n3703, new_n3702, new_n3701);
not_3  g03327(new_n3704, new_n3703);
xnor_3 g03328(new_n3705, new_n3704, new_n3700);
not_3  g03329(new_n3706, new_n3705);
nor_4  g03330(new_n3707, new_n3706, new_n3608);
not_3  g03331(new_n3708, new_n3608);
nor_4  g03332(new_n3709, new_n3705, new_n3708);
nor_4  g03333(new_n3710, new_n3709, new_n3707);
nor_4  g03334(new_n3711, new_n3627_1, new_n3609);
nor_4  g03335(new_n3712, new_n3635, new_n3711);
xnor_3 g03336(new_n3713, new_n3712, new_n3710);
xnor_3 g03337(new_n3714, new_n3713, new_n3679);
nand_4 g03338(new_n3715, new_n3714, new_n3645);
nand_4 g03339(new_n3716, new_n3715, new_n3640);
xnor_3 g03340(new_n3717, new_n3716, new_n3503);
nand_4 g03341(new_n3718, n7236, n6359);
not_3  g03342(new_n3719_1, new_n3718);
nand_4 g03343(new_n3720, n6358, n4086);
not_3  g03344(new_n3721, new_n3720);
not_3  g03345(new_n3722, new_n3657);
not_3  g03346(new_n3723, new_n3658);
nor_4  g03347(new_n3724, new_n3723, new_n3722);
not_3  g03348(new_n3725, new_n3656);
nor_4  g03349(new_n3726, new_n3659, new_n3725);
nor_4  g03350(new_n3727, new_n3726, new_n3724);
xnor_3 g03351(new_n3728, new_n3727, new_n3721);
nand_4 g03352(new_n3729, n5198, n405);
nand_4 g03353(new_n3730, n8433, n1471);
xnor_3 g03354(new_n3731, new_n3730, new_n3729);
xnor_3 g03355(new_n3732, new_n3731, new_n3728);
not_3  g03356(new_n3733, new_n3732);
nand_4 g03357(new_n3734, n8384, n217);
nand_4 g03358(new_n3735, n6611, n3992);
xor_3  g03359(new_n3736, new_n3735, new_n3734);
xnor_3 g03360(new_n3737, new_n3736, new_n3733);
not_3  g03361(new_n3738, new_n3737);
and_4  g03362(new_n3739, new_n3654_1, new_n3648);
nor_4  g03363(new_n3740, new_n3660, new_n3655);
nor_4  g03364(new_n3741, new_n3740, new_n3739);
xnor_3 g03365(new_n3742, new_n3741, new_n3738);
not_3  g03366(new_n3743, new_n3662);
nand_4 g03367(new_n3744, new_n3672, new_n3743);
xnor_3 g03368(new_n3745, new_n3744, new_n3742);
xnor_3 g03369(new_n3746, new_n3745, new_n3719_1);
nor_4  g03370(new_n3747, new_n3746, new_n3677_1);
nand_4 g03371(new_n3748, new_n3746, new_n3677_1);
not_3  g03372(new_n3749, new_n3748);
nor_4  g03373(new_n3750, new_n3749, new_n3747);
nand_4 g03374(new_n3751, n4805, n503);
not_3  g03375(new_n3752, new_n3751);
nand_4 g03376(new_n3753, n4826, n137);
nand_4 g03377(new_n3754_1, n7733, n6294);
nand_4 g03378(new_n3755, n12925, n6797);
xnor_3 g03379(new_n3756, new_n3755, new_n3754_1);
nor_4  g03380(new_n3757, new_n3756, new_n3753);
not_3  g03381(new_n3758, new_n3753);
not_3  g03382(new_n3759, new_n3756);
nor_4  g03383(new_n3760, new_n3759, new_n3758);
nor_4  g03384(new_n3761, new_n3760, new_n3757);
and_4  g03385(new_n3762, new_n3692, new_n3691);
not_3  g03386(new_n3763, new_n3690);
nor_4  g03387(new_n3764, new_n3693, new_n3763);
nor_4  g03388(new_n3765, new_n3764, new_n3762);
xnor_3 g03389(new_n3766, new_n3765, new_n3761);
nand_4 g03390(new_n3767, n11478, n4970);
nand_4 g03391(new_n3768, n7610, n5283);
xor_3  g03392(new_n3769, new_n3768, new_n3767);
xnor_3 g03393(new_n3770, new_n3769, new_n3766);
nand_4 g03394(new_n3771, new_n3688, new_n3682);
not_3  g03395(new_n3772, new_n3771);
nor_4  g03396(new_n3773, new_n3694, new_n3689);
nor_4  g03397(new_n3774, new_n3773, new_n3772);
not_3  g03398(new_n3775, new_n3774);
xnor_3 g03399(new_n3776, new_n3775, new_n3770);
not_3  g03400(new_n3777, new_n3696);
nand_4 g03401(new_n3778, new_n3704, new_n3700);
nand_4 g03402(new_n3779, new_n3778, new_n3777);
xnor_3 g03403(new_n3780, new_n3779, new_n3776);
xnor_3 g03404(new_n3781, new_n3780, new_n3752);
xnor_3 g03405(new_n3782, new_n3781, new_n3709);
xnor_3 g03406(new_n3783, new_n3782, new_n3750);
nor_4  g03407(new_n3784, new_n3712, new_n3710);
not_3  g03408(new_n3785, new_n3784);
not_3  g03409(new_n3786, new_n3679);
not_3  g03410(new_n3787, new_n3713);
nand_4 g03411(new_n3788, new_n3787, new_n3786);
nand_4 g03412(new_n3789, new_n3788, new_n3785);
xnor_3 g03413(new_n3790, new_n3789, new_n3783);
xnor_3 g03414(new_n3791, new_n3790, new_n3717);
not_3  g03415(new_n3792, new_n3791);
nor_4  g03416(new_n3793, new_n3792, new_n3411);
nor_4  g03417(new_n3794, new_n3791, new_n3410);
xor_3  g03418(new_n3795, new_n3403, new_n3402);
nand_4 g03419(new_n3796, new_n3645, new_n3640);
xnor_3 g03420(new_n3797, new_n3796, new_n3714);
nand_4 g03421(new_n3798, new_n3797, new_n3795);
not_3  g03422(new_n3799, new_n3798);
nor_4  g03423(new_n3800, new_n3797, new_n3795);
nor_4  g03424(new_n3801, new_n3800, new_n3799);
not_3  g03425(new_n3802, new_n3401);
xor_3  g03426(new_n3803, new_n3802, new_n3396);
nand_4 g03427(new_n3804, new_n3589, new_n3588);
xnor_3 g03428(new_n3805, new_n3804, new_n3636);
nor_4  g03429(new_n3806, new_n3805, new_n3803);
not_3  g03430(new_n3807, new_n3806);
not_3  g03431(new_n3808, new_n3584);
nor_4  g03432(new_n3809, new_n3808, new_n3570);
nor_4  g03433(new_n3810, new_n3809, new_n3585);
not_3  g03434(new_n3811, new_n3391);
nand_4 g03435(new_n3812, n9956, n7862);
not_3  g03436(new_n3813, new_n3812);
nor_4  g03437(new_n3814, new_n3813, new_n3336);
not_3  g03438(new_n3815, new_n3814);
nand_4 g03439(new_n3816, new_n3815, new_n3811);
nand_4 g03440(new_n3817, new_n3814, new_n3335);
nand_4 g03441(new_n3818, new_n3817, new_n3816);
not_3  g03442(new_n3819, new_n3818);
nor_4  g03443(new_n3820, new_n3819, new_n3810);
not_3  g03444(new_n3821, new_n3810);
nor_4  g03445(new_n3822, new_n3818, new_n3821);
nor_4  g03446(new_n3823, new_n3822, new_n3820);
not_3  g03447(new_n3824, new_n3823);
xor_3  g03448(new_n3825, new_n3579, new_n3434);
nor_4  g03449(new_n3826, new_n3825, new_n3812);
xor_3  g03450(new_n3827, new_n3393, new_n3392);
nor_4  g03451(new_n3828, new_n3827, new_n3826);
xor_3  g03452(new_n3829, new_n3582, new_n3580);
xnor_3 g03453(new_n3830, new_n3827, new_n3826);
nor_4  g03454(new_n3831, new_n3830, new_n3829);
nor_4  g03455(new_n3832, new_n3831, new_n3828);
nor_4  g03456(new_n3833, new_n3832, new_n3824);
nor_4  g03457(new_n3834, new_n3833, new_n3820);
not_3  g03458(new_n3835, new_n3803);
not_3  g03459(new_n3836, new_n3805);
nor_4  g03460(new_n3837, new_n3836, new_n3835);
nor_4  g03461(new_n3838, new_n3837, new_n3806);
nand_4 g03462(new_n3839, new_n3838, new_n3834);
nand_4 g03463(new_n3840, new_n3839, new_n3807);
nand_4 g03464(new_n3841, new_n3840, new_n3801);
nand_4 g03465(new_n3842_1, new_n3841, new_n3798);
nor_4  g03466(new_n3843, new_n3842_1, new_n3794);
nor_4  g03467(new_n3844, new_n3843, new_n3793);
nor_4  g03468(new_n3845, new_n3844, new_n3408);
not_3  g03469(new_n3846, new_n3408);
not_3  g03470(new_n3847, new_n3844);
nor_4  g03471(new_n3848, new_n3847, new_n3846);
nor_4  g03472(new_n3849_1, new_n3848, new_n3845);
nor_4  g03473(new_n3850, new_n3500, new_n3492);
not_3  g03474(new_n3851, new_n3850);
not_3  g03475(new_n3852, new_n3471);
nand_4 g03476(new_n3853, new_n3478, new_n3475);
nand_4 g03477(new_n3854, new_n3853, new_n3852);
nand_4 g03478(new_n3855, n9400, n8065);
not_3  g03479(new_n3856, new_n3855);
nand_4 g03480(new_n3857, n10439, n2464);
nand_4 g03481(new_n3858, n10391, n6877);
xor_3  g03482(new_n3859, new_n3858, new_n3857);
xnor_3 g03483(new_n3860, new_n3859, new_n3856);
xnor_3 g03484(new_n3861, new_n3860, new_n3854);
not_3  g03485(new_n3862, new_n3861);
nor_4  g03486(new_n3863, new_n3469, new_n3468);
nand_4 g03487(new_n3864, n11311, n8595);
not_3  g03488(new_n3865_1, new_n3864);
xor_3  g03489(new_n3866, new_n3865_1, new_n3863);
nand_4 g03490(new_n3867, n4203, n3602);
not_3  g03491(new_n3868, new_n3867);
nand_4 g03492(new_n3869, n6126, n4187);
nand_4 g03493(new_n3870, n12753, n3719);
xnor_3 g03494(new_n3871, new_n3870, new_n3869);
xnor_3 g03495(new_n3872, new_n3871, new_n3868);
xnor_3 g03496(new_n3873, new_n3872, new_n3866);
not_3  g03497(new_n3874, new_n3873);
xor_3  g03498(new_n3875, new_n3874, new_n3862);
nor_4  g03499(new_n3876, new_n3484, new_n3480);
nor_4  g03500(new_n3877, new_n3482, new_n3481);
not_3  g03501(new_n3878, new_n3877);
not_3  g03502(new_n3879, new_n3485);
not_3  g03503(new_n3880, new_n3491);
nand_4 g03504(new_n3881, new_n3880, new_n3879);
nor_4  g03505(new_n3882, new_n3881, new_n3878);
nor_4  g03506(new_n3883, new_n3491, new_n3485);
nor_4  g03507(new_n3884, new_n3883, new_n3877);
nor_4  g03508(new_n3885, new_n3884, new_n3882);
nor_4  g03509(new_n3886, new_n3885, new_n3876);
xnor_3 g03510(new_n3887, new_n3886, new_n3875);
xnor_3 g03511(new_n3888, new_n3887, new_n3851);
nand_4 g03512(new_n3889, new_n3501, new_n3466);
not_3  g03513(new_n3890, new_n3889);
nor_4  g03514(new_n3891, new_n3502, new_n3464);
nor_4  g03515(new_n3892, new_n3891, new_n3890);
xnor_3 g03516(new_n3893, new_n3892, new_n3888);
not_3  g03517(new_n3894, new_n3779);
nor_4  g03518(new_n3895, new_n3894, new_n3776);
not_3  g03519(new_n3896, new_n3895);
nand_4 g03520(new_n3897, n10965, n4805);
not_3  g03521(new_n3898, new_n3897);
nand_4 g03522(new_n3899, n5283, n4970);
nand_4 g03523(new_n3900, n11478, n503);
not_3  g03524(new_n3901, new_n3900);
xor_3  g03525(new_n3902, new_n3901, new_n3899);
xnor_3 g03526(new_n3903, new_n3902, new_n3898);
not_3  g03527(new_n3904, new_n3757);
nand_4 g03528(new_n3905, new_n3765, new_n3761);
nand_4 g03529(new_n3906, new_n3905, new_n3904);
xnor_3 g03530(new_n3907, new_n3906, new_n3903);
nor_4  g03531(new_n3908, new_n3755, new_n3754_1);
nand_4 g03532(new_n3909, n7610, n137);
not_3  g03533(new_n3910, new_n3909);
xor_3  g03534(new_n3911, new_n3910, new_n3908);
nand_4 g03535(new_n3912, n7733, n6797);
nand_4 g03536(new_n3913, n6294, n4826);
not_3  g03537(new_n3914, new_n3913);
nand_4 g03538(new_n3915, n12925, n3146);
not_3  g03539(new_n3916, new_n3915);
nor_4  g03540(new_n3917, new_n3916, new_n3914);
nor_4  g03541(new_n3918, new_n3915, new_n3913);
nor_4  g03542(new_n3919, new_n3918, new_n3917);
xor_3  g03543(new_n3920, new_n3919, new_n3912);
xnor_3 g03544(new_n3921, new_n3920, new_n3911);
xnor_3 g03545(new_n3922, new_n3921, new_n3907);
not_3  g03546(new_n3923, new_n3766);
nand_4 g03547(new_n3924, new_n3769, new_n3923);
nor_4  g03548(new_n3925, new_n3768, new_n3767);
nand_4 g03549(new_n3926, new_n3775, new_n3770);
not_3  g03550(new_n3927, new_n3926);
xnor_3 g03551(new_n3928, new_n3927, new_n3925);
nand_4 g03552(new_n3929, new_n3928, new_n3924);
xnor_3 g03553(new_n3930, new_n3929, new_n3922);
xnor_3 g03554(new_n3931, new_n3930, new_n3896);
nor_4  g03555(new_n3932_1, new_n3780, new_n3752);
not_3  g03556(new_n3933, new_n3932_1);
not_3  g03557(new_n3934, new_n3709);
not_3  g03558(new_n3935, new_n3780);
nor_4  g03559(new_n3936, new_n3935, new_n3751);
nor_4  g03560(new_n3937, new_n3932_1, new_n3936);
nand_4 g03561(new_n3938, new_n3937, new_n3934);
nand_4 g03562(new_n3939, new_n3938, new_n3933);
xnor_3 g03563(new_n3940, new_n3939, new_n3931);
not_3  g03564(new_n3941, new_n3742);
not_3  g03565(new_n3942, new_n3744);
nor_4  g03566(new_n3943, new_n3942, new_n3941);
nand_4 g03567(new_n3944, n11296, n7236);
nand_4 g03568(new_n3945, n8384, n6611);
nand_4 g03569(new_n3946, n6359, n3992);
not_3  g03570(new_n3947, new_n3946);
xor_3  g03571(new_n3948, new_n3947, new_n3945);
xnor_3 g03572(new_n3949, new_n3948, new_n3944);
nand_4 g03573(new_n3950, new_n3727, new_n3721);
not_3  g03574(new_n3951, new_n3728);
not_3  g03575(new_n3952, new_n3731);
nand_4 g03576(new_n3953, new_n3952, new_n3951);
nand_4 g03577(new_n3954, new_n3953, new_n3950);
xnor_3 g03578(new_n3955, new_n3954, new_n3949);
nor_4  g03579(new_n3956, new_n3730, new_n3729);
not_3  g03580(new_n3957, new_n3956);
nand_4 g03581(new_n3958, n6358, n217);
xor_3  g03582(new_n3959, new_n3958, new_n3957);
nand_4 g03583(new_n3960, n1471, n405);
not_3  g03584(new_n3961, new_n3960);
nand_4 g03585(new_n3962, n5198, n4086);
nand_4 g03586(new_n3963, n8433, n7646);
xor_3  g03587(new_n3964, new_n3963, new_n3962);
xnor_3 g03588(new_n3965, new_n3964, new_n3961);
xnor_3 g03589(new_n3966, new_n3965, new_n3959);
xnor_3 g03590(new_n3967, new_n3966, new_n3955);
nand_4 g03591(new_n3968, new_n3736, new_n3733);
nor_4  g03592(new_n3969, new_n3735, new_n3734);
nor_4  g03593(new_n3970, new_n3741, new_n3737);
xnor_3 g03594(new_n3971, new_n3970, new_n3969);
nand_4 g03595(new_n3972, new_n3971, new_n3968);
xnor_3 g03596(new_n3973, new_n3972, new_n3967);
xnor_3 g03597(new_n3974, new_n3973, new_n3943);
nand_4 g03598(new_n3975, new_n3745, new_n3718);
nand_4 g03599(new_n3976, new_n3748, new_n3975);
xnor_3 g03600(new_n3977, new_n3976, new_n3974);
xnor_3 g03601(new_n3978, new_n3977, new_n3940);
not_3  g03602(new_n3979, new_n3782);
nand_4 g03603(new_n3980, new_n3979, new_n3750);
nand_4 g03604(new_n3981, new_n3789, new_n3783);
nand_4 g03605(new_n3982, new_n3981, new_n3980);
xnor_3 g03606(new_n3983, new_n3982, new_n3978);
xnor_3 g03607(new_n3984, new_n3983, new_n3893);
not_3  g03608(new_n3985, new_n3984);
not_3  g03609(new_n3986_1, new_n3716);
nand_4 g03610(new_n3987, new_n3986_1, new_n3503);
not_3  g03611(new_n3988, new_n3790);
nand_4 g03612(new_n3989, new_n3988, new_n3717);
nand_4 g03613(new_n3990, new_n3989, new_n3987);
xnor_3 g03614(new_n3991, new_n3990, new_n3985);
xnor_3 g03615(n844, new_n3991, new_n3849_1);
nand_4 g03616(new_n3993, n7456, n6687);
not_3  g03617(new_n3994, new_n3993);
nand_4 g03618(new_n3995, n12591, n6687);
not_3  g03619(new_n3996, new_n3995);
nand_4 g03620(new_n3997, n4189, n1798);
not_3  g03621(new_n3998, new_n3997);
nor_4  g03622(new_n3999, new_n3998, new_n3996);
nor_4  g03623(new_n4000, new_n3997, new_n3995);
nand_4 g03624(new_n4001, n3932, n2564);
not_3  g03625(new_n4002, new_n4001);
nor_4  g03626(new_n4003, new_n4002, new_n4000);
nor_4  g03627(new_n4004, new_n4003, new_n3999);
nand_4 g03628(new_n4005_1, new_n4004, new_n3994);
not_3  g03629(new_n4006, new_n4005_1);
nor_4  g03630(new_n4007, new_n4004, new_n3994);
nor_4  g03631(new_n4008, new_n4007, new_n4006);
nand_4 g03632(new_n4009, n4189, n3932);
nand_4 g03633(new_n4010, n12591, n2564);
not_3  g03634(new_n4011, new_n4010);
nand_4 g03635(new_n4012, n6770, n1798);
not_3  g03636(new_n4013, new_n4012);
nor_4  g03637(new_n4014, new_n4013, new_n4011);
nor_4  g03638(new_n4015, new_n4012, new_n4010);
nor_4  g03639(new_n4016, new_n4015, new_n4014);
xnor_3 g03640(new_n4017, new_n4016, new_n4009);
xor_3  g03641(new_n4018, new_n4017, new_n4008);
not_3  g03642(new_n4019, new_n4018);
nand_4 g03643(new_n4020, n6687, n1798);
not_3  g03644(new_n4021, new_n4020);
nor_4  g03645(new_n4022, new_n4021, new_n4001);
nor_4  g03646(new_n4023, new_n4000, new_n3999);
nor_4  g03647(new_n4024, new_n4023, new_n4022);
not_3  g03648(new_n4025, new_n4024);
nor_4  g03649(new_n4026, new_n4025, new_n4001);
not_3  g03650(new_n4027, new_n4026);
xor_3  g03651(new_n4028, new_n4027, new_n4019);
not_3  g03652(new_n4029, new_n4028);
nand_4 g03653(new_n4030, n8336, n6703);
nand_4 g03654(new_n4031, n11876, n11222);
not_3  g03655(new_n4032, new_n4031);
nand_4 g03656(new_n4033, n12069, n5645);
xor_3  g03657(new_n4034, new_n4033, new_n4032);
nor_4  g03658(new_n4035, new_n4034, new_n4030);
nand_4 g03659(new_n4036, n9640, n8336);
nand_4 g03660(new_n4037, n10928, n6703);
not_3  g03661(new_n4038, new_n4037);
xor_3  g03662(new_n4039, new_n4038, new_n4036);
not_3  g03663(new_n4040, new_n4039);
nand_4 g03664(new_n4041, new_n4040, new_n4035);
not_3  g03665(new_n4042, new_n4041);
nor_4  g03666(new_n4043, new_n4033, new_n4031);
not_3  g03667(new_n4044, new_n4043);
nand_4 g03668(new_n4045, n12391, n5645);
nand_4 g03669(new_n4046, n12069, n1067);
xnor_3 g03670(new_n4047, new_n4046, new_n4045);
nor_4  g03671(new_n4048, new_n4047, new_n4044);
not_3  g03672(new_n4049, new_n4047);
nor_4  g03673(new_n4050, new_n4049, new_n4043);
nor_4  g03674(new_n4051, new_n4050, new_n4048);
not_3  g03675(new_n4052, new_n4051);
nand_4 g03676(new_n4053, n11222, n10898);
nand_4 g03677(new_n4054, n11876, n11153);
xor_3  g03678(new_n4055, new_n4054, new_n4053);
xnor_3 g03679(new_n4056, new_n4055, new_n4052);
not_3  g03680(new_n4057, new_n4056);
not_3  g03681(new_n4058, new_n4035);
xor_3  g03682(new_n4059, new_n4040, new_n4058);
nor_4  g03683(new_n4060, new_n4059, new_n4057);
nor_4  g03684(new_n4061, new_n4060, new_n4042);
not_3  g03685(new_n4062, new_n4030);
nand_4 g03686(new_n4063, n10928, n9640);
nor_4  g03687(new_n4064, new_n4063, new_n4062);
nand_4 g03688(new_n4065, n6986, n6703);
nand_4 g03689(new_n4066, n8336, n3022);
nand_4 g03690(new_n4067, new_n4066, new_n4065);
and_4  g03691(new_n4068, new_n4067, new_n4064);
nor_4  g03692(new_n4069, new_n4066, new_n4065);
nor_4  g03693(new_n4070, new_n4067, new_n4064);
nor_4  g03694(new_n4071, new_n4070, new_n4069);
not_3  g03695(new_n4072, new_n4071);
nor_4  g03696(new_n4073, new_n4072, new_n4068);
not_3  g03697(new_n4074, new_n4073);
xnor_3 g03698(new_n4075, new_n4074, new_n4061);
nor_4  g03699(new_n4076, new_n4046, new_n4045);
nand_4 g03700(new_n4077, n12069, n8665);
not_3  g03701(new_n4078, new_n4077);
nand_4 g03702(new_n4079, n12391, n1067);
nand_4 g03703(new_n4080, n7891, n5645);
xnor_3 g03704(new_n4081, new_n4080, new_n4079);
xor_3  g03705(new_n4082, new_n4081, new_n4078);
not_3  g03706(new_n4083, new_n4082);
xor_3  g03707(new_n4084, new_n4083, new_n4076);
nor_4  g03708(new_n4085, new_n4055, new_n4052);
nor_4  g03709(new_n4086_1, new_n4085, new_n4050);
nand_4 g03710(new_n4087, n11876, n5314);
nand_4 g03711(new_n4088_1, n11222, n3754);
nor_4  g03712(new_n4089, new_n4088_1, new_n4087);
nand_4 g03713(new_n4090, new_n4088_1, new_n4087);
nand_4 g03714(new_n4091, n11153, n10898);
nor_4  g03715(new_n4092, new_n4091, new_n4032);
nor_4  g03716(new_n4093, new_n4092, new_n4090);
nor_4  g03717(new_n4094_1, new_n4093, new_n4089);
not_3  g03718(new_n4095, new_n4094_1);
not_3  g03719(new_n4096, new_n4090);
not_3  g03720(new_n4097, new_n4092);
nor_4  g03721(new_n4098, new_n4097, new_n4096);
nor_4  g03722(new_n4099, new_n4098, new_n4095);
xnor_3 g03723(new_n4100, new_n4099, new_n4086_1);
xnor_3 g03724(new_n4101, new_n4100, new_n4084);
xnor_3 g03725(new_n4102, new_n4101, new_n4075);
not_3  g03726(new_n4103, new_n3999);
nand_4 g03727(new_n4104, new_n4022, new_n4103);
nand_4 g03728(new_n4105, new_n4104, new_n4025);
not_3  g03729(new_n4106, new_n4105);
nand_4 g03730(new_n4107, new_n4106, new_n4102);
xor_3  g03731(new_n4108, new_n4033, new_n4031);
xor_3  g03732(new_n4109, new_n4108, new_n4062);
nand_4 g03733(new_n4110, new_n4109, new_n4021);
not_3  g03734(new_n4111, new_n4110);
nand_4 g03735(new_n4112, n2564, n1798);
nand_4 g03736(new_n4113, n6687, n3932);
xor_3  g03737(new_n4114, new_n4113, new_n4112);
nor_4  g03738(new_n4115, new_n4114, new_n4111);
and_4  g03739(new_n4116, new_n4059, new_n4057);
nor_4  g03740(new_n4117, new_n4116, new_n4060);
not_3  g03741(new_n4118, new_n4114);
xor_3  g03742(new_n4119, new_n4118, new_n4111);
nor_4  g03743(new_n4120, new_n4119, new_n4117);
nor_4  g03744(new_n4121, new_n4120, new_n4115);
xnor_3 g03745(new_n4122, new_n4105, new_n4102);
nand_4 g03746(new_n4123, new_n4122, new_n4121);
nand_4 g03747(new_n4124, new_n4123, new_n4107);
xnor_3 g03748(new_n4125, new_n4124, new_n4029);
not_3  g03749(new_n4126, new_n4076);
nor_4  g03750(new_n4127, new_n4082, new_n4126);
nand_4 g03751(new_n4128, n12069, n11922);
not_3  g03752(new_n4129, new_n4128);
not_3  g03753(new_n4130, new_n4079);
not_3  g03754(new_n4131, new_n4080);
nor_4  g03755(new_n4132, new_n4131, new_n4130);
nor_4  g03756(new_n4133, new_n4081, new_n4078);
nor_4  g03757(new_n4134, new_n4133, new_n4132);
xnor_3 g03758(new_n4135, new_n4134, new_n4129);
nand_4 g03759(new_n4136, n7160, n5645);
nand_4 g03760(new_n4137, n7891, n1067);
nand_4 g03761(new_n4138, n12391, n8665);
nand_4 g03762(new_n4139, new_n4138, new_n4137);
nor_4  g03763(new_n4140, new_n4138, new_n4137);
not_3  g03764(new_n4141_1, new_n4140);
nand_4 g03765(new_n4142, new_n4141_1, new_n4139);
xnor_3 g03766(new_n4143, new_n4142, new_n4136);
xnor_3 g03767(new_n4144, new_n4143, new_n4135);
xnor_3 g03768(new_n4145, new_n4144, new_n4127);
nand_4 g03769(new_n4146, n11222, n2749);
not_3  g03770(new_n4147, new_n4146);
not_3  g03771(new_n4148, new_n4091);
nor_4  g03772(new_n4149, new_n4148, new_n4089);
nor_4  g03773(new_n4150, new_n4149, new_n4096);
xnor_3 g03774(new_n4151, new_n4150, new_n4147);
nand_4 g03775(new_n4152, n10898, n5314);
nand_4 g03776(new_n4153, n11153, n3754);
not_3  g03777(new_n4154, new_n4153);
nand_4 g03778(new_n4155_1, n11876, n996);
not_3  g03779(new_n4156, new_n4155_1);
nor_4  g03780(new_n4157, new_n4156, new_n4154);
nor_4  g03781(new_n4158, new_n4155_1, new_n4153);
nor_4  g03782(new_n4159_1, new_n4158, new_n4157);
xnor_3 g03783(new_n4160, new_n4159_1, new_n4152);
not_3  g03784(new_n4161, new_n4160);
xnor_3 g03785(new_n4162, new_n4161, new_n4151);
nor_4  g03786(new_n4163, new_n4094_1, new_n4091);
not_3  g03787(new_n4164, new_n4163);
nor_4  g03788(new_n4165, new_n4164, new_n4162);
not_3  g03789(new_n4166, new_n4162);
nor_4  g03790(new_n4167, new_n4163, new_n4166);
nor_4  g03791(new_n4168, new_n4167, new_n4165);
nor_4  g03792(new_n4169, new_n4168, new_n4145);
not_3  g03793(new_n4170, new_n4144);
xnor_3 g03794(new_n4171, new_n4170, new_n4127);
not_3  g03795(new_n4172, new_n4168);
nor_4  g03796(new_n4173, new_n4172, new_n4171);
nor_4  g03797(new_n4174, new_n4173, new_n4169);
nor_4  g03798(new_n4175, new_n4099, new_n4086_1);
nor_4  g03799(new_n4176, new_n4100, new_n4084);
nor_4  g03800(new_n4177, new_n4176, new_n4175);
not_3  g03801(new_n4178, new_n4177);
nor_4  g03802(new_n4179, new_n4178, new_n4174);
nand_4 g03803(new_n4180, new_n4178, new_n4174);
not_3  g03804(new_n4181, new_n4180);
nor_4  g03805(new_n4182, new_n4181, new_n4179);
not_3  g03806(new_n4183, new_n4182);
nand_4 g03807(new_n4184, n11023, n8336);
not_3  g03808(new_n4185, new_n4069);
not_3  g03809(new_n4186, new_n4063);
nand_4 g03810(new_n4187_1, new_n4067, new_n4186);
nand_4 g03811(new_n4188, new_n4187_1, new_n4185);
not_3  g03812(new_n4189_1, new_n4188);
xor_3  g03813(new_n4190_1, new_n4189_1, new_n4184);
nand_4 g03814(new_n4191, n9640, n6986);
not_3  g03815(new_n4192, new_n4191);
nand_4 g03816(new_n4193, n10928, n3022);
not_3  g03817(new_n4194, new_n4193);
nand_4 g03818(new_n4195, n6703, n2226);
not_3  g03819(new_n4196, new_n4195);
nor_4  g03820(new_n4197, new_n4196, new_n4194);
nor_4  g03821(new_n4198, new_n4195, new_n4193);
nor_4  g03822(new_n4199, new_n4198, new_n4197);
xor_3  g03823(new_n4200, new_n4199, new_n4192);
xnor_3 g03824(new_n4201, new_n4200, new_n4190_1);
not_3  g03825(new_n4202, new_n4201);
nor_4  g03826(new_n4203_1, new_n4071, new_n4063);
xor_3  g03827(new_n4204, new_n4203_1, new_n4202);
nand_4 g03828(new_n4205, new_n4074, new_n4061);
not_3  g03829(new_n4206, new_n4205);
nor_4  g03830(new_n4207, new_n4101, new_n4075);
nor_4  g03831(new_n4208, new_n4207, new_n4206);
nand_4 g03832(new_n4209, new_n4208, new_n4204);
not_3  g03833(new_n4210, new_n4209);
nor_4  g03834(new_n4211, new_n4208, new_n4204);
nor_4  g03835(new_n4212, new_n4211, new_n4210);
nor_4  g03836(new_n4213, new_n4212, new_n4183);
nand_4 g03837(new_n4214, new_n4212, new_n4183);
not_3  g03838(new_n4215, new_n4214);
nor_4  g03839(new_n4216, new_n4215, new_n4213);
xor_3  g03840(n911, new_n4216, new_n4125);
nand_4 g03841(new_n4218, n9956, n4189);
nand_4 g03842(new_n4219, n11917, n6687);
nand_4 g03843(new_n4220, new_n4219, new_n4218);
nor_4  g03844(new_n4221, new_n4219, new_n4218);
not_3  g03845(new_n4222, new_n4221);
and_4  g03846(new_n4223, new_n4222, new_n4220);
nand_4 g03847(new_n4224, n9956, n2564);
nand_4 g03848(new_n4225, n6687, n4921);
nor_4  g03849(new_n4226_1, new_n4225, new_n4224);
not_3  g03850(new_n4227, new_n4226_1);
nor_4  g03851(new_n4228, new_n4227, new_n4223);
not_3  g03852(new_n4229, new_n4228);
nand_4 g03853(new_n4230_1, n6687, n3842);
nand_4 g03854(new_n4231, n4921, n2564);
not_3  g03855(new_n4232, new_n4231);
nand_4 g03856(new_n4233, new_n4232, new_n4220);
nand_4 g03857(new_n4234, new_n4233, new_n4222);
not_3  g03858(new_n4235, new_n4234);
xor_3  g03859(new_n4236, new_n4235, new_n4230_1);
nand_4 g03860(new_n4237, n4921, n4189);
not_3  g03861(new_n4238, new_n4237);
nand_4 g03862(new_n4239, n11917, n2564);
not_3  g03863(new_n4240, new_n4239);
nand_4 g03864(new_n4241, n9956, n6770);
not_3  g03865(new_n4242, new_n4241);
nor_4  g03866(new_n4243, new_n4242, new_n4240);
nor_4  g03867(new_n4244, new_n4241, new_n4239);
nor_4  g03868(new_n4245, new_n4244, new_n4243);
xor_3  g03869(new_n4246, new_n4245, new_n4238);
xnor_3 g03870(new_n4247, new_n4246, new_n4236);
nor_4  g03871(new_n4248, new_n4247, new_n4229);
not_3  g03872(new_n4249, new_n4248);
nand_4 g03873(new_n4250, n6687, n2577);
nor_4  g03874(new_n4251, new_n4235, new_n4230_1);
not_3  g03875(new_n4252, new_n4251);
nand_4 g03876(new_n4253, new_n4246, new_n4236);
nand_4 g03877(new_n4254, new_n4253, new_n4252);
not_3  g03878(new_n4255, new_n4254);
xor_3  g03879(new_n4256, new_n4255, new_n4250);
nand_4 g03880(new_n4257, n3842, n2564);
nor_4  g03881(new_n4258, new_n4244, new_n4238);
nor_4  g03882(new_n4259, new_n4258, new_n4243);
xor_3  g03883(new_n4260, new_n4259, new_n4257);
not_3  g03884(new_n4261, new_n4260);
nand_4 g03885(new_n4262, n6770, n4921);
nand_4 g03886(new_n4263, n11917, n4189);
nand_4 g03887(new_n4264, n9956, n9920);
not_3  g03888(new_n4265, new_n4264);
xor_3  g03889(new_n4266, new_n4265, new_n4263);
xnor_3 g03890(new_n4267, new_n4266, new_n4262);
not_3  g03891(new_n4268, new_n4267);
xor_3  g03892(new_n4269, new_n4268, new_n4261);
xnor_3 g03893(new_n4270, new_n4269, new_n4256);
xnor_3 g03894(new_n4271, new_n4270, new_n4249);
not_3  g03895(new_n4272, new_n4247);
xor_3  g03896(new_n4273, new_n4272, new_n4229);
not_3  g03897(new_n4274, new_n4273);
nand_4 g03898(new_n4275, n8595, n8336);
not_3  g03899(new_n4276, new_n4275);
nand_4 g03900(new_n4277, n8336, n6126);
not_3  g03901(new_n4278, new_n4277);
nand_4 g03902(new_n4279, n6986, n3719);
not_3  g03903(new_n4280, new_n4279);
nor_4  g03904(new_n4281, new_n4280, new_n4278);
nor_4  g03905(new_n4282, new_n4279, new_n4277);
nand_4 g03906(new_n4283, n10928, n3602);
not_3  g03907(new_n4284, new_n4283);
nor_4  g03908(new_n4285, new_n4284, new_n4282);
nor_4  g03909(new_n4286, new_n4285, new_n4281);
nand_4 g03910(new_n4287, new_n4286, new_n4276);
not_3  g03911(new_n4288, new_n4287);
nor_4  g03912(new_n4289, new_n4286, new_n4276);
nor_4  g03913(new_n4290, new_n4289, new_n4288);
nand_4 g03914(new_n4291, n6986, n3602);
not_3  g03915(new_n4292, new_n4291);
nand_4 g03916(new_n4293, n10928, n6126);
nand_4 g03917(new_n4294, n3719, n2226);
not_3  g03918(new_n4295, new_n4294);
xor_3  g03919(new_n4296, new_n4295, new_n4293);
xnor_3 g03920(new_n4297, new_n4296, new_n4292);
nand_4 g03921(new_n4298, new_n4297, new_n4290);
not_3  g03922(new_n4299, new_n4290);
xnor_3 g03923(new_n4300_1, new_n4296, new_n4291);
nand_4 g03924(new_n4301, new_n4300_1, new_n4299);
nand_4 g03925(new_n4302, new_n4301, new_n4298);
nand_4 g03926(new_n4303, n8336, n3719);
not_3  g03927(new_n4304, new_n4303);
nor_4  g03928(new_n4305, new_n4304, new_n4283);
nor_4  g03929(new_n4306, new_n4282, new_n4281);
nor_4  g03930(new_n4307, new_n4306, new_n4305);
not_3  g03931(new_n4308, new_n4307);
nor_4  g03932(new_n4309, new_n4308, new_n4283);
xnor_3 g03933(new_n4310, new_n4309, new_n4302);
nand_4 g03934(new_n4311, n12925, n7891);
nand_4 g03935(new_n4312_1, n12069, n4826);
nand_4 g03936(new_n4313, new_n4312_1, new_n4311);
not_3  g03937(new_n4314, new_n4313);
not_3  g03938(new_n4315, new_n4311);
not_3  g03939(new_n4316, new_n4312_1);
nand_4 g03940(new_n4317, new_n4316, new_n4315);
not_3  g03941(new_n4318, new_n4317);
nor_4  g03942(new_n4319, new_n4318, new_n4314);
nand_4 g03943(new_n4320, n12069, n7733);
nand_4 g03944(new_n4321, n12925, n12391);
nor_4  g03945(new_n4322, new_n4321, new_n4320);
not_3  g03946(new_n4323, new_n4322);
nor_4  g03947(new_n4324, new_n4323, new_n4319);
not_3  g03948(new_n4325, new_n4324);
nand_4 g03949(new_n4326_1, n12069, n7610);
nand_4 g03950(new_n4327, n12391, n7733);
not_3  g03951(new_n4328, new_n4327);
nand_4 g03952(new_n4329, new_n4328, new_n4313);
nand_4 g03953(new_n4330, new_n4329, new_n4317);
not_3  g03954(new_n4331, new_n4330);
xnor_3 g03955(new_n4332, new_n4331, new_n4326_1);
nand_4 g03956(new_n4333_1, n12925, n7160);
not_3  g03957(new_n4334, new_n4333_1);
nand_4 g03958(new_n4335, n12391, n4826);
not_3  g03959(new_n4336, new_n4335);
nand_4 g03960(new_n4337, n7891, n7733);
not_3  g03961(new_n4338, new_n4337);
nor_4  g03962(new_n4339, new_n4338, new_n4336);
nor_4  g03963(new_n4340, new_n4337, new_n4335);
nor_4  g03964(new_n4341, new_n4340, new_n4339);
xnor_3 g03965(new_n4342, new_n4341, new_n4334);
xnor_3 g03966(new_n4343, new_n4342, new_n4332);
nor_4  g03967(new_n4344, new_n4343, new_n4325);
not_3  g03968(new_n4345, new_n4343);
nor_4  g03969(new_n4346, new_n4345, new_n4324);
nor_4  g03970(new_n4347, new_n4346, new_n4344);
nand_4 g03971(new_n4348, n11222, n217);
not_3  g03972(new_n4349, new_n4348);
nand_4 g03973(new_n4350, n8433, n5314);
not_3  g03974(new_n4351, new_n4350);
nand_4 g03975(new_n4352, n11222, n4086);
not_3  g03976(new_n4353, new_n4352);
nor_4  g03977(new_n4354, new_n4353, new_n4351);
nor_4  g03978(new_n4355, new_n4352, new_n4350);
nand_4 g03979(new_n4356, n11153, n405);
not_3  g03980(new_n4357, new_n4356);
nor_4  g03981(new_n4358, new_n4357, new_n4355);
nor_4  g03982(new_n4359, new_n4358, new_n4354);
xnor_3 g03983(new_n4360, new_n4359, new_n4349);
nand_4 g03984(new_n4361, n5314, n405);
nand_4 g03985(new_n4362, n8433, n996);
nand_4 g03986(new_n4363, n11153, n4086);
xnor_3 g03987(new_n4364, new_n4363, new_n4362);
xnor_3 g03988(new_n4365, new_n4364, new_n4361);
xnor_3 g03989(new_n4366, new_n4365, new_n4360);
not_3  g03990(new_n4367, new_n4355);
nand_4 g03991(new_n4368, n11222, n8433);
nand_4 g03992(new_n4369, new_n4368, new_n4357);
nand_4 g03993(new_n4370_1, new_n4369, new_n4354);
nand_4 g03994(new_n4371, new_n4370_1, new_n4367);
not_3  g03995(new_n4372, new_n4371);
nor_4  g03996(new_n4373, new_n4372, new_n4356);
not_3  g03997(new_n4374, new_n4373);
nor_4  g03998(new_n4375, new_n4374, new_n4366);
not_3  g03999(new_n4376, new_n4366);
nor_4  g04000(new_n4377, new_n4373, new_n4376);
nor_4  g04001(new_n4378_1, new_n4377, new_n4375);
not_3  g04002(new_n4379, new_n4378_1);
xnor_3 g04003(new_n4380, new_n4379, new_n4347);
nand_4 g04004(new_n4381, n12925, n12069);
nor_4  g04005(new_n4382, new_n4381, new_n4368);
not_3  g04006(new_n4383, new_n4382);
nand_4 g04007(new_n4384, n11153, n8433);
nand_4 g04008(new_n4385, n11222, n405);
xnor_3 g04009(new_n4386, new_n4385, new_n4384);
nand_4 g04010(new_n4387, new_n4386, new_n4383);
not_3  g04011(new_n4388, new_n4387);
nor_4  g04012(new_n4389, new_n4386, new_n4383);
nor_4  g04013(new_n4390, new_n4389, new_n4388);
xnor_3 g04014(new_n4391, new_n4321, new_n4320);
nand_4 g04015(new_n4392, new_n4391, new_n4390);
nand_4 g04016(new_n4393, new_n4392, new_n4387);
not_3  g04017(new_n4394, new_n4393);
nor_4  g04018(new_n4395, new_n4369, new_n4354);
nor_4  g04019(new_n4396, new_n4395, new_n4371);
nor_4  g04020(new_n4397_1, new_n4396, new_n4394);
not_3  g04021(new_n4398, new_n4397_1);
not_3  g04022(new_n4399, new_n4396);
nor_4  g04023(new_n4400, new_n4399, new_n4393);
nor_4  g04024(new_n4401, new_n4400, new_n4397_1);
not_3  g04025(new_n4402, new_n4319);
not_3  g04026(new_n4403, new_n4381);
nor_4  g04027(new_n4404, new_n4403, new_n4327);
not_3  g04028(new_n4405, new_n4404);
nand_4 g04029(new_n4406, new_n4405, new_n4402);
nand_4 g04030(new_n4407, new_n4404, new_n4313);
nand_4 g04031(new_n4408, new_n4407, new_n4406);
nand_4 g04032(new_n4409, new_n4408, new_n4401);
nand_4 g04033(new_n4410, new_n4409, new_n4398);
xnor_3 g04034(new_n4411, new_n4410, new_n4380);
xnor_3 g04035(new_n4412, new_n4411, new_n4310);
xnor_3 g04036(new_n4413, new_n4408, new_n4401);
not_3  g04037(new_n4414, new_n4413);
not_3  g04038(new_n4415, new_n4281);
nand_4 g04039(new_n4416, new_n4305, new_n4415);
nand_4 g04040(new_n4417, new_n4416, new_n4308);
nor_4  g04041(new_n4418, new_n4417, new_n4414);
xnor_3 g04042(new_n4419, new_n4417, new_n4414);
xnor_3 g04043(new_n4420, new_n4391, new_n4390);
not_3  g04044(new_n4421, new_n4420);
nand_4 g04045(new_n4422, n10928, n3719);
nand_4 g04046(new_n4423, n8336, n3602);
not_3  g04047(new_n4424, new_n4423);
xor_3  g04048(new_n4425, new_n4424, new_n4422);
nor_4  g04049(new_n4426, new_n4425, new_n4421);
xor_3  g04050(new_n4427, new_n4381, new_n4368);
nand_4 g04051(new_n4428, new_n4427, new_n4304);
xnor_3 g04052(new_n4429, new_n4425, new_n4421);
nor_4  g04053(new_n4430, new_n4429, new_n4428);
nor_4  g04054(new_n4431, new_n4430, new_n4426);
nor_4  g04055(new_n4432, new_n4431, new_n4419);
nor_4  g04056(new_n4433, new_n4432, new_n4418);
xnor_3 g04057(new_n4434, new_n4433, new_n4412);
not_3  g04058(new_n4435, new_n4434);
nand_4 g04059(new_n4436_1, new_n4435, new_n4274);
nand_4 g04060(new_n4437, new_n4434, new_n4273);
xnor_3 g04061(new_n4438, new_n4431, new_n4419);
not_3  g04062(new_n4439, new_n4438);
not_3  g04063(new_n4440, new_n4223);
nand_4 g04064(new_n4441, n9956, n6687);
not_3  g04065(new_n4442, new_n4441);
nor_4  g04066(new_n4443, new_n4442, new_n4231);
not_3  g04067(new_n4444, new_n4443);
nand_4 g04068(new_n4445, new_n4444, new_n4440);
nand_4 g04069(new_n4446, new_n4443, new_n4220);
nand_4 g04070(new_n4447, new_n4446, new_n4445);
not_3  g04071(new_n4448, new_n4447);
nor_4  g04072(new_n4449, new_n4448, new_n4439);
xnor_3 g04073(new_n4450, new_n4447, new_n4438);
not_3  g04074(new_n4451, new_n4428);
nor_4  g04075(new_n4452, new_n4427, new_n4304);
nor_4  g04076(new_n4453, new_n4452, new_n4451);
nand_4 g04077(new_n4454, new_n4453, new_n4442);
not_3  g04078(new_n4455, new_n4454);
xor_3  g04079(new_n4456, new_n4225, new_n4224);
nor_4  g04080(new_n4457, new_n4456, new_n4455);
not_3  g04081(new_n4458, new_n4429);
nor_4  g04082(new_n4459, new_n4458, new_n4451);
nor_4  g04083(new_n4460, new_n4459, new_n4430);
xnor_3 g04084(new_n4461, new_n4456, new_n4455);
nor_4  g04085(new_n4462, new_n4461, new_n4460);
nor_4  g04086(new_n4463, new_n4462, new_n4457);
nor_4  g04087(new_n4464, new_n4463, new_n4450);
nor_4  g04088(new_n4465, new_n4464, new_n4449);
nand_4 g04089(new_n4466, new_n4465, new_n4437);
nand_4 g04090(new_n4467, new_n4466, new_n4436_1);
xnor_3 g04091(new_n4468, new_n4467, new_n4271);
not_3  g04092(new_n4469, new_n4309);
nor_4  g04093(new_n4470, new_n4469, new_n4302);
nand_4 g04094(new_n4471, n10439, n8336);
not_3  g04095(new_n4472, new_n4471);
nand_4 g04096(new_n4473, new_n4298, new_n4287);
xnor_3 g04097(new_n4474, new_n4473, new_n4472);
nand_4 g04098(new_n4475, n10928, n8595);
not_3  g04099(new_n4476, new_n4475);
not_3  g04100(new_n4477, new_n4293);
nor_4  g04101(new_n4478, new_n4295, new_n4477);
nor_4  g04102(new_n4479, new_n4294, new_n4293);
nor_4  g04103(new_n4480, new_n4479, new_n4292);
nor_4  g04104(new_n4481, new_n4480, new_n4478);
xor_3  g04105(new_n4482, new_n4481, new_n4476);
not_3  g04106(new_n4483, new_n4482);
nand_4 g04107(new_n4484, n3602, n2226);
not_3  g04108(new_n4485, new_n4484);
nand_4 g04109(new_n4486, n6986, n6126);
nand_4 g04110(new_n4487, n3719, n1094);
xnor_3 g04111(new_n4488, new_n4487, new_n4486);
xor_3  g04112(new_n4489, new_n4488, new_n4485);
not_3  g04113(new_n4490, new_n4489);
xor_3  g04114(new_n4491, new_n4490, new_n4483);
nor_4  g04115(new_n4492, new_n4491, new_n4474);
xnor_3 g04116(new_n4493, new_n4473, new_n4471);
not_3  g04117(new_n4494, new_n4491);
nor_4  g04118(new_n4495, new_n4494, new_n4493);
nor_4  g04119(new_n4496, new_n4495, new_n4492);
xnor_3 g04120(new_n4497, new_n4496, new_n4470);
not_3  g04121(new_n4498, new_n4375);
nand_4 g04122(new_n4499_1, n11222, n6611);
not_3  g04123(new_n4500, new_n4499_1);
nand_4 g04124(new_n4501, n11153, n217);
nand_4 g04125(new_n4502, n996, n405);
nand_4 g04126(new_n4503, n5314, n4086);
not_3  g04127(new_n4504, new_n4503);
nand_4 g04128(new_n4505, n8433, n5767);
not_3  g04129(new_n4506, new_n4505);
nor_4  g04130(new_n4507, new_n4506, new_n4504);
nor_4  g04131(new_n4508, new_n4505, new_n4503);
nor_4  g04132(new_n4509, new_n4508, new_n4507);
xnor_3 g04133(new_n4510, new_n4509, new_n4502);
xnor_3 g04134(new_n4511, new_n4510, new_n4501);
not_3  g04135(new_n4512, new_n4511);
and_4  g04136(new_n4513, new_n4363, new_n4362);
not_3  g04137(new_n4514, new_n4361);
nor_4  g04138(new_n4515, new_n4363, new_n4362);
nor_4  g04139(new_n4516_1, new_n4515, new_n4514);
nor_4  g04140(new_n4517, new_n4516_1, new_n4513);
xnor_3 g04141(new_n4518, new_n4517, new_n4512);
nand_4 g04142(new_n4519, new_n4518, new_n4500);
xnor_3 g04143(new_n4520, new_n4517, new_n4511);
nand_4 g04144(new_n4521, new_n4520, new_n4499_1);
nand_4 g04145(new_n4522, new_n4521, new_n4519);
nand_4 g04146(new_n4523, new_n4359, new_n4349);
not_3  g04147(new_n4524, new_n4523);
nor_4  g04148(new_n4525, new_n4365, new_n4360);
nor_4  g04149(new_n4526, new_n4525, new_n4524);
xnor_3 g04150(new_n4527, new_n4526, new_n4522);
nor_4  g04151(new_n4528, new_n4527, new_n4498);
not_3  g04152(new_n4529, new_n4527);
nor_4  g04153(new_n4530, new_n4529, new_n4375);
nor_4  g04154(new_n4531, new_n4530, new_n4528);
not_3  g04155(new_n4532, new_n4344);
nand_4 g04156(new_n4533, n12069, n4970);
nand_4 g04157(new_n4534, n12391, n7610);
not_3  g04158(new_n4535, new_n4534);
nor_4  g04159(new_n4536, new_n4340, new_n4334);
nor_4  g04160(new_n4537, new_n4536, new_n4339);
xnor_3 g04161(new_n4538, new_n4537, new_n4535);
nand_4 g04162(new_n4539, n7733, n7160);
nand_4 g04163(new_n4540, n7891, n4826);
nand_4 g04164(new_n4541, n12925, n4828);
xnor_3 g04165(new_n4542, new_n4541, new_n4540);
xnor_3 g04166(new_n4543, new_n4542, new_n4539);
xnor_3 g04167(new_n4544, new_n4543, new_n4538);
xnor_3 g04168(new_n4545, new_n4544, new_n4533);
nor_4  g04169(new_n4546, new_n4331, new_n4326_1);
nor_4  g04170(new_n4547, new_n4342, new_n4332);
nor_4  g04171(new_n4548, new_n4547, new_n4546);
xnor_3 g04172(new_n4549, new_n4548, new_n4545);
xnor_3 g04173(new_n4550, new_n4549, new_n4532);
nor_4  g04174(new_n4551, new_n4378_1, new_n4347);
not_3  g04175(new_n4552, new_n4551);
nand_4 g04176(new_n4553_1, new_n4410, new_n4380);
nand_4 g04177(new_n4554, new_n4553_1, new_n4552);
xnor_3 g04178(new_n4555, new_n4554, new_n4550);
xnor_3 g04179(new_n4556, new_n4555, new_n4531);
not_3  g04180(new_n4557, new_n4556);
xnor_3 g04181(new_n4558, new_n4557, new_n4497);
nand_4 g04182(new_n4559, new_n4411, new_n4310);
not_3  g04183(new_n4560, new_n4412);
not_3  g04184(new_n4561, new_n4433);
nand_4 g04185(new_n4562, new_n4561, new_n4560);
nand_4 g04186(new_n4563, new_n4562, new_n4559);
xnor_3 g04187(new_n4564, new_n4563, new_n4558);
xor_3  g04188(n992, new_n4564, new_n4468);
nand_4 g04189(new_n4566, n7265, n6687);
not_3  g04190(new_n4567, new_n4566);
nand_4 g04191(new_n4568, n8336, n7946);
not_3  g04192(new_n4569, new_n4568);
nand_4 g04193(new_n4570, n11222, n9763);
nand_4 g04194(new_n4571, n12069, n2558);
xor_3  g04195(new_n4572, new_n4571, new_n4570);
xor_3  g04196(new_n4573, new_n4572, new_n4569);
xor_3  g04197(n1020, new_n4573, new_n4567);
not_3  g04198(new_n4575, new_n2193);
xnor_3 g04199(n1136, new_n4575, new_n2191);
and_4  g04200(new_n4577, new_n4437, new_n4436_1);
xor_3  g04201(n1138, new_n4577, new_n4465);
nand_4 g04202(new_n4579, n12591, n11757);
nand_4 g04203(new_n4580, n5240, n3932);
nand_4 g04204(new_n4581, n11821, n1798);
xnor_3 g04205(new_n4582, new_n4581, new_n4580);
nor_4  g04206(new_n4583, new_n4582, new_n4579);
not_3  g04207(new_n4584, new_n4579);
not_3  g04208(new_n4585, new_n4582);
nor_4  g04209(new_n4586, new_n4585, new_n4584);
nor_4  g04210(new_n4587, new_n4586, new_n4583);
nand_4 g04211(new_n4588, n5240, n1798);
not_3  g04212(new_n4589, new_n4588);
nand_4 g04213(new_n4590, n12591, n3172);
not_3  g04214(new_n4591, new_n4590);
nor_4  g04215(new_n4592, new_n4591, new_n4589);
nor_4  g04216(new_n4593, new_n4590, new_n4588);
nand_4 g04217(new_n4594, n11757, n3932);
not_3  g04218(new_n4595, new_n4594);
nor_4  g04219(new_n4596, new_n4595, new_n4593);
nor_4  g04220(new_n4597, new_n4596, new_n4592);
xnor_3 g04221(new_n4598, new_n4597, new_n4587);
nand_4 g04222(new_n4599, n7456, n1333);
not_3  g04223(new_n4600, new_n4599);
nand_4 g04224(new_n4601, n11757, n1798);
not_3  g04225(new_n4602, new_n4601);
nand_4 g04226(new_n4603, n12591, n1333);
not_3  g04227(new_n4604, new_n4603);
nor_4  g04228(new_n4605, new_n4604, new_n4602);
nor_4  g04229(new_n4606, new_n4603, new_n4601);
nand_4 g04230(new_n4607, n3932, n3172);
not_3  g04231(new_n4608, new_n4607);
nor_4  g04232(new_n4609, new_n4608, new_n4606);
nor_4  g04233(new_n4610, new_n4609, new_n4605);
nand_4 g04234(new_n4611, new_n4610, new_n4600);
xnor_3 g04235(new_n4612, new_n4610, new_n4599);
nor_4  g04236(new_n4613, new_n4593, new_n4592);
xnor_3 g04237(new_n4614, new_n4613, new_n4594);
nand_4 g04238(new_n4615, new_n4614, new_n4612);
nand_4 g04239(new_n4616, new_n4615, new_n4611);
nand_4 g04240(new_n4617, n11662, n1333);
nand_4 g04241(new_n4618, n7456, n3172);
xor_3  g04242(new_n4619, new_n4618, new_n4617);
xnor_3 g04243(new_n4620, new_n4619, new_n4616);
xnor_3 g04244(new_n4621, new_n4620, new_n4598);
nand_4 g04245(new_n4622, n11662, n7862);
not_3  g04246(new_n4623, new_n4622);
xnor_3 g04247(new_n4624, new_n4614, new_n4612);
not_3  g04248(new_n4625, new_n4624);
nor_4  g04249(new_n4626, new_n4625, new_n4623);
not_3  g04250(new_n4627, new_n4626);
nor_4  g04251(new_n4628, new_n4624, new_n4622);
nor_4  g04252(new_n4629, new_n4628, new_n4626);
nand_4 g04253(new_n4630, n7862, n7456);
nand_4 g04254(new_n4631, n3172, n1798);
not_3  g04255(new_n4632, new_n4631);
nand_4 g04256(new_n4633, n12591, n7862);
not_3  g04257(new_n4634_1, new_n4633);
nand_4 g04258(new_n4635, new_n4634_1, new_n4632);
nand_4 g04259(new_n4636, new_n4633, new_n4631);
nand_4 g04260(new_n4637, n3932, n1333);
not_3  g04261(new_n4638, new_n4637);
nand_4 g04262(new_n4639, new_n4638, new_n4636);
nand_4 g04263(new_n4640, new_n4639, new_n4635);
not_3  g04264(new_n4641, new_n4640);
nor_4  g04265(new_n4642, new_n4641, new_n4630);
xnor_3 g04266(new_n4643, new_n4641, new_n4630);
nor_4  g04267(new_n4644, new_n4606, new_n4605);
xnor_3 g04268(new_n4645, new_n4644, new_n4608);
nor_4  g04269(new_n4646, new_n4645, new_n4643);
nor_4  g04270(new_n4647, new_n4646, new_n4642);
nand_4 g04271(new_n4648, new_n4647, new_n4629);
nand_4 g04272(new_n4649, new_n4648, new_n4627);
nor_4  g04273(new_n4650, new_n4649, new_n4621);
not_3  g04274(new_n4651, new_n4650);
not_3  g04275(new_n4652, new_n4587);
not_3  g04276(new_n4653, new_n4597);
nor_4  g04277(new_n4654, new_n4653, new_n4652);
nor_4  g04278(new_n4655, new_n4654, new_n4583);
not_3  g04279(new_n4656, new_n4655);
nand_4 g04280(new_n4657, n10327, n1333);
nand_4 g04281(new_n4658, n11662, n3172);
nand_4 g04282(new_n4659, n9583, n7862);
not_3  g04283(new_n4660, new_n4659);
xor_3  g04284(new_n4661, new_n4660, new_n4658);
xnor_3 g04285(new_n4662, new_n4661, new_n4657);
xnor_3 g04286(new_n4663, new_n4662, new_n4656);
nor_4  g04287(new_n4664, new_n4581, new_n4580);
nand_4 g04288(new_n4665, n11757, n7456);
not_3  g04289(new_n4666, new_n4665);
xor_3  g04290(new_n4667, new_n4666, new_n4664);
not_3  g04291(new_n4668, new_n4667);
nand_4 g04292(new_n4669, n11821, n3932);
nand_4 g04293(new_n4670, n12591, n5240);
nand_4 g04294(new_n4671, n9080, n1798);
not_3  g04295(new_n4672, new_n4671);
xor_3  g04296(new_n4673, new_n4672, new_n4670);
xnor_3 g04297(new_n4674, new_n4673, new_n4669);
not_3  g04298(new_n4675, new_n4674);
xor_3  g04299(new_n4676, new_n4675, new_n4668);
xnor_3 g04300(new_n4677, new_n4676, new_n4663);
not_3  g04301(new_n4678, new_n4677);
nand_4 g04302(new_n4679, new_n4619, new_n4616);
nor_4  g04303(new_n4680, new_n4618, new_n4617);
nor_4  g04304(new_n4681, new_n4620, new_n4598);
xnor_3 g04305(new_n4682, new_n4681, new_n4680);
nand_4 g04306(new_n4683, new_n4682, new_n4679);
xnor_3 g04307(new_n4684, new_n4683, new_n4678);
xnor_3 g04308(new_n4685, new_n4684, new_n4651);
nand_4 g04309(new_n4686_1, n10327, n7862);
xnor_3 g04310(new_n4687, new_n4649, new_n4621);
nor_4  g04311(new_n4688, new_n4687, new_n4686_1);
not_3  g04312(new_n4689_1, new_n4688);
and_4  g04313(new_n4690, new_n4636, new_n4635);
nand_4 g04314(new_n4691, n1798, n1333);
nand_4 g04315(new_n4692, n7862, n3932);
nor_4  g04316(new_n4693, new_n4692, new_n4691);
not_3  g04317(new_n4694, new_n4693);
nor_4  g04318(new_n4695, new_n4694, new_n4690);
xor_3  g04319(new_n4696, new_n4645, new_n4643);
nand_4 g04320(new_n4697, new_n4696, new_n4695);
not_3  g04321(new_n4698, new_n4648);
nor_4  g04322(new_n4699, new_n4647, new_n4629);
nor_4  g04323(new_n4700, new_n4699, new_n4698);
nor_4  g04324(new_n4701, new_n4700, new_n4697);
not_3  g04325(new_n4702, new_n4686_1);
not_3  g04326(new_n4703, new_n4687);
nor_4  g04327(new_n4704, new_n4703, new_n4702);
nor_4  g04328(new_n4705, new_n4704, new_n4688);
nand_4 g04329(new_n4706, new_n4705, new_n4701);
nand_4 g04330(new_n4707, new_n4706, new_n4689_1);
xnor_3 g04331(new_n4708, new_n4707, new_n4685);
nand_4 g04332(new_n4709, n11311, n3022);
not_3  g04333(new_n4710, new_n4709);
nand_4 g04334(new_n4711, n9640, n4187);
nand_4 g04335(new_n4712, n6703, n4203);
not_3  g04336(new_n4713, new_n4712);
xor_3  g04337(new_n4714, new_n4713, new_n4711);
xnor_3 g04338(new_n4715, new_n4714, new_n4710);
not_3  g04339(new_n4716, new_n4715);
nand_4 g04340(new_n4717, n6703, n4187);
not_3  g04341(new_n4718, new_n4717);
nand_4 g04342(new_n4719, n3022, n2464);
not_3  g04343(new_n4720, new_n4719);
nor_4  g04344(new_n4721, new_n4720, new_n4718);
nor_4  g04345(new_n4722_1, new_n4719, new_n4717);
nand_4 g04346(new_n4723, n11311, n9640);
not_3  g04347(new_n4724, new_n4723);
nor_4  g04348(new_n4725, new_n4724, new_n4722_1);
nor_4  g04349(new_n4726, new_n4725, new_n4721);
xor_3  g04350(new_n4727, new_n4726, new_n4716);
nand_4 g04351(new_n4728, n10451, n9400);
nand_4 g04352(new_n4729, n11023, n2464);
xor_3  g04353(new_n4730, new_n4729, new_n4728);
xnor_3 g04354(new_n4731, new_n4730, new_n4727);
nand_4 g04355(new_n4732, n11023, n9400);
not_3  g04356(new_n4733_1, new_n4732);
nand_4 g04357(new_n4734, n11311, n6703);
not_3  g04358(new_n4735, new_n4734);
nand_4 g04359(new_n4736, n9400, n3022);
not_3  g04360(new_n4737, new_n4736);
nor_4  g04361(new_n4738, new_n4737, new_n4735);
nor_4  g04362(new_n4739, new_n4736, new_n4734);
nand_4 g04363(new_n4740, n9640, n2464);
not_3  g04364(new_n4741, new_n4740);
nor_4  g04365(new_n4742, new_n4741, new_n4739);
nor_4  g04366(new_n4743, new_n4742, new_n4738);
and_4  g04367(new_n4744, new_n4743, new_n4733_1);
xnor_3 g04368(new_n4745, new_n4743, new_n4733_1);
nor_4  g04369(new_n4746, new_n4722_1, new_n4721);
xnor_3 g04370(new_n4747, new_n4746, new_n4724);
nor_4  g04371(new_n4748, new_n4747, new_n4745);
nor_4  g04372(new_n4749, new_n4748, new_n4744);
xnor_3 g04373(new_n4750, new_n4749, new_n4731);
nand_4 g04374(new_n4751, n10451, n6877);
not_3  g04375(new_n4752, new_n4751);
xnor_3 g04376(new_n4753, new_n4747, new_n4745);
not_3  g04377(new_n4754, new_n4753);
nand_4 g04378(new_n4755, new_n4754, new_n4752);
nand_4 g04379(new_n4756, n11023, n6877);
not_3  g04380(new_n4757_1, new_n4756);
nand_4 g04381(new_n4758, n6703, n2464);
not_3  g04382(new_n4759, new_n4758);
nand_4 g04383(new_n4760, n6877, n3022);
not_3  g04384(new_n4761, new_n4760);
nor_4  g04385(new_n4762, new_n4761, new_n4759);
nor_4  g04386(new_n4763, new_n4760, new_n4758);
nand_4 g04387(new_n4764, n9640, n9400);
not_3  g04388(new_n4765, new_n4764);
nor_4  g04389(new_n4766, new_n4765, new_n4763);
nor_4  g04390(new_n4767, new_n4766, new_n4762);
and_4  g04391(new_n4768, new_n4767, new_n4757_1);
not_3  g04392(new_n4769, new_n4768);
xor_3  g04393(new_n4770, new_n4767, new_n4756);
not_3  g04394(new_n4771, new_n4770);
nor_4  g04395(new_n4772, new_n4739, new_n4738);
xor_3  g04396(new_n4773, new_n4772, new_n4740);
not_3  g04397(new_n4774, new_n4773);
nand_4 g04398(new_n4775, new_n4774, new_n4771);
nand_4 g04399(new_n4776, new_n4775, new_n4769);
xor_3  g04400(new_n4777, new_n4754, new_n4752);
nand_4 g04401(new_n4778, new_n4777, new_n4776);
nand_4 g04402(new_n4779, new_n4778, new_n4755);
nand_4 g04403(new_n4780, new_n4779, new_n4750);
not_3  g04404(new_n4781, new_n4714);
nand_4 g04405(new_n4782, new_n4781, new_n4710);
nand_4 g04406(new_n4783, new_n4726, new_n4715);
nand_4 g04407(new_n4784, new_n4783, new_n4782);
nand_4 g04408(new_n4785, n10278, n9400);
not_3  g04409(new_n4786, new_n4785);
nand_4 g04410(new_n4787, n10451, n2464);
not_3  g04411(new_n4788, new_n4787);
nand_4 g04412(new_n4789, n11423, n6877);
not_3  g04413(new_n4790, new_n4789);
nand_4 g04414(new_n4791, new_n4790, new_n4788);
nand_4 g04415(new_n4792, new_n4789, new_n4787);
nand_4 g04416(new_n4793, new_n4792, new_n4791);
xor_3  g04417(new_n4794, new_n4793, new_n4786);
xnor_3 g04418(new_n4795, new_n4794, new_n4784);
nor_4  g04419(new_n4796, new_n4712, new_n4711);
nand_4 g04420(new_n4797, n11311, n11023);
not_3  g04421(new_n4798, new_n4797);
xor_3  g04422(new_n4799, new_n4798, new_n4796);
nand_4 g04423(new_n4800, n9640, n4203);
not_3  g04424(new_n4801, new_n4800);
nand_4 g04425(new_n4802, n4187, n3022);
not_3  g04426(new_n4803, new_n4802);
nand_4 g04427(new_n4804, n12753, n6703);
not_3  g04428(new_n4805_1, new_n4804);
nor_4  g04429(new_n4806, new_n4805_1, new_n4803);
nor_4  g04430(new_n4807, new_n4804, new_n4802);
nor_4  g04431(new_n4808, new_n4807, new_n4806);
xor_3  g04432(new_n4809, new_n4808, new_n4801);
not_3  g04433(new_n4810, new_n4809);
xnor_3 g04434(new_n4811, new_n4810, new_n4799);
xnor_3 g04435(new_n4812, new_n4811, new_n4795);
not_3  g04436(new_n4813, new_n4730);
nor_4  g04437(new_n4814, new_n4813, new_n4727);
not_3  g04438(new_n4815, new_n4814);
nor_4  g04439(new_n4816, new_n4729, new_n4728);
not_3  g04440(new_n4817_1, new_n4816);
not_3  g04441(new_n4818, new_n4749);
nand_4 g04442(new_n4819, new_n4818, new_n4731);
xnor_3 g04443(new_n4820, new_n4819, new_n4817_1);
nand_4 g04444(new_n4821, new_n4820, new_n4815);
not_3  g04445(new_n4822, new_n4821);
xnor_3 g04446(new_n4823, new_n4822, new_n4812);
xnor_3 g04447(new_n4824, new_n4823, new_n4780);
nand_4 g04448(new_n4825, n10278, n6877);
xnor_3 g04449(new_n4826_1, new_n4779, new_n4750);
nor_4  g04450(new_n4827, new_n4826_1, new_n4825);
xnor_3 g04451(new_n4828_1, new_n4773, new_n4770);
not_3  g04452(new_n4829, new_n4762);
nand_4 g04453(new_n4830, n6877, n6703);
not_3  g04454(new_n4831, new_n4830);
nor_4  g04455(new_n4832, new_n4831, new_n4764);
nor_4  g04456(new_n4833, new_n4832, new_n4829);
nor_4  g04457(new_n4834, new_n4833, new_n4763);
nor_4  g04458(new_n4835, new_n4834, new_n4764);
not_3  g04459(new_n4836, new_n4835);
nor_4  g04460(new_n4837, new_n4836, new_n4828_1);
not_3  g04461(new_n4838, new_n4837);
xnor_3 g04462(new_n4839, new_n4777, new_n4776);
nor_4  g04463(new_n4840, new_n4839, new_n4838);
not_3  g04464(new_n4841, new_n4840);
xnor_3 g04465(new_n4842, new_n4826_1, new_n4825);
nor_4  g04466(new_n4843, new_n4842, new_n4841);
nor_4  g04467(new_n4844, new_n4843, new_n4827);
xnor_3 g04468(new_n4845, new_n4844, new_n4824);
nand_4 g04469(new_n4846, n12826, n4805);
nand_4 g04470(new_n4847, n8665, n137);
nand_4 g04471(new_n4848, n6294, n1067);
nand_4 g04472(new_n4849, n6797, n5645);
xnor_3 g04473(new_n4850, new_n4849, new_n4848);
nor_4  g04474(new_n4851, new_n4850, new_n4847);
not_3  g04475(new_n4852, new_n4847);
not_3  g04476(new_n4853, new_n4850);
nor_4  g04477(new_n4854, new_n4853, new_n4852);
nor_4  g04478(new_n4855, new_n4854, new_n4851);
nand_4 g04479(new_n4856, n6294, n5645);
nand_4 g04480(new_n4857, n8665, n5283);
and_4  g04481(new_n4858, new_n4857, new_n4856);
nand_4 g04482(new_n4859, n1067, n137);
not_3  g04483(new_n4860, new_n4859);
xnor_3 g04484(new_n4861, new_n4857, new_n4856);
nor_4  g04485(new_n4862, new_n4861, new_n4860);
nor_4  g04486(new_n4863, new_n4862, new_n4858);
xnor_3 g04487(new_n4864, new_n4863, new_n4855);
nand_4 g04488(new_n4865, n11922, n11478);
not_3  g04489(new_n4866, new_n4865);
nand_4 g04490(new_n4867, n11478, n8665);
not_3  g04491(new_n4868, new_n4867);
nand_4 g04492(new_n4869, n5283, n1067);
not_3  g04493(new_n4870, new_n4869);
nor_4  g04494(new_n4871, new_n4870, new_n4868);
nor_4  g04495(new_n4872, new_n4869, new_n4867);
nand_4 g04496(new_n4873, n5645, n137);
not_3  g04497(new_n4874, new_n4873);
nor_4  g04498(new_n4875, new_n4874, new_n4872);
nor_4  g04499(new_n4876, new_n4875, new_n4871);
nand_4 g04500(new_n4877, new_n4876, new_n4866);
xnor_3 g04501(new_n4878, new_n4861, new_n4859);
not_3  g04502(new_n4879, new_n4878);
xnor_3 g04503(new_n4880, new_n4876, new_n4865);
nand_4 g04504(new_n4881, new_n4880, new_n4879);
nand_4 g04505(new_n4882, new_n4881, new_n4877);
nand_4 g04506(new_n4883, n11478, n2551);
nand_4 g04507(new_n4884, n11922, n5283);
xor_3  g04508(new_n4885, new_n4884, new_n4883);
xnor_3 g04509(new_n4886, new_n4885, new_n4882);
xnor_3 g04510(new_n4887, new_n4886, new_n4864);
nand_4 g04511(new_n4888, n4805, n2551);
not_3  g04512(new_n4889, new_n4888);
nand_4 g04513(new_n4890, n11922, n4805);
not_3  g04514(new_n4891, new_n4890);
nand_4 g04515(new_n4892, n5645, n5283);
not_3  g04516(new_n4893, new_n4892);
nand_4 g04517(new_n4894, n8665, n4805);
not_3  g04518(new_n4895, new_n4894);
nand_4 g04519(new_n4896, new_n4895, new_n4893);
nand_4 g04520(new_n4897, n11478, n1067);
not_3  g04521(new_n4898, new_n4897);
nand_4 g04522(new_n4899, new_n4894, new_n4892);
nand_4 g04523(new_n4900, new_n4899, new_n4898);
nand_4 g04524(new_n4901, new_n4900, new_n4896);
nand_4 g04525(new_n4902, new_n4901, new_n4891);
not_3  g04526(new_n4903_1, new_n4902);
nor_4  g04527(new_n4904, new_n4901, new_n4891);
nor_4  g04528(new_n4905, new_n4904, new_n4903_1);
xnor_3 g04529(new_n4906, new_n4869, new_n4867);
xnor_3 g04530(new_n4907, new_n4906, new_n4873);
not_3  g04531(new_n4908, new_n4907);
nand_4 g04532(new_n4909, new_n4908, new_n4905);
nand_4 g04533(new_n4910, new_n4909, new_n4902);
nor_4  g04534(new_n4911, new_n4910, new_n4889);
xnor_3 g04535(new_n4912, new_n4880, new_n4878);
xnor_3 g04536(new_n4913, new_n4910, new_n4889);
nor_4  g04537(new_n4914, new_n4913, new_n4912);
nor_4  g04538(new_n4915, new_n4914, new_n4911);
not_3  g04539(new_n4916, new_n4915);
xnor_3 g04540(new_n4917, new_n4916, new_n4887);
nor_4  g04541(new_n4918, new_n4917, new_n4846);
nand_4 g04542(new_n4919, new_n4899, new_n4896);
nand_4 g04543(new_n4920, n4805, n1067);
nand_4 g04544(new_n4921_1, n11478, n5645);
nor_4  g04545(new_n4922, new_n4921_1, new_n4920);
nand_4 g04546(new_n4923, new_n4922, new_n4919);
xnor_3 g04547(new_n4924, new_n4908, new_n4905);
nor_4  g04548(new_n4925, new_n4924, new_n4923);
not_3  g04549(new_n4926, new_n4925);
not_3  g04550(new_n4927, new_n4912);
xnor_3 g04551(new_n4928_1, new_n4913, new_n4927);
nor_4  g04552(new_n4929, new_n4928_1, new_n4926);
not_3  g04553(new_n4930, new_n4929);
xnor_3 g04554(new_n4931, new_n4917, new_n4846);
nor_4  g04555(new_n4932, new_n4931, new_n4930);
nor_4  g04556(new_n4933, new_n4932, new_n4918);
nor_4  g04557(new_n4934, new_n4916, new_n4887);
not_3  g04558(new_n4935, new_n4851);
nand_4 g04559(new_n4936, new_n4863, new_n4855);
nand_4 g04560(new_n4937, new_n4936, new_n4935);
nand_4 g04561(new_n4938_1, n12826, n11478);
not_3  g04562(new_n4939, new_n4938_1);
nand_4 g04563(new_n4940, n5283, n2551);
nand_4 g04564(new_n4941, n4805, n4094);
nand_4 g04565(new_n4942, new_n4941, new_n4940);
not_3  g04566(new_n4943, new_n4940);
not_3  g04567(new_n4944, new_n4941);
nand_4 g04568(new_n4945, new_n4944, new_n4943);
nand_4 g04569(new_n4946, new_n4945, new_n4942);
xor_3  g04570(new_n4947, new_n4946, new_n4939);
xnor_3 g04571(new_n4948, new_n4947, new_n4937);
nor_4  g04572(new_n4949, new_n4849, new_n4848);
nand_4 g04573(new_n4950, n11922, n137);
not_3  g04574(new_n4951, new_n4950);
xor_3  g04575(new_n4952, new_n4951, new_n4949);
not_3  g04576(new_n4953, new_n4952);
nand_4 g04577(new_n4954, n6797, n1067);
not_3  g04578(new_n4955, new_n4954);
nand_4 g04579(new_n4956, n8665, n6294);
nand_4 g04580(new_n4957, n5645, n3146);
not_3  g04581(new_n4958, new_n4957);
xor_3  g04582(new_n4959, new_n4958, new_n4956);
xnor_3 g04583(new_n4960, new_n4959, new_n4955);
xnor_3 g04584(new_n4961, new_n4960, new_n4953);
xnor_3 g04585(new_n4962, new_n4961, new_n4948);
nand_4 g04586(new_n4963, new_n4885, new_n4882);
nor_4  g04587(new_n4964, new_n4884, new_n4883);
nor_4  g04588(new_n4965, new_n4886, new_n4864);
xnor_3 g04589(new_n4966, new_n4965, new_n4964);
nand_4 g04590(new_n4967, new_n4966, new_n4963);
xnor_3 g04591(new_n4968, new_n4967, new_n4962);
xnor_3 g04592(new_n4969, new_n4968, new_n4934);
xnor_3 g04593(new_n4970_1, new_n4969, new_n4933);
nand_4 g04594(new_n4971_1, n3992, n2749);
not_3  g04595(new_n4972, new_n4971_1);
nand_4 g04596(new_n4973, n11876, n6358);
not_3  g04597(new_n4974, new_n4973);
nand_4 g04598(new_n4975, n3992, n3754);
not_3  g04599(new_n4976, new_n4975);
nor_4  g04600(new_n4977, new_n4976, new_n4974);
nor_4  g04601(new_n4978, new_n4975, new_n4973);
nand_4 g04602(new_n4979, n10898, n8384);
not_3  g04603(new_n4980, new_n4979);
nor_4  g04604(new_n4981, new_n4980, new_n4978);
nor_4  g04605(new_n4982, new_n4981, new_n4977);
nand_4 g04606(new_n4983, new_n4982, new_n4972);
xnor_3 g04607(new_n4984, new_n4982, new_n4971_1);
nand_4 g04608(new_n4985, n10898, n6358);
not_3  g04609(new_n4986, new_n4985);
nand_4 g04610(new_n4987, n8384, n3754);
nand_4 g04611(new_n4988, n11876, n5198);
xnor_3 g04612(new_n4989, new_n4988, new_n4987);
xnor_3 g04613(new_n4990, new_n4989, new_n4986);
nand_4 g04614(new_n4991, new_n4990, new_n4984);
nand_4 g04615(new_n4992, new_n4991, new_n4983);
nand_4 g04616(new_n4993, n8384, n2749);
nand_4 g04617(new_n4994, n3992, n159);
xor_3  g04618(new_n4995, new_n4994, new_n4993);
xnor_3 g04619(new_n4996, new_n4995, new_n4992);
nand_4 g04620(new_n4997, n6358, n3754);
not_3  g04621(new_n4998, new_n4997);
nand_4 g04622(new_n4999, n10898, n5198);
nand_4 g04623(new_n5000, n11876, n1471);
xnor_3 g04624(new_n5001, new_n5000, new_n4999);
not_3  g04625(new_n5002, new_n5001);
nor_4  g04626(new_n5003, new_n5002, new_n4998);
nor_4  g04627(new_n5004, new_n5001, new_n4997);
nor_4  g04628(new_n5005, new_n5004, new_n5003);
not_3  g04629(new_n5006, new_n5005);
and_4  g04630(new_n5007, new_n4988, new_n4987);
nor_4  g04631(new_n5008, new_n4989, new_n4986);
nor_4  g04632(new_n5009, new_n5008, new_n5007);
nor_4  g04633(new_n5010, new_n5009, new_n5006);
not_3  g04634(new_n5011, new_n5009);
nor_4  g04635(new_n5012, new_n5011, new_n5005);
nor_4  g04636(new_n5013, new_n5012, new_n5010);
xnor_3 g04637(new_n5014, new_n5013, new_n4996);
nand_4 g04638(new_n5015, n7236, n159);
not_3  g04639(new_n5016, new_n5015);
nand_4 g04640(new_n5017, n7236, n2749);
not_3  g04641(new_n5018, new_n5017);
nand_4 g04642(new_n5019, n11876, n8384);
not_3  g04643(new_n5020, new_n5019);
nand_4 g04644(new_n5021, n7236, n3754);
not_3  g04645(new_n5022, new_n5021);
nor_4  g04646(new_n5023, new_n5022, new_n5020);
nand_4 g04647(new_n5024, n11876, n7236);
nor_4  g04648(new_n5025, new_n5024, new_n4987);
nand_4 g04649(new_n5026, n10898, n3992);
not_3  g04650(new_n5027, new_n5026);
nor_4  g04651(new_n5028, new_n5027, new_n5025);
nor_4  g04652(new_n5029, new_n5028, new_n5023);
nand_4 g04653(new_n5030_1, new_n5029, new_n5018);
not_3  g04654(new_n5031, new_n5030_1);
nor_4  g04655(new_n5032, new_n5029, new_n5018);
nor_4  g04656(new_n5033, new_n5032, new_n5031);
xnor_3 g04657(new_n5034_1, new_n4975, new_n4973);
xnor_3 g04658(new_n5035, new_n5034_1, new_n4979);
not_3  g04659(new_n5036, new_n5035);
nand_4 g04660(new_n5037, new_n5036, new_n5033);
nand_4 g04661(new_n5038, new_n5037, new_n5030_1);
nor_4  g04662(new_n5039, new_n5038, new_n5016);
not_3  g04663(new_n5040, new_n5039);
xnor_3 g04664(new_n5041, new_n4990, new_n4984);
not_3  g04665(new_n5042, new_n5038);
nor_4  g04666(new_n5043, new_n5042, new_n5015);
nor_4  g04667(new_n5044, new_n5043, new_n5039);
nand_4 g04668(new_n5045, new_n5044, new_n5041);
nand_4 g04669(new_n5046, new_n5045, new_n5040);
nor_4  g04670(new_n5047, new_n5046, new_n5014);
not_3  g04671(new_n5048, new_n5047);
nor_4  g04672(new_n5049, new_n5000, new_n4999);
not_3  g04673(new_n5050, new_n5049);
nand_4 g04674(new_n5051, n6358, n2749);
xor_3  g04675(new_n5052, new_n5051, new_n5050);
nand_4 g04676(new_n5053, n10898, n1471);
nand_4 g04677(new_n5054, n5198, n3754);
nand_4 g04678(new_n5055, n11876, n7646);
not_3  g04679(new_n5056, new_n5055);
xor_3  g04680(new_n5057, new_n5056, new_n5054);
xnor_3 g04681(new_n5058, new_n5057, new_n5053);
xnor_3 g04682(new_n5059, new_n5058, new_n5052);
nor_4  g04683(new_n5060, new_n5010, new_n5003);
nand_4 g04684(new_n5061, n3992, n1510);
nand_4 g04685(new_n5062, n8384, n159);
nand_4 g04686(new_n5063, n12247, n7236);
not_3  g04687(new_n5064, new_n5063);
xor_3  g04688(new_n5065, new_n5064, new_n5062);
xnor_3 g04689(new_n5066, new_n5065, new_n5061);
xnor_3 g04690(new_n5067, new_n5066, new_n5060);
xnor_3 g04691(new_n5068, new_n5067, new_n5059);
nand_4 g04692(new_n5069_1, new_n4995, new_n4992);
nor_4  g04693(new_n5070, new_n4994, new_n4993);
nor_4  g04694(new_n5071, new_n5013, new_n4996);
xnor_3 g04695(new_n5072, new_n5071, new_n5070);
nand_4 g04696(new_n5073, new_n5072, new_n5069_1);
xnor_3 g04697(new_n5074, new_n5073, new_n5068);
xnor_3 g04698(new_n5075, new_n5074, new_n5048);
nand_4 g04699(new_n5076, n7236, n1510);
not_3  g04700(new_n5077, new_n5076);
not_3  g04701(new_n5078, new_n5046);
xnor_3 g04702(new_n5079, new_n5078, new_n5014);
nand_4 g04703(new_n5080, new_n5079, new_n5077);
nor_4  g04704(new_n5081, new_n5025, new_n5023);
nand_4 g04705(new_n5082, n11876, n3992);
nand_4 g04706(new_n5083, n10898, n7236);
nor_4  g04707(new_n5084, new_n5083, new_n5082);
not_3  g04708(new_n5085, new_n5084);
nor_4  g04709(new_n5086, new_n5085, new_n5081);
not_3  g04710(new_n5087, new_n5086);
xnor_3 g04711(new_n5088, new_n5036, new_n5033);
nor_4  g04712(new_n5089, new_n5088, new_n5087);
xnor_3 g04713(new_n5090, new_n5044, new_n5041);
nand_4 g04714(new_n5091, new_n5090, new_n5089);
not_3  g04715(new_n5092, new_n5091);
xnor_3 g04716(new_n5093, new_n5079, new_n5076);
nand_4 g04717(new_n5094_1, new_n5093, new_n5092);
nand_4 g04718(new_n5095, new_n5094_1, new_n5080);
xnor_3 g04719(new_n5096, new_n5095, new_n5075);
xnor_3 g04720(new_n5097, new_n5096, new_n4970_1);
not_3  g04721(new_n5098, new_n4846);
xnor_3 g04722(new_n5099, new_n4917, new_n5098);
nor_4  g04723(new_n5100, new_n5099, new_n4929);
nor_4  g04724(new_n5101, new_n5100, new_n4932);
not_3  g04725(new_n5102, new_n5101);
xnor_3 g04726(new_n5103, new_n5093, new_n5092);
nand_4 g04727(new_n5104, new_n5103, new_n5102);
xnor_3 g04728(new_n5105_1, new_n5103, new_n5101);
nor_4  g04729(new_n5106, new_n5090, new_n5089);
nor_4  g04730(new_n5107, new_n5106, new_n5092);
not_3  g04731(new_n5108, new_n4923);
not_3  g04732(new_n5109, new_n4924);
nor_4  g04733(new_n5110, new_n5109, new_n5108);
nor_4  g04734(new_n5111, new_n5110, new_n4925);
not_3  g04735(new_n5112, new_n5088);
nor_4  g04736(new_n5113, new_n5112, new_n5086);
nor_4  g04737(new_n5114, new_n5113, new_n5089);
nor_4  g04738(new_n5115, new_n5114, new_n5111);
not_3  g04739(new_n5116, new_n5115);
xnor_3 g04740(new_n5117, new_n5083, new_n5082);
xnor_3 g04741(new_n5118, new_n4921_1, new_n4920);
nand_4 g04742(new_n5119, new_n5118, new_n5117);
not_3  g04743(new_n5120, new_n5119);
nand_4 g04744(new_n5121, n5645, n4805);
nor_4  g04745(new_n5122, new_n5121, new_n5024);
xnor_3 g04746(new_n5123, new_n5118, new_n5117);
nor_4  g04747(new_n5124, new_n5123, new_n5122);
nor_4  g04748(new_n5125, new_n5124, new_n5120);
not_3  g04749(new_n5126, new_n5121);
nor_4  g04750(new_n5127, new_n5126, new_n4897);
not_3  g04751(new_n5128, new_n5127);
nand_4 g04752(new_n5129, new_n5128, new_n4919);
nand_4 g04753(new_n5130, new_n5127, new_n4899);
nand_4 g04754(new_n5131, new_n5130, new_n5129);
not_3  g04755(new_n5132_1, new_n5131);
nor_4  g04756(new_n5133, new_n5132_1, new_n5125);
xnor_3 g04757(new_n5134, new_n5132_1, new_n5125);
not_3  g04758(new_n5135, new_n5024);
nor_4  g04759(new_n5136, new_n5026, new_n5135);
nor_4  g04760(new_n5137, new_n5136, new_n5081);
not_3  g04761(new_n5138, new_n5136);
nor_4  g04762(new_n5139, new_n5138, new_n5023);
nor_4  g04763(new_n5140, new_n5139, new_n5137);
nor_4  g04764(new_n5141, new_n5140, new_n5134);
nor_4  g04765(new_n5142, new_n5141, new_n5133);
xnor_3 g04766(new_n5143, new_n5114, new_n5111);
nor_4  g04767(new_n5144, new_n5143, new_n5142);
not_3  g04768(new_n5145, new_n5144);
nand_4 g04769(new_n5146, new_n5145, new_n5116);
not_3  g04770(new_n5147, new_n5146);
nor_4  g04771(new_n5148, new_n5147, new_n5107);
not_3  g04772(new_n5149, new_n5148);
not_3  g04773(new_n5150, new_n4928_1);
xor_3  g04774(new_n5151, new_n5150, new_n4926);
xnor_3 g04775(new_n5152, new_n5146, new_n5107);
nand_4 g04776(new_n5153_1, new_n5152, new_n5151);
nand_4 g04777(new_n5154, new_n5153_1, new_n5149);
nand_4 g04778(new_n5155, new_n5154, new_n5105_1);
nand_4 g04779(new_n5156, new_n5155, new_n5104);
xnor_3 g04780(new_n5157, new_n5156, new_n5097);
nand_4 g04781(new_n5158, new_n5157, new_n4845);
not_3  g04782(new_n5159, new_n4824);
xnor_3 g04783(new_n5160, new_n4844, new_n5159);
not_3  g04784(new_n5161, new_n4918);
nand_4 g04785(new_n5162, new_n5099, new_n4929);
nand_4 g04786(new_n5163, new_n5162, new_n5161);
xnor_3 g04787(new_n5164, new_n4969, new_n5163);
xnor_3 g04788(new_n5165, new_n5096, new_n5164);
xnor_3 g04789(new_n5166, new_n5156, new_n5165);
nand_4 g04790(new_n5167, new_n5166, new_n5160);
nand_4 g04791(new_n5168, new_n5167, new_n5158);
xnor_3 g04792(new_n5169, new_n4842, new_n4840);
xnor_3 g04793(new_n5170, new_n5154, new_n5105_1);
nand_4 g04794(new_n5171, new_n5170, new_n5169);
xnor_3 g04795(new_n5172, new_n4842, new_n4841);
xor_3  g04796(new_n5173, new_n5150, new_n4925);
not_3  g04797(new_n5174, new_n5152);
nor_4  g04798(new_n5175, new_n5174, new_n5173);
nor_4  g04799(new_n5176, new_n5175, new_n5148);
xnor_3 g04800(new_n5177, new_n5176, new_n5105_1);
nand_4 g04801(new_n5178, new_n5177, new_n5172);
not_3  g04802(new_n5179, new_n4839);
nor_4  g04803(new_n5180, new_n5179, new_n4837);
nor_4  g04804(new_n5181, new_n5180, new_n4840);
not_3  g04805(new_n5182, new_n4828_1);
xor_3  g04806(new_n5183, new_n4835, new_n5182);
xnor_3 g04807(new_n5184, new_n5143, new_n5142);
nand_4 g04808(new_n5185, new_n5184, new_n5183);
not_3  g04809(new_n5186, new_n5184);
xnor_3 g04810(new_n5187, new_n5186, new_n5183);
xnor_3 g04811(new_n5188, new_n5140, new_n5134);
not_3  g04812(new_n5189, new_n4834);
not_3  g04813(new_n5190, new_n4832);
nor_4  g04814(new_n5191_1, new_n5190, new_n4762);
nor_4  g04815(new_n5192, new_n5191_1, new_n5189);
nand_4 g04816(new_n5193, new_n5192, new_n5188);
not_3  g04817(new_n5194, new_n5193);
nor_4  g04818(new_n5195, new_n5192, new_n5188);
nor_4  g04819(new_n5196, new_n5195, new_n5194);
not_3  g04820(new_n5197, new_n5123);
xor_3  g04821(new_n5198_1, new_n5197, new_n5122);
nand_4 g04822(new_n5199, n9400, n6703);
nand_4 g04823(new_n5200, n9640, n6877);
xor_3  g04824(new_n5201, new_n5200, new_n5199);
nand_4 g04825(new_n5202, new_n5201, new_n5198_1);
xor_3  g04826(new_n5203, new_n5126, new_n5024);
nor_4  g04827(new_n5204, new_n5203, new_n4830);
not_3  g04828(new_n5205, new_n5202);
nor_4  g04829(new_n5206, new_n5201, new_n5198_1);
nor_4  g04830(new_n5207, new_n5206, new_n5205);
nand_4 g04831(new_n5208, new_n5207, new_n5204);
nand_4 g04832(new_n5209, new_n5208, new_n5202);
nand_4 g04833(new_n5210, new_n5209, new_n5196);
nand_4 g04834(new_n5211, new_n5210, new_n5193);
nand_4 g04835(new_n5212_1, new_n5211, new_n5187);
nand_4 g04836(new_n5213, new_n5212_1, new_n5185);
nor_4  g04837(new_n5214, new_n5213, new_n5181);
xnor_3 g04838(new_n5215, new_n5174, new_n5173);
xnor_3 g04839(new_n5216, new_n5213, new_n5181);
nor_4  g04840(new_n5217, new_n5216, new_n5215);
nor_4  g04841(new_n5218, new_n5217, new_n5214);
nand_4 g04842(new_n5219, new_n5218, new_n5178);
nand_4 g04843(new_n5220, new_n5219, new_n5171);
xnor_3 g04844(new_n5221, new_n5220, new_n5168);
not_3  g04845(new_n5222, new_n5221);
nand_4 g04846(new_n5223, new_n5222, new_n4708);
not_3  g04847(new_n5224, new_n4708);
nand_4 g04848(new_n5225, new_n5221, new_n5224);
xor_3  g04849(new_n5226, new_n4705, new_n4701);
not_3  g04850(new_n5227, new_n5226);
nand_4 g04851(new_n5228, new_n5178, new_n5171);
xnor_3 g04852(new_n5229, new_n5228, new_n5218);
not_3  g04853(new_n5230, new_n5229);
nand_4 g04854(new_n5231, new_n5230, new_n5227);
nand_4 g04855(new_n5232, new_n5229, new_n5226);
not_3  g04856(new_n5233, new_n4697);
xor_3  g04857(new_n5234, new_n4700, new_n5233);
not_3  g04858(new_n5235, new_n5215);
xnor_3 g04859(new_n5236, new_n5216, new_n5235);
nand_4 g04860(new_n5237, new_n5236, new_n5234);
not_3  g04861(new_n5238, new_n5237);
nor_4  g04862(new_n5239, new_n5236, new_n5234);
nor_4  g04863(new_n5240_1, new_n5239, new_n5238);
not_3  g04864(new_n5241, new_n4696);
xor_3  g04865(new_n5242, new_n5241, new_n4695);
not_3  g04866(new_n5243, new_n5242);
xnor_3 g04867(new_n5244, new_n5211, new_n5187);
not_3  g04868(new_n5245, new_n5244);
nor_4  g04869(new_n5246, new_n5245, new_n5243);
not_3  g04870(new_n5247, new_n5246);
xnor_3 g04871(new_n5248, new_n5209, new_n5196);
not_3  g04872(new_n5249, new_n4690);
nand_4 g04873(new_n5250, n7862, n1798);
not_3  g04874(new_n5251, new_n5250);
nor_4  g04875(new_n5252, new_n5251, new_n4637);
not_3  g04876(new_n5253, new_n5252);
nand_4 g04877(new_n5254, new_n5253, new_n5249);
nand_4 g04878(new_n5255, new_n5252, new_n4636);
nand_4 g04879(new_n5256, new_n5255, new_n5254);
nand_4 g04880(new_n5257_1, new_n5256, new_n5248);
not_3  g04881(new_n5258, new_n5257_1);
nor_4  g04882(new_n5259, new_n5256, new_n5248);
nor_4  g04883(new_n5260, new_n5259, new_n5258);
xor_3  g04884(new_n5261, new_n5203, new_n4830);
nand_4 g04885(new_n5262, new_n5261, new_n5251);
not_3  g04886(new_n5263, new_n5262);
xor_3  g04887(new_n5264, new_n4692, new_n4691);
or_4   g04888(new_n5265, new_n5264, new_n5263);
xnor_3 g04889(new_n5266, new_n5207, new_n5204);
xor_3  g04890(new_n5267, new_n5264, new_n5263);
nand_4 g04891(new_n5268, new_n5267, new_n5266);
nand_4 g04892(new_n5269, new_n5268, new_n5265);
nand_4 g04893(new_n5270, new_n5269, new_n5260);
nand_4 g04894(new_n5271, new_n5270, new_n5257_1);
nor_4  g04895(new_n5272, new_n5244, new_n5242);
nor_4  g04896(new_n5273, new_n5272, new_n5246);
nand_4 g04897(new_n5274, new_n5273, new_n5271);
nand_4 g04898(new_n5275, new_n5274, new_n5247);
nand_4 g04899(new_n5276, new_n5275, new_n5240_1);
nand_4 g04900(new_n5277, new_n5276, new_n5237);
nand_4 g04901(new_n5278, new_n5277, new_n5232);
nand_4 g04902(new_n5279, new_n5278, new_n5231);
nand_4 g04903(new_n5280, new_n5279, new_n5225);
nand_4 g04904(new_n5281, new_n5280, new_n5223);
nand_4 g04905(new_n5282, new_n4662, new_n4655);
nand_4 g04906(new_n5283_1, new_n4676, new_n4663);
nand_4 g04907(new_n5284, new_n5283_1, new_n5282);
not_3  g04908(new_n5285, new_n4658);
nor_4  g04909(new_n5286, new_n4660, new_n5285);
not_3  g04910(new_n5287, new_n4657);
nor_4  g04911(new_n5288, new_n4661, new_n5287);
nor_4  g04912(new_n5289, new_n5288, new_n5286);
xor_3  g04913(new_n5290, new_n5289, new_n5284);
xnor_3 g04914(new_n5291, new_n5290, new_n5281);
nor_4  g04915(new_n5292, new_n4823, new_n4780);
nor_4  g04916(new_n5293, new_n4844, new_n4824);
nor_4  g04917(new_n5294, new_n5293, new_n5292);
nand_4 g04918(new_n5295, new_n4968, new_n4934);
not_3  g04919(new_n5296, new_n4969);
nand_4 g04920(new_n5297, new_n5296, new_n5163);
nand_4 g04921(new_n5298, new_n5297, new_n5295);
xnor_3 g04922(new_n5299, new_n5298, new_n5294);
nand_4 g04923(new_n5300, n10327, n3172);
nand_4 g04924(new_n5301, n4203, n3022);
xor_3  g04925(new_n5302, new_n5301, new_n5300);
or_4   g04926(new_n5303, new_n4806, new_n4800);
not_3  g04927(new_n5304, new_n5303);
nor_4  g04928(new_n5305_1, new_n5304, new_n4807);
nand_4 g04929(new_n5306, n10278, n2464);
not_3  g04930(new_n5307, new_n5306);
nand_4 g04931(new_n5308, n11023, n4187);
nand_4 g04932(new_n5309, n11311, n10451);
xor_3  g04933(new_n5310, new_n5309, new_n5308);
xor_3  g04934(new_n5311, new_n5310, new_n5307);
xnor_3 g04935(new_n5312, new_n5311, new_n5305_1);
nand_4 g04936(new_n5313, new_n4798, new_n4796);
nand_4 g04937(new_n5314_1, new_n4809, new_n4799);
nand_4 g04938(new_n5315, new_n5314_1, new_n5313);
nand_4 g04939(new_n5316, n11423, n9400);
not_3  g04940(new_n5317, new_n5316);
xor_3  g04941(new_n5318, new_n5317, new_n5315);
xnor_3 g04942(new_n5319_1, new_n5318, new_n5312);
xnor_3 g04943(new_n5320_1, new_n5319_1, new_n5302);
not_3  g04944(new_n5321, new_n4794);
nor_4  g04945(new_n5322, new_n5321, new_n4784);
not_3  g04946(new_n5323, new_n4795);
nor_4  g04947(new_n5324, new_n4811, new_n5323);
nor_4  g04948(new_n5325, new_n5324, new_n5322);
nand_4 g04949(new_n5326, new_n5074, new_n5047);
nand_4 g04950(new_n5327, new_n5095, new_n5075);
nand_4 g04951(new_n5328, new_n5327, new_n5326);
xnor_3 g04952(new_n5329, new_n5328, new_n5325);
xnor_3 g04953(new_n5330, new_n5329, new_n5320_1);
xnor_3 g04954(new_n5331_1, new_n5330, new_n5299);
nand_4 g04955(new_n5332, new_n5220, new_n5158);
nand_4 g04956(new_n5333, new_n5332, new_n5167);
xnor_3 g04957(new_n5334, new_n5333, new_n5331_1);
nand_4 g04958(new_n5335, new_n4666, new_n4664);
nor_4  g04959(new_n5336, new_n4674, new_n4668);
not_3  g04960(new_n5337, new_n5336);
nand_4 g04961(new_n5338, new_n5337, new_n5335);
nand_4 g04962(new_n5339, n12591, n11821);
nand_4 g04963(new_n5340, n9080, n3932);
xor_3  g04964(new_n5341, new_n5340, new_n5339);
nand_4 g04965(new_n5342, n10174, n6703);
nand_4 g04966(new_n5343, n12753, n9640);
not_3  g04967(new_n5344, new_n5343);
xor_3  g04968(new_n5345, new_n5344, new_n5342);
nand_4 g04969(new_n5346, n9583, n1333);
nand_4 g04970(new_n5347, n6877, n2278);
xor_3  g04971(new_n5348, new_n5347, new_n5346);
xor_3  g04972(new_n5349, new_n5348, new_n5345);
xnor_3 g04973(new_n5350, new_n5349, new_n5341);
xnor_3 g04974(new_n5351, new_n5350, new_n5338);
nand_4 g04975(new_n5352, new_n4684, new_n4650);
nand_4 g04976(new_n5353, new_n4707, new_n4685);
nand_4 g04977(new_n5354, new_n5353, new_n5352);
nand_4 g04978(new_n5355, new_n4965, new_n4964);
not_3  g04979(new_n5356, new_n4962);
nand_4 g04980(new_n5357, new_n4967, new_n5356);
nand_4 g04981(new_n5358, new_n5357, new_n5355);
nand_4 g04982(new_n5359, n11922, n6294);
nand_4 g04983(new_n5360, new_n4951, new_n4949);
nand_4 g04984(new_n5361, new_n4960, new_n4952);
nand_4 g04985(new_n5362, new_n5361, new_n5360);
nand_4 g04986(new_n5363, n11478, n4094);
not_3  g04987(new_n5364, new_n5363);
xnor_3 g04988(new_n5365, new_n5364, new_n5362);
nor_4  g04989(new_n5366, new_n5051, new_n5050);
not_3  g04990(new_n5367, new_n5052);
nor_4  g04991(new_n5368, new_n5058, new_n5367);
nor_4  g04992(new_n5369, new_n5368, new_n5366);
not_3  g04993(new_n5370, new_n5062);
nor_4  g04994(new_n5371, new_n5064, new_n5370);
not_3  g04995(new_n5372, new_n5061);
nor_4  g04996(new_n5373, new_n5065, new_n5372);
nor_4  g04997(new_n5374, new_n5373, new_n5371);
nand_4 g04998(new_n5375, n12247, n3992);
nand_4 g04999(new_n5376, n8384, n1510);
not_3  g05000(new_n5377, new_n5376);
xor_3  g05001(new_n5378, new_n5377, new_n5375);
xnor_3 g05002(new_n5379, new_n5378, new_n5374);
xnor_3 g05003(new_n5380, new_n5379, new_n5369);
xnor_3 g05004(new_n5381, new_n5380, new_n5365);
xnor_3 g05005(new_n5382, new_n5381, new_n5359);
xnor_3 g05006(new_n5383, new_n5382, new_n5358);
xnor_3 g05007(new_n5384, new_n5383, new_n5354);
nand_4 g05008(new_n5385, new_n5071, new_n5070);
not_3  g05009(new_n5386, new_n5068);
nand_4 g05010(new_n5387, new_n5073, new_n5386);
nand_4 g05011(new_n5388, new_n5387, new_n5385);
not_3  g05012(new_n5389, new_n5060);
nand_4 g05013(new_n5390, new_n5066, new_n5389);
not_3  g05014(new_n5391, new_n5059);
nand_4 g05015(new_n5392, new_n5067, new_n5391);
nand_4 g05016(new_n5393, new_n5392, new_n5390);
not_3  g05017(new_n5394, new_n4947);
nor_4  g05018(new_n5395, new_n5394, new_n4937);
not_3  g05019(new_n5396, new_n4948);
nor_4  g05020(new_n5397, new_n4961, new_n5396);
nor_4  g05021(new_n5398, new_n5397, new_n5395);
xnor_3 g05022(new_n5399, new_n5398, new_n5393);
xnor_3 g05023(new_n5400, new_n5399, new_n5388);
not_3  g05024(new_n5401, new_n4956);
nor_4  g05025(new_n5402, new_n4958, new_n5401);
nor_4  g05026(new_n5403, new_n4959, new_n4955);
nor_4  g05027(new_n5404, new_n5403, new_n5402);
nand_4 g05028(new_n5405, n7862, n753);
nand_4 g05029(new_n5406, n12511, n7236);
not_3  g05030(new_n5407, new_n5406);
xor_3  g05031(new_n5408, new_n5407, new_n5405);
xnor_3 g05032(new_n5409, new_n5408, new_n5404);
nand_4 g05033(new_n5410, new_n4792, new_n4786);
nand_4 g05034(new_n5411_1, new_n5410, new_n4791);
nand_4 g05035(new_n5412, n10898, n7646);
nand_4 g05036(new_n5413, n6826, n1798);
xor_3  g05037(new_n5414, new_n5413, new_n5412);
nand_4 g05038(new_n5415, n11876, n4722);
nand_4 g05039(new_n5416, n3754, n1471);
xor_3  g05040(new_n5417, new_n5416, new_n5415);
xnor_3 g05041(new_n5418, new_n5417, new_n5414);
xnor_3 g05042(new_n5419, new_n5418, new_n5411_1);
xnor_3 g05043(new_n5420, new_n5419, new_n5409);
nand_4 g05044(new_n5421, n3146, n1067);
nand_4 g05045(new_n5422, n2551, n137);
xor_3  g05046(new_n5423, new_n5422, new_n5421);
nand_4 g05047(new_n5424, n8665, n6797);
nand_4 g05048(new_n5425, n12826, n5283);
xor_3  g05049(new_n5426, new_n5425, new_n5424);
xnor_3 g05050(new_n5427, new_n5426, new_n5423);
nand_4 g05051(new_n5428, new_n4942, new_n4939);
nand_4 g05052(new_n5429, new_n5428, new_n4945);
nand_4 g05053(new_n5430, n10685, n4805);
nand_4 g05054(new_n5431, n5645, n4938);
xor_3  g05055(new_n5432, new_n5431, new_n5430);
xnor_3 g05056(new_n5433, new_n5432, new_n5429);
xnor_3 g05057(new_n5434, new_n5433, new_n5427);
not_3  g05058(new_n5435_1, new_n5054);
nor_4  g05059(new_n5436, new_n5056, new_n5435_1);
not_3  g05060(new_n5437, new_n5053);
nor_4  g05061(new_n5438, new_n5057, new_n5437);
nor_4  g05062(new_n5439, new_n5438, new_n5436);
nand_4 g05063(new_n5440, n6358, n159);
nand_4 g05064(new_n5441, n5198, n2749);
xor_3  g05065(new_n5442, new_n5441, new_n5440);
xnor_3 g05066(new_n5443, new_n5442, new_n5439);
xnor_3 g05067(new_n5444, new_n5443, new_n5434);
xnor_3 g05068(new_n5445, new_n5444, new_n5420);
nand_4 g05069(new_n5446, new_n4681, new_n4680);
nand_4 g05070(new_n5447, new_n4683, new_n4677);
nand_4 g05071(new_n5448, new_n5447, new_n5446);
xnor_3 g05072(new_n5449, new_n5448, new_n5445);
xnor_3 g05073(new_n5450, new_n5449, new_n5400);
xnor_3 g05074(new_n5451, new_n5450, new_n5384);
xnor_3 g05075(new_n5452, new_n5451, new_n5351);
nor_4  g05076(new_n5453, new_n4819, new_n4817_1);
nor_4  g05077(new_n5454, new_n4822, new_n4812);
nor_4  g05078(new_n5455, new_n5454, new_n5453);
nand_4 g05079(new_n5456, new_n5096, new_n4970_1);
nand_4 g05080(new_n5457, new_n5156, new_n5165);
nand_4 g05081(new_n5458, new_n5457, new_n5456);
xnor_3 g05082(new_n5459, new_n5458, new_n5455);
xnor_3 g05083(new_n5460, new_n5459, new_n5452);
nor_4  g05084(new_n5461, new_n4671, new_n4670);
not_3  g05085(new_n5462, new_n4670);
nor_4  g05086(new_n5463, new_n4672, new_n5462);
or_4   g05087(new_n5464, new_n5463, new_n4669);
not_3  g05088(new_n5465, new_n5464);
or_4   g05089(new_n5466, new_n5465, new_n5461);
nand_4 g05090(new_n5467, n11757, n11662);
nand_4 g05091(new_n5468, n7456, n5240);
xor_3  g05092(new_n5469, new_n5468, new_n5467);
xor_3  g05093(new_n5470, new_n5469, new_n5466);
not_3  g05094(new_n5471, new_n5470);
xnor_3 g05095(new_n5472, new_n5471, new_n5460);
xnor_3 g05096(new_n5473, new_n5472, new_n5334);
nand_4 g05097(new_n5474, new_n5473, new_n5291);
not_3  g05098(new_n5475, new_n5290);
xnor_3 g05099(new_n5476, new_n5475, new_n5281);
xnor_3 g05100(new_n5477, new_n5470, new_n5460);
xnor_3 g05101(new_n5478, new_n5477, new_n5334);
nand_4 g05102(new_n5479, new_n5478, new_n5476);
nand_4 g05103(n1269, new_n5479, new_n5474);
nand_4 g05104(new_n5481, n10223, n4312);
not_3  g05105(new_n5482, new_n5481);
nand_4 g05106(new_n5483, n12705, n7265);
nand_4 g05107(new_n5484, n4312, n2879);
not_3  g05108(new_n5485, new_n5484);
nand_4 g05109(new_n5486, n10223, n1097);
xnor_3 g05110(new_n5487, new_n5486, new_n5483);
nor_4  g05111(new_n5488, new_n5487, new_n5485);
nor_4  g05112(new_n5489, new_n5488, new_n5483);
nor_4  g05113(new_n5490, new_n5489, new_n5482);
nor_4  g05114(new_n5491, new_n5489, new_n1087);
nor_4  g05115(new_n5492, new_n5491, new_n5481);
nor_4  g05116(new_n5493, new_n5492, new_n5490);
nand_4 g05117(new_n5494, n12025, n7265);
nand_4 g05118(new_n5495, n12705, n2879);
xor_3  g05119(new_n5496, new_n5495, new_n5494);
xnor_3 g05120(new_n5497, new_n5496, new_n5493);
not_3  g05121(new_n5498, new_n5497);
nand_4 g05122(new_n5499, n9195, n5964);
nand_4 g05123(new_n5500, n4634, n1097);
xor_3  g05124(new_n5501, new_n5500, new_n5499);
xnor_3 g05125(new_n5502, new_n5501, new_n5498);
nand_4 g05126(new_n5503, n5964, n4634);
not_3  g05127(new_n5504, new_n5503);
not_3  g05128(new_n5505, new_n1088);
not_3  g05129(new_n5506, new_n1089);
nor_4  g05130(new_n5507, new_n5506, new_n5505);
nor_4  g05131(new_n5508, new_n1089, new_n1088);
nor_4  g05132(new_n5509, new_n5508, new_n1087);
nor_4  g05133(new_n5510, new_n5509, new_n5507);
and_4  g05134(new_n5511, new_n5510, new_n5504);
xor_3  g05135(new_n5512, new_n5487, new_n5485);
xor_3  g05136(new_n5513, new_n5510, new_n5503);
nor_4  g05137(new_n5514, new_n5513, new_n5512);
nor_4  g05138(new_n5515, new_n5514, new_n5511);
xnor_3 g05139(new_n5516, new_n5515, new_n5502);
not_3  g05140(new_n5517, new_n5516);
nand_4 g05141(new_n5518, n9195, n5305);
not_3  g05142(new_n5519, new_n5518);
nand_4 g05143(new_n5520, new_n1091, new_n1085);
nand_4 g05144(new_n5521, new_n5520, new_n1082);
nor_4  g05145(new_n5522, new_n5521, new_n5519);
xor_3  g05146(new_n5523, new_n5510, new_n5504);
xnor_3 g05147(new_n5524, new_n5523, new_n5512);
xnor_3 g05148(new_n5525, new_n5521, new_n5519);
nor_4  g05149(new_n5526, new_n5525, new_n5524);
nor_4  g05150(new_n5527, new_n5526, new_n5522);
nand_4 g05151(new_n5528, new_n5527, new_n5517);
not_3  g05152(new_n5529, new_n5492);
nand_4 g05153(new_n5530, new_n5496, new_n5493);
nand_4 g05154(new_n5531, new_n5530, new_n5529);
nand_4 g05155(new_n5532, n5964, n2253);
nand_4 g05156(new_n5533, n9195, n1097);
nand_4 g05157(new_n5534, n5305, n3865);
not_3  g05158(new_n5535, new_n5534);
xor_3  g05159(new_n5536, new_n5535, new_n5533);
xnor_3 g05160(new_n5537, new_n5536, new_n5532);
xnor_3 g05161(new_n5538, new_n5537, new_n5531);
nor_4  g05162(new_n5539, new_n5495, new_n5494);
not_3  g05163(new_n5540, new_n5539);
nand_4 g05164(new_n5541, n4634, n4312);
xor_3  g05165(new_n5542, new_n5541, new_n5540);
nand_4 g05166(new_n5543, n12025, n2879);
nand_4 g05167(new_n5544, n11257, n7265);
nand_4 g05168(new_n5545, n12705, n10223);
not_3  g05169(new_n5546, new_n5545);
xor_3  g05170(new_n5547, new_n5546, new_n5544);
xnor_3 g05171(new_n5548, new_n5547, new_n5543);
xnor_3 g05172(new_n5549, new_n5548, new_n5542);
xnor_3 g05173(new_n5550, new_n5549, new_n5538);
nand_4 g05174(new_n5551, new_n5501, new_n5498);
nor_4  g05175(new_n5552, new_n5500, new_n5499);
nor_4  g05176(new_n5553, new_n5515, new_n5502);
xnor_3 g05177(new_n5554, new_n5553, new_n5552);
nand_4 g05178(new_n5555, new_n5554, new_n5551);
xnor_3 g05179(new_n5556, new_n5555, new_n5550);
xnor_3 g05180(new_n5557, new_n5556, new_n5528);
not_3  g05181(new_n5558, new_n5557);
nand_4 g05182(new_n5559, n5305, n2253);
not_3  g05183(new_n5560, new_n5559);
xnor_3 g05184(new_n5561, new_n5527, new_n5516);
nand_4 g05185(new_n5562, new_n5561, new_n5560);
nor_4  g05186(new_n5563, new_n1101, new_n1093);
not_3  g05187(new_n5564, new_n5563);
not_3  g05188(new_n5565, new_n5525);
xnor_3 g05189(new_n5566, new_n5565, new_n5524);
nor_4  g05190(new_n5567, new_n5566, new_n5564);
xnor_3 g05191(new_n5568, new_n5561, new_n5559);
nand_4 g05192(new_n5569, new_n5568, new_n5567);
nand_4 g05193(new_n5570, new_n5569, new_n5562);
xor_3  g05194(new_n5571, new_n5570, new_n5558);
not_3  g05195(new_n5572, new_n5569);
nor_4  g05196(new_n5573, new_n5568, new_n5567);
nor_4  g05197(new_n5574, new_n5573, new_n5572);
not_3  g05198(new_n5575, new_n5574);
nor_4  g05199(new_n5576, new_n1229, new_n1226);
not_3  g05200(new_n5577, new_n5576);
nand_4 g05201(new_n5578, n12145, n8759);
not_3  g05202(new_n5579_1, new_n1216);
nand_4 g05203(new_n5580, new_n1217, new_n5579_1);
nand_4 g05204(new_n5581, new_n1225, new_n1218);
nand_4 g05205(new_n5582, new_n5581, new_n5580);
not_3  g05206(new_n5583, new_n5582);
xnor_3 g05207(new_n5584, new_n5583, new_n5578);
nand_4 g05208(new_n5585, n6776, n2522);
not_3  g05209(new_n5586, new_n1222);
not_3  g05210(new_n5587, new_n1223);
nor_4  g05211(new_n5588, new_n5587, new_n5586);
nor_4  g05212(new_n5589, new_n1223, new_n1222);
nor_4  g05213(new_n5590, new_n5589, new_n1221);
nor_4  g05214(new_n5591, new_n5590, new_n5588);
xnor_3 g05215(new_n5592, new_n5591, new_n5585);
nand_4 g05216(new_n5593, n7436, n2024);
not_3  g05217(new_n5594, new_n5593);
nand_4 g05218(new_n5595, n12299, n9189);
nand_4 g05219(new_n5596, n8276, n7946);
xnor_3 g05220(new_n5597, new_n5596, new_n5595);
xnor_3 g05221(new_n5598, new_n5597, new_n5594);
xnor_3 g05222(new_n5599, new_n5598, new_n5592);
not_3  g05223(new_n5600, new_n5599);
xor_3  g05224(new_n5601, new_n5600, new_n5584);
nor_4  g05225(new_n5602, new_n5601, new_n5577);
not_3  g05226(new_n5603, new_n5602);
nand_4 g05227(new_n5604, n12221, n8759);
not_3  g05228(new_n5605, new_n5585);
nand_4 g05229(new_n5606, new_n5591, new_n5605);
nand_4 g05230(new_n5607, new_n5598, new_n5592);
nand_4 g05231(new_n5608, new_n5607, new_n5606);
nand_4 g05232(new_n5609, n12145, n6776);
nand_4 g05233(new_n5610, n12299, n2522);
xor_3  g05234(new_n5611, new_n5610, new_n5609);
xnor_3 g05235(new_n5612, new_n5611, new_n5608);
nand_4 g05236(new_n5613, n9189, n7436);
not_3  g05237(new_n5614, new_n5613);
nor_4  g05238(new_n5615, new_n5597, new_n5594);
nor_4  g05239(new_n5616, new_n5615, new_n5596);
nor_4  g05240(new_n5617, new_n5616, new_n5614);
nor_4  g05241(new_n5618, new_n5616, new_n1221);
nor_4  g05242(new_n5619, new_n5618, new_n5613);
nor_4  g05243(new_n5620, new_n5619, new_n5617);
nand_4 g05244(new_n5621, n8276, n2024);
nand_4 g05245(new_n5622, n9241, n7946);
xor_3  g05246(new_n5623, new_n5622, new_n5621);
xnor_3 g05247(new_n5624, new_n5623, new_n5620);
xnor_3 g05248(new_n5625, new_n5624, new_n5612);
nor_4  g05249(new_n5626, new_n5583, new_n5578);
nor_4  g05250(new_n5627, new_n5599, new_n5584);
nor_4  g05251(new_n5628, new_n5627, new_n5626);
xnor_3 g05252(new_n5629, new_n5628, new_n5625);
nor_4  g05253(new_n5630, new_n5629, new_n5604);
not_3  g05254(new_n5631, new_n5604);
not_3  g05255(new_n5632, new_n5629);
nor_4  g05256(new_n5633, new_n5632, new_n5631);
nor_4  g05257(new_n5634, new_n5633, new_n5630);
xnor_3 g05258(new_n5635, new_n5634, new_n5603);
xnor_3 g05259(new_n5636, new_n5601, new_n5576);
nand_4 g05260(new_n5637, n6016, n5331);
nand_4 g05261(new_n5638, n8476, n521);
not_3  g05262(new_n5639, new_n5638);
not_3  g05263(new_n5640, new_n1241);
nor_4  g05264(new_n5641_1, new_n1247, new_n5640);
nor_4  g05265(new_n5642, new_n5641_1, new_n1246);
xnor_3 g05266(new_n5643, new_n5642, new_n5639);
nand_4 g05267(new_n5644, n12648, n2498);
not_3  g05268(new_n5645_1, new_n5644);
nand_4 g05269(new_n5646, n5579, n2530);
not_3  g05270(new_n5647, new_n5646);
nand_4 g05271(new_n5648, n10545, n2558);
not_3  g05272(new_n5649, new_n5648);
nor_4  g05273(new_n5650, new_n5649, new_n5647);
nor_4  g05274(new_n5651, new_n5648, new_n5646);
nor_4  g05275(new_n5652, new_n5651, new_n5650);
xnor_3 g05276(new_n5653, new_n5652, new_n5645_1);
xnor_3 g05277(new_n5654, new_n5653, new_n5643);
nor_4  g05278(new_n5655, new_n5654, new_n5637);
not_3  g05279(new_n5656, new_n5637);
not_3  g05280(new_n5657, new_n5654);
nor_4  g05281(new_n5658, new_n5657, new_n5656);
nor_4  g05282(new_n5659, new_n5658, new_n5655);
nor_4  g05283(new_n5660, new_n1239, new_n1235);
nor_4  g05284(new_n5661, new_n1250, new_n1240);
nor_4  g05285(new_n5662, new_n5661, new_n5660);
not_3  g05286(new_n5663, new_n5662);
xnor_3 g05287(new_n5664, new_n5663, new_n5659);
xnor_3 g05288(new_n5665, new_n5664, new_n1255);
not_3  g05289(new_n5666, new_n1277);
nand_4 g05290(new_n5667, n7965, n7270);
nand_4 g05291(new_n5668, n7388, n806);
not_3  g05292(new_n5669, new_n5668);
not_3  g05293(new_n5670_1, new_n1263);
nor_4  g05294(new_n5671, new_n1269_1, new_n5670_1);
nor_4  g05295(new_n5672, new_n5671, new_n1268);
xnor_3 g05296(new_n5673, new_n5672, new_n5669);
nand_4 g05297(new_n5674, n9111, n2393);
not_3  g05298(new_n5675, new_n5674);
nand_4 g05299(new_n5676, n11892, n3342);
not_3  g05300(new_n5677, new_n5676);
nand_4 g05301(new_n5678, n9763, n5860);
not_3  g05302(new_n5679, new_n5678);
nor_4  g05303(new_n5680, new_n5679, new_n5677);
nor_4  g05304(new_n5681, new_n5678, new_n5676);
nor_4  g05305(new_n5682, new_n5681, new_n5680);
xnor_3 g05306(new_n5683, new_n5682, new_n5675);
xnor_3 g05307(new_n5684, new_n5683, new_n5673);
nor_4  g05308(new_n5685, new_n5684, new_n5667);
not_3  g05309(new_n5686, new_n5667);
not_3  g05310(new_n5687, new_n5684);
nor_4  g05311(new_n5688, new_n5687, new_n5686);
nor_4  g05312(new_n5689, new_n5688, new_n5685);
nor_4  g05313(new_n5690, new_n1261, new_n1259);
nor_4  g05314(new_n5691, new_n1272, new_n1262);
nor_4  g05315(new_n5692, new_n5691, new_n5690);
not_3  g05316(new_n5693_1, new_n5692);
xnor_3 g05317(new_n5694_1, new_n5693_1, new_n5689);
nor_4  g05318(new_n5695, new_n5694_1, new_n5666);
not_3  g05319(new_n5696, new_n5694_1);
nor_4  g05320(new_n5697, new_n5696, new_n1277);
nor_4  g05321(new_n5698, new_n5697, new_n5695);
xnor_3 g05322(new_n5699, new_n5698, new_n5665);
nor_4  g05323(new_n5700, new_n1280, new_n1258);
nor_4  g05324(new_n5701, new_n1287, new_n5700);
xnor_3 g05325(new_n5702, new_n5701, new_n5699);
nor_4  g05326(new_n5703, new_n5702, new_n5636);
not_3  g05327(new_n5704, new_n5703);
nand_4 g05328(new_n5705, new_n5702, new_n5636);
nor_4  g05329(new_n5706, new_n1233, new_n1230);
nor_4  g05330(new_n5707, new_n1288, new_n1234);
nor_4  g05331(new_n5708, new_n5707, new_n5706);
nand_4 g05332(new_n5709, new_n5708, new_n5705);
nand_4 g05333(new_n5710, new_n5709, new_n5704);
xnor_3 g05334(new_n5711, new_n5710, new_n5635);
not_3  g05335(new_n5712, new_n1255);
nor_4  g05336(new_n5713, new_n5664, new_n5712);
nand_4 g05337(new_n5714, n5798, n5331);
nand_4 g05338(new_n5715, n12648, n5579);
nand_4 g05339(new_n5716, n10545, n2498);
nand_4 g05340(new_n5717, n7690, n2558);
xnor_3 g05341(new_n5718, new_n5717, new_n5716);
nor_4  g05342(new_n5719, new_n5718, new_n5715);
not_3  g05343(new_n5720, new_n5715);
not_3  g05344(new_n5721, new_n5718);
nor_4  g05345(new_n5722, new_n5721, new_n5720);
nor_4  g05346(new_n5723, new_n5722, new_n5719);
nor_4  g05347(new_n5724, new_n5651, new_n5645_1);
nor_4  g05348(new_n5725, new_n5724, new_n5650);
xnor_3 g05349(new_n5726, new_n5725, new_n5723);
nand_4 g05350(new_n5727, n8476, n6016);
nand_4 g05351(new_n5728, n2530, n521);
xor_3  g05352(new_n5729, new_n5728, new_n5727);
xnor_3 g05353(new_n5730, new_n5729, new_n5726);
and_4  g05354(new_n5731, new_n5642, new_n5639);
nor_4  g05355(new_n5732, new_n5653, new_n5643);
nor_4  g05356(new_n5733, new_n5732, new_n5731);
xnor_3 g05357(new_n5734, new_n5733, new_n5730);
not_3  g05358(new_n5735, new_n5655);
nand_4 g05359(new_n5736, new_n5663, new_n5659);
nand_4 g05360(new_n5737, new_n5736, new_n5735);
xnor_3 g05361(new_n5738, new_n5737, new_n5734);
nor_4  g05362(new_n5739, new_n5738, new_n5714);
not_3  g05363(new_n5740, new_n5714);
not_3  g05364(new_n5741, new_n5738);
nor_4  g05365(new_n5742, new_n5741, new_n5740);
nor_4  g05366(new_n5743, new_n5742, new_n5739);
xnor_3 g05367(new_n5744, new_n5743, new_n5713);
not_3  g05368(new_n5745, new_n5695);
nand_4 g05369(new_n5746, n7965, n5153);
nand_4 g05370(new_n5747, n3342, n2393);
nand_4 g05371(new_n5748, n9763, n3986);
nand_4 g05372(new_n5749, n9111, n5860);
xnor_3 g05373(new_n5750, new_n5749, new_n5748);
nor_4  g05374(new_n5751, new_n5750, new_n5747);
not_3  g05375(new_n5752, new_n5747);
not_3  g05376(new_n5753, new_n5750);
nor_4  g05377(new_n5754, new_n5753, new_n5752);
nor_4  g05378(new_n5755, new_n5754, new_n5751);
nor_4  g05379(new_n5756, new_n5681, new_n5675);
nor_4  g05380(new_n5757, new_n5756, new_n5680);
xnor_3 g05381(new_n5758, new_n5757, new_n5755);
nand_4 g05382(new_n5759, n7388, n7270);
nand_4 g05383(new_n5760_1, n11892, n806);
xor_3  g05384(new_n5761, new_n5760_1, new_n5759);
xnor_3 g05385(new_n5762, new_n5761, new_n5758);
and_4  g05386(new_n5763, new_n5672, new_n5669);
nor_4  g05387(new_n5764, new_n5683, new_n5673);
nor_4  g05388(new_n5765, new_n5764, new_n5763);
xnor_3 g05389(new_n5766, new_n5765, new_n5762);
not_3  g05390(new_n5767_1, new_n5685);
nand_4 g05391(new_n5768, new_n5693_1, new_n5689);
nand_4 g05392(new_n5769, new_n5768, new_n5767_1);
xnor_3 g05393(new_n5770, new_n5769, new_n5766);
nor_4  g05394(new_n5771, new_n5770, new_n5746);
not_3  g05395(new_n5772, new_n5746);
not_3  g05396(new_n5773, new_n5770);
nor_4  g05397(new_n5774, new_n5773, new_n5772);
nor_4  g05398(new_n5775, new_n5774, new_n5771);
nor_4  g05399(new_n5776, new_n5775, new_n5745);
xnor_3 g05400(new_n5777, new_n5770, new_n5746);
nor_4  g05401(new_n5778, new_n5777, new_n5695);
nor_4  g05402(new_n5779, new_n5778, new_n5776);
not_3  g05403(new_n5780, new_n5779);
xnor_3 g05404(new_n5781, new_n5780, new_n5744);
nor_4  g05405(new_n5782, new_n5698, new_n5665);
nor_4  g05406(new_n5783, new_n5701, new_n5699);
nor_4  g05407(new_n5784, new_n5783, new_n5782);
not_3  g05408(new_n5785, new_n5784);
xnor_3 g05409(new_n5786, new_n5785, new_n5781);
xnor_3 g05410(new_n5787, new_n5786, new_n5711);
nor_4  g05411(new_n5788, new_n5787, new_n5575);
not_3  g05412(new_n5789, new_n5787);
nor_4  g05413(new_n5790, new_n5789, new_n5574);
xor_3  g05414(new_n5791, new_n5566, new_n5563);
not_3  g05415(new_n5792, new_n5708);
nand_4 g05416(new_n5793, new_n5705, new_n5704);
xnor_3 g05417(new_n5794, new_n5793, new_n5792);
not_3  g05418(new_n5795, new_n5794);
nor_4  g05419(new_n5796, new_n5795, new_n5791);
not_3  g05420(new_n5797, new_n5791);
nor_4  g05421(new_n5798_1, new_n5794, new_n5797);
nand_4 g05422(new_n5799, new_n1214, new_n1102);
not_3  g05423(new_n5800, new_n5799);
nor_4  g05424(new_n5801, new_n1289, new_n1215);
nor_4  g05425(new_n5802, new_n5801, new_n5800);
nor_4  g05426(new_n5803, new_n5802, new_n5798_1);
nor_4  g05427(new_n5804, new_n5803, new_n5796);
nor_4  g05428(new_n5805, new_n5804, new_n5790);
nor_4  g05429(new_n5806, new_n5805, new_n5788);
xnor_3 g05430(new_n5807, new_n5806, new_n5571);
not_3  g05431(new_n5808, new_n5630);
nand_4 g05432(new_n5809, new_n5634, new_n5602);
nand_4 g05433(new_n5810, new_n5809, new_n5808);
nor_4  g05434(new_n5811, new_n5628, new_n5625);
not_3  g05435(new_n5812, new_n5619);
nand_4 g05436(new_n5813, new_n5623, new_n5620);
nand_4 g05437(new_n5814_1, new_n5813, new_n5812);
nand_4 g05438(new_n5815, n12221, n6776);
nand_4 g05439(new_n5816, n12299, n12145);
nand_4 g05440(new_n5817, n10217, n8759);
not_3  g05441(new_n5818, new_n5817);
xor_3  g05442(new_n5819, new_n5818, new_n5816);
xnor_3 g05443(new_n5820, new_n5819, new_n5815);
xnor_3 g05444(new_n5821, new_n5820, new_n5814_1);
nor_4  g05445(new_n5822, new_n5622, new_n5621);
nand_4 g05446(new_n5823, n7436, n2522);
not_3  g05447(new_n5824, new_n5823);
xor_3  g05448(new_n5825, new_n5824, new_n5822);
nand_4 g05449(new_n5826, n9241, n2024);
nand_4 g05450(new_n5827, n10510, n7946);
nand_4 g05451(new_n5828, n9189, n8276);
nand_4 g05452(new_n5829, new_n5828, new_n5827);
not_3  g05453(new_n5830, new_n5827);
not_3  g05454(new_n5831, new_n5828);
nand_4 g05455(new_n5832, new_n5831, new_n5830);
nand_4 g05456(new_n5833, new_n5832, new_n5829);
xor_3  g05457(new_n5834, new_n5833, new_n5826);
xnor_3 g05458(new_n5835, new_n5834, new_n5825);
xnor_3 g05459(new_n5836, new_n5835, new_n5821);
nand_4 g05460(new_n5837, new_n5611, new_n5608);
nor_4  g05461(new_n5838, new_n5610, new_n5609);
nor_4  g05462(new_n5839, new_n5624, new_n5612);
xnor_3 g05463(new_n5840, new_n5839, new_n5838);
nand_4 g05464(new_n5841, new_n5840, new_n5837);
xnor_3 g05465(new_n5842, new_n5841, new_n5836);
not_3  g05466(new_n5843, new_n5842);
xor_3  g05467(new_n5844, new_n5843, new_n5811);
xnor_3 g05468(new_n5845, new_n5844, new_n5810);
not_3  g05469(new_n5846, new_n5710);
nand_4 g05470(new_n5847, new_n5846, new_n5635);
nand_4 g05471(new_n5848, new_n5786, new_n5711);
nand_4 g05472(new_n5849, new_n5848, new_n5847);
xnor_3 g05473(new_n5850, new_n5849, new_n5845);
not_3  g05474(new_n5851, new_n5734);
not_3  g05475(new_n5852, new_n5737);
nor_4  g05476(new_n5853, new_n5852, new_n5851);
not_3  g05477(new_n5854, new_n5719);
nand_4 g05478(new_n5855, new_n5725, new_n5723);
nand_4 g05479(new_n5856, new_n5855, new_n5854);
nand_4 g05480(new_n5857_1, n8476, n5798);
nand_4 g05481(new_n5858, n6016, n2530);
nand_4 g05482(new_n5859, n5331, n2347);
xnor_3 g05483(new_n5860_1, new_n5859, new_n5858);
xnor_3 g05484(new_n5861, new_n5860_1, new_n5857_1);
xnor_3 g05485(new_n5862, new_n5861, new_n5856);
nor_4  g05486(new_n5863, new_n5717, new_n5716);
nand_4 g05487(new_n5864, n12648, n521);
xnor_3 g05488(new_n5865, new_n5864, new_n5863);
nand_4 g05489(new_n5866, n7690, n2498);
not_3  g05490(new_n5867, new_n5866);
nand_4 g05491(new_n5868, n10545, n5579);
nand_4 g05492(new_n5869, n3616, n2558);
xnor_3 g05493(new_n5870, new_n5869, new_n5868);
xnor_3 g05494(new_n5871, new_n5870, new_n5867);
not_3  g05495(new_n5872, new_n5871);
xor_3  g05496(new_n5873, new_n5872, new_n5865);
xnor_3 g05497(new_n5874, new_n5873, new_n5862);
not_3  g05498(new_n5875, new_n5874);
not_3  g05499(new_n5876, new_n5726);
nand_4 g05500(new_n5877, new_n5729, new_n5876);
nor_4  g05501(new_n5878, new_n5728, new_n5727);
not_3  g05502(new_n5879, new_n5730);
nor_4  g05503(new_n5880, new_n5733, new_n5879);
xnor_3 g05504(new_n5881, new_n5880, new_n5878);
nand_4 g05505(new_n5882, new_n5881, new_n5877);
xnor_3 g05506(new_n5883, new_n5882, new_n5875);
xnor_3 g05507(new_n5884, new_n5883, new_n5853);
not_3  g05508(new_n5885, new_n5739);
nand_4 g05509(new_n5886, new_n5743, new_n5713);
nand_4 g05510(new_n5887, new_n5886, new_n5885);
xnor_3 g05511(new_n5888, new_n5887, new_n5884);
not_3  g05512(new_n5889, new_n5888);
not_3  g05513(new_n5890, new_n5766);
not_3  g05514(new_n5891, new_n5769);
nor_4  g05515(new_n5892, new_n5891, new_n5890);
not_3  g05516(new_n5893, new_n5892);
not_3  g05517(new_n5894, new_n5751);
nand_4 g05518(new_n5895, new_n5757, new_n5755);
nand_4 g05519(new_n5896, new_n5895, new_n5894);
nand_4 g05520(new_n5897, n7388, n5153);
nand_4 g05521(new_n5898, n11892, n7270);
nand_4 g05522(new_n5899, n7965, n2507);
xnor_3 g05523(new_n5900, new_n5899, new_n5898);
xnor_3 g05524(new_n5901, new_n5900, new_n5897);
xnor_3 g05525(new_n5902, new_n5901, new_n5896);
nor_4  g05526(new_n5903, new_n5749, new_n5748);
nand_4 g05527(new_n5904, n2393, n806);
xnor_3 g05528(new_n5905, new_n5904, new_n5903);
nand_4 g05529(new_n5906, n9111, n3986);
not_3  g05530(new_n5907, new_n5906);
nand_4 g05531(new_n5908, n5860, n3342);
nand_4 g05532(new_n5909, n9763, n5857);
xnor_3 g05533(new_n5910, new_n5909, new_n5908);
xnor_3 g05534(new_n5911, new_n5910, new_n5907);
not_3  g05535(new_n5912, new_n5911);
xor_3  g05536(new_n5913, new_n5912, new_n5905);
not_3  g05537(new_n5914, new_n5913);
xor_3  g05538(new_n5915, new_n5914, new_n5902);
not_3  g05539(new_n5916, new_n5915);
not_3  g05540(new_n5917, new_n5758);
nand_4 g05541(new_n5918, new_n5761, new_n5917);
nor_4  g05542(new_n5919, new_n5760_1, new_n5759);
not_3  g05543(new_n5920, new_n5762);
nor_4  g05544(new_n5921, new_n5765, new_n5920);
xnor_3 g05545(new_n5922, new_n5921, new_n5919);
nand_4 g05546(new_n5923, new_n5922, new_n5918);
xnor_3 g05547(new_n5924, new_n5923, new_n5916);
xnor_3 g05548(new_n5925, new_n5924, new_n5893);
nor_4  g05549(new_n5926, new_n5778, new_n5774);
not_3  g05550(new_n5927, new_n5926);
xnor_3 g05551(new_n5928, new_n5927, new_n5925);
not_3  g05552(new_n5929, new_n5928);
nor_4  g05553(new_n5930, new_n5929, new_n5889);
nor_4  g05554(new_n5931, new_n5928, new_n5888);
nor_4  g05555(new_n5932, new_n5931, new_n5930);
not_3  g05556(new_n5933, new_n5932);
nor_4  g05557(new_n5934_1, new_n5779, new_n5744);
not_3  g05558(new_n5935, new_n5934_1);
nand_4 g05559(new_n5936, new_n5784, new_n5781);
nand_4 g05560(new_n5937, new_n5936, new_n5935);
nor_4  g05561(new_n5938, new_n5937, new_n5933);
not_3  g05562(new_n5939, new_n5937);
nor_4  g05563(new_n5940, new_n5939, new_n5932);
nor_4  g05564(new_n5941, new_n5940, new_n5938);
xnor_3 g05565(new_n5942, new_n5941, new_n5850);
xnor_3 g05566(n1523, new_n5942, new_n5807);
nand_4 g05567(new_n5944, n7265, n4189);
nand_4 g05568(new_n5945, n10223, n6687);
nand_4 g05569(new_n5946, new_n5945, new_n5944);
not_3  g05570(new_n5947, new_n5944);
not_3  g05571(new_n5948, new_n5945);
nand_4 g05572(new_n5949, new_n5948, new_n5947);
and_4  g05573(new_n5950, new_n5949, new_n5946);
nand_4 g05574(new_n5951, n6687, n2879);
nand_4 g05575(new_n5952, n7265, n2564);
nor_4  g05576(new_n5953, new_n5952, new_n5951);
not_3  g05577(new_n5954, new_n5953);
nor_4  g05578(new_n5955, new_n5954, new_n5950);
nand_4 g05579(new_n5956, n6687, n4634);
not_3  g05580(new_n5957, new_n5956);
nand_4 g05581(new_n5958, n2879, n2564);
not_3  g05582(new_n5959, new_n5958);
nand_4 g05583(new_n5960, new_n5959, new_n5946);
nand_4 g05584(new_n5961, new_n5960, new_n5949);
xor_3  g05585(new_n5962, new_n5961, new_n5957);
nand_4 g05586(new_n5963, n4189, n2879);
nand_4 g05587(new_n5964_1, n10223, n2564);
nand_4 g05588(new_n5965, n7265, n6770);
xnor_3 g05589(new_n5966, new_n5965, new_n5964_1);
xor_3  g05590(new_n5967, new_n5966, new_n5963);
nand_4 g05591(new_n5968, new_n5967, new_n5962);
not_3  g05592(new_n5969, new_n5968);
nor_4  g05593(new_n5970, new_n5967, new_n5962);
nor_4  g05594(new_n5971, new_n5970, new_n5969);
nand_4 g05595(new_n5972, new_n5971, new_n5955);
not_3  g05596(new_n5973, new_n5972);
nand_4 g05597(new_n5974, n9195, n6687);
nand_4 g05598(new_n5975, n4634, n2564);
nand_4 g05599(new_n5976, n6770, n2879);
nand_4 g05600(new_n5977, n10223, n4189);
nand_4 g05601(new_n5978, n9920, n7265);
xnor_3 g05602(new_n5979, new_n5978, new_n5977);
xnor_3 g05603(new_n5980, new_n5979, new_n5976);
xnor_3 g05604(new_n5981, new_n5980, new_n5975);
nand_4 g05605(new_n5982, new_n5965, new_n5964_1);
not_3  g05606(new_n5983, new_n5982);
not_3  g05607(new_n5984, new_n5963);
nor_4  g05608(new_n5985, new_n5966, new_n5984);
nor_4  g05609(new_n5986, new_n5985, new_n5983);
xnor_3 g05610(new_n5987, new_n5986, new_n5981);
not_3  g05611(new_n5988, new_n5987);
nor_4  g05612(new_n5989, new_n5988, new_n5974);
not_3  g05613(new_n5990, new_n5974);
nor_4  g05614(new_n5991, new_n5987, new_n5990);
nor_4  g05615(new_n5992, new_n5991, new_n5989);
not_3  g05616(new_n5993, new_n5961);
nor_4  g05617(new_n5994, new_n5993, new_n5956);
not_3  g05618(new_n5995, new_n5994);
nand_4 g05619(new_n5996, new_n5968, new_n5995);
nand_4 g05620(new_n5997, new_n5996, new_n5992);
not_3  g05621(new_n5998, new_n5997);
nor_4  g05622(new_n5999, new_n5996, new_n5992);
nor_4  g05623(new_n6000, new_n5999, new_n5998);
xor_3  g05624(new_n6001, new_n6000, new_n5973);
nand_4 g05625(new_n6002, n8336, n2522);
nand_4 g05626(new_n6003, n9189, n8336);
not_3  g05627(new_n6004, new_n6003);
nand_4 g05628(new_n6005, n7946, n6986);
not_3  g05629(new_n6006, new_n6005);
nor_4  g05630(new_n6007, new_n6006, new_n6004);
nand_4 g05631(new_n6008, n10928, n2024);
not_3  g05632(new_n6009, new_n6008);
nor_4  g05633(new_n6010, new_n6005, new_n6003);
nor_4  g05634(new_n6011, new_n6010, new_n6009);
nor_4  g05635(new_n6012, new_n6011, new_n6007);
xor_3  g05636(new_n6013, new_n6012, new_n6002);
nand_4 g05637(new_n6014, n6986, n2024);
nand_4 g05638(new_n6015, n10928, n9189);
not_3  g05639(new_n6016_1, new_n6015);
nand_4 g05640(new_n6017, n7946, n2226);
not_3  g05641(new_n6018, new_n6017);
nor_4  g05642(new_n6019, new_n6018, new_n6016_1);
nor_4  g05643(new_n6020, new_n6017, new_n6015);
nor_4  g05644(new_n6021, new_n6020, new_n6019);
xor_3  g05645(new_n6022, new_n6021, new_n6014);
xnor_3 g05646(new_n6023, new_n6022, new_n6013);
not_3  g05647(new_n6024, new_n6007);
nor_4  g05648(new_n6025, new_n6008, new_n4569);
nor_4  g05649(new_n6026, new_n6025, new_n6024);
nor_4  g05650(new_n6027, new_n6026, new_n6010);
nor_4  g05651(new_n6028, new_n6027, new_n6008);
not_3  g05652(new_n6029, new_n6028);
nor_4  g05653(new_n6030, new_n6029, new_n6023);
not_3  g05654(new_n6031, new_n6030);
nand_4 g05655(new_n6032, n12145, n8336);
not_3  g05656(new_n6033, new_n6032);
nand_4 g05657(new_n6034, n10928, n2522);
not_3  g05658(new_n6035, new_n6014);
nor_4  g05659(new_n6036, new_n6020, new_n6035);
nor_4  g05660(new_n6037, new_n6036, new_n6019);
xor_3  g05661(new_n6038_1, new_n6037, new_n6034);
nand_4 g05662(new_n6039, n2226, n2024);
not_3  g05663(new_n6040, new_n6039);
nand_4 g05664(new_n6041, n9189, n6986);
nand_4 g05665(new_n6042, n7946, n1094);
xnor_3 g05666(new_n6043, new_n6042, new_n6041);
xor_3  g05667(new_n6044, new_n6043, new_n6040);
xnor_3 g05668(new_n6045, new_n6044, new_n6038_1);
not_3  g05669(new_n6046, new_n6045);
xor_3  g05670(new_n6047, new_n6046, new_n6033);
not_3  g05671(new_n6048, new_n6002);
and_4  g05672(new_n6049, new_n6012, new_n6048);
not_3  g05673(new_n6050, new_n6049);
nor_4  g05674(new_n6051, new_n6022, new_n6013);
not_3  g05675(new_n6052, new_n6051);
nand_4 g05676(new_n6053, new_n6052, new_n6050);
xnor_3 g05677(new_n6054, new_n6053, new_n6047);
xnor_3 g05678(new_n6055, new_n6054, new_n6031);
not_3  g05679(new_n6056, new_n6023);
xor_3  g05680(new_n6057, new_n6028, new_n6056);
nand_4 g05681(new_n6058, n7891, n2558);
nand_4 g05682(new_n6059, n12069, n5579);
nand_4 g05683(new_n6060, new_n6059, new_n6058);
not_3  g05684(new_n6061, new_n6060);
not_3  g05685(new_n6062, new_n6058);
not_3  g05686(new_n6063, new_n6059);
nand_4 g05687(new_n6064, new_n6063, new_n6062);
not_3  g05688(new_n6065, new_n6064);
nor_4  g05689(new_n6066, new_n6065, new_n6061);
nand_4 g05690(new_n6067, n12391, n2558);
nand_4 g05691(new_n6068, n12069, n2498);
nor_4  g05692(new_n6069, new_n6068, new_n6067);
not_3  g05693(new_n6070, new_n6069);
nor_4  g05694(new_n6071, new_n6070, new_n6066);
not_3  g05695(new_n6072, new_n6071);
nand_4 g05696(new_n6073, n12069, n521);
nand_4 g05697(new_n6074, n12391, n2498);
not_3  g05698(new_n6075, new_n6074);
nand_4 g05699(new_n6076, new_n6075, new_n6060);
nand_4 g05700(new_n6077, new_n6076, new_n6064);
not_3  g05701(new_n6078, new_n6077);
xnor_3 g05702(new_n6079, new_n6078, new_n6073);
nand_4 g05703(new_n6080, n7891, n2498);
not_3  g05704(new_n6081, new_n6080);
nand_4 g05705(new_n6082, n12391, n5579);
not_3  g05706(new_n6083, new_n6082);
nand_4 g05707(new_n6084, n7160, n2558);
not_3  g05708(new_n6085, new_n6084);
nor_4  g05709(new_n6086, new_n6085, new_n6083);
nor_4  g05710(new_n6087, new_n6084, new_n6082);
nor_4  g05711(new_n6088, new_n6087, new_n6086);
xnor_3 g05712(new_n6089_1, new_n6088, new_n6081);
xnor_3 g05713(new_n6090, new_n6089_1, new_n6079);
nor_4  g05714(new_n6091, new_n6090, new_n6072);
not_3  g05715(new_n6092, new_n6090);
nor_4  g05716(new_n6093, new_n6092, new_n6071);
nor_4  g05717(new_n6094, new_n6093, new_n6091);
nand_4 g05718(new_n6095, n11222, n806);
not_3  g05719(new_n6096, new_n6095);
nand_4 g05720(new_n6097, n11222, n3342);
nand_4 g05721(new_n6098, n9763, n5314);
nand_4 g05722(new_n6099, new_n6098, new_n6097);
not_3  g05723(new_n6100, new_n6099);
nand_4 g05724(new_n6101, n11153, n9111);
not_3  g05725(new_n6102, new_n6101);
nor_4  g05726(new_n6103, new_n6098, new_n6097);
nor_4  g05727(new_n6104, new_n6103, new_n6102);
nor_4  g05728(new_n6105, new_n6104, new_n6100);
nand_4 g05729(new_n6106, new_n6105, new_n6096);
not_3  g05730(new_n6107, new_n6106);
nor_4  g05731(new_n6108, new_n6105, new_n6096);
nor_4  g05732(new_n6109, new_n6108, new_n6107);
nand_4 g05733(new_n6110, n9111, n5314);
nand_4 g05734(new_n6111, n11153, n3342);
nand_4 g05735(new_n6112, n9763, n996);
xnor_3 g05736(new_n6113, new_n6112, new_n6111);
xnor_3 g05737(new_n6114, new_n6113, new_n6110);
not_3  g05738(new_n6115, new_n6114);
xnor_3 g05739(new_n6116, new_n6115, new_n6109);
not_3  g05740(new_n6117, new_n4570);
nor_4  g05741(new_n6118, new_n6101, new_n6117);
nor_4  g05742(new_n6119, new_n6118, new_n6099);
nor_4  g05743(new_n6120, new_n6119, new_n6103);
nor_4  g05744(new_n6121, new_n6120, new_n6101);
not_3  g05745(new_n6122, new_n6121);
nor_4  g05746(new_n6123, new_n6122, new_n6116);
not_3  g05747(new_n6124, new_n6116);
nor_4  g05748(new_n6125, new_n6121, new_n6124);
nor_4  g05749(new_n6126_1, new_n6125, new_n6123);
xnor_3 g05750(new_n6127, new_n6126_1, new_n6094);
not_3  g05751(new_n6128, new_n6127);
nor_4  g05752(new_n6129, new_n4571, new_n4570);
xnor_3 g05753(new_n6130, new_n6068, new_n6067);
not_3  g05754(new_n6131, new_n6130);
nor_4  g05755(new_n6132, new_n6131, new_n6129);
not_3  g05756(new_n6133, new_n6132);
not_3  g05757(new_n6134, new_n6129);
nor_4  g05758(new_n6135, new_n6130, new_n6134);
nor_4  g05759(new_n6136, new_n6135, new_n6132);
nand_4 g05760(new_n6137, n11153, n9763);
nand_4 g05761(new_n6138, n11222, n9111);
xnor_3 g05762(new_n6139, new_n6138, new_n6137);
nand_4 g05763(new_n6140, new_n6139, new_n6136);
nand_4 g05764(new_n6141, new_n6140, new_n6133);
not_3  g05765(new_n6142, new_n6141);
not_3  g05766(new_n6143, new_n6118);
nor_4  g05767(new_n6144, new_n6143, new_n6100);
not_3  g05768(new_n6145, new_n6144);
nand_4 g05769(new_n6146, new_n6145, new_n6120);
not_3  g05770(new_n6147, new_n6146);
nor_4  g05771(new_n6148, new_n6147, new_n6142);
xnor_3 g05772(new_n6149, new_n6146, new_n6141);
not_3  g05773(new_n6150, new_n4571);
nor_4  g05774(new_n6151, new_n6074, new_n6150);
not_3  g05775(new_n6152, new_n6151);
nor_4  g05776(new_n6153, new_n6152, new_n6060);
not_3  g05777(new_n6154, new_n6066);
nor_4  g05778(new_n6155, new_n6151, new_n6154);
nor_4  g05779(new_n6156, new_n6155, new_n6153);
not_3  g05780(new_n6157, new_n6156);
nor_4  g05781(new_n6158, new_n6157, new_n6149);
nor_4  g05782(new_n6159, new_n6158, new_n6148);
not_3  g05783(new_n6160, new_n6159);
nor_4  g05784(new_n6161, new_n6160, new_n6128);
nor_4  g05785(new_n6162, new_n6159, new_n6127);
nor_4  g05786(new_n6163, new_n6162, new_n6161);
not_3  g05787(new_n6164, new_n6163);
nand_4 g05788(new_n6165, new_n6164, new_n6057);
xnor_3 g05789(new_n6166, new_n6163, new_n6057);
xnor_3 g05790(new_n6167, new_n6157, new_n6149);
not_3  g05791(new_n6168, new_n6027);
not_3  g05792(new_n6169, new_n6025);
nor_4  g05793(new_n6170, new_n6169, new_n6007);
nor_4  g05794(new_n6171, new_n6170, new_n6168);
nand_4 g05795(new_n6172, new_n6171, new_n6167);
xnor_3 g05796(new_n6173, new_n6171, new_n6167);
not_3  g05797(new_n6174, new_n6173);
xnor_3 g05798(new_n6175, new_n6139, new_n6136);
not_3  g05799(new_n6176, new_n6175);
nand_4 g05800(new_n6177, n10928, n7946);
nand_4 g05801(new_n6178, n8336, n2024);
xor_3  g05802(new_n6179, new_n6178, new_n6177);
not_3  g05803(new_n6180, new_n6179);
nor_4  g05804(new_n6181, new_n6180, new_n6176);
nand_4 g05805(new_n6182, new_n4572, new_n4569);
xnor_3 g05806(new_n6183, new_n6179, new_n6175);
nor_4  g05807(new_n6184, new_n6183, new_n6182);
nor_4  g05808(new_n6185, new_n6184, new_n6181);
not_3  g05809(new_n6186, new_n6185);
nand_4 g05810(new_n6187, new_n6186, new_n6174);
nand_4 g05811(new_n6188, new_n6187, new_n6172);
nand_4 g05812(new_n6189, new_n6188, new_n6166);
nand_4 g05813(new_n6190, new_n6189, new_n6165);
xnor_3 g05814(new_n6191, new_n6190, new_n6055);
nand_4 g05815(new_n6192_1, n12069, n6016);
nand_4 g05816(new_n6193, n12391, n521);
not_3  g05817(new_n6194, new_n6193);
nor_4  g05818(new_n6195, new_n6087, new_n6081);
nor_4  g05819(new_n6196, new_n6195, new_n6086);
xnor_3 g05820(new_n6197, new_n6196, new_n6194);
nand_4 g05821(new_n6198, n7160, n2498);
nand_4 g05822(new_n6199, n7891, n5579);
nand_4 g05823(new_n6200, n4828, n2558);
xnor_3 g05824(new_n6201, new_n6200, new_n6199);
not_3  g05825(new_n6202, new_n6201);
nor_4  g05826(new_n6203, new_n6202, new_n6198);
not_3  g05827(new_n6204, new_n6198);
nor_4  g05828(new_n6205, new_n6201, new_n6204);
nor_4  g05829(new_n6206, new_n6205, new_n6203);
xnor_3 g05830(new_n6207, new_n6206, new_n6197);
xnor_3 g05831(new_n6208, new_n6207, new_n6192_1);
nor_4  g05832(new_n6209, new_n6078, new_n6073);
nor_4  g05833(new_n6210, new_n6089_1, new_n6079);
nor_4  g05834(new_n6211, new_n6210, new_n6209);
xnor_3 g05835(new_n6212, new_n6211, new_n6208);
not_3  g05836(new_n6213, new_n6212);
xor_3  g05837(new_n6214, new_n6213, new_n6091);
nand_4 g05838(new_n6215, n11222, n7270);
nand_4 g05839(new_n6216, n11153, n806);
not_3  g05840(new_n6217, new_n6216);
not_3  g05841(new_n6218, new_n6111);
not_3  g05842(new_n6219, new_n6112);
nor_4  g05843(new_n6220, new_n6219, new_n6218);
not_3  g05844(new_n6221, new_n6110);
nor_4  g05845(new_n6222, new_n6112, new_n6111);
nor_4  g05846(new_n6223, new_n6222, new_n6221);
nor_4  g05847(new_n6224, new_n6223, new_n6220);
xnor_3 g05848(new_n6225, new_n6224, new_n6217);
nand_4 g05849(new_n6226, n9111, n996);
not_3  g05850(new_n6227, new_n6226);
nand_4 g05851(new_n6228, n5314, n3342);
not_3  g05852(new_n6229, new_n6228);
nand_4 g05853(new_n6230, n9763, n5767);
not_3  g05854(new_n6231, new_n6230);
nor_4  g05855(new_n6232, new_n6231, new_n6229);
nor_4  g05856(new_n6233, new_n6230, new_n6228);
nor_4  g05857(new_n6234, new_n6233, new_n6232);
xnor_3 g05858(new_n6235, new_n6234, new_n6227);
xnor_3 g05859(new_n6236, new_n6235, new_n6225);
nor_4  g05860(new_n6237, new_n6236, new_n6215);
not_3  g05861(new_n6238, new_n6215);
not_3  g05862(new_n6239, new_n6236);
nor_4  g05863(new_n6240, new_n6239, new_n6238);
nor_4  g05864(new_n6241, new_n6240, new_n6237);
nand_4 g05865(new_n6242, new_n6115, new_n6109);
nand_4 g05866(new_n6243, new_n6242, new_n6106);
xnor_3 g05867(new_n6244, new_n6243, new_n6241);
not_3  g05868(new_n6245, new_n6244);
nor_4  g05869(new_n6246, new_n6245, new_n6123);
not_3  g05870(new_n6247, new_n6123);
nor_4  g05871(new_n6248, new_n6244, new_n6247);
nor_4  g05872(new_n6249, new_n6248, new_n6246);
xnor_3 g05873(new_n6250, new_n6249, new_n6214);
nor_4  g05874(new_n6251, new_n6126_1, new_n6094);
nor_4  g05875(new_n6252, new_n6162, new_n6251);
xnor_3 g05876(new_n6253, new_n6252, new_n6250);
xnor_3 g05877(new_n6254_1, new_n6253, new_n6191);
xnor_3 g05878(new_n6255, new_n6254_1, new_n6001);
not_3  g05879(new_n6256, new_n6255);
xor_3  g05880(new_n6257, new_n5971, new_n5955);
not_3  g05881(new_n6258, new_n6257);
xnor_3 g05882(new_n6259, new_n6188, new_n6166);
nand_4 g05883(new_n6260, new_n6259, new_n6258);
xnor_3 g05884(new_n6261, new_n6185, new_n6173);
not_3  g05885(new_n6262, new_n6261);
not_3  g05886(new_n6263, new_n5950);
nor_4  g05887(new_n6264, new_n5958, new_n4567);
not_3  g05888(new_n6265, new_n6264);
nand_4 g05889(new_n6266, new_n6265, new_n6263);
nand_4 g05890(new_n6267, new_n6264, new_n5946);
nand_4 g05891(new_n6268, new_n6267, new_n6266);
not_3  g05892(new_n6269, new_n6268);
nor_4  g05893(new_n6270, new_n6269, new_n6262);
not_3  g05894(new_n6271, new_n6270);
xor_3  g05895(new_n6272, new_n6269, new_n6262);
nand_4 g05896(new_n6273_1, new_n4573, new_n4567);
xor_3  g05897(new_n6274, new_n5952, new_n5951);
not_3  g05898(new_n6275, new_n6274);
nand_4 g05899(new_n6276, new_n6275, new_n6273_1);
not_3  g05900(new_n6277, new_n6183);
xor_3  g05901(new_n6278, new_n6277, new_n6182);
not_3  g05902(new_n6279, new_n6273_1);
xor_3  g05903(new_n6280, new_n6274, new_n6279);
nand_4 g05904(new_n6281, new_n6280, new_n6278);
nand_4 g05905(new_n6282, new_n6281, new_n6276);
nand_4 g05906(new_n6283, new_n6282, new_n6272);
nand_4 g05907(new_n6284, new_n6283, new_n6271);
xnor_3 g05908(new_n6285, new_n6259, new_n6257);
nand_4 g05909(new_n6286, new_n6285, new_n6284);
nand_4 g05910(new_n6287, new_n6286, new_n6260);
xor_3  g05911(n1658, new_n6287, new_n6256);
nand_4 g05912(new_n6289, n7862, n4634);
nand_4 g05913(new_n6290, n10223, n7862);
not_3  g05914(new_n6291, new_n6290);
nand_4 g05915(new_n6292, n7265, n3172);
not_3  g05916(new_n6293, new_n6292);
nor_4  g05917(new_n6294_1, new_n6293, new_n6291);
nor_4  g05918(new_n6295, new_n6292, new_n6290);
nand_4 g05919(new_n6296, n2879, n1333);
not_3  g05920(new_n6297, new_n6296);
nor_4  g05921(new_n6298, new_n6297, new_n6295);
nor_4  g05922(new_n6299, new_n6298, new_n6294_1);
xor_3  g05923(new_n6300, new_n6299, new_n6289);
nand_4 g05924(new_n6301, n3172, n2879);
nand_4 g05925(new_n6302, n10223, n1333);
not_3  g05926(new_n6303, new_n6302);
nand_4 g05927(new_n6304, n11757, n7265);
not_3  g05928(new_n6305, new_n6304);
nor_4  g05929(new_n6306, new_n6305, new_n6303);
nor_4  g05930(new_n6307, new_n6304, new_n6302);
nor_4  g05931(new_n6308, new_n6307, new_n6306);
xor_3  g05932(new_n6309, new_n6308, new_n6301);
xnor_3 g05933(new_n6310, new_n6309, new_n6300);
not_3  g05934(new_n6311, new_n6310);
nand_4 g05935(new_n6312, n7862, n7265);
not_3  g05936(new_n6313, new_n6312);
nor_4  g05937(new_n6314, new_n6313, new_n6296);
nor_4  g05938(new_n6315, new_n6295, new_n6294_1);
nor_4  g05939(new_n6316, new_n6315, new_n6314);
not_3  g05940(new_n6317, new_n6316);
nor_4  g05941(new_n6318, new_n6317, new_n6296);
xor_3  g05942(new_n6319, new_n6318, new_n6311);
nand_4 g05943(new_n6320, n6877, n2522);
nand_4 g05944(new_n6321, n2464, n2024);
nand_4 g05945(new_n6322, n9400, n9189);
nand_4 g05946(new_n6323, n11311, n7946);
xnor_3 g05947(new_n6324, new_n6323, new_n6322);
not_3  g05948(new_n6325, new_n6324);
nor_4  g05949(new_n6326, new_n6325, new_n6321);
not_3  g05950(new_n6327, new_n6321);
nor_4  g05951(new_n6328, new_n6324, new_n6327);
nor_4  g05952(new_n6329, new_n6328, new_n6326);
xnor_3 g05953(new_n6330, new_n6329, new_n6320);
nand_4 g05954(new_n6331, n9189, n6877);
not_3  g05955(new_n6332, new_n6331);
nand_4 g05956(new_n6333, n7946, n2464);
not_3  g05957(new_n6334, new_n6333);
nor_4  g05958(new_n6335, new_n6334, new_n6332);
nor_4  g05959(new_n6336, new_n6333, new_n6331);
nand_4 g05960(new_n6337, n9400, n2024);
not_3  g05961(new_n6338, new_n6337);
nor_4  g05962(new_n6339, new_n6338, new_n6336);
nor_4  g05963(new_n6340, new_n6339, new_n6335);
not_3  g05964(new_n6341, new_n6340);
nor_4  g05965(new_n6342, new_n6341, new_n6330);
not_3  g05966(new_n6343, new_n6330);
nor_4  g05967(new_n6344, new_n6340, new_n6343);
nor_4  g05968(new_n6345, new_n6344, new_n6342);
not_3  g05969(new_n6346, new_n6345);
nand_4 g05970(new_n6347, n7946, n6877);
not_3  g05971(new_n6348, new_n6347);
nor_4  g05972(new_n6349, new_n6348, new_n6337);
nor_4  g05973(new_n6350, new_n6336, new_n6335);
nor_4  g05974(new_n6351, new_n6350, new_n6349);
not_3  g05975(new_n6352, new_n6351);
nor_4  g05976(new_n6353, new_n6352, new_n6337);
not_3  g05977(new_n6354, new_n6353);
nor_4  g05978(new_n6355, new_n6354, new_n6346);
nor_4  g05979(new_n6356, new_n6353, new_n6345);
nor_4  g05980(new_n6357, new_n6356, new_n6355);
not_3  g05981(new_n6358_1, new_n6357);
nand_4 g05982(new_n6359_1, n4805, n2558);
nand_4 g05983(new_n6360, n9763, n7236);
xnor_3 g05984(new_n6361, new_n6360, new_n6359_1);
nor_4  g05985(new_n6362, new_n6361, new_n6347);
not_3  g05986(new_n6363, new_n6362);
nand_4 g05987(new_n6364, n9400, n7946);
nand_4 g05988(new_n6365, n6877, n2024);
not_3  g05989(new_n6366, new_n6365);
xnor_3 g05990(new_n6367, new_n6366, new_n6364);
not_3  g05991(new_n6368, new_n6367);
nor_4  g05992(new_n6369, new_n6368, new_n6363);
not_3  g05993(new_n6370, new_n6369);
nor_4  g05994(new_n6371, new_n6360, new_n6359_1);
nand_4 g05995(new_n6372, n9111, n7236);
nand_4 g05996(new_n6373, n9763, n3992);
xnor_3 g05997(new_n6374, new_n6373, new_n6372);
xnor_3 g05998(new_n6375, new_n6374, new_n6371);
nand_4 g05999(new_n6376, n4805, n2498);
nand_4 g06000(new_n6377, n11478, n2558);
not_3  g06001(new_n6378, new_n6377);
xnor_3 g06002(new_n6379, new_n6378, new_n6376);
not_3  g06003(new_n6380, new_n6379);
xnor_3 g06004(new_n6381, new_n6380, new_n6375);
nor_4  g06005(new_n6382, new_n6367, new_n6362);
nor_4  g06006(new_n6383, new_n6382, new_n6369);
nand_4 g06007(new_n6384, new_n6383, new_n6381);
nand_4 g06008(new_n6385, new_n6384, new_n6370);
not_3  g06009(new_n6386, new_n6335);
nand_4 g06010(new_n6387, new_n6349, new_n6386);
nand_4 g06011(new_n6388, new_n6387, new_n6352);
not_3  g06012(new_n6389, new_n6388);
nor_4  g06013(new_n6390, new_n6389, new_n6385);
not_3  g06014(new_n6391, new_n6390);
not_3  g06015(new_n6392, new_n6374);
nor_4  g06016(new_n6393, new_n6392, new_n6371);
not_3  g06017(new_n6394, new_n6393);
nand_4 g06018(new_n6395, new_n6380, new_n6375);
nand_4 g06019(new_n6396, new_n6395, new_n6394);
not_3  g06020(new_n6397, new_n6359_1);
nand_4 g06021(new_n6398, n11478, n2498);
nor_4  g06022(new_n6399, new_n6398, new_n6397);
not_3  g06023(new_n6400, new_n6399);
nand_4 g06024(new_n6401, n5283, n2558);
nand_4 g06025(new_n6402, n5579, n4805);
nand_4 g06026(new_n6403, new_n6402, new_n6401);
not_3  g06027(new_n6404, new_n6403);
nor_4  g06028(new_n6405, new_n6404, new_n6400);
not_3  g06029(new_n6406, new_n6405);
not_3  g06030(new_n6407, new_n6401);
not_3  g06031(new_n6408, new_n6402);
nand_4 g06032(new_n6409, new_n6408, new_n6407);
not_3  g06033(new_n6410, new_n6409);
nor_4  g06034(new_n6411, new_n6403, new_n6399);
nor_4  g06035(new_n6412, new_n6411, new_n6410);
nand_4 g06036(new_n6413, new_n6412, new_n6406);
xnor_3 g06037(new_n6414, new_n6413, new_n6396);
not_3  g06038(new_n6415, new_n6360);
nand_4 g06039(new_n6416, n9111, n3992);
nor_4  g06040(new_n6417, new_n6416, new_n6415);
not_3  g06041(new_n6418, new_n6417);
nand_4 g06042(new_n6419, n9763, n8384);
nand_4 g06043(new_n6420, n7236, n3342);
nand_4 g06044(new_n6421, new_n6420, new_n6419);
nor_4  g06045(new_n6422, new_n6421, new_n6418);
not_3  g06046(new_n6423, new_n6421);
not_3  g06047(new_n6424, new_n6419);
not_3  g06048(new_n6425, new_n6420);
nand_4 g06049(new_n6426, new_n6425, new_n6424);
not_3  g06050(new_n6427, new_n6426);
nor_4  g06051(new_n6428, new_n6427, new_n6423);
not_3  g06052(new_n6429_1, new_n6428);
nor_4  g06053(new_n6430, new_n6429_1, new_n6417);
nor_4  g06054(new_n6431_1, new_n6430, new_n6422);
not_3  g06055(new_n6432, new_n6431_1);
nor_4  g06056(new_n6433, new_n6432, new_n6414);
not_3  g06057(new_n6434, new_n6414);
nor_4  g06058(new_n6435, new_n6431_1, new_n6434);
nor_4  g06059(new_n6436, new_n6435, new_n6433);
not_3  g06060(new_n6437, new_n6385);
nor_4  g06061(new_n6438, new_n6388, new_n6437);
nor_4  g06062(new_n6439, new_n6438, new_n6390);
nand_4 g06063(new_n6440, new_n6439, new_n6436);
nand_4 g06064(new_n6441_1, new_n6440, new_n6391);
nor_4  g06065(new_n6442, new_n6441_1, new_n6358_1);
not_3  g06066(new_n6443, new_n6441_1);
nor_4  g06067(new_n6444, new_n6443, new_n6357);
nor_4  g06068(new_n6445_1, new_n6444, new_n6442);
nand_4 g06069(new_n6446, n4805, n521);
not_3  g06070(new_n6447, new_n6398);
nand_4 g06071(new_n6448, new_n6403, new_n6447);
nand_4 g06072(new_n6449, new_n6448, new_n6409);
not_3  g06073(new_n6450, new_n6449);
nor_4  g06074(new_n6451, new_n6450, new_n6446);
not_3  g06075(new_n6452, new_n6446);
nor_4  g06076(new_n6453, new_n6449, new_n6452);
nor_4  g06077(new_n6454, new_n6453, new_n6451);
nand_4 g06078(new_n6455, n5283, n2498);
nand_4 g06079(new_n6456, n2558, n137);
nand_4 g06080(new_n6457, n11478, n5579);
xnor_3 g06081(new_n6458, new_n6457, new_n6456);
xnor_3 g06082(new_n6459, new_n6458, new_n6455);
not_3  g06083(new_n6460, new_n6459);
xnor_3 g06084(new_n6461, new_n6460, new_n6454);
not_3  g06085(new_n6462, new_n6461);
nor_4  g06086(new_n6463, new_n6412, new_n6398);
nor_4  g06087(new_n6464, new_n6463, new_n6462);
not_3  g06088(new_n6465, new_n6463);
nor_4  g06089(new_n6466, new_n6465, new_n6461);
nor_4  g06090(new_n6467, new_n6466, new_n6464);
nand_4 g06091(new_n6468, n7236, n806);
not_3  g06092(new_n6469, new_n6416);
nand_4 g06093(new_n6470, new_n6421, new_n6469);
nand_4 g06094(new_n6471, new_n6470, new_n6426);
not_3  g06095(new_n6472, new_n6471);
nor_4  g06096(new_n6473, new_n6472, new_n6468);
not_3  g06097(new_n6474, new_n6468);
nor_4  g06098(new_n6475, new_n6471, new_n6474);
nor_4  g06099(new_n6476, new_n6475, new_n6473);
nand_4 g06100(new_n6477, n9111, n8384);
nand_4 g06101(new_n6478, n9763, n6358);
nand_4 g06102(new_n6479, n3992, n3342);
xnor_3 g06103(new_n6480, new_n6479, new_n6478);
xnor_3 g06104(new_n6481, new_n6480, new_n6477);
not_3  g06105(new_n6482, new_n6481);
xnor_3 g06106(new_n6483, new_n6482, new_n6476);
not_3  g06107(new_n6484, new_n6483);
nor_4  g06108(new_n6485, new_n6373, new_n6372);
not_3  g06109(new_n6486, new_n6485);
nor_4  g06110(new_n6487, new_n6428, new_n6486);
nor_4  g06111(new_n6488, new_n6487, new_n6484);
not_3  g06112(new_n6489, new_n6487);
nor_4  g06113(new_n6490, new_n6489, new_n6483);
nor_4  g06114(new_n6491, new_n6490, new_n6488);
xnor_3 g06115(new_n6492, new_n6491, new_n6467);
and_4  g06116(new_n6493, new_n6413, new_n6396);
nor_4  g06117(new_n6494, new_n6433, new_n6493);
xnor_3 g06118(new_n6495, new_n6494, new_n6492);
nor_4  g06119(new_n6496, new_n6495, new_n6445_1);
nand_4 g06120(new_n6497, new_n6495, new_n6445_1);
not_3  g06121(new_n6498, new_n6497);
nor_4  g06122(new_n6499, new_n6498, new_n6496);
nor_4  g06123(new_n6500, new_n6499, new_n6319);
not_3  g06124(new_n6501, new_n6500);
nand_4 g06125(new_n6502, new_n6499, new_n6319);
nand_4 g06126(new_n6503, new_n6502, new_n6501);
not_3  g06127(new_n6504, new_n6440);
nor_4  g06128(new_n6505, new_n6439, new_n6436);
nor_4  g06129(new_n6506, new_n6505, new_n6504);
not_3  g06130(new_n6507, new_n6314);
nor_4  g06131(new_n6508, new_n6507, new_n6294_1);
or_4   g06132(new_n6509, new_n6508, new_n6316);
nor_4  g06133(new_n6510, new_n6509, new_n6506);
xor_3  g06134(new_n6511, new_n6361, new_n6347);
nand_4 g06135(new_n6512, new_n6511, new_n6313);
not_3  g06136(new_n6513, new_n6512);
nand_4 g06137(new_n6514, n7265, n1333);
nand_4 g06138(new_n6515, n7862, n2879);
xor_3  g06139(new_n6516, new_n6515, new_n6514);
nor_4  g06140(new_n6517, new_n6516, new_n6513);
not_3  g06141(new_n6518, new_n6517);
not_3  g06142(new_n6519, new_n6381);
xor_3  g06143(new_n6520, new_n6383, new_n6519);
xor_3  g06144(new_n6521, new_n6516, new_n6513);
nand_4 g06145(new_n6522, new_n6521, new_n6520);
nand_4 g06146(new_n6523, new_n6522, new_n6518);
xnor_3 g06147(new_n6524, new_n6509, new_n6506);
nor_4  g06148(new_n6525, new_n6524, new_n6523);
nor_4  g06149(new_n6526, new_n6525, new_n6510);
xor_3  g06150(n1847, new_n6526, new_n6503);
nand_4 g06151(new_n6528, n5305, n1798);
nand_4 g06152(new_n6529, n8759, n6703);
not_3  g06153(new_n6530, new_n6529);
nand_4 g06154(new_n6531, n5645, n5331);
nand_4 g06155(new_n6532, n11876, n7965);
xor_3  g06156(new_n6533, new_n6532, new_n6531);
not_3  g06157(new_n6534, new_n6533);
xor_3  g06158(new_n6535, new_n6534, new_n6530);
nor_4  g06159(new_n6536, new_n6535, new_n6528);
nand_4 g06160(new_n6537, n5305, n3932);
nand_4 g06161(new_n6538, n5964, n1798);
xor_3  g06162(new_n6539, new_n6538, new_n6537);
xor_3  g06163(new_n6540, new_n6539, new_n6536);
nor_4  g06164(new_n6541, new_n6534, new_n6529);
nand_4 g06165(new_n6542, n9640, n8759);
nand_4 g06166(new_n6543, n6776, n6703);
xor_3  g06167(new_n6544, new_n6543, new_n6542);
xnor_3 g06168(new_n6545, new_n6544, new_n6541);
nor_4  g06169(new_n6546, new_n6532, new_n6531);
not_3  g06170(new_n6547, new_n6546);
nand_4 g06171(new_n6548, n10898, n7965);
nand_4 g06172(new_n6549, n11876, n7388);
xnor_3 g06173(new_n6550, new_n6549, new_n6548);
nor_4  g06174(new_n6551, new_n6550, new_n6547);
not_3  g06175(new_n6552, new_n6550);
nor_4  g06176(new_n6553, new_n6552, new_n6546);
nor_4  g06177(new_n6554, new_n6553, new_n6551);
nand_4 g06178(new_n6555, n5331, n1067);
nand_4 g06179(new_n6556, n8476, n5645);
xor_3  g06180(new_n6557, new_n6556, new_n6555);
xnor_3 g06181(new_n6558, new_n6557, new_n6554);
nor_4  g06182(new_n6559, new_n6558, new_n6545);
and_4  g06183(new_n6560, new_n6558, new_n6545);
nor_4  g06184(new_n6561, new_n6560, new_n6559);
xor_3  g06185(n2096, new_n6561, new_n6540);
xor_3  g06186(n2131, new_n3840, new_n3801);
nand_4 g06187(new_n6564, n7456, n2564);
not_3  g06188(new_n6565, new_n6564);
not_3  g06189(new_n6566, new_n4009);
nor_4  g06190(new_n6567, new_n4015, new_n6566);
nor_4  g06191(new_n6568, new_n6567, new_n4014);
nand_4 g06192(new_n6569, new_n6568, new_n6565);
xnor_3 g06193(new_n6570, new_n6568, new_n6564);
nand_4 g06194(new_n6571, n6770, n3932);
nand_4 g06195(new_n6572, n12591, n4189);
not_3  g06196(new_n6573, new_n6572);
nand_4 g06197(new_n6574, n9920, n1798);
not_3  g06198(new_n6575, new_n6574);
nor_4  g06199(new_n6576, new_n6575, new_n6573);
nor_4  g06200(new_n6577, new_n6574, new_n6572);
nor_4  g06201(new_n6578_1, new_n6577, new_n6576);
xnor_3 g06202(new_n6579, new_n6578_1, new_n6571);
nand_4 g06203(new_n6580, new_n6579, new_n6570);
nand_4 g06204(new_n6581, new_n6580, new_n6569);
nand_4 g06205(new_n6582, n11662, n2564);
nand_4 g06206(new_n6583, n7456, n4189);
xor_3  g06207(new_n6584, new_n6583, new_n6582);
xnor_3 g06208(new_n6585, new_n6584, new_n6581);
nand_4 g06209(new_n6586, n12591, n6770);
not_3  g06210(new_n6587, new_n6586);
nand_4 g06211(new_n6588, n3627, n1798);
nand_4 g06212(new_n6589, n9920, n3932);
xor_3  g06213(new_n6590, new_n6589, new_n6588);
xnor_3 g06214(new_n6591, new_n6590, new_n6587);
not_3  g06215(new_n6592, new_n6591);
not_3  g06216(new_n6593, new_n6571);
nor_4  g06217(new_n6594, new_n6577, new_n6593);
nor_4  g06218(new_n6595, new_n6594, new_n6576);
not_3  g06219(new_n6596, new_n6595);
xor_3  g06220(new_n6597, new_n6596, new_n6592);
xnor_3 g06221(new_n6598, new_n6597, new_n6585);
not_3  g06222(new_n6599, new_n6598);
nand_4 g06223(new_n6600, n11662, n6687);
not_3  g06224(new_n6601, new_n6600);
nand_4 g06225(new_n6602, new_n4017, new_n4008);
nand_4 g06226(new_n6603, new_n6602, new_n4005_1);
nor_4  g06227(new_n6604_1, new_n6603, new_n6601);
not_3  g06228(new_n6605, new_n6604_1);
not_3  g06229(new_n6606, new_n6570);
xor_3  g06230(new_n6607, new_n6579, new_n6606);
not_3  g06231(new_n6608, new_n6603);
nor_4  g06232(new_n6609, new_n6608, new_n6600);
nor_4  g06233(new_n6610, new_n6609, new_n6604_1);
nand_4 g06234(new_n6611_1, new_n6610, new_n6607);
nand_4 g06235(new_n6612, new_n6611_1, new_n6605);
not_3  g06236(new_n6613, new_n6612);
nand_4 g06237(new_n6614, new_n6613, new_n6599);
nand_4 g06238(new_n6615, new_n6590, new_n6587);
not_3  g06239(new_n6616, new_n6615);
nor_4  g06240(new_n6617, new_n6596, new_n6591);
nor_4  g06241(new_n6618, new_n6617, new_n6616);
not_3  g06242(new_n6619, new_n6618);
nand_4 g06243(new_n6620, n10327, n2564);
nand_4 g06244(new_n6621, n11662, n4189);
nand_4 g06245(new_n6622, n9583, n6687);
not_3  g06246(new_n6623, new_n6622);
xor_3  g06247(new_n6624, new_n6623, new_n6621);
xnor_3 g06248(new_n6625, new_n6624, new_n6620);
xnor_3 g06249(new_n6626, new_n6625, new_n6619);
nor_4  g06250(new_n6627, new_n6589, new_n6588);
nand_4 g06251(new_n6628, n7456, n6770);
not_3  g06252(new_n6629, new_n6628);
xor_3  g06253(new_n6630, new_n6629, new_n6627);
nand_4 g06254(new_n6631, n3932, n3627);
nand_4 g06255(new_n6632, n12591, n9920);
nand_4 g06256(new_n6633, n4516, n1798);
nand_4 g06257(new_n6634, new_n6633, new_n6632);
not_3  g06258(new_n6635, new_n6632);
not_3  g06259(new_n6636, new_n6633);
nand_4 g06260(new_n6637, new_n6636, new_n6635);
nand_4 g06261(new_n6638, new_n6637, new_n6634);
xor_3  g06262(new_n6639, new_n6638, new_n6631);
xnor_3 g06263(new_n6640, new_n6639, new_n6630);
not_3  g06264(new_n6641, new_n6640);
xnor_3 g06265(new_n6642, new_n6641, new_n6626);
nand_4 g06266(new_n6643, new_n6584, new_n6581);
nor_4  g06267(new_n6644, new_n6583, new_n6582);
nor_4  g06268(new_n6645_1, new_n6597, new_n6585);
xnor_3 g06269(new_n6646, new_n6645_1, new_n6644);
nand_4 g06270(new_n6647, new_n6646, new_n6643);
xnor_3 g06271(new_n6648, new_n6647, new_n6642);
xnor_3 g06272(new_n6649, new_n6648, new_n6614);
nand_4 g06273(new_n6650, n10327, n6687);
not_3  g06274(new_n6651, new_n6650);
xnor_3 g06275(new_n6652, new_n6612, new_n6598);
not_3  g06276(new_n6653, new_n6652);
nand_4 g06277(new_n6654, new_n6653, new_n6651);
nor_4  g06278(new_n6655, new_n4027, new_n4019);
not_3  g06279(new_n6656, new_n6655);
not_3  g06280(new_n6657, new_n6611_1);
nor_4  g06281(new_n6658, new_n6610, new_n6607);
nor_4  g06282(new_n6659, new_n6658, new_n6657);
nor_4  g06283(new_n6660, new_n6659, new_n6656);
nor_4  g06284(new_n6661, new_n6652, new_n6650);
nor_4  g06285(new_n6662, new_n6653, new_n6651);
nor_4  g06286(new_n6663, new_n6662, new_n6661);
nand_4 g06287(new_n6664, new_n6663, new_n6660);
nand_4 g06288(new_n6665, new_n6664, new_n6654);
xnor_3 g06289(new_n6666, new_n6665, new_n6649);
nand_4 g06290(new_n6667, n3022, n2226);
nand_4 g06291(new_n6668, n9640, n1094);
nand_4 g06292(new_n6669, n10678, n6703);
xnor_3 g06293(new_n6670, new_n6669, new_n6668);
nor_4  g06294(new_n6671, new_n6670, new_n6667);
not_3  g06295(new_n6672, new_n6667);
not_3  g06296(new_n6673, new_n6670);
nor_4  g06297(new_n6674, new_n6673, new_n6672);
nor_4  g06298(new_n6675, new_n6674, new_n6671);
nand_4 g06299(new_n6676, n6986, n3022);
not_3  g06300(new_n6677, new_n6676);
nand_4 g06301(new_n6678, n6703, n1094);
not_3  g06302(new_n6679, new_n6678);
nor_4  g06303(new_n6680, new_n6679, new_n6677);
nor_4  g06304(new_n6681, new_n6678, new_n6676);
nand_4 g06305(new_n6682, n9640, n2226);
not_3  g06306(new_n6683, new_n6682);
nor_4  g06307(new_n6684, new_n6683, new_n6681);
nor_4  g06308(new_n6685, new_n6684, new_n6680);
xnor_3 g06309(new_n6686, new_n6685, new_n6675);
nand_4 g06310(new_n6687_1, n10928, n10451);
nand_4 g06311(new_n6688, n11023, n6986);
xor_3  g06312(new_n6689_1, new_n6688, new_n6687_1);
xnor_3 g06313(new_n6690, new_n6689_1, new_n6686);
nand_4 g06314(new_n6691, n11023, n10928);
not_3  g06315(new_n6692, new_n6691);
nor_4  g06316(new_n6693, new_n4198, new_n4192);
nor_4  g06317(new_n6694, new_n6693, new_n4197);
nand_4 g06318(new_n6695, new_n6694, new_n6692);
xor_3  g06319(new_n6696, new_n6694, new_n6692);
nor_4  g06320(new_n6697, new_n6681, new_n6680);
xor_3  g06321(new_n6698, new_n6697, new_n6683);
nand_4 g06322(new_n6699, new_n6698, new_n6696);
nand_4 g06323(new_n6700, new_n6699, new_n6695);
xnor_3 g06324(new_n6701, new_n6700, new_n6690);
not_3  g06325(new_n6702, new_n6701);
nand_4 g06326(new_n6703_1, n10451, n8336);
not_3  g06327(new_n6704, new_n6703_1);
xor_3  g06328(new_n6705, new_n6694, new_n6691);
xor_3  g06329(new_n6706, new_n6697, new_n6682);
nor_4  g06330(new_n6707, new_n6706, new_n6705);
nor_4  g06331(new_n6708, new_n6698, new_n6696);
nor_4  g06332(new_n6709, new_n6708, new_n6707);
nand_4 g06333(new_n6710, new_n6709, new_n6704);
nor_4  g06334(new_n6711, new_n4189_1, new_n4184);
not_3  g06335(new_n6712, new_n6711);
nand_4 g06336(new_n6713, new_n4200, new_n4190_1);
nand_4 g06337(new_n6714, new_n6713, new_n6712);
xnor_3 g06338(new_n6715, new_n6706, new_n6705);
xnor_3 g06339(new_n6716, new_n6715, new_n6704);
nand_4 g06340(new_n6717, new_n6716, new_n6714);
nand_4 g06341(new_n6718, new_n6717, new_n6710);
nand_4 g06342(new_n6719, new_n6718, new_n6702);
nand_4 g06343(new_n6720, new_n6685, new_n6675);
not_3  g06344(new_n6721, new_n6720);
nor_4  g06345(new_n6722, new_n6721, new_n6671);
not_3  g06346(new_n6723, new_n6722);
nand_4 g06347(new_n6724, n10928, n10278);
nand_4 g06348(new_n6725, n10451, n6986);
nand_4 g06349(new_n6726, n11423, n8336);
not_3  g06350(new_n6727, new_n6726);
xor_3  g06351(new_n6728, new_n6727, new_n6725);
xnor_3 g06352(new_n6729, new_n6728, new_n6724);
xnor_3 g06353(new_n6730, new_n6729, new_n6723);
nor_4  g06354(new_n6731, new_n6669, new_n6668);
not_3  g06355(new_n6732, new_n6731);
nand_4 g06356(new_n6733, n11023, n2226);
xor_3  g06357(new_n6734, new_n6733, new_n6732);
not_3  g06358(new_n6735, new_n6734);
nand_4 g06359(new_n6736, n10678, n9640);
nand_4 g06360(new_n6737, n3022, n1094);
nand_4 g06361(new_n6738, n7320, n6703);
not_3  g06362(new_n6739, new_n6738);
xor_3  g06363(new_n6740, new_n6739, new_n6737);
xnor_3 g06364(new_n6741, new_n6740, new_n6736);
xnor_3 g06365(new_n6742_1, new_n6741, new_n6735);
xnor_3 g06366(new_n6743, new_n6742_1, new_n6730);
not_3  g06367(new_n6744, new_n6743);
not_3  g06368(new_n6745, new_n6686);
nand_4 g06369(new_n6746, new_n6689_1, new_n6745);
nor_4  g06370(new_n6747, new_n6688, new_n6687_1);
nand_4 g06371(new_n6748, new_n6700, new_n6690);
not_3  g06372(new_n6749, new_n6748);
xnor_3 g06373(new_n6750, new_n6749, new_n6747);
nand_4 g06374(new_n6751, new_n6750, new_n6746);
xnor_3 g06375(new_n6752, new_n6751, new_n6744);
xnor_3 g06376(new_n6753, new_n6752, new_n6719);
nand_4 g06377(new_n6754, n10278, n8336);
not_3  g06378(new_n6755, new_n6754);
xnor_3 g06379(new_n6756, new_n6718, new_n6701);
nor_4  g06380(new_n6757, new_n6756, new_n6755);
not_3  g06381(new_n6758, new_n4203_1);
nor_4  g06382(new_n6759, new_n6758, new_n4201);
not_3  g06383(new_n6760, new_n6759);
xnor_3 g06384(new_n6761, new_n6716, new_n6714);
nor_4  g06385(new_n6762, new_n6761, new_n6760);
not_3  g06386(new_n6763, new_n6756);
xor_3  g06387(new_n6764, new_n6763, new_n6755);
nor_4  g06388(new_n6765, new_n6764, new_n6762);
nor_4  g06389(new_n6766, new_n6765, new_n6757);
not_3  g06390(new_n6767, new_n6766);
xnor_3 g06391(new_n6768, new_n6767, new_n6753);
nand_4 g06392(new_n6769, n8665, n7160);
nand_4 g06393(new_n6770_1, n4828, n1067);
nand_4 g06394(new_n6771, n5645, n2515);
xnor_3 g06395(new_n6772, new_n6771, new_n6770_1);
nor_4  g06396(new_n6773, new_n6772, new_n6769);
not_3  g06397(new_n6774, new_n6769);
not_3  g06398(new_n6775, new_n6772);
nor_4  g06399(new_n6776_1, new_n6775, new_n6774);
nor_4  g06400(new_n6777, new_n6776_1, new_n6773);
nand_4 g06401(new_n6778, n8665, n7891);
nand_4 g06402(new_n6779, n5645, n4828);
and_4  g06403(new_n6780, new_n6779, new_n6778);
nand_4 g06404(new_n6781, n7160, n1067);
not_3  g06405(new_n6782, new_n6781);
xnor_3 g06406(new_n6783, new_n6779, new_n6778);
nor_4  g06407(new_n6784, new_n6783, new_n6782);
nor_4  g06408(new_n6785, new_n6784, new_n6780);
xnor_3 g06409(new_n6786, new_n6785, new_n6777);
nand_4 g06410(new_n6787, n12391, n2551);
nand_4 g06411(new_n6788, n11922, n7891);
not_3  g06412(new_n6789, new_n6788);
xor_3  g06413(new_n6790, new_n6789, new_n6787);
xnor_3 g06414(new_n6791, new_n6790, new_n6786);
nand_4 g06415(new_n6792, n12391, n11922);
not_3  g06416(new_n6793, new_n4136);
nand_4 g06417(new_n6794, new_n4139, new_n6793);
nand_4 g06418(new_n6795, new_n6794, new_n4141_1);
not_3  g06419(new_n6796, new_n6795);
nor_4  g06420(new_n6797_1, new_n6796, new_n6792);
xnor_3 g06421(new_n6798, new_n6783, new_n6781);
xnor_3 g06422(new_n6799, new_n6796, new_n6792);
nor_4  g06423(new_n6800, new_n6799, new_n6798);
nor_4  g06424(new_n6801, new_n6800, new_n6797_1);
xnor_3 g06425(new_n6802, new_n6801, new_n6791);
nand_4 g06426(new_n6803, n12069, n2551);
xnor_3 g06427(new_n6804, new_n6799, new_n6798);
nor_4  g06428(new_n6805, new_n6804, new_n6803);
not_3  g06429(new_n6806_1, new_n6805);
nand_4 g06430(new_n6807, new_n6804, new_n6803);
nand_4 g06431(new_n6808, new_n4134, new_n4129);
nor_4  g06432(new_n6809_1, new_n4143, new_n4135);
not_3  g06433(new_n6810, new_n6809_1);
nand_4 g06434(new_n6811, new_n6810, new_n6808);
nand_4 g06435(new_n6812, new_n6811, new_n6807);
nand_4 g06436(new_n6813, new_n6812, new_n6806_1);
not_3  g06437(new_n6814, new_n6813);
nor_4  g06438(new_n6815, new_n6814, new_n6802);
not_3  g06439(new_n6816, new_n6815);
nand_4 g06440(new_n6817, new_n6785, new_n6777);
not_3  g06441(new_n6818, new_n6817);
nor_4  g06442(new_n6819, new_n6818, new_n6773);
not_3  g06443(new_n6820, new_n6819);
nand_4 g06444(new_n6821, n12826, n12391);
nand_4 g06445(new_n6822_1, n7891, n2551);
nand_4 g06446(new_n6823, n12069, n4094);
not_3  g06447(new_n6824, new_n6823);
xor_3  g06448(new_n6825, new_n6824, new_n6822_1);
xnor_3 g06449(new_n6826_1, new_n6825, new_n6821);
xnor_3 g06450(new_n6827, new_n6826_1, new_n6820);
nor_4  g06451(new_n6828, new_n6771, new_n6770_1);
not_3  g06452(new_n6829, new_n6828);
nand_4 g06453(new_n6830, n11922, n7160);
xor_3  g06454(new_n6831, new_n6830, new_n6829);
nand_4 g06455(new_n6832, n2515, n1067);
not_3  g06456(new_n6833, new_n6832);
nand_4 g06457(new_n6834, n8665, n4828);
nand_4 g06458(new_n6835, n5645, n1199);
xor_3  g06459(new_n6836, new_n6835, new_n6834);
xnor_3 g06460(new_n6837, new_n6836, new_n6833);
xnor_3 g06461(new_n6838, new_n6837, new_n6831);
xnor_3 g06462(new_n6839, new_n6838, new_n6827);
not_3  g06463(new_n6840, new_n6786);
not_3  g06464(new_n6841, new_n6790);
nand_4 g06465(new_n6842, new_n6841, new_n6840);
nor_4  g06466(new_n6843, new_n6788, new_n6787);
nor_4  g06467(new_n6844, new_n6801, new_n6791);
xnor_3 g06468(new_n6845, new_n6844, new_n6843);
nand_4 g06469(new_n6846, new_n6845, new_n6842);
xnor_3 g06470(new_n6847, new_n6846, new_n6839);
xnor_3 g06471(new_n6848, new_n6847, new_n6816);
nand_4 g06472(new_n6849, n12826, n12069);
not_3  g06473(new_n6850, new_n6849);
not_3  g06474(new_n6851, new_n6802);
nor_4  g06475(new_n6852, new_n6813, new_n6851);
nor_4  g06476(new_n6853, new_n6852, new_n6815);
nor_4  g06477(new_n6854, new_n6853, new_n6850);
nand_4 g06478(new_n6855, new_n4170, new_n4127);
not_3  g06479(new_n6856, new_n6807);
nor_4  g06480(new_n6857, new_n6856, new_n6805);
xnor_3 g06481(new_n6858, new_n6857, new_n6811);
nor_4  g06482(new_n6859, new_n6858, new_n6855);
xnor_3 g06483(new_n6860_1, new_n6853, new_n6850);
nor_4  g06484(new_n6861, new_n6860_1, new_n6859);
nor_4  g06485(new_n6862, new_n6861, new_n6854);
xnor_3 g06486(new_n6863, new_n6862, new_n6848);
nand_4 g06487(new_n6864, n3754, n996);
nand_4 g06488(new_n6865, n10898, n5767);
nand_4 g06489(new_n6866, n11876, n5319);
xnor_3 g06490(new_n6867, new_n6866, new_n6865);
nor_4  g06491(new_n6868, new_n6867, new_n6864);
not_3  g06492(new_n6869, new_n6864);
not_3  g06493(new_n6870, new_n6867);
nor_4  g06494(new_n6871, new_n6870, new_n6869);
nor_4  g06495(new_n6872, new_n6871, new_n6868);
nand_4 g06496(new_n6873, n5314, n3754);
nand_4 g06497(new_n6874, n10898, n996);
and_4  g06498(new_n6875, new_n6874, new_n6873);
nand_4 g06499(new_n6876, n11876, n5767);
not_3  g06500(new_n6877_1, new_n6876);
xnor_3 g06501(new_n6878, new_n6874, new_n6873);
nor_4  g06502(new_n6879, new_n6878, new_n6877_1);
nor_4  g06503(new_n6880, new_n6879, new_n6875);
xnor_3 g06504(new_n6881, new_n6880, new_n6872);
nand_4 g06505(new_n6882, n11153, n159);
nand_4 g06506(new_n6883, n5314, n2749);
not_3  g06507(new_n6884, new_n6883);
xor_3  g06508(new_n6885, new_n6884, new_n6882);
xnor_3 g06509(new_n6886, new_n6885, new_n6881);
nand_4 g06510(new_n6887, n11153, n2749);
not_3  g06511(new_n6888, new_n6887);
not_3  g06512(new_n6889, new_n4152);
nor_4  g06513(new_n6890, new_n4158, new_n6889);
nor_4  g06514(new_n6891, new_n6890, new_n4157);
and_4  g06515(new_n6892, new_n6891, new_n6888);
xnor_3 g06516(new_n6893, new_n6891, new_n6887);
not_3  g06517(new_n6894, new_n6893);
xnor_3 g06518(new_n6895, new_n6878, new_n6876);
nor_4  g06519(new_n6896, new_n6895, new_n6894);
nor_4  g06520(new_n6897, new_n6896, new_n6892);
xnor_3 g06521(new_n6898, new_n6897, new_n6886);
nand_4 g06522(new_n6899, n11222, n159);
xnor_3 g06523(new_n6900, new_n6895, new_n6894);
nor_4  g06524(new_n6901, new_n6900, new_n6899);
not_3  g06525(new_n6902, new_n6901);
nand_4 g06526(new_n6903, new_n6900, new_n6899);
nand_4 g06527(new_n6904, new_n4150, new_n4147);
not_3  g06528(new_n6905, new_n6904);
nor_4  g06529(new_n6906, new_n4161, new_n4151);
nor_4  g06530(new_n6907, new_n6906, new_n6905);
not_3  g06531(new_n6908, new_n6907);
nand_4 g06532(new_n6909, new_n6908, new_n6903);
nand_4 g06533(new_n6910, new_n6909, new_n6902);
not_3  g06534(new_n6911, new_n6910);
nor_4  g06535(new_n6912, new_n6911, new_n6898);
not_3  g06536(new_n6913, new_n6881);
not_3  g06537(new_n6914, new_n6885);
nand_4 g06538(new_n6915, new_n6914, new_n6913);
nor_4  g06539(new_n6916, new_n6883, new_n6882);
nor_4  g06540(new_n6917, new_n6897, new_n6886);
xnor_3 g06541(new_n6918, new_n6917, new_n6916);
nand_4 g06542(new_n6919, new_n6918, new_n6915);
not_3  g06543(new_n6920, new_n6868);
nand_4 g06544(new_n6921, new_n6880, new_n6872);
nand_4 g06545(new_n6922, new_n6921, new_n6920);
nand_4 g06546(new_n6923, n11153, n1510);
not_3  g06547(new_n6924, new_n6923);
nand_4 g06548(new_n6925, n5314, n159);
nand_4 g06549(new_n6926, n12247, n11222);
not_3  g06550(new_n6927, new_n6926);
xor_3  g06551(new_n6928, new_n6927, new_n6925);
xnor_3 g06552(new_n6929, new_n6928, new_n6924);
not_3  g06553(new_n6930, new_n6929);
xnor_3 g06554(new_n6931, new_n6930, new_n6922);
nor_4  g06555(new_n6932, new_n6866, new_n6865);
nand_4 g06556(new_n6933, n2749, n996);
not_3  g06557(new_n6934, new_n6933);
xor_3  g06558(new_n6935, new_n6934, new_n6932);
not_3  g06559(new_n6936, new_n6935);
nand_4 g06560(new_n6937, n10898, n5319);
not_3  g06561(new_n6938, new_n6937);
nand_4 g06562(new_n6939, n11876, n9457);
nand_4 g06563(new_n6940, n5767, n3754);
not_3  g06564(new_n6941, new_n6940);
xor_3  g06565(new_n6942, new_n6941, new_n6939);
xnor_3 g06566(new_n6943, new_n6942, new_n6938);
xnor_3 g06567(new_n6944, new_n6943, new_n6936);
not_3  g06568(new_n6945, new_n6944);
xnor_3 g06569(new_n6946, new_n6945, new_n6931);
xnor_3 g06570(new_n6947, new_n6946, new_n6919);
xnor_3 g06571(new_n6948, new_n6947, new_n6912);
nand_4 g06572(new_n6949, n11222, n1510);
not_3  g06573(new_n6950, new_n6949);
not_3  g06574(new_n6951, new_n6898);
nor_4  g06575(new_n6952, new_n6910, new_n6951);
nor_4  g06576(new_n6953, new_n6952, new_n6912);
nor_4  g06577(new_n6954, new_n6953, new_n6950);
not_3  g06578(new_n6955, new_n4165);
nand_4 g06579(new_n6956, new_n6903, new_n6902);
xnor_3 g06580(new_n6957, new_n6956, new_n6908);
not_3  g06581(new_n6958, new_n6957);
nor_4  g06582(new_n6959, new_n6958, new_n6955);
xnor_3 g06583(new_n6960, new_n6953, new_n6950);
nor_4  g06584(new_n6961, new_n6960, new_n6959);
nor_4  g06585(new_n6962, new_n6961, new_n6954);
xnor_3 g06586(new_n6963, new_n6962, new_n6948);
xnor_3 g06587(new_n6964, new_n6960, new_n6959);
xnor_3 g06588(new_n6965, new_n6860_1, new_n6859);
nor_4  g06589(new_n6966, new_n6965, new_n6964);
not_3  g06590(new_n6967, new_n6966);
not_3  g06591(new_n6968, new_n6959);
xnor_3 g06592(new_n6969, new_n6960, new_n6968);
not_3  g06593(new_n6970, new_n6859);
xnor_3 g06594(new_n6971, new_n6860_1, new_n6970);
nor_4  g06595(new_n6972, new_n6971, new_n6969);
xnor_3 g06596(new_n6973, new_n6858, new_n6855);
not_3  g06597(new_n6974, new_n6973);
not_3  g06598(new_n6975, new_n4169);
nand_4 g06599(new_n6976, new_n4180, new_n6975);
not_3  g06600(new_n6977, new_n6976);
nand_4 g06601(new_n6978, new_n6977, new_n6974);
nand_4 g06602(new_n6979, new_n6976, new_n6973);
nor_4  g06603(new_n6980, new_n6957, new_n4165);
nor_4  g06604(new_n6981, new_n6980, new_n6959);
nand_4 g06605(new_n6982, new_n6981, new_n6979);
nand_4 g06606(new_n6983, new_n6982, new_n6978);
nor_4  g06607(new_n6984, new_n6983, new_n6972);
not_3  g06608(new_n6985, new_n6984);
nand_4 g06609(new_n6986_1, new_n6985, new_n6967);
xnor_3 g06610(new_n6987, new_n6986_1, new_n6963);
xnor_3 g06611(new_n6988, new_n6987, new_n6863);
xnor_3 g06612(new_n6989, new_n6988, new_n6768);
not_3  g06613(new_n6990, new_n6762);
not_3  g06614(new_n6991, new_n6764);
nor_4  g06615(new_n6992, new_n6991, new_n6990);
nor_4  g06616(new_n6993, new_n6992, new_n6765);
not_3  g06617(new_n6994, new_n6993);
not_3  g06618(new_n6995, new_n6761);
xor_3  g06619(new_n6996, new_n6995, new_n6760);
not_3  g06620(new_n6997, new_n6996);
not_3  g06621(new_n6998, new_n6981);
xnor_3 g06622(new_n6999, new_n6976, new_n6974);
xnor_3 g06623(new_n7000, new_n6999, new_n6998);
nand_4 g06624(new_n7001, new_n7000, new_n6997);
xnor_3 g06625(new_n7002, new_n6999, new_n6981);
nand_4 g06626(new_n7003, new_n7002, new_n6996);
nand_4 g06627(new_n7004, new_n4214, new_n4209);
nand_4 g06628(new_n7005, new_n7004, new_n7003);
nand_4 g06629(new_n7006, new_n7005, new_n7001);
nand_4 g06630(new_n7007, new_n7006, new_n6994);
xnor_3 g06631(new_n7008, new_n7006, new_n6993);
not_3  g06632(new_n7009, new_n6972);
nand_4 g06633(new_n7010, new_n7009, new_n6967);
xnor_3 g06634(new_n7011, new_n7010, new_n6983);
nand_4 g06635(new_n7012, new_n7011, new_n7008);
nand_4 g06636(new_n7013, new_n7012, new_n7007);
xnor_3 g06637(new_n7014, new_n7013, new_n6989);
nand_4 g06638(new_n7015, new_n7014, new_n6666);
not_3  g06639(new_n7016, new_n6666);
not_3  g06640(new_n7017, new_n7014);
nand_4 g06641(new_n7018, new_n7017, new_n7016);
nand_4 g06642(new_n7019, new_n7018, new_n7015);
not_3  g06643(new_n7020, new_n6663);
xor_3  g06644(new_n7021, new_n7020, new_n6660);
not_3  g06645(new_n7022, new_n7021);
xnor_3 g06646(new_n7023, new_n7011, new_n7008);
not_3  g06647(new_n7024, new_n7023);
nand_4 g06648(new_n7025, new_n7024, new_n7022);
nand_4 g06649(new_n7026, new_n7023, new_n7021);
xor_3  g06650(new_n7027, new_n6659, new_n6655);
not_3  g06651(new_n7028, new_n7027);
nand_4 g06652(new_n7029, new_n7003, new_n7001);
xnor_3 g06653(new_n7030, new_n7029, new_n7004);
nor_4  g06654(new_n7031, new_n7030, new_n7028);
nand_4 g06655(new_n7032, new_n4124, new_n4028);
nand_4 g06656(new_n7033, new_n4216, new_n4125);
nand_4 g06657(new_n7034, new_n7033, new_n7032);
xnor_3 g06658(new_n7035, new_n7030, new_n7028);
nor_4  g06659(new_n7036, new_n7035, new_n7034);
nor_4  g06660(new_n7037, new_n7036, new_n7031);
nand_4 g06661(new_n7038, new_n7037, new_n7026);
nand_4 g06662(new_n7039, new_n7038, new_n7025);
xnor_3 g06663(n2301, new_n7039, new_n7019);
xor_3  g06664(n2316, new_n4122, new_n4121);
nand_4 g06665(new_n7042, n4634, n1333);
not_3  g06666(new_n7043, new_n7042);
not_3  g06667(new_n7044, new_n6301);
nor_4  g06668(new_n7045, new_n6307, new_n7044);
nor_4  g06669(new_n7046, new_n7045, new_n6306);
nand_4 g06670(new_n7047, new_n7046, new_n7043);
xnor_3 g06671(new_n7048, new_n7046, new_n7042);
nand_4 g06672(new_n7049, n11757, n2879);
not_3  g06673(new_n7050, new_n7049);
nand_4 g06674(new_n7051, n10223, n3172);
not_3  g06675(new_n7052, new_n7051);
nand_4 g06676(new_n7053, n7265, n5240);
not_3  g06677(new_n7054, new_n7053);
nor_4  g06678(new_n7055, new_n7054, new_n7052);
not_3  g06679(new_n7056, new_n7055);
nor_4  g06680(new_n7057, new_n7053, new_n7051);
not_3  g06681(new_n7058, new_n7057);
nand_4 g06682(new_n7059, new_n7058, new_n7056);
xnor_3 g06683(new_n7060, new_n7059, new_n7050);
nand_4 g06684(new_n7061, new_n7060, new_n7048);
nand_4 g06685(new_n7062, new_n7061, new_n7047);
nand_4 g06686(new_n7063, n4634, n3172);
nand_4 g06687(new_n7064, n9195, n1333);
xor_3  g06688(new_n7065, new_n7064, new_n7063);
xnor_3 g06689(new_n7066, new_n7065, new_n7062);
nand_4 g06690(new_n7067, n11757, n10223);
not_3  g06691(new_n7068, new_n7067);
nand_4 g06692(new_n7069, n5240, n2879);
nand_4 g06693(new_n7070, n11821, n7265);
xnor_3 g06694(new_n7071, new_n7070, new_n7069);
not_3  g06695(new_n7072, new_n7071);
nor_4  g06696(new_n7073, new_n7072, new_n7068);
nor_4  g06697(new_n7074, new_n7071, new_n7067);
nor_4  g06698(new_n7075, new_n7074, new_n7073);
nor_4  g06699(new_n7076, new_n7057, new_n7050);
nor_4  g06700(new_n7077, new_n7076, new_n7055);
not_3  g06701(new_n7078, new_n7077);
xor_3  g06702(new_n7079, new_n7078, new_n7075);
xnor_3 g06703(new_n7080, new_n7079, new_n7066);
not_3  g06704(new_n7081, new_n7080);
nand_4 g06705(new_n7082, n9195, n7862);
xnor_3 g06706(new_n7083, new_n7060, new_n7048);
nor_4  g06707(new_n7084, new_n7083, new_n7082);
not_3  g06708(new_n7085, new_n7084);
not_3  g06709(new_n7086, new_n6289);
nand_4 g06710(new_n7087, new_n6299, new_n7086);
xor_3  g06711(new_n7088, new_n6299, new_n7086);
xor_3  g06712(new_n7089, new_n6308, new_n7044);
nand_4 g06713(new_n7090, new_n7089, new_n7088);
nand_4 g06714(new_n7091, new_n7090, new_n7087);
not_3  g06715(new_n7092, new_n7082);
not_3  g06716(new_n7093, new_n7083);
nor_4  g06717(new_n7094, new_n7093, new_n7092);
nor_4  g06718(new_n7095, new_n7094, new_n7084);
nand_4 g06719(new_n7096, new_n7095, new_n7091);
nand_4 g06720(new_n7097, new_n7096, new_n7085);
nand_4 g06721(new_n7098, new_n7097, new_n7081);
not_3  g06722(new_n7099, new_n7075);
nor_4  g06723(new_n7100, new_n7077, new_n7099);
nor_4  g06724(new_n7101, new_n7100, new_n7073);
nand_4 g06725(new_n7102, n2253, n1333);
nand_4 g06726(new_n7103, n9195, n3172);
nand_4 g06727(new_n7104, n7862, n3865);
xor_3  g06728(new_n7105, new_n7104, new_n7103);
xnor_3 g06729(new_n7106, new_n7105, new_n7102);
xnor_3 g06730(new_n7107, new_n7106, new_n7101);
nor_4  g06731(new_n7108, new_n7070, new_n7069);
nand_4 g06732(new_n7109, n11757, n4634);
not_3  g06733(new_n7110, new_n7109);
xor_3  g06734(new_n7111, new_n7110, new_n7108);
nand_4 g06735(new_n7112, n11821, n2879);
not_3  g06736(new_n7113, new_n7112);
nand_4 g06737(new_n7114, n10223, n5240);
nand_4 g06738(new_n7115, n9080, n7265);
xnor_3 g06739(new_n7116, new_n7115, new_n7114);
and_4  g06740(new_n7117, new_n7116, new_n7113);
nor_4  g06741(new_n7118, new_n7116, new_n7113);
nor_4  g06742(new_n7119, new_n7118, new_n7117);
xnor_3 g06743(new_n7120, new_n7119, new_n7111);
not_3  g06744(new_n7121, new_n7120);
xnor_3 g06745(new_n7122, new_n7121, new_n7107);
nand_4 g06746(new_n7123, new_n7065, new_n7062);
nor_4  g06747(new_n7124, new_n7064, new_n7063);
nor_4  g06748(new_n7125, new_n7079, new_n7066);
xnor_3 g06749(new_n7126, new_n7125, new_n7124);
nand_4 g06750(new_n7127, new_n7126, new_n7123);
xnor_3 g06751(new_n7128, new_n7127, new_n7122);
xnor_3 g06752(new_n7129, new_n7128, new_n7098);
nand_4 g06753(new_n7130, n7862, n2253);
not_3  g06754(new_n7131, new_n7130);
xnor_3 g06755(new_n7132, new_n7097, new_n7080);
nand_4 g06756(new_n7133, new_n7132, new_n7131);
not_3  g06757(new_n7134, new_n6318);
nor_4  g06758(new_n7135, new_n7134, new_n6310);
not_3  g06759(new_n7136, new_n7135);
xnor_3 g06760(new_n7137, new_n7095, new_n7091);
nor_4  g06761(new_n7138, new_n7137, new_n7136);
xnor_3 g06762(new_n7139, new_n7132, new_n7130);
nand_4 g06763(new_n7140, new_n7139, new_n7138);
nand_4 g06764(new_n7141, new_n7140, new_n7133);
xor_3  g06765(new_n7142, new_n7141, new_n7129);
not_3  g06766(new_n7143, new_n7142);
not_3  g06767(new_n7144, new_n7138);
xnor_3 g06768(new_n7145, new_n7139, new_n7144);
not_3  g06769(new_n7146, new_n7145);
not_3  g06770(new_n7147, new_n7137);
xor_3  g06771(new_n7148, new_n7147, new_n7136);
not_3  g06772(new_n7149, new_n6355);
nand_4 g06773(new_n7150, n12145, n6877);
nand_4 g06774(new_n7151, n9400, n2522);
not_3  g06775(new_n7152, new_n7151);
nand_4 g06776(new_n7153, n11311, n2024);
not_3  g06777(new_n7154, new_n7153);
nand_4 g06778(new_n7155, n9189, n2464);
nand_4 g06779(new_n7156, n7946, n4187);
xnor_3 g06780(new_n7157, new_n7156, new_n7155);
xnor_3 g06781(new_n7158, new_n7157, new_n7154);
xnor_3 g06782(new_n7159_1, new_n7158, new_n7152);
and_4  g06783(new_n7160_1, new_n6323, new_n6322);
nor_4  g06784(new_n7161, new_n6328, new_n7160_1);
xnor_3 g06785(new_n7162, new_n7161, new_n7159_1);
xnor_3 g06786(new_n7163, new_n7162, new_n7150);
nor_4  g06787(new_n7164, new_n6329, new_n6320);
nor_4  g06788(new_n7165, new_n6342, new_n7164);
not_3  g06789(new_n7166, new_n7165);
xnor_3 g06790(new_n7167, new_n7166, new_n7163);
nor_4  g06791(new_n7168, new_n7167, new_n7149);
not_3  g06792(new_n7169, new_n7167);
nor_4  g06793(new_n7170, new_n7169, new_n6355);
nor_4  g06794(new_n7171, new_n7170, new_n7168);
not_3  g06795(new_n7172, new_n6442);
nand_4 g06796(new_n7173, new_n6497, new_n7172);
xnor_3 g06797(new_n7174, new_n7173, new_n7171);
not_3  g06798(new_n7175, new_n6466);
nand_4 g06799(new_n7176, n11478, n521);
not_3  g06800(new_n7177, new_n7176);
not_3  g06801(new_n7178, new_n6456);
not_3  g06802(new_n7179, new_n6457);
nor_4  g06803(new_n7180, new_n7179, new_n7178);
not_3  g06804(new_n7181, new_n6455);
nor_4  g06805(new_n7182, new_n6457, new_n6456);
nor_4  g06806(new_n7183, new_n7182, new_n7181);
nor_4  g06807(new_n7184, new_n7183, new_n7180);
xnor_3 g06808(new_n7185, new_n7184, new_n7177);
nand_4 g06809(new_n7186, n2498, n137);
not_3  g06810(new_n7187, new_n7186);
nand_4 g06811(new_n7188, n5579, n5283);
not_3  g06812(new_n7189, new_n7188);
nand_4 g06813(new_n7190, n6294, n2558);
not_3  g06814(new_n7191, new_n7190);
nor_4  g06815(new_n7192, new_n7191, new_n7189);
not_3  g06816(new_n7193_1, new_n7192);
nor_4  g06817(new_n7194, new_n7190, new_n7188);
not_3  g06818(new_n7195, new_n7194);
nand_4 g06819(new_n7196, new_n7195, new_n7193_1);
xnor_3 g06820(new_n7197, new_n7196, new_n7187);
xnor_3 g06821(new_n7198, new_n7197, new_n7185);
not_3  g06822(new_n7199, new_n7198);
nand_4 g06823(new_n7200, n6016, n4805);
not_3  g06824(new_n7201, new_n7200);
not_3  g06825(new_n7202, new_n6451);
nand_4 g06826(new_n7203, new_n6460, new_n6454);
nand_4 g06827(new_n7204, new_n7203, new_n7202);
nor_4  g06828(new_n7205, new_n7204, new_n7201);
not_3  g06829(new_n7206, new_n7204);
nor_4  g06830(new_n7207, new_n7206, new_n7200);
nor_4  g06831(new_n7208, new_n7207, new_n7205);
nand_4 g06832(new_n7209, new_n7208, new_n7199);
not_3  g06833(new_n7210, new_n7209);
nor_4  g06834(new_n7211, new_n7208, new_n7199);
nor_4  g06835(new_n7212, new_n7211, new_n7210);
xnor_3 g06836(new_n7213, new_n7212, new_n7175);
not_3  g06837(new_n7214, new_n6490);
nand_4 g06838(new_n7215, n7270, n7236);
not_3  g06839(new_n7216, new_n7215);
not_3  g06840(new_n7217, new_n6473);
nand_4 g06841(new_n7218, new_n6482, new_n6476);
nand_4 g06842(new_n7219, new_n7218, new_n7217);
nor_4  g06843(new_n7220, new_n7219, new_n7216);
not_3  g06844(new_n7221, new_n7219);
nor_4  g06845(new_n7222, new_n7221, new_n7215);
nor_4  g06846(new_n7223, new_n7222, new_n7220);
nand_4 g06847(new_n7224, n3992, n806);
not_3  g06848(new_n7225, new_n7224);
not_3  g06849(new_n7226, new_n6478);
not_3  g06850(new_n7227, new_n6479);
nor_4  g06851(new_n7228, new_n7227, new_n7226);
not_3  g06852(new_n7229, new_n6477);
nor_4  g06853(new_n7230, new_n6479, new_n6478);
nor_4  g06854(new_n7231, new_n7230, new_n7229);
nor_4  g06855(new_n7232, new_n7231, new_n7228);
nand_4 g06856(new_n7233, new_n7232, new_n7225);
not_3  g06857(new_n7234, new_n7233);
nor_4  g06858(new_n7235, new_n7232, new_n7225);
nor_4  g06859(new_n7236_1, new_n7235, new_n7234);
not_3  g06860(new_n7237, new_n7236_1);
nand_4 g06861(new_n7238, n9111, n6358);
nand_4 g06862(new_n7239, n8384, n3342);
nand_4 g06863(new_n7240, n9763, n5198);
xnor_3 g06864(new_n7241, new_n7240, new_n7239);
xnor_3 g06865(new_n7242, new_n7241, new_n7238);
xnor_3 g06866(new_n7243, new_n7242, new_n7237);
nand_4 g06867(new_n7244, new_n7243, new_n7223);
not_3  g06868(new_n7245, new_n7244);
nor_4  g06869(new_n7246, new_n7243, new_n7223);
nor_4  g06870(new_n7247, new_n7246, new_n7245);
xnor_3 g06871(new_n7248, new_n7247, new_n7214);
xnor_3 g06872(new_n7249, new_n7248, new_n7213);
nor_4  g06873(new_n7250, new_n6491, new_n6467);
nor_4  g06874(new_n7251, new_n6494, new_n6492);
nor_4  g06875(new_n7252, new_n7251, new_n7250);
xnor_3 g06876(new_n7253, new_n7252, new_n7249);
xnor_3 g06877(new_n7254, new_n7253, new_n7174);
not_3  g06878(new_n7255, new_n7254);
nand_4 g06879(new_n7256, new_n7255, new_n7148);
xnor_3 g06880(new_n7257, new_n7254, new_n7148);
nand_4 g06881(new_n7258, new_n6526, new_n6502);
nand_4 g06882(new_n7259, new_n7258, new_n6501);
nand_4 g06883(new_n7260, new_n7259, new_n7257);
nand_4 g06884(new_n7261, new_n7260, new_n7256);
nand_4 g06885(new_n7262, new_n7261, new_n7146);
nor_4  g06886(new_n7263, new_n7247, new_n7214);
not_3  g06887(new_n7264, new_n7263);
nand_4 g06888(new_n7265_1, n7236, n5153);
nand_4 g06889(new_n7266, n6358, n3342);
nand_4 g06890(new_n7267, n9111, n5198);
nand_4 g06891(new_n7268, n9763, n1471);
xnor_3 g06892(new_n7269, new_n7268, new_n7267);
nor_4  g06893(new_n7270_1, new_n7269, new_n7266);
not_3  g06894(new_n7271, new_n7266);
not_3  g06895(new_n7272, new_n7269);
nor_4  g06896(new_n7273, new_n7272, new_n7271);
nor_4  g06897(new_n7274, new_n7273, new_n7270_1);
and_4  g06898(new_n7275, new_n7240, new_n7239);
not_3  g06899(new_n7276, new_n7238);
nor_4  g06900(new_n7277, new_n7241, new_n7276);
nor_4  g06901(new_n7278, new_n7277, new_n7275);
xnor_3 g06902(new_n7279, new_n7278, new_n7274);
nand_4 g06903(new_n7280, n7270, n3992);
nand_4 g06904(new_n7281, n8384, n806);
not_3  g06905(new_n7282, new_n7281);
xor_3  g06906(new_n7283, new_n7282, new_n7280);
xnor_3 g06907(new_n7284, new_n7283, new_n7279);
nor_4  g06908(new_n7285, new_n7242, new_n7237);
nor_4  g06909(new_n7286, new_n7285, new_n7234);
xnor_3 g06910(new_n7287, new_n7286, new_n7284);
not_3  g06911(new_n7288, new_n7220);
nand_4 g06912(new_n7289, new_n7244, new_n7288);
xnor_3 g06913(new_n7290, new_n7289, new_n7287);
xnor_3 g06914(new_n7291, new_n7290, new_n7265_1);
xnor_3 g06915(new_n7292, new_n7291, new_n7264);
nor_4  g06916(new_n7293, new_n7212, new_n7175);
nand_4 g06917(new_n7294_1, n5798, n4805);
nand_4 g06918(new_n7295, n5579, n137);
nand_4 g06919(new_n7296, n6797, n2558);
nand_4 g06920(new_n7297, n6294, n2498);
xnor_3 g06921(new_n7298, new_n7297, new_n7296);
nor_4  g06922(new_n7299, new_n7298, new_n7295);
not_3  g06923(new_n7300, new_n7295);
not_3  g06924(new_n7301, new_n7298);
nor_4  g06925(new_n7302, new_n7301, new_n7300);
nor_4  g06926(new_n7303, new_n7302, new_n7299);
nor_4  g06927(new_n7304, new_n7194, new_n7187);
nor_4  g06928(new_n7305, new_n7304, new_n7192);
xnor_3 g06929(new_n7306, new_n7305, new_n7303);
nand_4 g06930(new_n7307, n11478, n6016);
nand_4 g06931(new_n7308, n5283, n521);
xor_3  g06932(new_n7309, new_n7308, new_n7307);
xnor_3 g06933(new_n7310, new_n7309, new_n7306);
and_4  g06934(new_n7311, new_n7184, new_n7177);
not_3  g06935(new_n7312, new_n7197);
nor_4  g06936(new_n7313, new_n7312, new_n7185);
nor_4  g06937(new_n7314, new_n7313, new_n7311);
xnor_3 g06938(new_n7315, new_n7314, new_n7310);
not_3  g06939(new_n7316, new_n7205);
nand_4 g06940(new_n7317, new_n7209, new_n7316);
xnor_3 g06941(new_n7318, new_n7317, new_n7315);
not_3  g06942(new_n7319, new_n7318);
nand_4 g06943(new_n7320_1, new_n7319, new_n7294_1);
not_3  g06944(new_n7321, new_n7294_1);
nand_4 g06945(new_n7322, new_n7318, new_n7321);
nand_4 g06946(new_n7323, new_n7322, new_n7320_1);
xnor_3 g06947(new_n7324, new_n7323, new_n7293);
xnor_3 g06948(new_n7325, new_n7324, new_n7292);
nand_4 g06949(new_n7326, new_n7248, new_n7213);
not_3  g06950(new_n7327, new_n7326);
nor_4  g06951(new_n7328, new_n7252, new_n7249);
nor_4  g06952(new_n7329, new_n7328, new_n7327);
not_3  g06953(new_n7330, new_n7329);
nand_4 g06954(new_n7331, new_n7330, new_n7325);
not_3  g06955(new_n7332, new_n7331);
nor_4  g06956(new_n7333, new_n7330, new_n7325);
nor_4  g06957(new_n7334, new_n7333, new_n7332);
nor_4  g06958(new_n7335, new_n7173, new_n7171);
not_3  g06959(new_n7336, new_n7335);
not_3  g06960(new_n7337, new_n7174);
not_3  g06961(new_n7338, new_n7253);
nand_4 g06962(new_n7339, new_n7338, new_n7337);
nand_4 g06963(new_n7340, new_n7339, new_n7336);
not_3  g06964(new_n7341, new_n7340);
nand_4 g06965(new_n7342, n12221, n6877);
not_3  g06966(new_n7343, new_n7342);
not_3  g06967(new_n7344, new_n7150);
nand_4 g06968(new_n7345, new_n7162, new_n7344);
nand_4 g06969(new_n7346, new_n7166, new_n7163);
nand_4 g06970(new_n7347, new_n7346, new_n7345);
nor_4  g06971(new_n7348, new_n7158, new_n7152);
nor_4  g06972(new_n7349, new_n7161, new_n7159_1);
nor_4  g06973(new_n7350, new_n7349, new_n7348);
not_3  g06974(new_n7351, new_n7350);
nand_4 g06975(new_n7352, n11311, n9189);
not_3  g06976(new_n7353, new_n7352);
nand_4 g06977(new_n7354_1, n4187, n2024);
nand_4 g06978(new_n7355, n7946, n4203);
not_3  g06979(new_n7356, new_n7355);
xor_3  g06980(new_n7357, new_n7356, new_n7354_1);
xnor_3 g06981(new_n7358, new_n7357, new_n7353);
and_4  g06982(new_n7359, new_n7156, new_n7155);
nor_4  g06983(new_n7360, new_n7156, new_n7155);
nor_4  g06984(new_n7361, new_n7360, new_n7154);
nor_4  g06985(new_n7362, new_n7361, new_n7359);
not_3  g06986(new_n7363, new_n7362);
xnor_3 g06987(new_n7364, new_n7363, new_n7358);
nand_4 g06988(new_n7365, n12145, n9400);
nand_4 g06989(new_n7366, n2522, n2464);
xor_3  g06990(new_n7367, new_n7366, new_n7365);
xnor_3 g06991(new_n7368, new_n7367, new_n7364);
xnor_3 g06992(new_n7369, new_n7368, new_n7351);
xnor_3 g06993(new_n7370, new_n7369, new_n7347);
xnor_3 g06994(new_n7371, new_n7370, new_n7343);
xnor_3 g06995(new_n7372, new_n7371, new_n7168);
xnor_3 g06996(new_n7373, new_n7372, new_n7341);
xnor_3 g06997(new_n7374, new_n7373, new_n7334);
xnor_3 g06998(new_n7375, new_n7261, new_n7145);
nand_4 g06999(new_n7376, new_n7375, new_n7374);
nand_4 g07000(new_n7377, new_n7376, new_n7262);
nand_4 g07001(new_n7378, new_n7377, new_n7143);
xnor_3 g07002(new_n7379, new_n7377, new_n7142);
xnor_3 g07003(new_n7380, new_n7368, new_n7350);
nand_4 g07004(new_n7381, new_n7380, new_n7347);
nand_4 g07005(new_n7382, new_n7357, new_n7352);
nand_4 g07006(new_n7383, new_n7363, new_n7358);
nand_4 g07007(new_n7384, new_n7383, new_n7382);
nand_4 g07008(new_n7385, n12221, n9400);
not_3  g07009(new_n7386, new_n7385);
nand_4 g07010(new_n7387, n12145, n2464);
nand_4 g07011(new_n7388_1, n10217, n6877);
not_3  g07012(new_n7389, new_n7388_1);
xor_3  g07013(new_n7390, new_n7389, new_n7387);
xnor_3 g07014(new_n7391, new_n7390, new_n7386);
xnor_3 g07015(new_n7392, new_n7391, new_n7384);
nor_4  g07016(new_n7393, new_n7355, new_n7354_1);
nand_4 g07017(new_n7394, n11311, n2522);
not_3  g07018(new_n7395, new_n7394);
xor_3  g07019(new_n7396, new_n7395, new_n7393);
nand_4 g07020(new_n7397, n4203, n2024);
nand_4 g07021(new_n7398, n9189, n4187);
not_3  g07022(new_n7399, new_n7398);
nand_4 g07023(new_n7400, n12753, n7946);
not_3  g07024(new_n7401, new_n7400);
nand_4 g07025(new_n7402, new_n7401, new_n7399);
nand_4 g07026(new_n7403, new_n7400, new_n7398);
nand_4 g07027(new_n7404, new_n7403, new_n7402);
xor_3  g07028(new_n7405, new_n7404, new_n7397);
xnor_3 g07029(new_n7406, new_n7405, new_n7396);
xnor_3 g07030(new_n7407, new_n7406, new_n7392);
nand_4 g07031(new_n7408, new_n7367, new_n7364);
nor_4  g07032(new_n7409, new_n7366, new_n7365);
nor_4  g07033(new_n7410, new_n7367, new_n7364);
nor_4  g07034(new_n7411, new_n7410, new_n7351);
xnor_3 g07035(new_n7412, new_n7411, new_n7409);
nand_4 g07036(new_n7413, new_n7412, new_n7408);
xnor_3 g07037(new_n7414, new_n7413, new_n7407);
xnor_3 g07038(new_n7415, new_n7414, new_n7381);
xnor_3 g07039(new_n7416, new_n7380, new_n7347);
nor_4  g07040(new_n7417, new_n7416, new_n7342);
not_3  g07041(new_n7418, new_n7168);
nor_4  g07042(new_n7419, new_n7371, new_n7418);
nor_4  g07043(new_n7420, new_n7419, new_n7417);
xnor_3 g07044(new_n7421, new_n7420, new_n7415);
not_3  g07045(new_n7422, new_n7317);
nand_4 g07046(new_n7423, new_n7422, new_n7315);
nand_4 g07047(new_n7424, n4805, n2347);
nand_4 g07048(new_n7425, n6016, n5283);
nand_4 g07049(new_n7426, n11478, n5798);
not_3  g07050(new_n7427, new_n7426);
xor_3  g07051(new_n7428, new_n7427, new_n7425);
xnor_3 g07052(new_n7429, new_n7428, new_n7424);
nand_4 g07053(new_n7430, new_n7305, new_n7303);
not_3  g07054(new_n7431, new_n7430);
nor_4  g07055(new_n7432, new_n7431, new_n7299);
not_3  g07056(new_n7433, new_n7432);
xnor_3 g07057(new_n7434, new_n7433, new_n7429);
nor_4  g07058(new_n7435, new_n7297, new_n7296);
nand_4 g07059(new_n7436_1, n521, n137);
xor_3  g07060(new_n7437, new_n7436_1, new_n7435);
nand_4 g07061(new_n7438, n6797, n2498);
nand_4 g07062(new_n7439, n6294, n5579);
nand_4 g07063(new_n7440, n3146, n2558);
not_3  g07064(new_n7441, new_n7440);
xor_3  g07065(new_n7442, new_n7441, new_n7439);
xnor_3 g07066(new_n7443, new_n7442, new_n7438);
xnor_3 g07067(new_n7444, new_n7443, new_n7437);
xnor_3 g07068(new_n7445, new_n7444, new_n7434);
not_3  g07069(new_n7446, new_n7306);
nand_4 g07070(new_n7447, new_n7309, new_n7446);
nor_4  g07071(new_n7448, new_n7308, new_n7307);
not_3  g07072(new_n7449, new_n7310);
nor_4  g07073(new_n7450, new_n7314, new_n7449);
xnor_3 g07074(new_n7451, new_n7450, new_n7448);
nand_4 g07075(new_n7452, new_n7451, new_n7447);
xnor_3 g07076(new_n7453, new_n7452, new_n7445);
xnor_3 g07077(new_n7454, new_n7453, new_n7423);
nand_4 g07078(new_n7455, new_n7320_1, new_n7293);
nand_4 g07079(new_n7456_1, new_n7455, new_n7322);
xnor_3 g07080(new_n7457, new_n7456_1, new_n7454);
nor_4  g07081(new_n7458, new_n7289, new_n7287);
not_3  g07082(new_n7459, new_n7458);
not_3  g07083(new_n7460, new_n7279);
not_3  g07084(new_n7461, new_n7283);
nand_4 g07085(new_n7462, new_n7461, new_n7460);
nor_4  g07086(new_n7463, new_n7281, new_n7280);
nor_4  g07087(new_n7464, new_n7286, new_n7284);
xnor_3 g07088(new_n7465, new_n7464, new_n7463);
nand_4 g07089(new_n7466, new_n7465, new_n7462);
nor_4  g07090(new_n7467, new_n7268, new_n7267);
nand_4 g07091(new_n7468, n6358, n806);
not_3  g07092(new_n7469, new_n7468);
xor_3  g07093(new_n7470, new_n7469, new_n7467);
nand_4 g07094(new_n7471, n9111, n1471);
nand_4 g07095(new_n7472, n5198, n3342);
nand_4 g07096(new_n7473, n9763, n7646);
nand_4 g07097(new_n7474, new_n7473, new_n7472);
not_3  g07098(new_n7475, new_n7472);
not_3  g07099(new_n7476, new_n7473);
nand_4 g07100(new_n7477, new_n7476, new_n7475);
nand_4 g07101(new_n7478, new_n7477, new_n7474);
xor_3  g07102(new_n7479, new_n7478, new_n7471);
xnor_3 g07103(new_n7480, new_n7479, new_n7470);
not_3  g07104(new_n7481, new_n7480);
not_3  g07105(new_n7482, new_n7270_1);
nand_4 g07106(new_n7483, new_n7278, new_n7274);
nand_4 g07107(new_n7484, new_n7483, new_n7482);
nand_4 g07108(new_n7485, n5153, n3992);
nand_4 g07109(new_n7486, n8384, n7270);
nand_4 g07110(new_n7487, n7236, n2507);
not_3  g07111(new_n7488, new_n7487);
xor_3  g07112(new_n7489, new_n7488, new_n7486);
xnor_3 g07113(new_n7490, new_n7489, new_n7485);
xnor_3 g07114(new_n7491, new_n7490, new_n7484);
xnor_3 g07115(new_n7492, new_n7491, new_n7481);
xnor_3 g07116(new_n7493, new_n7492, new_n7466);
xnor_3 g07117(new_n7494, new_n7493, new_n7459);
nor_4  g07118(new_n7495, new_n7290, new_n7265_1);
not_3  g07119(new_n7496, new_n7495);
nand_4 g07120(new_n7497, new_n7290, new_n7265_1);
nand_4 g07121(new_n7498, new_n7497, new_n7263);
nand_4 g07122(new_n7499, new_n7498, new_n7496);
xnor_3 g07123(new_n7500_1, new_n7499, new_n7494);
xnor_3 g07124(new_n7501, new_n7500_1, new_n7457);
not_3  g07125(new_n7502, new_n7324);
nand_4 g07126(new_n7503, new_n7502, new_n7292);
nand_4 g07127(new_n7504, new_n7331, new_n7503);
xnor_3 g07128(new_n7505, new_n7504, new_n7501);
xnor_3 g07129(new_n7506, new_n7505, new_n7421);
nand_4 g07130(new_n7507, new_n7372, new_n7341);
not_3  g07131(new_n7508, new_n7334);
not_3  g07132(new_n7509, new_n7373);
nand_4 g07133(new_n7510, new_n7509, new_n7508);
nand_4 g07134(new_n7511, new_n7510, new_n7507);
xnor_3 g07135(new_n7512, new_n7511, new_n7506);
nand_4 g07136(new_n7513, new_n7512, new_n7379);
nand_4 g07137(new_n7514, new_n7513, new_n7378);
not_3  g07138(new_n7515, new_n7421);
nand_4 g07139(new_n7516, new_n7505, new_n7515);
nand_4 g07140(new_n7517, new_n7511, new_n7506);
nand_4 g07141(new_n7518, new_n7517, new_n7516);
nor_4  g07142(new_n7519, new_n7453, new_n7423);
not_3  g07143(new_n7520, new_n7456_1);
nor_4  g07144(new_n7521, new_n7520, new_n7454);
nor_4  g07145(new_n7522, new_n7521, new_n7519);
xnor_3 g07146(new_n7523_1, new_n7522, new_n7518);
not_3  g07147(new_n7524, new_n7457);
nand_4 g07148(new_n7525, new_n7500_1, new_n7524);
nand_4 g07149(new_n7526, new_n7504, new_n7501);
nand_4 g07150(new_n7527, new_n7526, new_n7525);
nand_4 g07151(new_n7528, new_n7432, new_n7429);
nand_4 g07152(new_n7529, new_n7444, new_n7434);
nand_4 g07153(new_n7530, new_n7529, new_n7528);
nand_4 g07154(new_n7531, n11478, n2347);
not_3  g07155(new_n7532, new_n7531);
xnor_3 g07156(new_n7533, new_n7532, new_n7530);
nand_4 g07157(new_n7534, n3342, n1471);
not_3  g07158(new_n7535, new_n7534);
not_3  g07159(new_n7536, new_n7435);
nor_4  g07160(new_n7537, new_n7436_1, new_n7536);
nor_4  g07161(new_n7538, new_n7443, new_n7437);
nor_4  g07162(new_n7539, new_n7538, new_n7537);
not_3  g07163(new_n7540, new_n7387);
nor_4  g07164(new_n7541, new_n7389, new_n7540);
nor_4  g07165(new_n7542, new_n7390, new_n7386);
nor_4  g07166(new_n7543, new_n7542, new_n7541);
nand_4 g07167(new_n7544, n7236, n6431);
not_3  g07168(new_n7545, new_n7544);
nand_4 g07169(new_n7546_1, n9111, n7646);
nand_4 g07170(new_n7547, n9763, n4722);
xor_3  g07171(new_n7548, new_n7547, new_n7546_1);
xnor_3 g07172(new_n7549, new_n7548, new_n7545);
xnor_3 g07173(new_n7550, new_n7549, new_n7543);
xnor_3 g07174(new_n7551, new_n7550, new_n7539);
xnor_3 g07175(new_n7552, new_n7551, new_n7535);
not_3  g07176(new_n7553, new_n7391);
nand_4 g07177(new_n7554, new_n7553, new_n7384);
nand_4 g07178(new_n7555, new_n7406, new_n7392);
nand_4 g07179(new_n7556, new_n7555, new_n7554);
nand_4 g07180(new_n7557, new_n7395, new_n7393);
nand_4 g07181(new_n7558, new_n7405, new_n7396);
nand_4 g07182(new_n7559, new_n7558, new_n7557);
nand_4 g07183(new_n7560, n10217, n9400);
not_3  g07184(new_n7561, new_n7560);
xnor_3 g07185(new_n7562, new_n7561, new_n7559);
nand_4 g07186(new_n7563, n9189, n4203);
not_3  g07187(new_n7564, new_n7563);
nand_4 g07188(new_n7565, n4187, n2522);
nand_4 g07189(new_n7566, n12145, n11311);
xor_3  g07190(new_n7567, new_n7566, new_n7565);
xnor_3 g07191(new_n7568_1, new_n7567, new_n7564);
nand_4 g07192(new_n7569, n7823, n6877);
nand_4 g07193(new_n7570, n12753, n2024);
not_3  g07194(new_n7571, new_n7570);
xor_3  g07195(new_n7572, new_n7571, new_n7569);
xnor_3 g07196(new_n7573, new_n7572, new_n7568_1);
not_3  g07197(new_n7574, new_n7397);
nand_4 g07198(new_n7575, new_n7403, new_n7574);
and_4  g07199(new_n7576, new_n7575, new_n7402);
nand_4 g07200(new_n7577, n10174, n7946);
nand_4 g07201(new_n7578, n12221, n2464);
xor_3  g07202(new_n7579, new_n7578, new_n7577);
xnor_3 g07203(new_n7580, new_n7579, new_n7576);
xnor_3 g07204(new_n7581, new_n7580, new_n7573);
xnor_3 g07205(new_n7582, new_n7581, new_n7562);
xnor_3 g07206(new_n7583, new_n7582, new_n7556);
xnor_3 g07207(new_n7584, new_n7583, new_n7552);
xnor_3 g07208(new_n7585, new_n7584, new_n7533);
nand_4 g07209(new_n7586, new_n7464, new_n7463);
not_3  g07210(new_n7587, new_n7492);
nand_4 g07211(new_n7588, new_n7587, new_n7466);
nand_4 g07212(new_n7589, new_n7588, new_n7586);
nand_4 g07213(new_n7590, new_n7411, new_n7409);
nand_4 g07214(new_n7591, new_n7413, new_n7407);
nand_4 g07215(new_n7592, new_n7591, new_n7590);
xnor_3 g07216(new_n7593, new_n7592, new_n7589);
xnor_3 g07217(new_n7594, new_n7593, new_n7585);
not_3  g07218(new_n7595, new_n7439);
nor_4  g07219(new_n7596, new_n7441, new_n7595);
not_3  g07220(new_n7597, new_n7438);
nor_4  g07221(new_n7598, new_n7442, new_n7597);
or_4   g07222(new_n7599, new_n7598, new_n7596);
nand_4 g07223(new_n7600, new_n7493, new_n7458);
nand_4 g07224(new_n7601, new_n7499, new_n7494);
nand_4 g07225(new_n7602, new_n7601, new_n7600);
xnor_3 g07226(new_n7603, new_n7602, new_n7599);
xnor_3 g07227(new_n7604, new_n7603, new_n7594);
xnor_3 g07228(new_n7605, new_n7604, new_n7527);
nor_4  g07229(new_n7606, new_n7414, new_n7381);
nor_4  g07230(new_n7607, new_n7420, new_n7415);
nor_4  g07231(new_n7608, new_n7607, new_n7606);
not_3  g07232(new_n7609, new_n7098);
nand_4 g07233(new_n7610_1, new_n7128, new_n7609);
nand_4 g07234(new_n7611, new_n7141, new_n7129);
nand_4 g07235(new_n7612, new_n7611, new_n7610_1);
nand_4 g07236(new_n7613, new_n7125, new_n7124);
not_3  g07237(new_n7614, new_n7122);
nand_4 g07238(new_n7615, new_n7127, new_n7614);
nand_4 g07239(new_n7616, new_n7615, new_n7613);
not_3  g07240(new_n7617, new_n7425);
nor_4  g07241(new_n7618, new_n7427, new_n7617);
not_3  g07242(new_n7619, new_n7424);
nor_4  g07243(new_n7620, new_n7428, new_n7619);
nor_4  g07244(new_n7621, new_n7620, new_n7618);
nor_4  g07245(new_n7622, new_n7106, new_n7101);
nor_4  g07246(new_n7623, new_n7120, new_n7107);
nor_4  g07247(new_n7624, new_n7623, new_n7622);
nand_4 g07248(new_n7625, n7862, n2512);
not_3  g07249(new_n7626, new_n7108);
nand_4 g07250(new_n7627, new_n7109, new_n7626);
nand_4 g07251(new_n7628, new_n7119, new_n7111);
nand_4 g07252(new_n7629, new_n7628, new_n7627);
xnor_3 g07253(new_n7630, new_n7629, new_n7625);
nor_4  g07254(new_n7631, new_n7104, new_n7103);
not_3  g07255(new_n7632, new_n7102);
nand_4 g07256(new_n7633, new_n7104, new_n7103);
nand_4 g07257(new_n7634, new_n7633, new_n7632);
not_3  g07258(new_n7635, new_n7634);
nor_4  g07259(new_n7636, new_n7635, new_n7631);
nand_4 g07260(new_n7637, n11821, n10223);
nand_4 g07261(new_n7638, n5240, n4634);
nand_4 g07262(new_n7639, n9080, n2879);
xnor_3 g07263(new_n7640, new_n7639, new_n7638);
and_4  g07264(new_n7641, new_n7640, new_n7637);
nor_4  g07265(new_n7642, new_n7640, new_n7637);
nor_4  g07266(new_n7643, new_n7642, new_n7641);
xnor_3 g07267(new_n7644, new_n7643, new_n7636);
and_4  g07268(new_n7645, new_n7115, new_n7114);
nor_4  g07269(new_n7646_1, new_n7118, new_n7645);
nand_4 g07270(new_n7647, n11757, n9195);
not_3  g07271(new_n7648, new_n7647);
nand_4 g07272(new_n7649, n3172, n2253);
nand_4 g07273(new_n7650, n3865, n1333);
xnor_3 g07274(new_n7651, new_n7650, new_n7649);
xnor_3 g07275(new_n7652, new_n7651, new_n7648);
xnor_3 g07276(new_n7653, new_n7652, new_n7646_1);
xnor_3 g07277(new_n7654, new_n7653, new_n7644);
xnor_3 g07278(new_n7655, new_n7654, new_n7630);
xnor_3 g07279(new_n7656, new_n7655, new_n7624);
xnor_3 g07280(new_n7657, new_n7656, new_n7621);
not_3  g07281(new_n7658, new_n7484);
nand_4 g07282(new_n7659, new_n7490, new_n7658);
nand_4 g07283(new_n7660, new_n7491, new_n7480);
nand_4 g07284(new_n7661, new_n7660, new_n7659);
nand_4 g07285(new_n7662, n5798, n5283);
nand_4 g07286(new_n7663, n7265, n6826);
nand_4 g07287(new_n7664, n6294, n521);
xor_3  g07288(new_n7665, new_n7664, new_n7663);
xor_3  g07289(new_n7666, new_n7665, new_n7662);
xnor_3 g07290(new_n7667, new_n7666, new_n7661);
xnor_3 g07291(new_n7668, new_n7667, new_n7657);
xnor_3 g07292(new_n7669, new_n7668, new_n7616);
xnor_3 g07293(new_n7670, new_n7669, new_n7612);
xnor_3 g07294(new_n7671, new_n7670, new_n7608);
nand_4 g07295(new_n7672, new_n7450, new_n7448);
nand_4 g07296(new_n7673, new_n7452, new_n7445);
nand_4 g07297(new_n7674, new_n7673, new_n7672);
nand_4 g07298(new_n7675, n6797, n5579);
not_3  g07299(new_n7676_1, new_n7675);
nand_4 g07300(new_n7677, new_n7469, new_n7467);
nand_4 g07301(new_n7678, new_n7479, new_n7470);
nand_4 g07302(new_n7679, new_n7678, new_n7677);
xor_3  g07303(new_n7680, new_n7679, new_n7676_1);
nand_4 g07304(new_n7681, n4805, n1576);
nand_4 g07305(new_n7682, n3992, n2507);
xor_3  g07306(new_n7683, new_n7682, new_n7681);
nand_4 g07307(new_n7684, n3146, n2498);
nand_4 g07308(new_n7685, n6016, n137);
xor_3  g07309(new_n7686, new_n7685, new_n7684);
xor_3  g07310(new_n7687, new_n7686, new_n7683);
nand_4 g07311(new_n7688, n8384, n5153);
nand_4 g07312(new_n7689, n7270, n6358);
xor_3  g07313(new_n7690_1, new_n7689, new_n7688);
not_3  g07314(new_n7691, new_n7471);
nand_4 g07315(new_n7692, new_n7474, new_n7691);
and_4  g07316(new_n7693, new_n7692, new_n7477);
xor_3  g07317(new_n7694, new_n7693, new_n7690_1);
xnor_3 g07318(new_n7695, new_n7694, new_n7687);
not_3  g07319(new_n7696, new_n7486);
nor_4  g07320(new_n7697, new_n7488, new_n7696);
not_3  g07321(new_n7698, new_n7485);
nor_4  g07322(new_n7699, new_n7489, new_n7698);
nor_4  g07323(new_n7700, new_n7699, new_n7697);
nand_4 g07324(new_n7701, n4938, n2558);
nand_4 g07325(new_n7702, n5198, n806);
xor_3  g07326(new_n7703, new_n7702, new_n7701);
xor_3  g07327(new_n7704, new_n7703, new_n7700);
xnor_3 g07328(new_n7705, new_n7704, new_n7695);
xnor_3 g07329(new_n7706, new_n7705, new_n7680);
xnor_3 g07330(new_n7707, new_n7706, new_n7674);
xnor_3 g07331(new_n7708, new_n7707, new_n7671);
xnor_3 g07332(new_n7709, new_n7708, new_n7605);
xnor_3 g07333(new_n7710, new_n7709, new_n7523_1);
xnor_3 g07334(n2383, new_n7710, new_n7514);
not_3  g07335(new_n7712, new_n6272);
xor_3  g07336(n2425, new_n6282, new_n7712);
not_3  g07337(new_n7714, new_n3043);
nor_4  g07338(new_n7715, new_n7714, new_n3041);
xnor_3 g07339(n2431, new_n7715, new_n3093);
xnor_3 g07340(n2434, new_n2187, new_n2186);
not_3  g07341(new_n7718, new_n5266);
xor_3  g07342(n2581, new_n5267, new_n7718);
nand_4 g07343(new_n7720, new_n7026, new_n7025);
xnor_3 g07344(n2624, new_n7720, new_n7037);
nand_4 g07345(new_n7722, n6126, n2226);
nand_4 g07346(new_n7723, n3602, n1094);
nand_4 g07347(new_n7724, n10678, n3719);
not_3  g07348(new_n7725, new_n7724);
xor_3  g07349(new_n7726, new_n7725, new_n7723);
xnor_3 g07350(new_n7727, new_n7726, new_n7722);
and_4  g07351(new_n7728, new_n4487, new_n4486);
nor_4  g07352(new_n7729, new_n4488, new_n4485);
nor_4  g07353(new_n7730_1, new_n7729, new_n7728);
xnor_3 g07354(new_n7731, new_n7730_1, new_n7727);
nand_4 g07355(new_n7732, n10928, n10439);
nand_4 g07356(new_n7733_1, n8595, n6986);
xor_3  g07357(new_n7734, new_n7733_1, new_n7732);
xnor_3 g07358(new_n7735, new_n7734, new_n7731);
and_4  g07359(new_n7736, new_n4481, new_n4476);
nor_4  g07360(new_n7737, new_n4489, new_n4483);
nor_4  g07361(new_n7738, new_n7737, new_n7736);
xnor_3 g07362(new_n7739, new_n7738, new_n7735);
nand_4 g07363(new_n7740, new_n4473, new_n4472);
nand_4 g07364(new_n7741, new_n4494, new_n4493);
nand_4 g07365(new_n7742, new_n7741, new_n7740);
not_3  g07366(new_n7743, new_n7742);
nor_4  g07367(new_n7744, new_n7743, new_n7739);
not_3  g07368(new_n7745, new_n7722);
not_3  g07369(new_n7746, new_n7726);
nor_4  g07370(new_n7747, new_n7746, new_n7745);
nor_4  g07371(new_n7748, new_n7730_1, new_n7727);
nor_4  g07372(new_n7749, new_n7748, new_n7747);
nand_4 g07373(new_n7750, n10928, n8065);
nand_4 g07374(new_n7751, n10439, n6986);
nand_4 g07375(new_n7752, n10391, n8336);
not_3  g07376(new_n7753, new_n7752);
xor_3  g07377(new_n7754, new_n7753, new_n7751);
xnor_3 g07378(new_n7755, new_n7754, new_n7750);
xnor_3 g07379(new_n7756, new_n7755, new_n7749);
nor_4  g07380(new_n7757, new_n7724, new_n7723);
nand_4 g07381(new_n7758, n8595, n2226);
not_3  g07382(new_n7759, new_n7758);
xor_3  g07383(new_n7760, new_n7759, new_n7757);
not_3  g07384(new_n7761, new_n7760);
nand_4 g07385(new_n7762, n10678, n3602);
nand_4 g07386(new_n7763, n6126, n1094);
nand_4 g07387(new_n7764, n7320, n3719);
not_3  g07388(new_n7765, new_n7764);
xor_3  g07389(new_n7766, new_n7765, new_n7763);
xnor_3 g07390(new_n7767, new_n7766, new_n7762);
not_3  g07391(new_n7768, new_n7767);
xor_3  g07392(new_n7769, new_n7768, new_n7761);
xnor_3 g07393(new_n7770, new_n7769, new_n7756);
not_3  g07394(new_n7771, new_n7770);
nand_4 g07395(new_n7772, new_n7734, new_n7731);
nor_4  g07396(new_n7773, new_n7733_1, new_n7732);
not_3  g07397(new_n7774, new_n7773);
not_3  g07398(new_n7775, new_n7734);
xnor_3 g07399(new_n7776, new_n7775, new_n7731);
not_3  g07400(new_n7777, new_n7738);
nand_4 g07401(new_n7778, new_n7777, new_n7776);
xnor_3 g07402(new_n7779, new_n7778, new_n7774);
nand_4 g07403(new_n7780, new_n7779, new_n7772);
xnor_3 g07404(new_n7781, new_n7780, new_n7771);
xnor_3 g07405(new_n7782, new_n7781, new_n7744);
nand_4 g07406(new_n7783, n8336, n8065);
xnor_3 g07407(new_n7784, new_n7743, new_n7739);
nand_4 g07408(new_n7785, new_n7784, new_n7783);
nand_4 g07409(new_n7786, new_n4496, new_n4470);
xnor_3 g07410(new_n7787, new_n7742, new_n7739);
xnor_3 g07411(new_n7788, new_n7787, new_n7783);
nand_4 g07412(new_n7789, new_n7788, new_n7786);
nand_4 g07413(new_n7790, new_n7789, new_n7785);
xnor_3 g07414(new_n7791, new_n7790, new_n7782);
nand_4 g07415(new_n7792, n7160, n4826);
nand_4 g07416(new_n7793, n7733, n4828);
nand_4 g07417(new_n7794, n12925, n2515);
xnor_3 g07418(new_n7795, new_n7794, new_n7793);
nor_4  g07419(new_n7796, new_n7795, new_n7792);
not_3  g07420(new_n7797, new_n7792);
not_3  g07421(new_n7798, new_n7795);
nor_4  g07422(new_n7799, new_n7798, new_n7797);
nor_4  g07423(new_n7800, new_n7799, new_n7796);
not_3  g07424(new_n7801, new_n4540);
not_3  g07425(new_n7802, new_n4541);
nor_4  g07426(new_n7803, new_n7802, new_n7801);
not_3  g07427(new_n7804, new_n4539);
nor_4  g07428(new_n7805, new_n4542, new_n7804);
nor_4  g07429(new_n7806, new_n7805, new_n7803);
xnor_3 g07430(new_n7807, new_n7806, new_n7800);
not_3  g07431(new_n7808, new_n7807);
nand_4 g07432(new_n7809, n12391, n4970);
nand_4 g07433(new_n7810, n7891, n7610);
xor_3  g07434(new_n7811, new_n7810, new_n7809);
xnor_3 g07435(new_n7812, new_n7811, new_n7808);
nand_4 g07436(new_n7813, new_n4537, new_n4535);
not_3  g07437(new_n7814, new_n7813);
nor_4  g07438(new_n7815, new_n4543, new_n4538);
nor_4  g07439(new_n7816, new_n7815, new_n7814);
xnor_3 g07440(new_n7817, new_n7816, new_n7812);
nor_4  g07441(new_n7818, new_n4544, new_n4533);
nor_4  g07442(new_n7819, new_n4548, new_n4545);
nor_4  g07443(new_n7820, new_n7819, new_n7818);
nor_4  g07444(new_n7821, new_n7820, new_n7817);
not_3  g07445(new_n7822, new_n7821);
not_3  g07446(new_n7823_1, new_n7796);
nand_4 g07447(new_n7824, new_n7806, new_n7800);
nand_4 g07448(new_n7825, new_n7824, new_n7823_1);
nand_4 g07449(new_n7826, n12391, n503);
not_3  g07450(new_n7827, new_n7826);
nand_4 g07451(new_n7828, n7891, n4970);
nand_4 g07452(new_n7829, n12069, n10965);
xnor_3 g07453(new_n7830, new_n7829, new_n7828);
xor_3  g07454(new_n7831, new_n7830, new_n7827);
xnor_3 g07455(new_n7832, new_n7831, new_n7825);
nor_4  g07456(new_n7833, new_n7794, new_n7793);
not_3  g07457(new_n7834, new_n7833);
nand_4 g07458(new_n7835, n7610, n7160);
xor_3  g07459(new_n7836, new_n7835, new_n7834);
nand_4 g07460(new_n7837, n7733, n2515);
not_3  g07461(new_n7838, new_n7837);
nand_4 g07462(new_n7839, n4828, n4826);
nand_4 g07463(new_n7840, n12925, n1199);
xnor_3 g07464(new_n7841, new_n7840, new_n7839);
xor_3  g07465(new_n7842, new_n7841, new_n7838);
xnor_3 g07466(new_n7843, new_n7842, new_n7836);
xnor_3 g07467(new_n7844, new_n7843, new_n7832);
nand_4 g07468(new_n7845, new_n7811, new_n7808);
nor_4  g07469(new_n7846, new_n7810, new_n7809);
xnor_3 g07470(new_n7847, new_n7811, new_n7807);
not_3  g07471(new_n7848, new_n7816);
nand_4 g07472(new_n7849, new_n7848, new_n7847);
not_3  g07473(new_n7850, new_n7849);
xnor_3 g07474(new_n7851, new_n7850, new_n7846);
nand_4 g07475(new_n7852, new_n7851, new_n7845);
xnor_3 g07476(new_n7853, new_n7852, new_n7844);
xnor_3 g07477(new_n7854, new_n7853, new_n7822);
nand_4 g07478(new_n7855, n12069, n503);
not_3  g07479(new_n7856, new_n7855);
not_3  g07480(new_n7857, new_n7817);
xnor_3 g07481(new_n7858, new_n7820, new_n7857);
nand_4 g07482(new_n7859, new_n7858, new_n7856);
nor_4  g07483(new_n7860, new_n4549, new_n4532);
xnor_3 g07484(new_n7861, new_n7858, new_n7855);
nand_4 g07485(new_n7862_1, new_n7861, new_n7860);
nand_4 g07486(new_n7863, new_n7862_1, new_n7859);
xnor_3 g07487(new_n7864, new_n7863, new_n7854);
nand_4 g07488(new_n7865, n11222, n6359);
not_3  g07489(new_n7866, new_n7865);
nand_4 g07490(new_n7867, n4086, n996);
nand_4 g07491(new_n7868, n5767, n405);
nand_4 g07492(new_n7869, n8433, n5319);
xnor_3 g07493(new_n7870, new_n7869, new_n7868);
nor_4  g07494(new_n7871, new_n7870, new_n7867);
not_3  g07495(new_n7872, new_n7867);
not_3  g07496(new_n7873, new_n7870);
nor_4  g07497(new_n7874, new_n7873, new_n7872);
nor_4  g07498(new_n7875, new_n7874, new_n7871);
not_3  g07499(new_n7876, new_n4502);
nor_4  g07500(new_n7877, new_n4508, new_n7876);
nor_4  g07501(new_n7878, new_n7877, new_n4507);
xnor_3 g07502(new_n7879, new_n7878, new_n7875);
nand_4 g07503(new_n7880, n11153, n6611);
nand_4 g07504(new_n7881, n5314, n217);
xor_3  g07505(new_n7882, new_n7881, new_n7880);
xnor_3 g07506(new_n7883, new_n7882, new_n7879);
not_3  g07507(new_n7884, new_n4501);
nand_4 g07508(new_n7885, new_n4510, new_n7884);
nand_4 g07509(new_n7886, new_n4517, new_n4511);
nand_4 g07510(new_n7887, new_n7886, new_n7885);
xnor_3 g07511(new_n7888, new_n7887, new_n7883);
not_3  g07512(new_n7889, new_n4526);
nand_4 g07513(new_n7890, new_n7889, new_n4521);
nand_4 g07514(new_n7891_1, new_n7890, new_n4519);
not_3  g07515(new_n7892, new_n7891_1);
nor_4  g07516(new_n7893, new_n7892, new_n7888);
not_3  g07517(new_n7894, new_n7888);
nor_4  g07518(new_n7895, new_n7891_1, new_n7894);
nor_4  g07519(new_n7896, new_n7895, new_n7893);
nand_4 g07520(new_n7897, new_n7896, new_n7866);
xnor_3 g07521(new_n7898, new_n7896, new_n7865);
nand_4 g07522(new_n7899, new_n7898, new_n4528);
nand_4 g07523(new_n7900, new_n7899, new_n7897);
nor_4  g07524(new_n7901, new_n7869, new_n7868);
nand_4 g07525(new_n7902, n996, n217);
not_3  g07526(new_n7903, new_n7902);
xor_3  g07527(new_n7904, new_n7903, new_n7901);
not_3  g07528(new_n7905, new_n7904);
nand_4 g07529(new_n7906, n5319, n405);
not_3  g07530(new_n7907, new_n7906);
nand_4 g07531(new_n7908, n5767, n4086);
nand_4 g07532(new_n7909, n9457, n8433);
xnor_3 g07533(new_n7910, new_n7909, new_n7908);
xor_3  g07534(new_n7911, new_n7910, new_n7907);
nor_4  g07535(new_n7912, new_n7911, new_n7905);
not_3  g07536(new_n7913, new_n7911);
nor_4  g07537(new_n7914, new_n7913, new_n7904);
nor_4  g07538(new_n7915, new_n7914, new_n7912);
nand_4 g07539(new_n7916, new_n7878, new_n7875);
not_3  g07540(new_n7917, new_n7916);
nor_4  g07541(new_n7918, new_n7917, new_n7871);
not_3  g07542(new_n7919, new_n7918);
nand_4 g07543(new_n7920, n11153, n6359);
not_3  g07544(new_n7921, new_n7920);
nand_4 g07545(new_n7922, n6611, n5314);
nand_4 g07546(new_n7923, n11296, n11222);
nand_4 g07547(new_n7924, new_n7923, new_n7922);
not_3  g07548(new_n7925, new_n7922);
not_3  g07549(new_n7926, new_n7923);
nand_4 g07550(new_n7927, new_n7926, new_n7925);
nand_4 g07551(new_n7928, new_n7927, new_n7924);
xor_3  g07552(new_n7929, new_n7928, new_n7921);
xnor_3 g07553(new_n7930, new_n7929, new_n7919);
xnor_3 g07554(new_n7931, new_n7930, new_n7915);
not_3  g07555(new_n7932, new_n7879);
nand_4 g07556(new_n7933, new_n7882, new_n7932);
nor_4  g07557(new_n7934, new_n7881, new_n7880);
nand_4 g07558(new_n7935, new_n7887, new_n7883);
not_3  g07559(new_n7936, new_n7935);
xnor_3 g07560(new_n7937, new_n7936, new_n7934);
nand_4 g07561(new_n7938, new_n7937, new_n7933);
xnor_3 g07562(new_n7939, new_n7938, new_n7931);
xnor_3 g07563(new_n7940, new_n7939, new_n7893);
xnor_3 g07564(new_n7941, new_n7940, new_n7900);
xnor_3 g07565(new_n7942, new_n7941, new_n7864);
xnor_3 g07566(new_n7943, new_n7861, new_n7860);
not_3  g07567(new_n7944, new_n7943);
not_3  g07568(new_n7945, new_n4528);
xnor_3 g07569(new_n7946_1, new_n7898, new_n7945);
nor_4  g07570(new_n7947, new_n7946_1, new_n7944);
not_3  g07571(new_n7948, new_n4550);
not_3  g07572(new_n7949, new_n4554);
nor_4  g07573(new_n7950, new_n7949, new_n7948);
nor_4  g07574(new_n7951, new_n4555, new_n4531);
nor_4  g07575(new_n7952, new_n7951, new_n7950);
xnor_3 g07576(new_n7953, new_n7946_1, new_n7944);
nor_4  g07577(new_n7954, new_n7953, new_n7952);
nor_4  g07578(new_n7955, new_n7954, new_n7947);
xnor_3 g07579(new_n7956, new_n7955, new_n7942);
nand_4 g07580(new_n7957, new_n7956, new_n7791);
xnor_3 g07581(new_n7958, new_n7956, new_n7791);
not_3  g07582(new_n7959, new_n7958);
not_3  g07583(new_n7960, new_n7783);
nand_4 g07584(new_n7961, new_n7787, new_n7960);
nand_4 g07585(new_n7962, new_n7961, new_n7785);
xnor_3 g07586(new_n7963, new_n7962, new_n7786);
xnor_3 g07587(new_n7964, new_n7953, new_n7952);
not_3  g07588(new_n7965_1, new_n7964);
nand_4 g07589(new_n7966_1, new_n7965_1, new_n7963);
xnor_3 g07590(new_n7967, new_n7964, new_n7963);
nor_4  g07591(new_n7968, new_n4557, new_n4497);
not_3  g07592(new_n7969, new_n4563);
nor_4  g07593(new_n7970, new_n7969, new_n4558);
nor_4  g07594(new_n7971, new_n7970, new_n7968);
nand_4 g07595(new_n7972, new_n7971, new_n7967);
nand_4 g07596(new_n7973, new_n7972, new_n7966_1);
nand_4 g07597(new_n7974, new_n7973, new_n7959);
nand_4 g07598(new_n7975, new_n7974, new_n7957);
nand_4 g07599(new_n7976, new_n7781, new_n7744);
not_3  g07600(new_n7977, new_n7976);
nor_4  g07601(new_n7978, new_n7790, new_n7782);
nor_4  g07602(new_n7979, new_n7978, new_n7977);
xnor_3 g07603(new_n7980, new_n7979, new_n7975);
not_3  g07604(new_n7981_1, new_n7941);
nand_4 g07605(new_n7982, new_n7981_1, new_n7864);
not_3  g07606(new_n7983, new_n7947);
not_3  g07607(new_n7984, new_n7952);
xnor_3 g07608(new_n7985, new_n7946_1, new_n7943);
nand_4 g07609(new_n7986, new_n7985, new_n7984);
nand_4 g07610(new_n7987, new_n7986, new_n7983);
nand_4 g07611(new_n7988, new_n7987, new_n7942);
nand_4 g07612(new_n7989, new_n7988, new_n7982);
nand_4 g07613(new_n7990, new_n7853, new_n7821);
nand_4 g07614(new_n7991, new_n7863, new_n7854);
nand_4 g07615(new_n7992, new_n7991, new_n7990);
and_4  g07616(new_n7993, new_n7909, new_n7908);
nor_4  g07617(new_n7994, new_n7910, new_n7907);
nor_4  g07618(new_n7995, new_n7994, new_n7993);
nand_4 g07619(new_n7996, n11296, n11153);
xor_3  g07620(new_n7997, new_n7996, new_n7995);
not_3  g07621(new_n7998, new_n7751);
nor_4  g07622(new_n7999, new_n7753, new_n7998);
not_3  g07623(new_n8000, new_n7750);
nor_4  g07624(new_n8001, new_n7754, new_n8000);
nor_4  g07625(new_n8002, new_n8001, new_n7999);
nand_4 g07626(new_n8003, n6611, n996);
nand_4 g07627(new_n8004, n6359, n5314);
xor_3  g07628(new_n8005, new_n8004, new_n8003);
nand_4 g07629(new_n8006, n12069, n7546);
nand_4 g07630(new_n8007, n12925, n6578);
xor_3  g07631(new_n8008, new_n8007, new_n8006);
xnor_3 g07632(new_n8009, new_n8008, new_n8005);
nand_4 g07633(new_n8010, n7733, n1199);
nand_4 g07634(new_n8011, n7160, n4970);
not_3  g07635(new_n8012, new_n8011);
xor_3  g07636(new_n8013, new_n8012, new_n8010);
xnor_3 g07637(new_n8014, new_n8013, new_n8009);
xnor_3 g07638(new_n8015, new_n8014, new_n8002);
nand_4 g07639(new_n8016, new_n7903, new_n7901);
nand_4 g07640(new_n8017, new_n7913, new_n7904);
nand_4 g07641(new_n8018, new_n8017, new_n8016);
nand_4 g07642(new_n8019, n5767, n217);
nand_4 g07643(new_n8020, new_n7924, new_n7921);
nand_4 g07644(new_n8021, new_n8020, new_n7927);
xor_3  g07645(new_n8022, new_n8021, new_n8019);
xor_3  g07646(new_n8023, new_n8022, new_n8018);
xnor_3 g07647(new_n8024, new_n8023, new_n8015);
xnor_3 g07648(new_n8025, new_n8024, new_n7997);
nand_4 g07649(new_n8026, new_n7929, new_n7918);
not_3  g07650(new_n8027, new_n7915);
nand_4 g07651(new_n8028_1, new_n7930, new_n8027);
nand_4 g07652(new_n8029, new_n8028_1, new_n8026);
nand_4 g07653(new_n8030, n7610, n4828);
nand_4 g07654(new_n8031, n4826, n2515);
not_3  g07655(new_n8032, new_n8031);
xor_3  g07656(new_n8033, new_n8032, new_n8030);
xnor_3 g07657(new_n8034, new_n8033, new_n8029);
nand_4 g07658(new_n8035, n4921, n4516);
nand_4 g07659(new_n8036, n2564, n1835);
xor_3  g07660(new_n8037, new_n8036, new_n8035);
xnor_3 g07661(new_n8038, new_n8037, new_n8034);
xnor_3 g07662(new_n8039, new_n8038, new_n8025);
xnor_3 g07663(new_n8040, new_n8039, new_n7992);
xnor_3 g07664(new_n8041, new_n8040, new_n7989);
nand_4 g07665(new_n8042, new_n7939, new_n7893);
not_3  g07666(new_n8043, new_n7940);
nand_4 g07667(new_n8044, new_n8043, new_n7900);
nand_4 g07668(new_n8045, new_n8044, new_n8042);
nand_4 g07669(new_n8046, new_n7850, new_n7846);
not_3  g07670(new_n8047, new_n7844);
nand_4 g07671(new_n8048, new_n7852, new_n8047);
nand_4 g07672(new_n8049, new_n8048, new_n8046);
nand_4 g07673(new_n8050, n4189, n2577);
not_3  g07674(new_n8051, new_n8050);
nand_4 g07675(new_n8052, n6687, n1835);
not_3  g07676(new_n8053, new_n8052);
nor_4  g07677(new_n8054, new_n8053, new_n8051);
nand_4 g07678(new_n8055, n9637, n2564);
not_3  g07679(new_n8056, new_n8055);
xor_3  g07680(new_n8057, new_n8053, new_n8050);
nor_4  g07681(new_n8058, new_n8057, new_n8056);
nor_4  g07682(new_n8059, new_n8058, new_n8054);
xnor_3 g07683(new_n8060, new_n8059, new_n8049);
nand_4 g07684(new_n8061, n11917, n6770);
not_3  g07685(new_n8062, new_n8061);
nand_4 g07686(new_n8063, n9920, n4921);
nand_4 g07687(new_n8064, n9956, n3627);
not_3  g07688(new_n8065_1, new_n8064);
xor_3  g07689(new_n8066, new_n8065_1, new_n8063);
not_3  g07690(new_n8067, new_n8066);
nor_4  g07691(new_n8068, new_n8067, new_n8062);
xor_3  g07692(new_n8069, new_n8067, new_n8062);
not_3  g07693(new_n8070, new_n8069);
not_3  g07694(new_n8071, new_n4263);
nor_4  g07695(new_n8072, new_n4265, new_n8071);
not_3  g07696(new_n8073, new_n4262);
nor_4  g07697(new_n8074, new_n4266, new_n8073);
nor_4  g07698(new_n8075, new_n8074, new_n8072);
nor_4  g07699(new_n8076, new_n8075, new_n8070);
nor_4  g07700(new_n8077, new_n8076, new_n8068);
xnor_3 g07701(new_n8078, new_n8057, new_n8055);
not_3  g07702(new_n8079, new_n8078);
nand_4 g07703(new_n8080, new_n8079, new_n8077);
nor_4  g07704(new_n8081, new_n8064, new_n8063);
nand_4 g07705(new_n8082, n6770, n3842);
xor_3  g07706(new_n8083, new_n8082, new_n8081);
nand_4 g07707(new_n8084, n4921, n3627);
nand_4 g07708(new_n8085, n11917, n9920);
nand_4 g07709(new_n8086, n9956, n4516);
not_3  g07710(new_n8087, new_n8086);
xor_3  g07711(new_n8088, new_n8087, new_n8085);
xnor_3 g07712(new_n8089, new_n8088, new_n8084);
not_3  g07713(new_n8090, new_n8089);
xor_3  g07714(new_n8091, new_n8090, new_n8083);
not_3  g07715(new_n8092, new_n8091);
xnor_3 g07716(new_n8093, new_n8078, new_n8077);
nand_4 g07717(new_n8094, new_n8093, new_n8092);
nand_4 g07718(new_n8095, new_n8094, new_n8080);
nand_4 g07719(new_n8096, n9920, n3842);
xnor_3 g07720(new_n8097, new_n8096, new_n8095);
xnor_3 g07721(new_n8098, new_n8097, new_n8060);
xnor_3 g07722(new_n8099, new_n8098, new_n8045);
nand_4 g07723(new_n8100_1, new_n7936, new_n7934);
not_3  g07724(new_n8101, new_n7931);
nand_4 g07725(new_n8102, new_n7938, new_n8101);
nand_4 g07726(new_n8103, new_n8102, new_n8100_1);
nand_4 g07727(new_n8104, new_n7759, new_n7757);
nand_4 g07728(new_n8105, new_n7768, new_n7760);
nand_4 g07729(new_n8106, new_n8105, new_n8104);
nand_4 g07730(new_n8107, n10439, n2226);
nand_4 g07731(new_n8108, n10678, n6126);
xor_3  g07732(new_n8109, new_n8108, new_n8107);
nand_4 g07733(new_n8110, n11222, n1357);
nand_4 g07734(new_n8111, n8433, n4817);
xor_3  g07735(new_n8112, new_n8111, new_n8110);
nand_4 g07736(new_n8113, n10928, n10391);
nand_4 g07737(new_n8114, n8595, n1094);
not_3  g07738(new_n8115, new_n8114);
xor_3  g07739(new_n8116, new_n8115, new_n8113);
xor_3  g07740(new_n8117, new_n8116, new_n8112);
xnor_3 g07741(new_n8118, new_n8117, new_n8109);
xnor_3 g07742(new_n8119, new_n8118, new_n8106);
not_3  g07743(new_n8120, new_n7763);
nor_4  g07744(new_n8121, new_n7765, new_n8120);
not_3  g07745(new_n8122, new_n7762);
nor_4  g07746(new_n8123, new_n7766, new_n8122);
nor_4  g07747(new_n8124, new_n8123, new_n8121);
nand_4 g07748(new_n8125, n9457, n405);
not_3  g07749(new_n8126, new_n8125);
xnor_3 g07750(new_n8127, new_n8126, new_n8124);
nand_4 g07751(new_n8128, n8065, n6986);
nand_4 g07752(new_n8129, n8336, n4190);
not_3  g07753(new_n8130, new_n8129);
xor_3  g07754(new_n8131, new_n8130, new_n8128);
nand_4 g07755(new_n8132, n7523, n3719);
nand_4 g07756(new_n8133, n7320, n3602);
xor_3  g07757(new_n8134, new_n8133, new_n8132);
xor_3  g07758(new_n8135, new_n8134, new_n8131);
xnor_3 g07759(new_n8136, new_n8135, new_n8127);
nand_4 g07760(new_n8137, n11536, n6687);
and_4  g07761(new_n8138_1, new_n7829, new_n7828);
nor_4  g07762(new_n8139, new_n7830, new_n7827);
nor_4  g07763(new_n8140, new_n8139, new_n8138_1);
xor_3  g07764(new_n8141, new_n8140, new_n8137);
xnor_3 g07765(new_n8142, new_n8141, new_n8136);
xnor_3 g07766(new_n8143, new_n8142, new_n8119);
xnor_3 g07767(new_n8144, new_n8143, new_n8103);
not_3  g07768(new_n8145, new_n7749);
nand_4 g07769(new_n8146, new_n7755, new_n8145);
nand_4 g07770(new_n8147, new_n7769, new_n7756);
nand_4 g07771(new_n8148, new_n8147, new_n8146);
not_3  g07772(new_n8149, new_n8082);
nor_4  g07773(new_n8150, new_n8149, new_n8081);
nor_4  g07774(new_n8151, new_n8090, new_n8083);
nor_4  g07775(new_n8152, new_n8151, new_n8150);
nand_4 g07776(new_n8153, n9637, n4189);
not_3  g07777(new_n8154, new_n8085);
nor_4  g07778(new_n8155, new_n8087, new_n8154);
not_3  g07779(new_n8156, new_n8084);
nor_4  g07780(new_n8157, new_n8088, new_n8156);
nor_4  g07781(new_n8158, new_n8157, new_n8155);
nand_4 g07782(new_n8159, n5319, n4086);
not_3  g07783(new_n8160, new_n8159);
nand_4 g07784(new_n8161, n6770, n2577);
nand_4 g07785(new_n8162, n11917, n3627);
xor_3  g07786(new_n8163, new_n8162, new_n8161);
xnor_3 g07787(new_n8164, new_n8163, new_n8160);
xnor_3 g07788(new_n8165, new_n8164, new_n8158);
xnor_3 g07789(new_n8166, new_n8165, new_n8153);
xnor_3 g07790(new_n8167, new_n8166, new_n8152);
nand_4 g07791(new_n8168, n9956, n2087);
nor_4  g07792(new_n8169, new_n7835, new_n7834);
not_3  g07793(new_n8170, new_n7836);
nor_4  g07794(new_n8171, new_n7842, new_n8170);
nor_4  g07795(new_n8172, new_n8171, new_n8169);
and_4  g07796(new_n8173, new_n7840, new_n7839);
nor_4  g07797(new_n8174, new_n7841, new_n7838);
nor_4  g07798(new_n8175, new_n8174, new_n8173);
nand_4 g07799(new_n8176, n12391, n10965);
nand_4 g07800(new_n8177, n7891, n503);
xor_3  g07801(new_n8178, new_n8177, new_n8176);
xnor_3 g07802(new_n8179, new_n8178, new_n8175);
xnor_3 g07803(new_n8180, new_n8179, new_n8172);
xnor_3 g07804(new_n8181, new_n8180, new_n8168);
xnor_3 g07805(new_n8182, new_n8181, new_n8167);
xnor_3 g07806(new_n8183, new_n8182, new_n8148);
not_3  g07807(new_n8184, new_n7778);
nand_4 g07808(new_n8185, new_n8184, new_n7773);
nand_4 g07809(new_n8186, new_n7780, new_n7770);
nand_4 g07810(new_n8187, new_n8186, new_n8185);
nand_4 g07811(new_n8188, n2577, n2564);
nand_4 g07812(new_n8189, n4189, n3842);
nor_4  g07813(new_n8190, new_n8189, new_n8188);
xnor_3 g07814(new_n8191, new_n8075, new_n8069);
not_3  g07815(new_n8192, new_n8191);
xor_3  g07816(new_n8193, new_n8189, new_n8188);
xnor_3 g07817(new_n8194, new_n8193, new_n8192);
not_3  g07818(new_n8195, new_n4257);
and_4  g07819(new_n8196, new_n4259, new_n8195);
nor_4  g07820(new_n8197, new_n4267, new_n4260);
nor_4  g07821(new_n8198, new_n8197, new_n8196);
nor_4  g07822(new_n8199, new_n8198, new_n8194);
nand_4 g07823(new_n8200, new_n8199, new_n8190);
xnor_3 g07824(new_n8201, new_n8093, new_n8091);
nand_4 g07825(new_n8202_1, new_n8193, new_n8192);
xnor_3 g07826(new_n8203, new_n8199, new_n8190);
nand_4 g07827(new_n8204, new_n8203, new_n8202_1);
nand_4 g07828(new_n8205, new_n8204, new_n8201);
nand_4 g07829(new_n8206, new_n8205, new_n8200);
xnor_3 g07830(new_n8207, new_n8206, new_n8187);
xnor_3 g07831(new_n8208, new_n8207, new_n8183);
xnor_3 g07832(new_n8209, new_n8208, new_n8144);
xnor_3 g07833(new_n8210, new_n8209, new_n8099);
xnor_3 g07834(new_n8211, new_n8210, new_n8041);
xnor_3 g07835(new_n8212, new_n8211, new_n7980);
xnor_3 g07836(new_n8213, new_n8198, new_n8194);
not_3  g07837(new_n8214, new_n4250);
nand_4 g07838(new_n8215, new_n4254, new_n8214);
nand_4 g07839(new_n8216, new_n4269, new_n4256);
nand_4 g07840(new_n8217, new_n8216, new_n8215);
not_3  g07841(new_n8218, new_n8217);
nor_4  g07842(new_n8219, new_n8218, new_n8213);
xnor_3 g07843(new_n8220, new_n8204, new_n8201);
xnor_3 g07844(new_n8221, new_n8220, new_n8219);
nand_4 g07845(new_n8222, n9637, n6687);
not_3  g07846(new_n8223, new_n8222);
not_3  g07847(new_n8224, new_n8213);
nor_4  g07848(new_n8225, new_n8217, new_n8224);
nor_4  g07849(new_n8226, new_n8225, new_n8219);
nand_4 g07850(new_n8227, new_n8226, new_n8223);
nor_4  g07851(new_n8228, new_n4270, new_n4249);
xnor_3 g07852(new_n8229, new_n8226, new_n8222);
nand_4 g07853(new_n8230, new_n8229, new_n8228);
nand_4 g07854(new_n8231, new_n8230, new_n8227);
xnor_3 g07855(new_n8232, new_n8231, new_n8221);
not_3  g07856(new_n8233, new_n8232);
xnor_3 g07857(new_n8234, new_n7973, new_n7958);
not_3  g07858(new_n8235, new_n8234);
nand_4 g07859(new_n8236_1, new_n8235, new_n8233);
nand_4 g07860(new_n8237, new_n8234, new_n8232);
not_3  g07861(new_n8238, new_n8229);
xnor_3 g07862(new_n8239, new_n8238, new_n8228);
not_3  g07863(new_n8240, new_n4271);
nand_4 g07864(new_n8241, new_n4467, new_n8240);
nand_4 g07865(new_n8242, new_n4564, new_n4468);
nand_4 g07866(new_n8243, new_n8242, new_n8241);
nor_4  g07867(new_n8244, new_n8243, new_n8239);
xnor_3 g07868(new_n8245, new_n7971, new_n7967);
xnor_3 g07869(new_n8246, new_n8243, new_n8239);
nor_4  g07870(new_n8247, new_n8246, new_n8245);
nor_4  g07871(new_n8248, new_n8247, new_n8244);
nand_4 g07872(new_n8249, new_n8248, new_n8237);
nand_4 g07873(new_n8250, new_n8249, new_n8236_1);
not_3  g07874(new_n8251, new_n8220);
nand_4 g07875(new_n8252, new_n8251, new_n8219);
nand_4 g07876(new_n8253, new_n8231, new_n8221);
nand_4 g07877(new_n8254, new_n8253, new_n8252);
not_3  g07878(new_n8255, new_n7831);
nor_4  g07879(new_n8256, new_n8255, new_n7825);
not_3  g07880(new_n8257, new_n7832);
nor_4  g07881(new_n8258, new_n7843, new_n8257);
nor_4  g07882(new_n8259, new_n8258, new_n8256);
xnor_3 g07883(new_n8260, new_n8259, new_n8254);
xnor_3 g07884(new_n8261, new_n8260, new_n8250);
xnor_3 g07885(n2679, new_n8261, new_n8212);
not_3  g07886(new_n8263, new_n6000);
nor_4  g07887(new_n8264, new_n8263, new_n5972);
nand_4 g07888(new_n8265, n6687, n2253);
not_3  g07889(new_n8266, new_n8265);
nand_4 g07890(new_n8267, n10223, n6770);
not_3  g07891(new_n8268, new_n8267);
nand_4 g07892(new_n8269, n9920, n2879);
nand_4 g07893(new_n8270, n7265, n3627);
xnor_3 g07894(new_n8271, new_n8270, new_n8269);
xnor_3 g07895(new_n8272, new_n8271, new_n8268);
not_3  g07896(new_n8273, new_n5977);
not_3  g07897(new_n8274, new_n5978);
nor_4  g07898(new_n8275, new_n8274, new_n8273);
not_3  g07899(new_n8276_1, new_n5976);
nor_4  g07900(new_n8277, new_n5979, new_n8276_1);
nor_4  g07901(new_n8278, new_n8277, new_n8275);
xnor_3 g07902(new_n8279, new_n8278, new_n8272);
not_3  g07903(new_n8280, new_n8279);
nand_4 g07904(new_n8281, n9195, n2564);
nand_4 g07905(new_n8282, n4634, n4189);
xor_3  g07906(new_n8283, new_n8282, new_n8281);
not_3  g07907(new_n8284, new_n8283);
xor_3  g07908(new_n8285, new_n8284, new_n8280);
nor_4  g07909(new_n8286, new_n5980, new_n5975);
not_3  g07910(new_n8287, new_n5986);
nor_4  g07911(new_n8288, new_n8287, new_n5981);
nor_4  g07912(new_n8289, new_n8288, new_n8286);
xnor_3 g07913(new_n8290, new_n8289, new_n8285);
not_3  g07914(new_n8291, new_n5989);
nand_4 g07915(new_n8292, new_n5997, new_n8291);
xnor_3 g07916(new_n8293, new_n8292, new_n8290);
xnor_3 g07917(new_n8294, new_n8293, new_n8266);
xor_3  g07918(new_n8295, new_n8294, new_n8264);
not_3  g07919(new_n8296, new_n6001);
nand_4 g07920(new_n8297, new_n6254_1, new_n8296);
nand_4 g07921(new_n8298, new_n6287, new_n6255);
nand_4 g07922(new_n8299, new_n8298, new_n8297);
xnor_3 g07923(new_n8300, new_n8299, new_n8295);
nor_4  g07924(new_n8301, new_n6054, new_n6031);
nand_4 g07925(new_n8302, n12221, n8336);
not_3  g07926(new_n8303_1, new_n8302);
nand_4 g07927(new_n8304, n9189, n2226);
nand_4 g07928(new_n8305, n2024, n1094);
nand_4 g07929(new_n8306, n10678, n7946);
xnor_3 g07930(new_n8307, new_n8306, new_n8305);
nor_4  g07931(new_n8308, new_n8307, new_n8304);
not_3  g07932(new_n8309, new_n8304);
not_3  g07933(new_n8310, new_n8307);
nor_4  g07934(new_n8311, new_n8310, new_n8309);
nor_4  g07935(new_n8312, new_n8311, new_n8308);
not_3  g07936(new_n8313, new_n6041);
not_3  g07937(new_n8314, new_n6042);
nor_4  g07938(new_n8315, new_n8314, new_n8313);
nor_4  g07939(new_n8316, new_n6043, new_n6040);
nor_4  g07940(new_n8317, new_n8316, new_n8315);
xnor_3 g07941(new_n8318, new_n8317, new_n8312);
not_3  g07942(new_n8319, new_n8318);
nand_4 g07943(new_n8320, n12145, n10928);
nand_4 g07944(new_n8321, n6986, n2522);
xor_3  g07945(new_n8322, new_n8321, new_n8320);
not_3  g07946(new_n8323, new_n8322);
xor_3  g07947(new_n8324, new_n8323, new_n8319);
not_3  g07948(new_n8325, new_n6034);
and_4  g07949(new_n8326, new_n6037, new_n8325);
nor_4  g07950(new_n8327, new_n6044, new_n6038_1);
nor_4  g07951(new_n8328, new_n8327, new_n8326);
xnor_3 g07952(new_n8329, new_n8328, new_n8324);
nand_4 g07953(new_n8330, new_n6046, new_n6033);
nand_4 g07954(new_n8331, new_n6053, new_n6047);
nand_4 g07955(new_n8332, new_n8331, new_n8330);
not_3  g07956(new_n8333, new_n8332);
nor_4  g07957(new_n8334, new_n8333, new_n8329);
not_3  g07958(new_n8335, new_n8329);
nor_4  g07959(new_n8336_1, new_n8332, new_n8335);
nor_4  g07960(new_n8337, new_n8336_1, new_n8334);
xnor_3 g07961(new_n8338, new_n8337, new_n8303_1);
xnor_3 g07962(new_n8339, new_n8338, new_n8301);
not_3  g07963(new_n8340, new_n6190);
nor_4  g07964(new_n8341, new_n8340, new_n6055);
not_3  g07965(new_n8342, new_n8341);
nand_4 g07966(new_n8343, new_n6253, new_n6191);
nand_4 g07967(new_n8344, new_n8343, new_n8342);
xnor_3 g07968(new_n8345, new_n8344, new_n8339);
not_3  g07969(new_n8346, new_n6091);
nor_4  g07970(new_n8347, new_n6212, new_n8346);
not_3  g07971(new_n8348, new_n8347);
nand_4 g07972(new_n8349, n12069, n5798);
nand_4 g07973(new_n8350, n7160, n5579);
not_3  g07974(new_n8351, new_n8350);
nor_4  g07975(new_n8352, new_n6205, new_n6200);
nor_4  g07976(new_n8353, new_n8352, new_n8351);
nor_4  g07977(new_n8354, new_n8352, new_n6081);
nor_4  g07978(new_n8355, new_n8354, new_n8350);
nor_4  g07979(new_n8356, new_n8355, new_n8353);
nand_4 g07980(new_n8357, n4828, n2498);
nand_4 g07981(new_n8358, n2558, n2515);
xor_3  g07982(new_n8359, new_n8358, new_n8357);
xnor_3 g07983(new_n8360, new_n8359, new_n8356);
nand_4 g07984(new_n8361, n12391, n6016);
nand_4 g07985(new_n8362, n7891, n521);
not_3  g07986(new_n8363, new_n8362);
xor_3  g07987(new_n8364, new_n8363, new_n8361);
xnor_3 g07988(new_n8365, new_n8364, new_n8360);
and_4  g07989(new_n8366, new_n6196, new_n6194);
nor_4  g07990(new_n8367, new_n6206, new_n6197);
nor_4  g07991(new_n8368, new_n8367, new_n8366);
xnor_3 g07992(new_n8369, new_n8368, new_n8365);
nor_4  g07993(new_n8370, new_n6207, new_n6192_1);
nor_4  g07994(new_n8371, new_n6211, new_n6208);
nor_4  g07995(new_n8372, new_n8371, new_n8370);
xnor_3 g07996(new_n8373, new_n8372, new_n8369);
xnor_3 g07997(new_n8374, new_n8373, new_n8349);
xnor_3 g07998(new_n8375, new_n8374, new_n8348);
not_3  g07999(new_n8376, new_n6248);
nand_4 g08000(new_n8377, n11222, n5153);
nand_4 g08001(new_n8378, n3342, n996);
nand_4 g08002(new_n8379, n9111, n5767);
nand_4 g08003(new_n8380, n9763, n5319);
xnor_3 g08004(new_n8381, new_n8380, new_n8379);
nor_4  g08005(new_n8382, new_n8381, new_n8378);
not_3  g08006(new_n8383, new_n8378);
not_3  g08007(new_n8384_1, new_n8381);
nor_4  g08008(new_n8385, new_n8384_1, new_n8383);
nor_4  g08009(new_n8386, new_n8385, new_n8382);
nor_4  g08010(new_n8387, new_n6233, new_n6227);
nor_4  g08011(new_n8388, new_n8387, new_n6232);
xnor_3 g08012(new_n8389, new_n8388, new_n8386);
not_3  g08013(new_n8390, new_n8389);
nand_4 g08014(new_n8391, n11153, n7270);
nand_4 g08015(new_n8392, n5314, n806);
xor_3  g08016(new_n8393, new_n8392, new_n8391);
xnor_3 g08017(new_n8394, new_n8393, new_n8390);
and_4  g08018(new_n8395, new_n6224, new_n6217);
nor_4  g08019(new_n8396, new_n6235, new_n6225);
nor_4  g08020(new_n8397, new_n8396, new_n8395);
xnor_3 g08021(new_n8398_1, new_n8397, new_n8394);
not_3  g08022(new_n8399, new_n6237);
nand_4 g08023(new_n8400, new_n6243, new_n6241);
nand_4 g08024(new_n8401, new_n8400, new_n8399);
not_3  g08025(new_n8402, new_n8401);
xnor_3 g08026(new_n8403, new_n8402, new_n8398_1);
xnor_3 g08027(new_n8404, new_n8403, new_n8377);
not_3  g08028(new_n8405, new_n8404);
nor_4  g08029(new_n8406, new_n8405, new_n8376);
nor_4  g08030(new_n8407, new_n8404, new_n6248);
nor_4  g08031(new_n8408, new_n8407, new_n8406);
nand_4 g08032(new_n8409, new_n8408, new_n8375);
not_3  g08033(new_n8410, new_n8375);
not_3  g08034(new_n8411, new_n8408);
nand_4 g08035(new_n8412, new_n8411, new_n8410);
nand_4 g08036(new_n8413, new_n8412, new_n8409);
nor_4  g08037(new_n8414, new_n6249, new_n6214);
nor_4  g08038(new_n8415, new_n6252, new_n6250);
nor_4  g08039(new_n8416, new_n8415, new_n8414);
xnor_3 g08040(new_n8417, new_n8416, new_n8413);
not_3  g08041(new_n8418, new_n8417);
xnor_3 g08042(new_n8419, new_n8418, new_n8345);
nor_4  g08043(new_n8420, new_n8419, new_n8300);
not_3  g08044(new_n8421, new_n8300);
not_3  g08045(new_n8422, new_n8419);
nor_4  g08046(new_n8423, new_n8422, new_n8421);
nor_4  g08047(n2708, new_n8423, new_n8420);
xor_3  g08048(n2818, new_n1050, new_n1049);
xnor_3 g08049(n2902, new_n2189, new_n2164);
nand_4 g08050(new_n8427, n11407, n5305);
not_3  g08051(new_n8428, new_n8427);
nand_4 g08052(new_n8429, n12709, n8759);
not_3  g08053(new_n8430, new_n8429);
nand_4 g08054(new_n8431, n12489, n5331);
nand_4 g08055(new_n8432, n10990, n7965);
not_3  g08056(new_n8433_1, new_n8432);
xor_3  g08057(new_n8434, new_n8433_1, new_n8431);
not_3  g08058(new_n8435, new_n8434);
xor_3  g08059(new_n8436, new_n8435, new_n8430);
xor_3  g08060(n3071, new_n8436, new_n8428);
not_3  g08061(new_n8438, new_n3084);
xor_3  g08062(n3124, new_n3087, new_n8438);
nand_4 g08063(new_n8440, new_n8436, new_n8428);
nand_4 g08064(new_n8441, n11407, n5964);
nand_4 g08065(new_n8442, n5305, n5212);
xor_3  g08066(new_n8443, new_n8442, new_n8441);
not_3  g08067(new_n8444, new_n8443);
nand_4 g08068(new_n8445, new_n8444, new_n8440);
nor_4  g08069(new_n8446, new_n8434, new_n8429);
nand_4 g08070(new_n8447, n11728, n8759);
nand_4 g08071(new_n8448, n12709, n6776);
not_3  g08072(new_n8449, new_n8448);
xor_3  g08073(new_n8450, new_n8449, new_n8447);
not_3  g08074(new_n8451, new_n8450);
nand_4 g08075(new_n8452, new_n8451, new_n8446);
not_3  g08076(new_n8453, new_n8452);
nor_4  g08077(new_n8454, new_n8451, new_n8446);
nor_4  g08078(new_n8455, new_n8454, new_n8453);
not_3  g08079(new_n8456, new_n8455);
nor_4  g08080(new_n8457, new_n8432, new_n8431);
nand_4 g08081(new_n8458, n7159, n5331);
nand_4 g08082(new_n8459, n12489, n8476);
not_3  g08083(new_n8460, new_n8459);
xor_3  g08084(new_n8461, new_n8460, new_n8458);
not_3  g08085(new_n8462, new_n8461);
xor_3  g08086(new_n8463, new_n8462, new_n8457);
nand_4 g08087(new_n8464, n7965, n5760);
nand_4 g08088(new_n8465, n10990, n7388);
xor_3  g08089(new_n8466, new_n8465, new_n8464);
not_3  g08090(new_n8467, new_n8466);
nor_4  g08091(new_n8468, new_n8467, new_n8463);
not_3  g08092(new_n8469, new_n8463);
nor_4  g08093(new_n8470, new_n8466, new_n8469);
nor_4  g08094(new_n8471, new_n8470, new_n8468);
xnor_3 g08095(new_n8472, new_n8471, new_n8456);
not_3  g08096(new_n8473, new_n8445);
nor_4  g08097(new_n8474, new_n8444, new_n8440);
nor_4  g08098(new_n8475, new_n8474, new_n8473);
nand_4 g08099(new_n8476_1, new_n8475, new_n8472);
nand_4 g08100(new_n8477, new_n8476_1, new_n8445);
nand_4 g08101(new_n8478, n5964, n5212);
nor_4  g08102(new_n8479, new_n8478, new_n8428);
nand_4 g08103(new_n8480, n11407, n1097);
nand_4 g08104(new_n8481, n11877, n5305);
nand_4 g08105(new_n8482, new_n8481, new_n8480);
nor_4  g08106(new_n8483, new_n8482, new_n8479);
nor_4  g08107(new_n8484, new_n8481, new_n8480);
nor_4  g08108(new_n8485, new_n8484, new_n8483);
not_3  g08109(new_n8486, new_n8485);
not_3  g08110(new_n8487, new_n8479);
not_3  g08111(new_n8488, new_n8482);
nor_4  g08112(new_n8489, new_n8488, new_n8487);
nor_4  g08113(new_n8490, new_n8489, new_n8486);
not_3  g08114(new_n8491, new_n8490);
nor_4  g08115(new_n8492, new_n8491, new_n8477);
not_3  g08116(new_n8493, new_n8477);
nor_4  g08117(new_n8494, new_n8490, new_n8493);
nor_4  g08118(new_n8495, new_n8494, new_n8492);
nor_4  g08119(new_n8496, new_n8471, new_n8456);
nor_4  g08120(new_n8497, new_n8496, new_n8453);
nand_4 g08121(new_n8498, n11728, n6776);
nor_4  g08122(new_n8499, new_n8498, new_n8430);
nand_4 g08123(new_n8500, n12709, n12299);
not_3  g08124(new_n8501, new_n8500);
nand_4 g08125(new_n8502, n8759, n6429);
not_3  g08126(new_n8503, new_n8502);
nand_4 g08127(new_n8504, new_n8503, new_n8501);
nand_4 g08128(new_n8505, new_n8502, new_n8500);
and_4  g08129(new_n8506, new_n8505, new_n8504);
nor_4  g08130(new_n8507, new_n8506, new_n8499);
not_3  g08131(new_n8508, new_n8498);
nand_4 g08132(new_n8509, new_n8505, new_n8508);
nor_4  g08133(new_n8510, new_n8509, new_n8430);
nor_4  g08134(new_n8511, new_n8510, new_n8507);
xnor_3 g08135(new_n8512, new_n8511, new_n8497);
not_3  g08136(new_n8513, new_n8431);
nand_4 g08137(new_n8514, n8476, n7159);
nor_4  g08138(new_n8515, new_n8514, new_n8513);
nand_4 g08139(new_n8516, n12489, n2530);
not_3  g08140(new_n8517, new_n8516);
nand_4 g08141(new_n8518, n12777, n5331);
not_3  g08142(new_n8519, new_n8518);
nor_4  g08143(new_n8520, new_n8519, new_n8517);
nor_4  g08144(new_n8521, new_n8518, new_n8516);
nor_4  g08145(new_n8522, new_n8521, new_n8520);
nor_4  g08146(new_n8523, new_n8522, new_n8515);
not_3  g08147(new_n8524, new_n8523);
not_3  g08148(new_n8525, new_n8520);
nand_4 g08149(new_n8526, new_n8525, new_n8515);
nand_4 g08150(new_n8527, new_n8526, new_n8524);
nand_4 g08151(new_n8528, n7388, n5760);
nor_4  g08152(new_n8529, new_n8528, new_n8433_1);
nand_4 g08153(new_n8530, n11892, n10990);
not_3  g08154(new_n8531, new_n8530);
nand_4 g08155(new_n8532, n7965, n1478);
not_3  g08156(new_n8533, new_n8532);
nor_4  g08157(new_n8534, new_n8533, new_n8531);
nor_4  g08158(new_n8535, new_n8532, new_n8530);
nor_4  g08159(new_n8536, new_n8535, new_n8534);
nor_4  g08160(new_n8537, new_n8536, new_n8529);
not_3  g08161(new_n8538, new_n8537);
not_3  g08162(new_n8539, new_n8534);
nand_4 g08163(new_n8540, new_n8539, new_n8529);
nand_4 g08164(new_n8541, new_n8540, new_n8538);
xor_3  g08165(new_n8542, new_n8541, new_n8527);
nor_4  g08166(new_n8543, new_n8462, new_n8457);
nor_4  g08167(new_n8544, new_n8470, new_n8543);
nand_4 g08168(new_n8545, new_n8544, new_n8542);
not_3  g08169(new_n8546, new_n8545);
nor_4  g08170(new_n8547, new_n8544, new_n8542);
nor_4  g08171(new_n8548, new_n8547, new_n8546);
nand_4 g08172(new_n8549, new_n8548, new_n8512);
not_3  g08173(new_n8550, new_n8549);
nor_4  g08174(new_n8551, new_n8548, new_n8512);
nor_4  g08175(new_n8552, new_n8551, new_n8550);
xor_3  g08176(n3214, new_n8552, new_n8495);
not_3  g08177(new_n8554, new_n5802);
nor_4  g08178(new_n8555, new_n5798_1, new_n5796);
xor_3  g08179(n3230, new_n8555, new_n8554);
not_3  g08180(new_n8557, new_n5279);
nand_4 g08181(new_n8558, new_n5225, new_n5223);
xnor_3 g08182(n3272, new_n8558, new_n8557);
nand_4 g08183(new_n8560, n5964, n4370);
not_3  g08184(new_n8561, new_n8560);
nand_4 g08185(new_n8562, n11407, n4312);
not_3  g08186(new_n8563, new_n8562);
nand_4 g08187(new_n8564, n11877, n5964);
not_3  g08188(new_n8565, new_n8564);
nor_4  g08189(new_n8566, new_n8565, new_n8563);
nor_4  g08190(new_n8567, new_n8564, new_n8562);
nand_4 g08191(new_n8568, n5212, n1097);
not_3  g08192(new_n8569, new_n8568);
nor_4  g08193(new_n8570, new_n8569, new_n8567);
nor_4  g08194(new_n8571, new_n8570, new_n8566);
nand_4 g08195(new_n8572, new_n8571, new_n8561);
xor_3  g08196(new_n8573, new_n8571, new_n8561);
nand_4 g08197(new_n8574, n5212, n4312);
not_3  g08198(new_n8575, new_n8574);
nand_4 g08199(new_n8576, n11877, n1097);
not_3  g08200(new_n8577, new_n8576);
nand_4 g08201(new_n8578, n12705, n11407);
not_3  g08202(new_n8579, new_n8578);
nor_4  g08203(new_n8580, new_n8579, new_n8577);
nor_4  g08204(new_n8581, new_n8578, new_n8576);
nor_4  g08205(new_n8582, new_n8581, new_n8580);
xor_3  g08206(new_n8583, new_n8582, new_n8575);
nand_4 g08207(new_n8584, new_n8583, new_n8573);
nand_4 g08208(new_n8585, new_n8584, new_n8572);
not_3  g08209(new_n8586, new_n8585);
nand_4 g08210(new_n8587, n5964, n5320);
nand_4 g08211(new_n8588, n4370, n1097);
xor_3  g08212(new_n8589, new_n8588, new_n8587);
not_3  g08213(new_n8590, new_n8589);
xor_3  g08214(new_n8591, new_n8590, new_n8586);
nand_4 g08215(new_n8592, n11877, n4312);
not_3  g08216(new_n8593, new_n8592);
nand_4 g08217(new_n8594, n12705, n5212);
nand_4 g08218(new_n8595_1, n12025, n11407);
xnor_3 g08219(new_n8596, new_n8595_1, new_n8594);
xnor_3 g08220(new_n8597, new_n8596, new_n8593);
nor_4  g08221(new_n8598, new_n8581, new_n8575);
nor_4  g08222(new_n8599, new_n8598, new_n8580);
xor_3  g08223(new_n8600, new_n8599, new_n8597);
xnor_3 g08224(new_n8601, new_n8600, new_n8591);
nand_4 g08225(new_n8602, n5320, n5305);
xnor_3 g08226(new_n8603, new_n8583, new_n8573);
nand_4 g08227(new_n8604, new_n8603, new_n8602);
not_3  g08228(new_n8605, new_n8602);
not_3  g08229(new_n8606, new_n8603);
xor_3  g08230(new_n8607, new_n8606, new_n8605);
nand_4 g08231(new_n8608, n5305, n4370);
not_3  g08232(new_n8609, new_n8608);
not_3  g08233(new_n8610, new_n8478);
nor_4  g08234(new_n8611, new_n8484, new_n8610);
nor_4  g08235(new_n8612, new_n8611, new_n8488);
and_4  g08236(new_n8613, new_n8612, new_n8609);
xor_3  g08237(new_n8614, new_n8612, new_n8608);
nor_4  g08238(new_n8615, new_n8567, new_n8566);
xor_3  g08239(new_n8616, new_n8615, new_n8568);
nor_4  g08240(new_n8617, new_n8616, new_n8614);
nor_4  g08241(new_n8618, new_n8617, new_n8613);
nand_4 g08242(new_n8619, new_n8618, new_n8607);
nand_4 g08243(new_n8620, new_n8619, new_n8604);
nor_4  g08244(new_n8621, new_n8620, new_n8601);
not_3  g08245(new_n8622, new_n8621);
nand_4 g08246(new_n8623, new_n8596, new_n8592);
not_3  g08247(new_n8624, new_n8599);
nand_4 g08248(new_n8625, new_n8624, new_n8597);
and_4  g08249(new_n8626, new_n8625, new_n8623);
nand_4 g08250(new_n8627, n12000, n5964);
nand_4 g08251(new_n8628, n5320, n1097);
nand_4 g08252(new_n8629, n9725, n5305);
not_3  g08253(new_n8630, new_n8629);
xor_3  g08254(new_n8631, new_n8630, new_n8628);
xnor_3 g08255(new_n8632, new_n8631, new_n8627);
xnor_3 g08256(new_n8633, new_n8632, new_n8626);
not_3  g08257(new_n8634, new_n8633);
nor_4  g08258(new_n8635, new_n8595_1, new_n8594);
nand_4 g08259(new_n8636, n4370, n4312);
xor_3  g08260(new_n8637, new_n8636, new_n8635);
nand_4 g08261(new_n8638, n12025, n5212);
nand_4 g08262(new_n8639, n12705, n11877);
nand_4 g08263(new_n8640, n11407, n11257);
not_3  g08264(new_n8641, new_n8640);
xor_3  g08265(new_n8642, new_n8641, new_n8639);
xnor_3 g08266(new_n8643, new_n8642, new_n8638);
xnor_3 g08267(new_n8644, new_n8643, new_n8637);
xnor_3 g08268(new_n8645, new_n8644, new_n8634);
nor_4  g08269(new_n8646, new_n8590, new_n8586);
nor_4  g08270(new_n8647, new_n8588, new_n8587);
nand_4 g08271(new_n8648, new_n8600, new_n8591);
xnor_3 g08272(new_n8649, new_n8648, new_n8647);
nor_4  g08273(new_n8650, new_n8649, new_n8646);
not_3  g08274(new_n8651, new_n8650);
xnor_3 g08275(new_n8652, new_n8651, new_n8645);
xnor_3 g08276(new_n8653, new_n8652, new_n8622);
nand_4 g08277(new_n8654, n12000, n5305);
xnor_3 g08278(new_n8655, new_n8620, new_n8601);
nor_4  g08279(new_n8656, new_n8655, new_n8654);
not_3  g08280(new_n8657, new_n8656);
xor_3  g08281(new_n8658, new_n8616, new_n8614);
nor_4  g08282(new_n8659, new_n8485, new_n8478);
nand_4 g08283(new_n8660, new_n8659, new_n8658);
not_3  g08284(new_n8661, new_n8619);
nor_4  g08285(new_n8662, new_n8618, new_n8607);
nor_4  g08286(new_n8663, new_n8662, new_n8661);
nor_4  g08287(new_n8664, new_n8663, new_n8660);
not_3  g08288(new_n8665_1, new_n8654);
not_3  g08289(new_n8666, new_n8655);
nor_4  g08290(new_n8667, new_n8666, new_n8665_1);
nor_4  g08291(new_n8668, new_n8667, new_n8656);
nand_4 g08292(new_n8669, new_n8668, new_n8664);
nand_4 g08293(new_n8670, new_n8669, new_n8657);
xnor_3 g08294(new_n8671, new_n8670, new_n8653);
not_3  g08295(new_n8672, new_n8671);
nand_4 g08296(new_n8673, n8759, n8717);
not_3  g08297(new_n8674, new_n8673);
nand_4 g08298(new_n8675, n7436, n6429);
not_3  g08299(new_n8676, new_n8675);
nand_4 g08300(new_n8677, n12709, n9241);
nand_4 g08301(new_n8678, n11728, n8276);
xnor_3 g08302(new_n8679, new_n8678, new_n8677);
xnor_3 g08303(new_n8680, new_n8679, new_n8676);
nand_4 g08304(new_n8681, n12299, n6429);
not_3  g08305(new_n8682, new_n8681);
nand_4 g08306(new_n8683, n12709, n8276);
not_3  g08307(new_n8684, new_n8683);
nor_4  g08308(new_n8685, new_n8684, new_n8682);
nor_4  g08309(new_n8686, new_n8683, new_n8681);
nand_4 g08310(new_n8687, n11728, n7436);
not_3  g08311(new_n8688, new_n8687);
nor_4  g08312(new_n8689, new_n8688, new_n8686);
nor_4  g08313(new_n8690, new_n8689, new_n8685);
xor_3  g08314(new_n8691, new_n8690, new_n8680);
nand_4 g08315(new_n8692, n6776, n2433);
nand_4 g08316(new_n8693, n12299, n8819);
xor_3  g08317(new_n8694, new_n8693, new_n8692);
xnor_3 g08318(new_n8695, new_n8694, new_n8691);
not_3  g08319(new_n8696, new_n8695);
nand_4 g08320(new_n8697, n8819, n6776);
not_3  g08321(new_n8698, new_n8697);
nand_4 g08322(new_n8699, n12709, n7436);
not_3  g08323(new_n8700, new_n8699);
nand_4 g08324(new_n8701, n6776, n6429);
not_3  g08325(new_n8702, new_n8701);
nor_4  g08326(new_n8703, new_n8702, new_n8700);
nor_4  g08327(new_n8704, new_n8701, new_n8699);
nand_4 g08328(new_n8705, n12299, n11728);
not_3  g08329(new_n8706, new_n8705);
nor_4  g08330(new_n8707, new_n8706, new_n8704);
nor_4  g08331(new_n8708, new_n8707, new_n8703);
and_4  g08332(new_n8709, new_n8708, new_n8698);
xor_3  g08333(new_n8710, new_n8708, new_n8697);
nor_4  g08334(new_n8711, new_n8686, new_n8685);
xor_3  g08335(new_n8712, new_n8711, new_n8687);
nor_4  g08336(new_n8713, new_n8712, new_n8710);
nor_4  g08337(new_n8714, new_n8713, new_n8709);
xnor_3 g08338(new_n8715, new_n8714, new_n8696);
nand_4 g08339(new_n8716, n8759, n2433);
xnor_3 g08340(new_n8717_1, new_n8712, new_n8710);
nand_4 g08341(new_n8718, new_n8717_1, new_n8716);
not_3  g08342(new_n8719, new_n8716);
not_3  g08343(new_n8720, new_n8717_1);
xor_3  g08344(new_n8721, new_n8720, new_n8719);
nand_4 g08345(new_n8722, n8819, n8759);
nand_4 g08346(new_n8723, new_n8509, new_n8504);
not_3  g08347(new_n8724, new_n8723);
nor_4  g08348(new_n8725, new_n8724, new_n8722);
xor_3  g08349(new_n8726, new_n8723, new_n8722);
nor_4  g08350(new_n8727, new_n8704, new_n8703);
xor_3  g08351(new_n8728, new_n8727, new_n8705);
nor_4  g08352(new_n8729, new_n8728, new_n8726);
nor_4  g08353(new_n8730, new_n8729, new_n8725);
nand_4 g08354(new_n8731, new_n8730, new_n8721);
nand_4 g08355(new_n8732, new_n8731, new_n8718);
xnor_3 g08356(new_n8733, new_n8732, new_n8715);
nand_4 g08357(new_n8734, new_n8733, new_n8674);
not_3  g08358(new_n8735, new_n8726);
not_3  g08359(new_n8736, new_n8728);
xor_3  g08360(new_n8737, new_n8736, new_n8735);
not_3  g08361(new_n8738, new_n8737);
not_3  g08362(new_n8739, new_n8507);
nor_4  g08363(new_n8740, new_n8739, new_n8498);
not_3  g08364(new_n8741, new_n8740);
nor_4  g08365(new_n8742, new_n8741, new_n8738);
xnor_3 g08366(new_n8743, new_n8730, new_n8721);
nand_4 g08367(new_n8744, new_n8743, new_n8742);
not_3  g08368(new_n8745, new_n8744);
xnor_3 g08369(new_n8746, new_n8733, new_n8673);
nand_4 g08370(new_n8747, new_n8746, new_n8745);
nand_4 g08371(new_n8748, new_n8747, new_n8734);
not_3  g08372(new_n8749, new_n8715);
nor_4  g08373(new_n8750, new_n8732, new_n8749);
nand_4 g08374(new_n8751, new_n8679, new_n8675);
not_3  g08375(new_n8752, new_n8690);
nand_4 g08376(new_n8753, new_n8752, new_n8680);
and_4  g08377(new_n8754, new_n8753, new_n8751);
nand_4 g08378(new_n8755, n8717, n6776);
not_3  g08379(new_n8756, new_n8755);
nand_4 g08380(new_n8757, n12299, n2433);
nand_4 g08381(new_n8758, n8759, n7730);
nor_4  g08382(new_n8759_1, new_n8758, new_n8757);
not_3  g08383(new_n8760, new_n8757);
not_3  g08384(new_n8761, new_n8758);
nor_4  g08385(new_n8762, new_n8761, new_n8760);
nor_4  g08386(new_n8763, new_n8762, new_n8759_1);
xnor_3 g08387(new_n8764, new_n8763, new_n8756);
xnor_3 g08388(new_n8765, new_n8764, new_n8754);
not_3  g08389(new_n8766, new_n8765);
nor_4  g08390(new_n8767, new_n8678, new_n8677);
nand_4 g08391(new_n8768, n8819, n7436);
xor_3  g08392(new_n8769, new_n8768, new_n8767);
nand_4 g08393(new_n8770, n11728, n9241);
nand_4 g08394(new_n8771, n8276, n6429);
nand_4 g08395(new_n8772, n12709, n10510);
not_3  g08396(new_n8773, new_n8772);
xor_3  g08397(new_n8774, new_n8773, new_n8771);
xnor_3 g08398(new_n8775, new_n8774, new_n8770);
xnor_3 g08399(new_n8776, new_n8775, new_n8769);
not_3  g08400(new_n8777, new_n8776);
xor_3  g08401(new_n8778, new_n8777, new_n8766);
nand_4 g08402(new_n8779, new_n8694, new_n8691);
nor_4  g08403(new_n8780, new_n8693, new_n8692);
nor_4  g08404(new_n8781, new_n8714, new_n8695);
xnor_3 g08405(new_n8782, new_n8781, new_n8780);
nand_4 g08406(new_n8783, new_n8782, new_n8779);
xnor_3 g08407(new_n8784, new_n8783, new_n8778);
xnor_3 g08408(new_n8785, new_n8784, new_n8750);
xnor_3 g08409(new_n8786, new_n8785, new_n8748);
nand_4 g08410(new_n8787, n2393, n1478);
nand_4 g08411(new_n8788, n5860, n5760);
nand_4 g08412(new_n8789, n10990, n3986);
xnor_3 g08413(new_n8790, new_n8789, new_n8788);
nor_4  g08414(new_n8791, new_n8790, new_n8787);
not_3  g08415(new_n8792, new_n8787);
not_3  g08416(new_n8793, new_n8790);
nor_4  g08417(new_n8794, new_n8793, new_n8792);
nor_4  g08418(new_n8795, new_n8794, new_n8791);
nand_4 g08419(new_n8796, n11892, n1478);
not_3  g08420(new_n8797, new_n8796);
nand_4 g08421(new_n8798, n10990, n5860);
not_3  g08422(new_n8799, new_n8798);
nor_4  g08423(new_n8800, new_n8799, new_n8797);
nor_4  g08424(new_n8801, new_n8798, new_n8796);
nand_4 g08425(new_n8802, n5760, n2393);
not_3  g08426(new_n8803, new_n8802);
nor_4  g08427(new_n8804, new_n8803, new_n8801);
nor_4  g08428(new_n8805, new_n8804, new_n8800);
xnor_3 g08429(new_n8806, new_n8805, new_n8795);
not_3  g08430(new_n8807, new_n8806);
nand_4 g08431(new_n8808, n12947, n7388);
nand_4 g08432(new_n8809, n11892, n11791);
xor_3  g08433(new_n8810, new_n8809, new_n8808);
xnor_3 g08434(new_n8811, new_n8810, new_n8807);
nand_4 g08435(new_n8812, n11791, n7388);
not_3  g08436(new_n8813, new_n8812);
nand_4 g08437(new_n8814, n10990, n2393);
not_3  g08438(new_n8815, new_n8814);
nand_4 g08439(new_n8816, n7388, n1478);
not_3  g08440(new_n8817, new_n8816);
nor_4  g08441(new_n8818, new_n8817, new_n8815);
nor_4  g08442(new_n8819_1, new_n8816, new_n8814);
nand_4 g08443(new_n8820, n11892, n5760);
not_3  g08444(new_n8821, new_n8820);
nor_4  g08445(new_n8822, new_n8821, new_n8819_1);
nor_4  g08446(new_n8823, new_n8822, new_n8818);
and_4  g08447(new_n8824, new_n8823, new_n8813);
xnor_3 g08448(new_n8825, new_n8823, new_n8813);
nor_4  g08449(new_n8826, new_n8801, new_n8800);
xnor_3 g08450(new_n8827, new_n8826, new_n8803);
nor_4  g08451(new_n8828, new_n8827, new_n8825);
nor_4  g08452(new_n8829, new_n8828, new_n8824);
xnor_3 g08453(new_n8830, new_n8829, new_n8811);
nand_4 g08454(new_n8831, n12947, n7965);
not_3  g08455(new_n8832, new_n8831);
nand_4 g08456(new_n8833, n11791, n7965);
not_3  g08457(new_n8834, new_n8833);
not_3  g08458(new_n8835, new_n8528);
nor_4  g08459(new_n8836, new_n8535, new_n8835);
nor_4  g08460(new_n8837, new_n8836, new_n8534);
nand_4 g08461(new_n8838, new_n8837, new_n8834);
xnor_3 g08462(new_n8839, new_n8837, new_n8833);
xnor_3 g08463(new_n8840, new_n8816, new_n8814);
xnor_3 g08464(new_n8841, new_n8840, new_n8820);
not_3  g08465(new_n8842, new_n8841);
nand_4 g08466(new_n8843, new_n8842, new_n8839);
nand_4 g08467(new_n8844, new_n8843, new_n8838);
nor_4  g08468(new_n8845, new_n8844, new_n8832);
not_3  g08469(new_n8846, new_n8845);
xnor_3 g08470(new_n8847, new_n8827, new_n8825);
not_3  g08471(new_n8848, new_n8844);
nor_4  g08472(new_n8849, new_n8848, new_n8831);
nor_4  g08473(new_n8850, new_n8849, new_n8845);
nand_4 g08474(new_n8851, new_n8850, new_n8847);
nand_4 g08475(new_n8852, new_n8851, new_n8846);
nor_4  g08476(new_n8853, new_n8852, new_n8830);
nor_4  g08477(new_n8854, new_n8789, new_n8788);
nand_4 g08478(new_n8855, n11791, n2393);
not_3  g08479(new_n8856, new_n8855);
xor_3  g08480(new_n8857, new_n8856, new_n8854);
not_3  g08481(new_n8858, new_n8857);
nand_4 g08482(new_n8859, n5760, n3986);
nand_4 g08483(new_n8860, n5860, n1478);
nand_4 g08484(new_n8861, n10990, n5857);
nand_4 g08485(new_n8862, new_n8861, new_n8860);
not_3  g08486(new_n8863, new_n8860);
not_3  g08487(new_n8864, new_n8861);
nand_4 g08488(new_n8865, new_n8864, new_n8863);
nand_4 g08489(new_n8866, new_n8865, new_n8862);
xor_3  g08490(new_n8867, new_n8866, new_n8859);
xnor_3 g08491(new_n8868, new_n8867, new_n8858);
nand_4 g08492(new_n8869, new_n8805, new_n8795);
not_3  g08493(new_n8870, new_n8869);
nor_4  g08494(new_n8871, new_n8870, new_n8791);
nand_4 g08495(new_n8872, n7388, n6441);
nand_4 g08496(new_n8873, n12947, n11892);
nand_4 g08497(new_n8874, n11999, n7965);
xor_3  g08498(new_n8875, new_n8874, new_n8873);
xnor_3 g08499(new_n8876, new_n8875, new_n8872);
xnor_3 g08500(new_n8877, new_n8876, new_n8871);
not_3  g08501(new_n8878, new_n8877);
nor_4  g08502(new_n8879, new_n8878, new_n8868);
xnor_3 g08503(new_n8880, new_n8867, new_n8857);
nor_4  g08504(new_n8881, new_n8877, new_n8880);
nor_4  g08505(new_n8882, new_n8881, new_n8879);
nand_4 g08506(new_n8883, new_n8810, new_n8807);
nor_4  g08507(new_n8884, new_n8809, new_n8808);
nor_4  g08508(new_n8885, new_n8829, new_n8811);
xnor_3 g08509(new_n8886, new_n8885, new_n8884);
nand_4 g08510(new_n8887, new_n8886, new_n8883);
xnor_3 g08511(new_n8888, new_n8887, new_n8882);
xnor_3 g08512(new_n8889, new_n8888, new_n8853);
nand_4 g08513(new_n8890, n7965, n6441);
not_3  g08514(new_n8891, new_n8890);
xnor_3 g08515(new_n8892, new_n8852, new_n8830);
not_3  g08516(new_n8893, new_n8892);
nand_4 g08517(new_n8894, new_n8893, new_n8891);
nand_4 g08518(new_n8895, new_n8892, new_n8890);
xor_3  g08519(new_n8896, new_n8841, new_n8839);
not_3  g08520(new_n8897, new_n8896);
nand_4 g08521(new_n8898, new_n8537, new_n8835);
not_3  g08522(new_n8899, new_n8898);
nand_4 g08523(new_n8900, new_n8899, new_n8897);
xnor_3 g08524(new_n8901, new_n8850, new_n8847);
not_3  g08525(new_n8902, new_n8901);
nor_4  g08526(new_n8903, new_n8902, new_n8900);
nand_4 g08527(new_n8904, new_n8903, new_n8895);
nand_4 g08528(new_n8905, new_n8904, new_n8894);
xnor_3 g08529(new_n8906, new_n8905, new_n8889);
nand_4 g08530(new_n8907, n12777, n12648);
nand_4 g08531(new_n8908, n10545, n7159);
nand_4 g08532(new_n8909, n12489, n7690);
xnor_3 g08533(new_n8910, new_n8909, new_n8908);
nor_4  g08534(new_n8911, new_n8910, new_n8907);
not_3  g08535(new_n8912, new_n8907);
not_3  g08536(new_n8913, new_n8910);
nor_4  g08537(new_n8914, new_n8913, new_n8912);
nor_4  g08538(new_n8915, new_n8914, new_n8911);
nand_4 g08539(new_n8916, n12777, n2530);
not_3  g08540(new_n8917, new_n8916);
nand_4 g08541(new_n8918, n12489, n10545);
not_3  g08542(new_n8919, new_n8918);
nor_4  g08543(new_n8920, new_n8919, new_n8917);
nor_4  g08544(new_n8921, new_n8918, new_n8916);
nand_4 g08545(new_n8922, n12648, n7159);
not_3  g08546(new_n8923, new_n8922);
nor_4  g08547(new_n8924, new_n8923, new_n8921);
nor_4  g08548(new_n8925, new_n8924, new_n8920);
xnor_3 g08549(new_n8926, new_n8925, new_n8915);
not_3  g08550(new_n8927, new_n8926);
nand_4 g08551(new_n8928, n11967, n8476);
nand_4 g08552(new_n8929, n6254, n2530);
xor_3  g08553(new_n8930, new_n8929, new_n8928);
xnor_3 g08554(new_n8931, new_n8930, new_n8927);
nand_4 g08555(new_n8932, n8476, n6254);
not_3  g08556(new_n8933, new_n8932);
nand_4 g08557(new_n8934, n12648, n12489);
not_3  g08558(new_n8935, new_n8934);
nand_4 g08559(new_n8936, n12777, n8476);
not_3  g08560(new_n8937, new_n8936);
nor_4  g08561(new_n8938, new_n8937, new_n8935);
nor_4  g08562(new_n8939, new_n8936, new_n8934);
nand_4 g08563(new_n8940, n7159, n2530);
not_3  g08564(new_n8941, new_n8940);
nor_4  g08565(new_n8942, new_n8941, new_n8939);
nor_4  g08566(new_n8943, new_n8942, new_n8938);
and_4  g08567(new_n8944, new_n8943, new_n8933);
xnor_3 g08568(new_n8945, new_n8943, new_n8933);
nor_4  g08569(new_n8946, new_n8921, new_n8920);
xnor_3 g08570(new_n8947, new_n8946, new_n8923);
nor_4  g08571(new_n8948, new_n8947, new_n8945);
nor_4  g08572(new_n8949, new_n8948, new_n8944);
xnor_3 g08573(new_n8950, new_n8949, new_n8931);
nand_4 g08574(new_n8951, n11967, n5331);
not_3  g08575(new_n8952, new_n8951);
xnor_3 g08576(new_n8953, new_n8947, new_n8945);
not_3  g08577(new_n8954, new_n8953);
nor_4  g08578(new_n8955, new_n8954, new_n8952);
not_3  g08579(new_n8956, new_n8955);
nor_4  g08580(new_n8957, new_n8953, new_n8951);
nor_4  g08581(new_n8958, new_n8957, new_n8955);
nand_4 g08582(new_n8959, n6254, n5331);
not_3  g08583(new_n8960, new_n8959);
not_3  g08584(new_n8961, new_n8514);
nor_4  g08585(new_n8962, new_n8521, new_n8961);
nor_4  g08586(new_n8963, new_n8962, new_n8520);
nand_4 g08587(new_n8964, new_n8963, new_n8960);
not_3  g08588(new_n8965, new_n8964);
xnor_3 g08589(new_n8966, new_n8963, new_n8960);
nor_4  g08590(new_n8967, new_n8939, new_n8938);
xnor_3 g08591(new_n8968, new_n8967, new_n8941);
nor_4  g08592(new_n8969, new_n8968, new_n8966);
nor_4  g08593(new_n8970, new_n8969, new_n8965);
nand_4 g08594(new_n8971, new_n8970, new_n8958);
nand_4 g08595(new_n8972, new_n8971, new_n8956);
nor_4  g08596(new_n8973, new_n8972, new_n8950);
not_3  g08597(new_n8974, new_n8973);
nand_4 g08598(new_n8975, n5331, n1353);
nand_4 g08599(new_n8976, n11967, n2530);
nand_4 g08600(new_n8977, n8476, n447);
not_3  g08601(new_n8978, new_n8977);
xor_3  g08602(new_n8979, new_n8978, new_n8976);
xnor_3 g08603(new_n8980, new_n8979, new_n8975);
nand_4 g08604(new_n8981, new_n8925, new_n8915);
not_3  g08605(new_n8982, new_n8981);
nor_4  g08606(new_n8983, new_n8982, new_n8911);
not_3  g08607(new_n8984, new_n8983);
xnor_3 g08608(new_n8985, new_n8984, new_n8980);
nor_4  g08609(new_n8986, new_n8909, new_n8908);
nand_4 g08610(new_n8987, n12648, n6254);
not_3  g08611(new_n8988, new_n8987);
xor_3  g08612(new_n8989, new_n8988, new_n8986);
not_3  g08613(new_n8990, new_n8989);
nand_4 g08614(new_n8991, n7690, n7159);
not_3  g08615(new_n8992, new_n8991);
nand_4 g08616(new_n8993, n12777, n10545);
nand_4 g08617(new_n8994, n12489, n3616);
not_3  g08618(new_n8995, new_n8994);
xor_3  g08619(new_n8996, new_n8995, new_n8993);
xnor_3 g08620(new_n8997, new_n8996, new_n8992);
xnor_3 g08621(new_n8998, new_n8997, new_n8990);
xnor_3 g08622(new_n8999, new_n8998, new_n8985);
nand_4 g08623(new_n9000, new_n8930, new_n8927);
nor_4  g08624(new_n9001, new_n8929, new_n8928);
nor_4  g08625(new_n9002, new_n8949, new_n8931);
xnor_3 g08626(new_n9003, new_n9002, new_n9001);
nand_4 g08627(new_n9004, new_n9003, new_n9000);
xnor_3 g08628(new_n9005, new_n9004, new_n8999);
xnor_3 g08629(new_n9006, new_n9005, new_n8974);
nand_4 g08630(new_n9007, n5331, n447);
not_3  g08631(new_n9008, new_n9007);
xnor_3 g08632(new_n9009, new_n8972, new_n8950);
not_3  g08633(new_n9010, new_n9009);
nand_4 g08634(new_n9011, new_n9010, new_n9008);
nand_4 g08635(new_n9012, new_n9009, new_n9007);
not_3  g08636(new_n9013, new_n8966);
xor_3  g08637(new_n9014, new_n8968, new_n9013);
nand_4 g08638(new_n9015, new_n8523, new_n8961);
nor_4  g08639(new_n9016, new_n9015, new_n9014);
xnor_3 g08640(new_n9017, new_n8970, new_n8958);
nand_4 g08641(new_n9018, new_n9017, new_n9016);
not_3  g08642(new_n9019, new_n9018);
nand_4 g08643(new_n9020, new_n9019, new_n9012);
nand_4 g08644(new_n9021, new_n9020, new_n9011);
xnor_3 g08645(new_n9022, new_n9021, new_n9006);
xnor_3 g08646(new_n9023, new_n9022, new_n8906);
nand_4 g08647(new_n9024, new_n8895, new_n8894);
xnor_3 g08648(new_n9025, new_n9024, new_n8903);
not_3  g08649(new_n9026, new_n9025);
nand_4 g08650(new_n9027, new_n9012, new_n9011);
xnor_3 g08651(new_n9028, new_n9027, new_n9019);
not_3  g08652(new_n9029, new_n9028);
nand_4 g08653(new_n9030, new_n9029, new_n9026);
nand_4 g08654(new_n9031, new_n9028, new_n9025);
xnor_3 g08655(new_n9032, new_n9017, new_n9016);
xnor_3 g08656(new_n9033, new_n8902, new_n8900);
nand_4 g08657(new_n9034, new_n9033, new_n9032);
xnor_3 g08658(new_n9035, new_n9033, new_n9032);
not_3  g08659(new_n9036, new_n9035);
xnor_3 g08660(new_n9037, new_n9015, new_n9014);
xor_3  g08661(new_n9038, new_n8898, new_n8897);
nor_4  g08662(new_n9039, new_n9038, new_n9037);
nor_4  g08663(new_n9040, new_n8541, new_n8527);
nor_4  g08664(new_n9041, new_n8546, new_n9040);
xnor_3 g08665(new_n9042, new_n9038, new_n9037);
nor_4  g08666(new_n9043, new_n9042, new_n9041);
nor_4  g08667(new_n9044, new_n9043, new_n9039);
nand_4 g08668(new_n9045, new_n9044, new_n9036);
nand_4 g08669(new_n9046, new_n9045, new_n9034);
nand_4 g08670(new_n9047, new_n9046, new_n9031);
nand_4 g08671(new_n9048, new_n9047, new_n9030);
xnor_3 g08672(new_n9049, new_n9048, new_n9023);
xnor_3 g08673(new_n9050, new_n9049, new_n8786);
not_3  g08674(new_n9051, new_n8747);
nor_4  g08675(new_n9052, new_n8746, new_n8745);
nor_4  g08676(new_n9053, new_n9052, new_n9051);
not_3  g08677(new_n9054, new_n9034);
not_3  g08678(new_n9055, new_n9014);
not_3  g08679(new_n9056, new_n9015);
nor_4  g08680(new_n9057, new_n9056, new_n9055);
nor_4  g08681(new_n9058, new_n9057, new_n9016);
xor_3  g08682(new_n9059, new_n8899, new_n8897);
nand_4 g08683(new_n9060, new_n9059, new_n9058);
not_3  g08684(new_n9061, new_n9041);
nor_4  g08685(new_n9062, new_n9059, new_n9058);
nor_4  g08686(new_n9063, new_n9062, new_n9039);
nand_4 g08687(new_n9064, new_n9063, new_n9061);
nand_4 g08688(new_n9065, new_n9064, new_n9060);
nor_4  g08689(new_n9066, new_n9065, new_n9035);
nor_4  g08690(new_n9067, new_n9066, new_n9054);
nand_4 g08691(new_n9068, new_n9031, new_n9030);
xnor_3 g08692(new_n9069, new_n9068, new_n9067);
nand_4 g08693(new_n9070, new_n9069, new_n9053);
not_3  g08694(new_n9071, new_n9053);
xnor_3 g08695(new_n9072, new_n9068, new_n9046);
nand_4 g08696(new_n9073, new_n9072, new_n9071);
xnor_3 g08697(new_n9074, new_n8743, new_n8742);
not_3  g08698(new_n9075, new_n9074);
xnor_3 g08699(new_n9076, new_n9065, new_n9035);
nand_4 g08700(new_n9077, new_n9076, new_n9075);
nor_4  g08701(new_n9078, new_n8740, new_n8737);
nor_4  g08702(new_n9079, new_n9078, new_n8742);
xnor_3 g08703(new_n9080_1, new_n9042, new_n9061);
nand_4 g08704(new_n9081, new_n9080_1, new_n9079);
not_3  g08705(new_n9082, new_n9079);
xnor_3 g08706(new_n9083, new_n9042, new_n9041);
nor_4  g08707(new_n9084, new_n9083, new_n9082);
nor_4  g08708(new_n9085, new_n9080_1, new_n9079);
nor_4  g08709(new_n9086, new_n9085, new_n9084);
not_3  g08710(new_n9087, new_n8511);
nor_4  g08711(new_n9088, new_n9087, new_n8497);
not_3  g08712(new_n9089, new_n9088);
nand_4 g08713(new_n9090, new_n8549, new_n9089);
nand_4 g08714(new_n9091, new_n9090, new_n9086);
nand_4 g08715(new_n9092, new_n9091, new_n9081);
xnor_3 g08716(new_n9093, new_n9076, new_n9074);
nand_4 g08717(new_n9094, new_n9093, new_n9092);
nand_4 g08718(new_n9095, new_n9094, new_n9077);
nand_4 g08719(new_n9096, new_n9095, new_n9073);
nand_4 g08720(new_n9097, new_n9096, new_n9070);
xnor_3 g08721(new_n9098, new_n9097, new_n9050);
nand_4 g08722(new_n9099, new_n9098, new_n8672);
xnor_3 g08723(new_n9100, new_n9098, new_n8671);
xnor_3 g08724(new_n9101, new_n8668, new_n8664);
not_3  g08725(new_n9102, new_n9077);
xnor_3 g08726(new_n9103, new_n9083, new_n9082);
not_3  g08727(new_n9104, new_n9090);
nor_4  g08728(new_n9105, new_n9104, new_n9103);
nor_4  g08729(new_n9106, new_n9105, new_n9084);
xnor_3 g08730(new_n9107, new_n9076, new_n9075);
nor_4  g08731(new_n9108, new_n9107, new_n9106);
nor_4  g08732(new_n9109, new_n9108, new_n9102);
nand_4 g08733(new_n9110, new_n9073, new_n9070);
xnor_3 g08734(new_n9111_1, new_n9110, new_n9109);
nand_4 g08735(new_n9112, new_n9111_1, new_n9101);
not_3  g08736(new_n9113, new_n9112);
not_3  g08737(new_n9114, new_n9101);
xnor_3 g08738(new_n9115, new_n9110, new_n9095);
nand_4 g08739(new_n9116, new_n9115, new_n9114);
nand_4 g08740(new_n9117, new_n9116, new_n9112);
not_3  g08741(new_n9118, new_n8660);
not_3  g08742(new_n9119, new_n8663);
nor_4  g08743(new_n9120, new_n9119, new_n9118);
nor_4  g08744(new_n9121, new_n9120, new_n8664);
not_3  g08745(new_n9122, new_n9121);
xnor_3 g08746(new_n9123, new_n9107, new_n9106);
nand_4 g08747(new_n9124, new_n9123, new_n9122);
not_3  g08748(new_n9125, new_n9124);
nor_4  g08749(new_n9126, new_n9093, new_n9092);
nor_4  g08750(new_n9127, new_n9126, new_n9108);
nand_4 g08751(new_n9128, new_n9127, new_n9121);
nand_4 g08752(new_n9129, new_n9128, new_n9124);
nor_4  g08753(new_n9130, new_n8659, new_n8658);
nor_4  g08754(new_n9131, new_n9130, new_n9118);
xnor_3 g08755(new_n9132, new_n9090, new_n9103);
nor_4  g08756(new_n9133, new_n9132, new_n9131);
not_3  g08757(new_n9134, new_n8492);
nand_4 g08758(new_n9135, new_n8552, new_n8495);
nand_4 g08759(new_n9136, new_n9135, new_n9134);
xnor_3 g08760(new_n9137_1, new_n9132, new_n9131);
nor_4  g08761(new_n9138, new_n9137_1, new_n9136);
nor_4  g08762(new_n9139, new_n9138, new_n9133);
nor_4  g08763(new_n9140, new_n9139, new_n9129);
nor_4  g08764(new_n9141, new_n9140, new_n9125);
nor_4  g08765(new_n9142, new_n9141, new_n9117);
nor_4  g08766(new_n9143, new_n9142, new_n9113);
nand_4 g08767(new_n9144, new_n9143, new_n9100);
nand_4 g08768(new_n9145, new_n9144, new_n9099);
nor_4  g08769(new_n9146, new_n9049, new_n8786);
nor_4  g08770(new_n9147, new_n9097, new_n9050);
nor_4  g08771(new_n9148, new_n9147, new_n9146);
not_3  g08772(new_n9149, new_n8906);
nand_4 g08773(new_n9150, new_n9022, new_n9149);
nand_4 g08774(new_n9151, new_n9048, new_n9023);
nand_4 g08775(new_n9152, new_n9151, new_n9150);
nand_4 g08776(new_n9153, new_n8888, new_n8853);
not_3  g08777(new_n9154, new_n8889);
nand_4 g08778(new_n9155, new_n8905, new_n9154);
nand_4 g08779(new_n9156, new_n9155, new_n9153);
nand_4 g08780(new_n9157, new_n8885, new_n8884);
not_3  g08781(new_n9158, new_n8882);
nand_4 g08782(new_n9159, new_n8887, new_n9158);
nand_4 g08783(new_n9160, new_n9159, new_n9157);
not_3  g08784(new_n9161, new_n8767);
nor_4  g08785(new_n9162, new_n8768, new_n9161);
nor_4  g08786(new_n9163, new_n8775, new_n8769);
nor_4  g08787(new_n9164, new_n9163, new_n9162);
nand_4 g08788(new_n9165, n9241, n6429);
nand_4 g08789(new_n9166, n12299, n8717);
xor_3  g08790(new_n9167, new_n9166, new_n9165);
nand_4 g08791(new_n9168, n7730, n6776);
nand_4 g08792(new_n9169, n8819, n8276);
xor_3  g08793(new_n9170, new_n9169, new_n9168);
xor_3  g08794(new_n9171, new_n9170, new_n9167);
not_3  g08795(new_n9172, new_n8771);
nor_4  g08796(new_n9173, new_n8773, new_n9172);
not_3  g08797(new_n9174, new_n8770);
nor_4  g08798(new_n9175, new_n8774, new_n9174);
nor_4  g08799(new_n9176, new_n9175, new_n9173);
nand_4 g08800(new_n9177, n7436, n2433);
xnor_3 g08801(new_n9178, new_n9177, new_n9176);
xnor_3 g08802(new_n9179, new_n9178, new_n9171);
xnor_3 g08803(new_n9180, new_n9179, new_n9164);
or_4   g08804(new_n9181, new_n8762, new_n8755);
not_3  g08805(new_n9182, new_n9181);
nor_4  g08806(new_n9183, new_n9182, new_n8759_1);
nand_4 g08807(new_n9184, n12777, n7690);
nand_4 g08808(new_n9185, n7159, n3616);
xor_3  g08809(new_n9186, new_n9185, new_n9184);
nand_4 g08810(new_n9187, n11999, n7388);
nand_4 g08811(new_n9188, n11892, n6441);
xor_3  g08812(new_n9189_1, new_n9188, new_n9187);
xnor_3 g08813(new_n9190, new_n9189_1, new_n9186);
nand_4 g08814(new_n9191, n10022, n7965);
nand_4 g08815(new_n9192, n10990, n45);
xor_3  g08816(new_n9193, new_n9192, new_n9191);
nand_4 g08817(new_n9194, n3986, n1478);
nand_4 g08818(new_n9195_1, n5857, n5760);
xor_3  g08819(new_n9196, new_n9195_1, new_n9194);
xnor_3 g08820(new_n9197, new_n9196, new_n9193);
xnor_3 g08821(new_n9198, new_n9197, new_n9190);
not_3  g08822(new_n9199, new_n8993);
nor_4  g08823(new_n9200, new_n8995, new_n9199);
nor_4  g08824(new_n9201, new_n8996, new_n8992);
nor_4  g08825(new_n9202, new_n9201, new_n9200);
nand_4 g08826(new_n9203, n8476, n1353);
not_3  g08827(new_n9204, new_n9203);
xnor_3 g08828(new_n9205, new_n9204, new_n9202);
xnor_3 g08829(new_n9206, new_n9205, new_n9198);
xnor_3 g08830(new_n9207, new_n9206, new_n9183);
xnor_3 g08831(new_n9208, new_n9207, new_n9180);
xnor_3 g08832(new_n9209, new_n9208, new_n9160);
xnor_3 g08833(new_n9210, new_n9209, new_n9156);
xnor_3 g08834(new_n9211, new_n9210, new_n9152);
xnor_3 g08835(new_n9212, new_n9211, new_n9148);
nand_4 g08836(new_n9213, new_n8784, new_n8750);
not_3  g08837(new_n9214, new_n8785);
nand_4 g08838(new_n9215, new_n9214, new_n8748);
nand_4 g08839(new_n9216, new_n9215, new_n9213);
nand_4 g08840(new_n9217, n2530, n447);
xnor_3 g08841(new_n9218, new_n9217, new_n9216);
nand_4 g08842(new_n9219, new_n8781, new_n8780);
not_3  g08843(new_n9220, new_n8778);
nand_4 g08844(new_n9221, new_n8783, new_n9220);
nand_4 g08845(new_n9222, new_n9221, new_n9219);
nand_4 g08846(new_n9223, n12648, n11967);
nand_4 g08847(new_n9224, n11791, n5860);
xor_3  g08848(new_n9225, new_n9224, new_n9223);
nand_4 g08849(new_n9226, n5331, n4436);
nand_4 g08850(new_n9227, n12489, n4499);
xor_3  g08851(new_n9228, new_n9227, new_n9226);
xor_3  g08852(new_n9229, new_n9228, new_n9225);
not_3  g08853(new_n9230, new_n8859);
nand_4 g08854(new_n9231, new_n8862, new_n9230);
nand_4 g08855(new_n9232, new_n9231, new_n8865);
nor_4  g08856(new_n9233, new_n8874, new_n8873);
not_3  g08857(new_n9234, new_n8872);
nand_4 g08858(new_n9235, new_n8874, new_n8873);
nand_4 g08859(new_n9236, new_n9235, new_n9234);
not_3  g08860(new_n9237, new_n9236);
nor_4  g08861(new_n9238, new_n9237, new_n9233);
xor_3  g08862(new_n9239, new_n9238, new_n9232);
xnor_3 g08863(new_n9240, new_n9239, new_n9229);
xnor_3 g08864(new_n9241_1, new_n9240, new_n9222);
not_3  g08865(new_n9242, new_n8647);
nor_4  g08866(new_n9243, new_n8648, new_n9242);
nor_4  g08867(new_n9244, new_n8650, new_n8645);
nor_4  g08868(new_n9245, new_n9244, new_n9243);
nand_4 g08869(new_n9246, n11257, n5212);
not_3  g08870(new_n9247, new_n8754);
nand_4 g08871(new_n9248, new_n8764, new_n9247);
nand_4 g08872(new_n9249, new_n8776, new_n8765);
nand_4 g08873(new_n9250, new_n9249, new_n9248);
nand_4 g08874(new_n9251, n12709, n10644);
not_3  g08875(new_n9252, new_n9251);
xnor_3 g08876(new_n9253, new_n9252, new_n9250);
nand_4 g08877(new_n9254, n11728, n10510);
not_3  g08878(new_n9255, new_n8626);
nand_4 g08879(new_n9256, new_n8632, new_n9255);
nand_4 g08880(new_n9257, new_n8644, new_n8633);
nand_4 g08881(new_n9258, new_n9257, new_n9256);
xnor_3 g08882(new_n9259, new_n9258, new_n9254);
xnor_3 g08883(new_n9260, new_n9259, new_n9253);
xnor_3 g08884(new_n9261, new_n9260, new_n9246);
xnor_3 g08885(new_n9262, new_n9261, new_n9245);
xnor_3 g08886(new_n9263, new_n9262, new_n9241_1);
nand_4 g08887(new_n9264, new_n9005, new_n8973);
nand_4 g08888(new_n9265, new_n9021, new_n9006);
nand_4 g08889(new_n9266, new_n9265, new_n9264);
nand_4 g08890(new_n9267, n12947, n2393);
not_3  g08891(new_n9268, new_n9267);
nand_4 g08892(new_n9269, new_n8856, new_n8854);
nand_4 g08893(new_n9270, new_n8867, new_n8857);
nand_4 g08894(new_n9271, new_n9270, new_n9269);
xor_3  g08895(new_n9272, new_n9271, new_n9268);
nand_4 g08896(new_n9273, new_n8983, new_n8980);
not_3  g08897(new_n9274, new_n8998);
nand_4 g08898(new_n9275, new_n9274, new_n8985);
nand_4 g08899(new_n9276, new_n9275, new_n9273);
nand_4 g08900(new_n9277, n10545, n6254);
nand_4 g08901(new_n9278, new_n8988, new_n8986);
nand_4 g08902(new_n9279, new_n8997, new_n8989);
nand_4 g08903(new_n9280, new_n9279, new_n9278);
nand_4 g08904(new_n9281, n8759, n1198);
not_3  g08905(new_n9282, new_n9281);
xnor_3 g08906(new_n9283, new_n9282, new_n9280);
xnor_3 g08907(new_n9284, new_n9283, new_n9277);
xnor_3 g08908(new_n9285, new_n9284, new_n9276);
nand_4 g08909(new_n9286, n12705, n4370);
not_3  g08910(new_n9287, new_n9286);
nand_4 g08911(new_n9288, n9725, n5964);
nand_4 g08912(new_n9289, n12000, n1097);
xor_3  g08913(new_n9290, new_n9289, new_n9288);
nand_4 g08914(new_n9291, n5320, n4312);
nand_4 g08915(new_n9292, n12025, n11877);
xor_3  g08916(new_n9293, new_n9292, new_n9291);
xnor_3 g08917(new_n9294, new_n9293, new_n9290);
xnor_3 g08918(new_n9295, new_n9294, new_n9287);
not_3  g08919(new_n9296, new_n8628);
nor_4  g08920(new_n9297, new_n8630, new_n9296);
not_3  g08921(new_n9298, new_n8627);
nor_4  g08922(new_n9299, new_n8631, new_n9298);
nor_4  g08923(new_n9300, new_n9299, new_n9297);
not_3  g08924(new_n9301, new_n8639);
nor_4  g08925(new_n9302, new_n8641, new_n9301);
not_3  g08926(new_n9303, new_n8638);
nor_4  g08927(new_n9304, new_n8642, new_n9303);
nor_4  g08928(new_n9305, new_n9304, new_n9302);
xnor_3 g08929(new_n9306, new_n9305, new_n9300);
xnor_3 g08930(new_n9307, new_n9306, new_n9295);
not_3  g08931(new_n9308, new_n8976);
nor_4  g08932(new_n9309, new_n8978, new_n9308);
not_3  g08933(new_n9310, new_n8975);
nor_4  g08934(new_n9311, new_n8979, new_n9310);
nor_4  g08935(new_n9312, new_n9311, new_n9309);
nand_4 g08936(new_n9313, n11407, n10547);
nand_4 g08937(new_n9314, n6604, n5305);
not_3  g08938(new_n9315, new_n9314);
xor_3  g08939(new_n9316, new_n9315, new_n9313);
xnor_3 g08940(new_n9317, new_n9316, new_n9312);
not_3  g08941(new_n9318, new_n8636);
or_4   g08942(new_n9319, new_n9318, new_n8635);
not_3  g08943(new_n9320, new_n8637);
nand_4 g08944(new_n9321, new_n8643, new_n9320);
nand_4 g08945(new_n9322, new_n9321, new_n9319);
xnor_3 g08946(new_n9323, new_n9322, new_n9317);
xnor_3 g08947(new_n9324, new_n9323, new_n9307);
xnor_3 g08948(new_n9325, new_n9324, new_n9285);
xnor_3 g08949(new_n9326, new_n9325, new_n9272);
xnor_3 g08950(new_n9327, new_n9326, new_n9266);
xnor_3 g08951(new_n9328, new_n9327, new_n9263);
nand_4 g08952(new_n9329, new_n8652, new_n8621);
nand_4 g08953(new_n9330, new_n8670, new_n8653);
nand_4 g08954(new_n9331, new_n9330, new_n9329);
nand_4 g08955(new_n9332, new_n9002, new_n9001);
not_3  g08956(new_n9333, new_n8999);
nand_4 g08957(new_n9334, new_n9004, new_n9333);
nand_4 g08958(new_n9335, new_n9334, new_n9332);
not_3  g08959(new_n9336, new_n8871);
nor_4  g08960(new_n9337, new_n8876, new_n9336);
nor_4  g08961(new_n9338, new_n8879, new_n9337);
xnor_3 g08962(new_n9339, new_n9338, new_n9335);
xnor_3 g08963(new_n9340, new_n9339, new_n9331);
xnor_3 g08964(new_n9341, new_n9340, new_n9328);
xnor_3 g08965(new_n9342, new_n9341, new_n9218);
xnor_3 g08966(new_n9343, new_n9342, new_n9212);
xnor_3 g08967(n3287, new_n9343, new_n9145);
xnor_3 g08968(n3339, new_n9141, new_n9117);
not_3  g08969(new_n9346, new_n4119);
xor_3  g08970(n3456, new_n9346, new_n4117);
nand_4 g08971(new_n9348, n6687, n4005);
not_3  g08972(new_n9349, new_n9348);
nand_4 g08973(new_n9350, n12720, n6770);
not_3  g08974(new_n9351, new_n9350);
nand_4 g08975(new_n9352, n9920, n2509);
nand_4 g08976(new_n9353, n6038, n3627);
xor_3  g08977(new_n9354, new_n9353, new_n9352);
xnor_3 g08978(new_n9355, new_n9354, new_n9351);
nand_4 g08979(new_n9356, n9920, n6038);
not_3  g08980(new_n9357, new_n9356);
nand_4 g08981(new_n9358, n12720, n4189);
not_3  g08982(new_n9359, new_n9358);
nor_4  g08983(new_n9360, new_n9359, new_n9357);
nand_4 g08984(new_n9361, n6770, n2509);
not_3  g08985(new_n9362, new_n9361);
xnor_3 g08986(new_n9363, new_n9358, new_n9356);
nor_4  g08987(new_n9364, new_n9363, new_n9362);
nor_4  g08988(new_n9365, new_n9364, new_n9360);
not_3  g08989(new_n9366, new_n9365);
xnor_3 g08990(new_n9367, new_n9366, new_n9355);
nand_4 g08991(new_n9368, n2564, n2508);
not_3  g08992(new_n9369, new_n9368);
nand_4 g08993(new_n9370, n6770, n6038);
not_3  g08994(new_n9371, new_n9370);
nand_4 g08995(new_n9372, n4189, n2509);
not_3  g08996(new_n9373, new_n9372);
nor_4  g08997(new_n9374, new_n9373, new_n9371);
nand_4 g08998(new_n9375, n12720, n2564);
not_3  g08999(new_n9376, new_n9375);
xnor_3 g09000(new_n9377, new_n9372, new_n9370);
nor_4  g09001(new_n9378, new_n9377, new_n9376);
nor_4  g09002(new_n9379, new_n9378, new_n9374);
nand_4 g09003(new_n9380, new_n9379, new_n9369);
xnor_3 g09004(new_n9381, new_n9363, new_n9362);
xnor_3 g09005(new_n9382, new_n9379, new_n9368);
nand_4 g09006(new_n9383, new_n9382, new_n9381);
nand_4 g09007(new_n9384, new_n9383, new_n9380);
nand_4 g09008(new_n9385, n2585, n2564);
nand_4 g09009(new_n9386, n4189, n2508);
xor_3  g09010(new_n9387_1, new_n9386, new_n9385);
xnor_3 g09011(new_n9388, new_n9387_1, new_n9384);
xnor_3 g09012(new_n9389, new_n9388, new_n9367);
nand_4 g09013(new_n9390, n6687, n2585);
not_3  g09014(new_n9391, new_n9390);
nand_4 g09015(new_n9392, n6687, n2508);
nand_4 g09016(new_n9393, new_n9359, new_n378);
nand_4 g09017(new_n9394, n6038, n4189);
nand_4 g09018(new_n9395, n12720, n6687);
nand_4 g09019(new_n9396, new_n9395, new_n9394);
nand_4 g09020(new_n9397, n2564, n2509);
not_3  g09021(new_n9398, new_n9397);
nand_4 g09022(new_n9399, new_n9398, new_n9396);
nand_4 g09023(new_n9400_1, new_n9399, new_n9393);
not_3  g09024(new_n9401, new_n9400_1);
nor_4  g09025(new_n9402, new_n9401, new_n9392);
not_3  g09026(new_n9403, new_n9402);
not_3  g09027(new_n9404, new_n9392);
xor_3  g09028(new_n9405, new_n9400_1, new_n9404);
xor_3  g09029(new_n9406, new_n9377, new_n9375);
nand_4 g09030(new_n9407, new_n9406, new_n9405);
nand_4 g09031(new_n9408, new_n9407, new_n9403);
nor_4  g09032(new_n9409, new_n9408, new_n9391);
not_3  g09033(new_n9410, new_n9409);
xor_3  g09034(new_n9411, new_n9382, new_n9381);
not_3  g09035(new_n9412, new_n9408);
xor_3  g09036(new_n9413, new_n9412, new_n9391);
nor_4  g09037(new_n9414, new_n9413, new_n9411);
not_3  g09038(new_n9415, new_n9414);
nand_4 g09039(new_n9416, new_n9415, new_n9410);
nor_4  g09040(new_n9417, new_n9416, new_n9389);
not_3  g09041(new_n9418, new_n9389);
nor_4  g09042(new_n9419, new_n9414, new_n9409);
nor_4  g09043(new_n9420, new_n9419, new_n9418);
nor_4  g09044(new_n9421, new_n9420, new_n9417);
nand_4 g09045(new_n9422, new_n9421, new_n9349);
not_3  g09046(new_n9423, new_n9393);
not_3  g09047(new_n9424, new_n9396);
nor_4  g09048(new_n9425, new_n9424, new_n9423);
nand_4 g09049(new_n9426, n6038, n2564);
nand_4 g09050(new_n9427, n6687, n2509);
nor_4  g09051(new_n9428, new_n9427, new_n9426);
not_3  g09052(new_n9429, new_n9428);
nor_4  g09053(new_n9430, new_n9429, new_n9425);
xor_3  g09054(new_n9431, new_n9406, new_n9405);
nand_4 g09055(new_n9432, new_n9431, new_n9430);
not_3  g09056(new_n9433, new_n9411);
not_3  g09057(new_n9434, new_n9413);
nor_4  g09058(new_n9435, new_n9434, new_n9433);
nor_4  g09059(new_n9436, new_n9435, new_n9414);
nor_4  g09060(new_n9437, new_n9436, new_n9432);
xnor_3 g09061(new_n9438, new_n9421, new_n9348);
nand_4 g09062(new_n9439, new_n9438, new_n9437);
nand_4 g09063(new_n9440, new_n9439, new_n9422);
nor_4  g09064(new_n9441, new_n9354, new_n9351);
not_3  g09065(new_n9442, new_n9441);
nor_4  g09066(new_n9443, new_n9365, new_n9355);
not_3  g09067(new_n9444, new_n9443);
nand_4 g09068(new_n9445, new_n9444, new_n9442);
nand_4 g09069(new_n9446, n4005, n2564);
nand_4 g09070(new_n9447, n4189, n2585);
nand_4 g09071(new_n9448, n12706, n6687);
not_3  g09072(new_n9449, new_n9448);
xor_3  g09073(new_n9450, new_n9449, new_n9447);
xnor_3 g09074(new_n9451, new_n9450, new_n9446);
not_3  g09075(new_n9452, new_n9451);
xnor_3 g09076(new_n9453, new_n9452, new_n9445);
nor_4  g09077(new_n9454, new_n9353, new_n9352);
nand_4 g09078(new_n9455, n6770, n2508);
not_3  g09079(new_n9456, new_n9455);
xor_3  g09080(new_n9457_1, new_n9456, new_n9454);
not_3  g09081(new_n9458, new_n9457_1);
nand_4 g09082(new_n9459, n3627, n2509);
not_3  g09083(new_n9460, new_n9459);
nand_4 g09084(new_n9461, n12720, n9920);
nand_4 g09085(new_n9462, n6038, n4516);
nand_4 g09086(new_n9463, new_n9462, new_n9461);
not_3  g09087(new_n9464, new_n9461);
not_3  g09088(new_n9465, new_n9462);
nand_4 g09089(new_n9466, new_n9465, new_n9464);
nand_4 g09090(new_n9467, new_n9466, new_n9463);
xor_3  g09091(new_n9468, new_n9467, new_n9460);
xnor_3 g09092(new_n9469, new_n9468, new_n9458);
xnor_3 g09093(new_n9470, new_n9469, new_n9453);
nand_4 g09094(new_n9471, new_n9387_1, new_n9384);
nor_4  g09095(new_n9472, new_n9386, new_n9385);
nor_4  g09096(new_n9473, new_n9388, new_n9367);
xnor_3 g09097(new_n9474, new_n9473, new_n9472);
nand_4 g09098(new_n9475, new_n9474, new_n9471);
xnor_3 g09099(new_n9476, new_n9475, new_n9470);
xnor_3 g09100(new_n9477, new_n9476, new_n9417);
xnor_3 g09101(new_n9478, new_n9477, new_n9440);
not_3  g09102(new_n9479, new_n9478);
nand_4 g09103(new_n9480, n8336, n1209);
nand_4 g09104(new_n9481, n7354, n6986);
nand_4 g09105(new_n9482, new_n9481, new_n9480);
not_3  g09106(new_n9483, new_n9482);
not_3  g09107(new_n9484, new_n9480);
not_3  g09108(new_n9485, new_n9481);
nand_4 g09109(new_n9486, new_n9485, new_n9484);
not_3  g09110(new_n9487, new_n9486);
nor_4  g09111(new_n9488, new_n9487, new_n9483);
nand_4 g09112(new_n9489, n10928, n7354);
nand_4 g09113(new_n9490, n8336, n7500);
nor_4  g09114(new_n9491, new_n9490, new_n9489);
not_3  g09115(new_n9492, new_n9491);
nor_4  g09116(new_n9493, new_n9492, new_n9488);
not_3  g09117(new_n9494, new_n9493);
nand_4 g09118(new_n9495, n8336, n5105);
not_3  g09119(new_n9496, new_n9495);
nand_4 g09120(new_n9497, n10928, n7500);
not_3  g09121(new_n9498, new_n9497);
nand_4 g09122(new_n9499, new_n9498, new_n9482);
nand_4 g09123(new_n9500, new_n9499, new_n9486);
xor_3  g09124(new_n9501, new_n9500, new_n9496);
nand_4 g09125(new_n9502, n7500, n6986);
not_3  g09126(new_n9503, new_n9502);
nand_4 g09127(new_n9504, n7354, n2226);
not_3  g09128(new_n9505, new_n9504);
nand_4 g09129(new_n9506, n10928, n1209);
not_3  g09130(new_n9507, new_n9506);
nor_4  g09131(new_n9508, new_n9507, new_n9505);
nor_4  g09132(new_n9509, new_n9506, new_n9504);
nor_4  g09133(new_n9510, new_n9509, new_n9508);
xor_3  g09134(new_n9511, new_n9510, new_n9503);
xnor_3 g09135(new_n9512, new_n9511, new_n9501);
nor_4  g09136(new_n9513, new_n9512, new_n9494);
nand_4 g09137(new_n9514, n8336, n4141);
not_3  g09138(new_n9515, new_n9514);
not_3  g09139(new_n9516, new_n9500);
nor_4  g09140(new_n9517, new_n9516, new_n9495);
not_3  g09141(new_n9518, new_n9517);
nand_4 g09142(new_n9519, new_n9511, new_n9501);
nand_4 g09143(new_n9520, new_n9519, new_n9518);
not_3  g09144(new_n9521, new_n9520);
xor_3  g09145(new_n9522, new_n9521, new_n9515);
nand_4 g09146(new_n9523, n10928, n5105);
not_3  g09147(new_n9524, new_n9523);
nor_4  g09148(new_n9525, new_n9509, new_n9503);
nor_4  g09149(new_n9526, new_n9525, new_n9508);
xor_3  g09150(new_n9527, new_n9526, new_n9524);
nand_4 g09151(new_n9528, n6986, n1209);
not_3  g09152(new_n9529, new_n9528);
nand_4 g09153(new_n9530, n7500, n2226);
nand_4 g09154(new_n9531, n7354, n1094);
xnor_3 g09155(new_n9532, new_n9531, new_n9530);
xor_3  g09156(new_n9533, new_n9532, new_n9529);
xnor_3 g09157(new_n9534, new_n9533, new_n9527);
xnor_3 g09158(new_n9535, new_n9534, new_n9522);
nand_4 g09159(new_n9536, new_n9535, new_n9513);
not_3  g09160(new_n9537, new_n9536);
nand_4 g09161(new_n9538, n8336, n4928);
not_3  g09162(new_n9539, new_n9538);
nand_4 g09163(new_n9540, n2226, n1209);
not_3  g09164(new_n9541, new_n9540);
not_3  g09165(new_n9542, new_n9530);
not_3  g09166(new_n9543, new_n9531);
nor_4  g09167(new_n9544, new_n9543, new_n9542);
nor_4  g09168(new_n9545, new_n9532, new_n9529);
nor_4  g09169(new_n9546, new_n9545, new_n9544);
xnor_3 g09170(new_n9547, new_n9546, new_n9541);
nand_4 g09171(new_n9548, n7500, n1094);
nand_4 g09172(new_n9549, n10678, n7354);
not_3  g09173(new_n9550, new_n9549);
xor_3  g09174(new_n9551, new_n9550, new_n9548);
xnor_3 g09175(new_n9552, new_n9551, new_n9547);
not_3  g09176(new_n9553, new_n9552);
nand_4 g09177(new_n9554, n10928, n4141);
nand_4 g09178(new_n9555, n6986, n5105);
xor_3  g09179(new_n9556, new_n9555, new_n9554);
not_3  g09180(new_n9557, new_n9556);
xor_3  g09181(new_n9558, new_n9557, new_n9553);
and_4  g09182(new_n9559, new_n9526, new_n9524);
not_3  g09183(new_n9560, new_n9527);
nor_4  g09184(new_n9561, new_n9533, new_n9560);
nor_4  g09185(new_n9562, new_n9561, new_n9559);
xnor_3 g09186(new_n9563, new_n9562, new_n9558);
not_3  g09187(new_n9564, new_n9563);
nor_4  g09188(new_n9565, new_n9520, new_n9515);
nor_4  g09189(new_n9566, new_n9534, new_n9522);
nor_4  g09190(new_n9567, new_n9566, new_n9565);
xnor_3 g09191(new_n9568, new_n9567, new_n9564);
xnor_3 g09192(new_n9569, new_n9568, new_n9539);
xnor_3 g09193(new_n9570, new_n9569, new_n9537);
nand_4 g09194(new_n9571_1, n8028, n5314);
not_3  g09195(new_n9572, new_n9571_1);
nand_4 g09196(new_n9573, n11222, n1980);
not_3  g09197(new_n9574, new_n9573);
nand_4 g09198(new_n9575, new_n9574, new_n9572);
nand_4 g09199(new_n9576, new_n9573, new_n9571_1);
nand_4 g09200(new_n9577, new_n9576, new_n9575);
nand_4 g09201(new_n9578_1, n11153, n8028);
nand_4 g09202(new_n9579, n11222, n10848);
nor_4  g09203(new_n9580, new_n9579, new_n9578_1);
and_4  g09204(new_n9581, new_n9580, new_n9577);
not_3  g09205(new_n9582, new_n9581);
nand_4 g09206(new_n9583_1, n11222, n7294);
nand_4 g09207(new_n9584, n11153, n10848);
not_3  g09208(new_n9585, new_n9584);
nand_4 g09209(new_n9586, new_n9585, new_n9576);
nand_4 g09210(new_n9587, new_n9586, new_n9575);
not_3  g09211(new_n9588, new_n9587);
xnor_3 g09212(new_n9589, new_n9588, new_n9583_1);
nand_4 g09213(new_n9590, n10848, n5314);
not_3  g09214(new_n9591, new_n9590);
nand_4 g09215(new_n9592, n8028, n996);
not_3  g09216(new_n9593, new_n9592);
nand_4 g09217(new_n9594, n11153, n1980);
not_3  g09218(new_n9595, new_n9594);
nor_4  g09219(new_n9596, new_n9595, new_n9593);
nor_4  g09220(new_n9597, new_n9594, new_n9592);
nor_4  g09221(new_n9598, new_n9597, new_n9596);
xnor_3 g09222(new_n9599, new_n9598, new_n9591);
xnor_3 g09223(new_n9600, new_n9599, new_n9589);
nor_4  g09224(new_n9601, new_n9600, new_n9582);
not_3  g09225(new_n9602, new_n9601);
nor_4  g09226(new_n9603, new_n9588, new_n9583_1);
nor_4  g09227(new_n9604, new_n9599, new_n9589);
nor_4  g09228(new_n9605, new_n9604, new_n9603);
nand_4 g09229(new_n9606, n12704, n11222);
not_3  g09230(new_n9607, new_n9606);
nand_4 g09231(new_n9608, n11153, n7294);
not_3  g09232(new_n9609, new_n9608);
nor_4  g09233(new_n9610, new_n9597, new_n9591);
nor_4  g09234(new_n9611, new_n9610, new_n9596);
xnor_3 g09235(new_n9612, new_n9611, new_n9609);
nand_4 g09236(new_n9613, n10848, n996);
not_3  g09237(new_n9614, new_n9613);
nand_4 g09238(new_n9615, n5314, n1980);
not_3  g09239(new_n9616, new_n9615);
nand_4 g09240(new_n9617, n8028, n5767);
not_3  g09241(new_n9618, new_n9617);
nor_4  g09242(new_n9619, new_n9618, new_n9616);
not_3  g09243(new_n9620, new_n9619);
nor_4  g09244(new_n9621, new_n9617, new_n9615);
not_3  g09245(new_n9622, new_n9621);
nand_4 g09246(new_n9623, new_n9622, new_n9620);
xnor_3 g09247(new_n9624, new_n9623, new_n9614);
xnor_3 g09248(new_n9625, new_n9624, new_n9612);
nor_4  g09249(new_n9626, new_n9625, new_n9607);
not_3  g09250(new_n9627, new_n9625);
nor_4  g09251(new_n9628, new_n9627, new_n9606);
nor_4  g09252(new_n9629, new_n9628, new_n9626);
xnor_3 g09253(new_n9630, new_n9629, new_n9605);
not_3  g09254(new_n9631, new_n9630);
nor_4  g09255(new_n9632, new_n9631, new_n9602);
nor_4  g09256(new_n9633, new_n9630, new_n9601);
nor_4  g09257(new_n9634, new_n9633, new_n9632);
nand_4 g09258(new_n9635, n7891, n1564);
nand_4 g09259(new_n9636, n12069, n533);
nand_4 g09260(new_n9637_1, new_n9636, new_n9635);
nor_4  g09261(new_n9638, new_n9636, new_n9635);
not_3  g09262(new_n9639, new_n9638);
nand_4 g09263(new_n9640_1, new_n9639, new_n9637_1);
not_3  g09264(new_n9641, new_n9640_1);
nand_4 g09265(new_n9642, n12391, n1564);
nand_4 g09266(new_n9643, n12069, n1512);
nor_4  g09267(new_n9644, new_n9643, new_n9642);
not_3  g09268(new_n9645, new_n9644);
nor_4  g09269(new_n9646, new_n9645, new_n9641);
not_3  g09270(new_n9647, new_n9646);
nand_4 g09271(new_n9648, n12069, n2802);
nand_4 g09272(new_n9649, n12391, n1512);
not_3  g09273(new_n9650, new_n9649);
nand_4 g09274(new_n9651, new_n9650, new_n9637_1);
nand_4 g09275(new_n9652, new_n9651, new_n9639);
not_3  g09276(new_n9653, new_n9652);
nor_4  g09277(new_n9654, new_n9653, new_n9648);
not_3  g09278(new_n9655, new_n9648);
nor_4  g09279(new_n9656, new_n9652, new_n9655);
nor_4  g09280(new_n9657, new_n9656, new_n9654);
nand_4 g09281(new_n9658, n7891, n1512);
nand_4 g09282(new_n9659, n7160, n1564);
nand_4 g09283(new_n9660, n12391, n533);
xnor_3 g09284(new_n9661, new_n9660, new_n9659);
xnor_3 g09285(new_n9662, new_n9661, new_n9658);
not_3  g09286(new_n9663, new_n9662);
xnor_3 g09287(new_n9664, new_n9663, new_n9657);
nor_4  g09288(new_n9665, new_n9664, new_n9647);
not_3  g09289(new_n9666, new_n9664);
nor_4  g09290(new_n9667, new_n9666, new_n9646);
nor_4  g09291(new_n9668, new_n9667, new_n9665);
not_3  g09292(new_n9669, new_n9600);
nor_4  g09293(new_n9670, new_n9669, new_n9581);
nor_4  g09294(new_n9671, new_n9670, new_n9601);
nor_4  g09295(new_n9672, new_n9671, new_n9668);
nand_4 g09296(new_n9673, new_n9650, new_n382);
nand_4 g09297(new_n9674, new_n9673, new_n9640_1);
not_3  g09298(new_n9675, new_n9651);
nand_4 g09299(new_n9676, new_n9675, new_n382);
nand_4 g09300(new_n9677, new_n9676, new_n9674);
not_3  g09301(new_n9678, new_n381_1);
nor_4  g09302(new_n9679, new_n9584, new_n9678);
not_3  g09303(new_n9680, new_n9679);
nand_4 g09304(new_n9681, new_n9680, new_n9577);
nand_4 g09305(new_n9682, new_n9679, new_n9576);
nand_4 g09306(new_n9683, new_n9682, new_n9681);
and_4  g09307(new_n9684, new_n9683, new_n9677);
nor_4  g09308(new_n9685, new_n382, new_n381_1);
xnor_3 g09309(new_n9686, new_n9579, new_n9578_1);
not_3  g09310(new_n9687, new_n9686);
nor_4  g09311(new_n9688, new_n9687, new_n9685);
xor_3  g09312(new_n9689, new_n9686, new_n9685);
xor_3  g09313(new_n9690, new_n9643, new_n9642);
nor_4  g09314(new_n9691, new_n9690, new_n9689);
nor_4  g09315(new_n9692, new_n9691, new_n9688);
xnor_3 g09316(new_n9693, new_n9683, new_n9677);
nor_4  g09317(new_n9694, new_n9693, new_n9692);
nor_4  g09318(new_n9695, new_n9694, new_n9684);
xnor_3 g09319(new_n9696, new_n9671, new_n9668);
nor_4  g09320(new_n9697, new_n9696, new_n9695);
nor_4  g09321(new_n9698, new_n9697, new_n9672);
nor_4  g09322(new_n9699, new_n9698, new_n9634);
nand_4 g09323(new_n9700, n12069, n6806);
nand_4 g09324(new_n9701, n12391, n2802);
not_3  g09325(new_n9702, new_n9701);
not_3  g09326(new_n9703, new_n9659);
not_3  g09327(new_n9704, new_n9660);
nor_4  g09328(new_n9705, new_n9704, new_n9703);
not_3  g09329(new_n9706_1, new_n9658);
nor_4  g09330(new_n9707, new_n9661, new_n9706_1);
nor_4  g09331(new_n9708, new_n9707, new_n9705);
xnor_3 g09332(new_n9709, new_n9708, new_n9702);
nand_4 g09333(new_n9710, n7891, n533);
nand_4 g09334(new_n9711, n4828, n1564);
nand_4 g09335(new_n9712, n7160, n1512);
xnor_3 g09336(new_n9713, new_n9712, new_n9711);
xnor_3 g09337(new_n9714, new_n9713, new_n9710);
xnor_3 g09338(new_n9715, new_n9714, new_n9709);
nand_4 g09339(new_n9716, new_n9715, new_n9700);
not_3  g09340(new_n9717, new_n9716);
nor_4  g09341(new_n9718, new_n9715, new_n9700);
nor_4  g09342(new_n9719, new_n9718, new_n9717);
not_3  g09343(new_n9720, new_n9654);
nand_4 g09344(new_n9721, new_n9663, new_n9657);
nand_4 g09345(new_n9722, new_n9721, new_n9720);
not_3  g09346(new_n9723, new_n9722);
xnor_3 g09347(new_n9724, new_n9723, new_n9719);
nand_4 g09348(new_n9725_1, new_n9724, new_n9665);
not_3  g09349(new_n9726, new_n9725_1);
nor_4  g09350(new_n9727, new_n9724, new_n9665);
nor_4  g09351(new_n9728, new_n9727, new_n9726);
xnor_3 g09352(new_n9729, new_n9698, new_n9634);
nor_4  g09353(new_n9730, new_n9729, new_n9728);
nor_4  g09354(new_n9731, new_n9730, new_n9699);
not_3  g09355(new_n9732, new_n9731);
nand_4 g09356(new_n9733, n11222, n5814);
nand_4 g09357(new_n9734, n1980, n996);
nand_4 g09358(new_n9735, n8028, n5319);
nand_4 g09359(new_n9736, n10848, n5767);
xnor_3 g09360(new_n9737, new_n9736, new_n9735);
nor_4  g09361(new_n9738, new_n9737, new_n9734);
not_3  g09362(new_n9739, new_n9734);
not_3  g09363(new_n9740, new_n9737);
nor_4  g09364(new_n9741, new_n9740, new_n9739);
nor_4  g09365(new_n9742, new_n9741, new_n9738);
nor_4  g09366(new_n9743, new_n9621, new_n9614);
nor_4  g09367(new_n9744, new_n9743, new_n9619);
xnor_3 g09368(new_n9745, new_n9744, new_n9742);
nand_4 g09369(new_n9746, n12704, n11153);
nand_4 g09370(new_n9747, n7294, n5314);
xor_3  g09371(new_n9748, new_n9747, new_n9746);
xnor_3 g09372(new_n9749, new_n9748, new_n9745);
and_4  g09373(new_n9750, new_n9611, new_n9609);
not_3  g09374(new_n9751, new_n9624);
nor_4  g09375(new_n9752, new_n9751, new_n9612);
nor_4  g09376(new_n9753, new_n9752, new_n9750);
xnor_3 g09377(new_n9754, new_n9753, new_n9749);
not_3  g09378(new_n9755, new_n9628);
nor_4  g09379(new_n9756_1, new_n9626, new_n9605);
not_3  g09380(new_n9757, new_n9756_1);
nand_4 g09381(new_n9758, new_n9757, new_n9755);
xnor_3 g09382(new_n9759, new_n9758, new_n9754);
xnor_3 g09383(new_n9760, new_n9759, new_n9733);
xnor_3 g09384(new_n9761, new_n9760, new_n9632);
nand_4 g09385(new_n9762, n12069, n5069);
nand_4 g09386(new_n9763_1, n7160, n533);
nand_4 g09387(new_n9764, n2515, n1564);
nand_4 g09388(new_n9765, n4828, n1512);
xnor_3 g09389(new_n9766, new_n9765, new_n9764);
nor_4  g09390(new_n9767_1, new_n9766, new_n9763_1);
not_3  g09391(new_n9768, new_n9763_1);
not_3  g09392(new_n9769, new_n9766);
nor_4  g09393(new_n9770, new_n9769, new_n9768);
nor_4  g09394(new_n9771, new_n9770, new_n9767_1);
and_4  g09395(new_n9772, new_n9712, new_n9711);
not_3  g09396(new_n9773, new_n9710);
nor_4  g09397(new_n9774, new_n9713, new_n9773);
nor_4  g09398(new_n9775, new_n9774, new_n9772);
xnor_3 g09399(new_n9776, new_n9775, new_n9771);
nand_4 g09400(new_n9777, n7891, n2802);
nand_4 g09401(new_n9778, n12391, n6806);
xor_3  g09402(new_n9779, new_n9778, new_n9777);
not_3  g09403(new_n9780, new_n9779);
nor_4  g09404(new_n9781, new_n9780, new_n9776);
not_3  g09405(new_n9782, new_n9776);
nor_4  g09406(new_n9783, new_n9779, new_n9782);
nor_4  g09407(new_n9784, new_n9783, new_n9781);
nand_4 g09408(new_n9785, new_n9708, new_n9702);
not_3  g09409(new_n9786, new_n9785);
nor_4  g09410(new_n9787, new_n9714, new_n9709);
nor_4  g09411(new_n9788, new_n9787, new_n9786);
not_3  g09412(new_n9789, new_n9788);
xnor_3 g09413(new_n9790, new_n9789, new_n9784);
nand_4 g09414(new_n9791, new_n9723, new_n9719);
nand_4 g09415(new_n9792, new_n9791, new_n9716);
xnor_3 g09416(new_n9793, new_n9792, new_n9790);
nand_4 g09417(new_n9794, new_n9793, new_n9762);
not_3  g09418(new_n9795, new_n9762);
not_3  g09419(new_n9796, new_n9792);
xnor_3 g09420(new_n9797, new_n9796, new_n9790);
nand_4 g09421(new_n9798, new_n9797, new_n9795);
nand_4 g09422(new_n9799, new_n9798, new_n9794);
xnor_3 g09423(new_n9800, new_n9799, new_n9725_1);
not_3  g09424(new_n9801, new_n9800);
nand_4 g09425(new_n9802, new_n9801, new_n9761);
not_3  g09426(new_n9803, new_n9761);
nand_4 g09427(new_n9804, new_n9800, new_n9803);
nand_4 g09428(new_n9805, new_n9804, new_n9802);
xnor_3 g09429(new_n9806, new_n9805, new_n9732);
nor_4  g09430(new_n9807, new_n9806, new_n9570);
xnor_3 g09431(new_n9808, new_n9806, new_n9570);
nor_4  g09432(new_n9809, new_n9535, new_n9513);
nor_4  g09433(new_n9810, new_n9809, new_n9537);
xnor_3 g09434(new_n9811, new_n9729, new_n9728);
nand_4 g09435(new_n9812, new_n9811, new_n9810);
not_3  g09436(new_n9813, new_n9812);
not_3  g09437(new_n9814, new_n9810);
not_3  g09438(new_n9815, new_n9728);
xnor_3 g09439(new_n9816, new_n9729, new_n9815);
nand_4 g09440(new_n9817, new_n9816, new_n9814);
nand_4 g09441(new_n9818, new_n9817, new_n9812);
not_3  g09442(new_n9819, new_n9512);
xor_3  g09443(new_n9820_1, new_n9819, new_n9494);
not_3  g09444(new_n9821, new_n9696);
xnor_3 g09445(new_n9822, new_n9821, new_n9695);
nor_4  g09446(new_n9823, new_n9822, new_n9820_1);
xnor_3 g09447(new_n9824, new_n9822, new_n9820_1);
xnor_3 g09448(new_n9825, new_n9693, new_n9692);
nor_4  g09449(new_n9826, new_n9497, new_n380);
not_3  g09450(new_n9827, new_n9826);
nor_4  g09451(new_n9828, new_n9827, new_n9482);
not_3  g09452(new_n9829, new_n9488);
nor_4  g09453(new_n9830, new_n9826, new_n9829);
nor_4  g09454(new_n9831, new_n9830, new_n9828);
not_3  g09455(new_n9832, new_n9831);
nor_4  g09456(new_n9833, new_n9832, new_n9825);
not_3  g09457(new_n9834, new_n9833);
not_3  g09458(new_n9835, new_n9825);
xor_3  g09459(new_n9836, new_n9831, new_n9835);
xnor_3 g09460(new_n9837, new_n9690, new_n9689);
xor_3  g09461(new_n9838, new_n9490, new_n9489);
nand_4 g09462(new_n9839, new_n9838, new_n9837);
not_3  g09463(new_n9840, new_n9839);
nor_4  g09464(new_n9841, new_n384, new_n379);
not_3  g09465(new_n9842, new_n9841);
xnor_3 g09466(new_n9843, new_n9838, new_n9837);
nor_4  g09467(new_n9844, new_n9843, new_n9842);
nor_4  g09468(new_n9845, new_n9844, new_n9840);
nand_4 g09469(new_n9846, new_n9845, new_n9836);
nand_4 g09470(new_n9847, new_n9846, new_n9834);
nor_4  g09471(new_n9848, new_n9847, new_n9824);
nor_4  g09472(new_n9849, new_n9848, new_n9823);
nor_4  g09473(new_n9850, new_n9849, new_n9818);
nor_4  g09474(new_n9851, new_n9850, new_n9813);
nor_4  g09475(new_n9852, new_n9851, new_n9808);
nor_4  g09476(new_n9853, new_n9852, new_n9807);
nand_4 g09477(new_n9854, new_n9567, new_n9564);
and_4  g09478(new_n9855, new_n9546, new_n9541);
nor_4  g09479(new_n9856, new_n9551, new_n9547);
nor_4  g09480(new_n9857, new_n9856, new_n9855);
nand_4 g09481(new_n9858, n10928, n4928);
nand_4 g09482(new_n9859, n6986, n4141);
nand_4 g09483(new_n9860, n8336, n8236);
xor_3  g09484(new_n9861, new_n9860, new_n9859);
not_3  g09485(new_n9862, new_n9861);
xor_3  g09486(new_n9863, new_n9862, new_n9858);
not_3  g09487(new_n9864, new_n9863);
xnor_3 g09488(new_n9865, new_n9864, new_n9857);
nor_4  g09489(new_n9866, new_n9549, new_n9548);
not_3  g09490(new_n9867, new_n9866);
nand_4 g09491(new_n9868, n5105, n2226);
xor_3  g09492(new_n9869, new_n9868, new_n9867);
nand_4 g09493(new_n9870, n10678, n7500);
nand_4 g09494(new_n9871, n7354, n7320);
nand_4 g09495(new_n9872, n1209, n1094);
not_3  g09496(new_n9873, new_n9872);
xor_3  g09497(new_n9874, new_n9873, new_n9871);
xnor_3 g09498(new_n9875, new_n9874, new_n9870);
xnor_3 g09499(new_n9876, new_n9875, new_n9869);
xnor_3 g09500(new_n9877, new_n9876, new_n9865);
nand_4 g09501(new_n9878, new_n9556, new_n9553);
nor_4  g09502(new_n9879, new_n9555, new_n9554);
nor_4  g09503(new_n9880, new_n9562, new_n9558);
xnor_3 g09504(new_n9881, new_n9880, new_n9879);
nand_4 g09505(new_n9882, new_n9881, new_n9878);
xnor_3 g09506(new_n9883, new_n9882, new_n9877);
xnor_3 g09507(new_n9884, new_n9883, new_n9854);
nand_4 g09508(new_n9885, new_n9568, new_n9538);
nand_4 g09509(new_n9886, new_n9569, new_n9536);
nand_4 g09510(new_n9887, new_n9886, new_n9885);
xnor_3 g09511(new_n9888, new_n9887, new_n9884);
not_3  g09512(new_n9889, new_n9888);
not_3  g09513(new_n9890, new_n9754);
not_3  g09514(new_n9891, new_n9758);
nor_4  g09515(new_n9892, new_n9891, new_n9890);
not_3  g09516(new_n9893, new_n9892);
nand_4 g09517(new_n9894, new_n9744, new_n9742);
not_3  g09518(new_n9895, new_n9894);
nor_4  g09519(new_n9896, new_n9895, new_n9738);
not_3  g09520(new_n9897, new_n9896);
nand_4 g09521(new_n9898, n11153, n5814);
nand_4 g09522(new_n9899, n12704, n5314);
nand_4 g09523(new_n9900, n11222, n4903);
not_3  g09524(new_n9901, new_n9900);
xor_3  g09525(new_n9902, new_n9901, new_n9899);
xnor_3 g09526(new_n9903, new_n9902, new_n9898);
xnor_3 g09527(new_n9904, new_n9903, new_n9897);
nor_4  g09528(new_n9905, new_n9736, new_n9735);
nand_4 g09529(new_n9906, n7294, n996);
not_3  g09530(new_n9907, new_n9906);
xor_3  g09531(new_n9908, new_n9907, new_n9905);
nand_4 g09532(new_n9909, n10848, n5319);
not_3  g09533(new_n9910, new_n9909);
nand_4 g09534(new_n9911, n5767, n1980);
nand_4 g09535(new_n9912, n9457, n8028);
not_3  g09536(new_n9913, new_n9912);
xor_3  g09537(new_n9914, new_n9913, new_n9911);
xnor_3 g09538(new_n9915, new_n9914, new_n9910);
xnor_3 g09539(new_n9916, new_n9915, new_n9908);
xnor_3 g09540(new_n9917, new_n9916, new_n9904);
not_3  g09541(new_n9918, new_n9917);
not_3  g09542(new_n9919, new_n9745);
nand_4 g09543(new_n9920_1, new_n9748, new_n9919);
nor_4  g09544(new_n9921, new_n9747, new_n9746);
not_3  g09545(new_n9922, new_n9749);
nor_4  g09546(new_n9923, new_n9753, new_n9922);
xnor_3 g09547(new_n9924, new_n9923, new_n9921);
nand_4 g09548(new_n9925, new_n9924, new_n9920_1);
xnor_3 g09549(new_n9926, new_n9925, new_n9918);
xnor_3 g09550(new_n9927, new_n9926, new_n9893);
not_3  g09551(new_n9928, new_n9733);
not_3  g09552(new_n9929, new_n9759);
nor_4  g09553(new_n9930, new_n9929, new_n9928);
nor_4  g09554(new_n9931, new_n9759, new_n9733);
nor_4  g09555(new_n9932, new_n9931, new_n9632);
nor_4  g09556(new_n9933, new_n9932, new_n9930);
xnor_3 g09557(new_n9934, new_n9933, new_n9927);
nor_4  g09558(new_n9935, new_n9792, new_n9790);
not_3  g09559(new_n9936, new_n9935);
not_3  g09560(new_n9937, new_n9781);
nor_4  g09561(new_n9938_1, new_n9778, new_n9777);
nand_4 g09562(new_n9939, new_n9789, new_n9784);
not_3  g09563(new_n9940, new_n9939);
xnor_3 g09564(new_n9941, new_n9940, new_n9938_1);
nand_4 g09565(new_n9942, new_n9941, new_n9937);
nor_4  g09566(new_n9943, new_n9765, new_n9764);
nand_4 g09567(new_n9944, n7160, n2802);
not_3  g09568(new_n9945, new_n9944);
xor_3  g09569(new_n9946, new_n9945, new_n9943);
nand_4 g09570(new_n9947, n2515, n1512);
not_3  g09571(new_n9948, new_n9947);
nand_4 g09572(new_n9949, n1564, n1199);
nand_4 g09573(new_n9950, n4828, n533);
nand_4 g09574(new_n9951, new_n9950, new_n9949);
not_3  g09575(new_n9952, new_n9949);
not_3  g09576(new_n9953, new_n9950);
nand_4 g09577(new_n9954, new_n9953, new_n9952);
nand_4 g09578(new_n9955, new_n9954, new_n9951);
xor_3  g09579(new_n9956_1, new_n9955, new_n9948);
not_3  g09580(new_n9957, new_n9956_1);
nor_4  g09581(new_n9958, new_n9957, new_n9946);
not_3  g09582(new_n9959, new_n9946);
nor_4  g09583(new_n9960, new_n9956_1, new_n9959);
nor_4  g09584(new_n9961, new_n9960, new_n9958);
not_3  g09585(new_n9962, new_n9767_1);
nand_4 g09586(new_n9963, new_n9775, new_n9771);
nand_4 g09587(new_n9964, new_n9963, new_n9962);
nand_4 g09588(new_n9965, n12391, n5069);
nand_4 g09589(new_n9966, n7891, n6806);
nand_4 g09590(new_n9967, n12069, n12044);
not_3  g09591(new_n9968, new_n9967);
xor_3  g09592(new_n9969, new_n9968, new_n9966);
xnor_3 g09593(new_n9970, new_n9969, new_n9965);
xnor_3 g09594(new_n9971, new_n9970, new_n9964);
xnor_3 g09595(new_n9972, new_n9971, new_n9961);
xnor_3 g09596(new_n9973, new_n9972, new_n9942);
xnor_3 g09597(new_n9974, new_n9973, new_n9936);
nand_4 g09598(new_n9975, new_n9794, new_n9726);
nand_4 g09599(new_n9976, new_n9975, new_n9798);
xnor_3 g09600(new_n9977, new_n9976, new_n9974);
nand_4 g09601(new_n9978, new_n9804, new_n9731);
nand_4 g09602(new_n9979, new_n9978, new_n9802);
xnor_3 g09603(new_n9980, new_n9979, new_n9977);
xnor_3 g09604(new_n9981, new_n9980, new_n9934);
nand_4 g09605(new_n9982, new_n9981, new_n9889);
not_3  g09606(new_n9983, new_n9934);
xnor_3 g09607(new_n9984, new_n9980, new_n9983);
nand_4 g09608(new_n9985, new_n9984, new_n9888);
nand_4 g09609(new_n9986, new_n9985, new_n9982);
xnor_3 g09610(new_n9987, new_n9986, new_n9853);
not_3  g09611(new_n9988, new_n9987);
nand_4 g09612(new_n9989, new_n9988, new_n9479);
nand_4 g09613(new_n9990, new_n9987, new_n9478);
not_3  g09614(new_n9991, new_n9439);
nor_4  g09615(new_n9992, new_n9438, new_n9437);
nor_4  g09616(new_n9993, new_n9992, new_n9991);
xnor_3 g09617(new_n9994, new_n9436, new_n9432);
not_3  g09618(new_n9995, new_n9994);
xnor_3 g09619(new_n9996, new_n9849, new_n9818);
not_3  g09620(new_n9997, new_n9996);
nand_4 g09621(new_n9998, new_n9997, new_n9995);
nand_4 g09622(new_n9999, new_n9996, new_n9994);
not_3  g09623(new_n10000, new_n9430);
xnor_3 g09624(new_n10001, new_n9431, new_n10000);
not_3  g09625(new_n10002, new_n9824);
xnor_3 g09626(new_n10003, new_n9847, new_n10002);
nor_4  g09627(new_n10004, new_n10003, new_n10001);
xnor_3 g09628(new_n10005, new_n10003, new_n10001);
xnor_3 g09629(new_n10006, new_n9845, new_n9836);
nor_4  g09630(new_n10007, new_n9397, new_n378);
nor_4  g09631(new_n10008, new_n10007, new_n9425);
not_3  g09632(new_n10009, new_n10007);
nor_4  g09633(new_n10010, new_n10009, new_n9424);
nor_4  g09634(new_n10011, new_n10010, new_n10008);
nor_4  g09635(new_n10012, new_n10011, new_n10006);
xnor_3 g09636(new_n10013, new_n10011, new_n10006);
not_3  g09637(new_n10014, new_n386);
nor_4  g09638(new_n10015, new_n10014, new_n377);
xor_3  g09639(new_n10016, new_n9427, new_n9426);
nor_4  g09640(new_n10017, new_n10016, new_n10015);
xnor_3 g09641(new_n10018, new_n9843, new_n9841);
xnor_3 g09642(new_n10019, new_n10016, new_n10015);
nor_4  g09643(new_n10020, new_n10019, new_n10018);
nor_4  g09644(new_n10021, new_n10020, new_n10017);
nor_4  g09645(new_n10022_1, new_n10021, new_n10013);
nor_4  g09646(new_n10023, new_n10022_1, new_n10012);
nor_4  g09647(new_n10024, new_n10023, new_n10005);
nor_4  g09648(new_n10025, new_n10024, new_n10004);
nand_4 g09649(new_n10026, new_n10025, new_n9999);
nand_4 g09650(new_n10027, new_n10026, new_n9998);
nor_4  g09651(new_n10028, new_n10027, new_n9993);
not_3  g09652(new_n10029, new_n9851);
xnor_3 g09653(new_n10030, new_n10029, new_n9808);
xnor_3 g09654(new_n10031, new_n10027, new_n9993);
nor_4  g09655(new_n10032, new_n10031, new_n10030);
nor_4  g09656(new_n10033, new_n10032, new_n10028);
nand_4 g09657(new_n10034, new_n10033, new_n9990);
nand_4 g09658(new_n10035, new_n10034, new_n9989);
nor_4  g09659(new_n10036, new_n9883, new_n9854);
nor_4  g09660(new_n10037, new_n9887, new_n9884);
nor_4  g09661(new_n10038, new_n10037, new_n10036);
nand_4 g09662(new_n10039, new_n9973, new_n9935);
nand_4 g09663(new_n10040, new_n9976, new_n9974);
nand_4 g09664(new_n10041, new_n10040, new_n10039);
nand_4 g09665(new_n10042, new_n9907, new_n9905);
nand_4 g09666(new_n10043, new_n9915, new_n9908);
nand_4 g09667(new_n10044, new_n10043, new_n10042);
nand_4 g09668(new_n10045, n10848, n9457);
nand_4 g09669(new_n10046, n11222, n1906);
not_3  g09670(new_n10047, new_n10046);
xor_3  g09671(new_n10048, new_n10047, new_n10045);
xor_3  g09672(new_n10049, new_n10048, new_n10044);
not_3  g09673(new_n10050, new_n9911);
nor_4  g09674(new_n10051, new_n9913, new_n10050);
nor_4  g09675(new_n10052, new_n9914, new_n9910);
nor_4  g09676(new_n10053, new_n10052, new_n10051);
nand_4 g09677(new_n10054, n8028, n4817);
not_3  g09678(new_n10055, new_n10054);
nand_4 g09679(new_n10056, n6578, n1564);
nand_4 g09680(new_n10057, n5814, n5314);
xor_3  g09681(new_n10058, new_n10057, new_n10056);
xor_3  g09682(new_n10059, new_n10058, new_n10055);
xnor_3 g09683(new_n10060, new_n10059, new_n10053);
not_3  g09684(new_n10061, new_n9899);
nor_4  g09685(new_n10062, new_n9901, new_n10061);
not_3  g09686(new_n10063, new_n9898);
nor_4  g09687(new_n10064, new_n9902, new_n10063);
nor_4  g09688(new_n10065, new_n10064, new_n10062);
nand_4 g09689(new_n10066, n7294, n5767);
nand_4 g09690(new_n10067, n12069, n5694);
nand_4 g09691(new_n10068, n11153, n4903);
xor_3  g09692(new_n10069, new_n10068, new_n10067);
xor_3  g09693(new_n10070, new_n10069, new_n10066);
xnor_3 g09694(new_n10071, new_n10070, new_n10065);
xnor_3 g09695(new_n10072, new_n10071, new_n10060);
xnor_3 g09696(new_n10073, new_n10072, new_n10049);
xnor_3 g09697(new_n10074, new_n10073, new_n10041);
xnor_3 g09698(new_n10075, new_n10074, new_n10038);
not_3  g09699(new_n10076, new_n9476);
nand_4 g09700(new_n10077, new_n10076, new_n9417);
nand_4 g09701(new_n10078, new_n9477, new_n9440);
nand_4 g09702(new_n10079, new_n10078, new_n10077);
nand_4 g09703(new_n10080, new_n9923, new_n9921);
nand_4 g09704(new_n10081, new_n9925, new_n9917);
nand_4 g09705(new_n10082, new_n10081, new_n10080);
nand_4 g09706(new_n10083, n5319, n1980);
xnor_3 g09707(new_n10084, new_n10083, new_n10082);
nand_4 g09708(new_n10085, n12720, n3627);
nand_4 g09709(new_n10086, n4516, n2509);
xor_3  g09710(new_n10087, new_n10086, new_n10085);
nand_4 g09711(new_n10088, new_n9463, new_n9460);
and_4  g09712(new_n10089, new_n10088, new_n9466);
xnor_3 g09713(new_n10090, new_n10089, new_n10087);
nand_4 g09714(new_n10091, n12706, n2564);
not_3  g09715(new_n10092, new_n10091);
nand_4 g09716(new_n10093, n9920, n2508);
nand_4 g09717(new_n10094, n4189, n4005);
xor_3  g09718(new_n10095, new_n10094, new_n10093);
xnor_3 g09719(new_n10096, new_n10095, new_n10092);
xnor_3 g09720(new_n10097, new_n10096, new_n10090);
not_3  g09721(new_n10098, new_n9447);
nor_4  g09722(new_n10099, new_n9449, new_n10098);
not_3  g09723(new_n10100, new_n9446);
nor_4  g09724(new_n10101, new_n9450, new_n10100);
nor_4  g09725(new_n10102, new_n10101, new_n10099);
or_4   g09726(new_n10103, new_n9456, new_n9454);
nand_4 g09727(new_n10104, new_n9468, new_n9457_1);
nand_4 g09728(new_n10105, new_n10104, new_n10103);
xnor_3 g09729(new_n10106, new_n10105, new_n10102);
xnor_3 g09730(new_n10107, new_n10106, new_n10097);
xnor_3 g09731(new_n10108, new_n10107, new_n10084);
nand_4 g09732(new_n10109, new_n9473, new_n9472);
nand_4 g09733(new_n10110, new_n9475, new_n9470);
nand_4 g09734(new_n10111, new_n10110, new_n10109);
nand_4 g09735(new_n10112, new_n9451, new_n9445);
nand_4 g09736(new_n10113, new_n9469, new_n9453);
nand_4 g09737(new_n10114, new_n10113, new_n10112);
nand_4 g09738(new_n10115, n6770, n2585);
nand_4 g09739(new_n10116, new_n9951, new_n9948);
and_4  g09740(new_n10117, new_n10116, new_n9954);
nand_4 g09741(new_n10118, n6687, n615);
nand_4 g09742(new_n10119, n6038, n2087);
xor_3  g09743(new_n10120, new_n10119, new_n10118);
xnor_3 g09744(new_n10121, new_n10120, new_n10117);
xnor_3 g09745(new_n10122, new_n10121, new_n10115);
xnor_3 g09746(new_n10123, new_n10122, new_n10114);
xnor_3 g09747(new_n10124, new_n10123, new_n10111);
xnor_3 g09748(new_n10125, new_n10124, new_n10108);
nand_4 g09749(new_n10126, new_n9940, new_n9938_1);
not_3  g09750(new_n10127, new_n9972);
nand_4 g09751(new_n10128, new_n10127, new_n9942);
nand_4 g09752(new_n10129, new_n10128, new_n10126);
not_3  g09753(new_n10130, new_n9964);
nand_4 g09754(new_n10131, new_n9970, new_n10130);
not_3  g09755(new_n10132, new_n9961);
nand_4 g09756(new_n10133, new_n9971, new_n10132);
nand_4 g09757(new_n10134, new_n10133, new_n10131);
nand_4 g09758(new_n10135, new_n9945, new_n9943);
not_3  g09759(new_n10136, new_n9960);
nand_4 g09760(new_n10137, new_n10136, new_n10135);
nand_4 g09761(new_n10138, n12391, n12044);
nand_4 g09762(new_n10139, n1512, n1199);
nand_4 g09763(new_n10140, n7160, n6806);
xor_3  g09764(new_n10141, new_n10140, new_n10139);
nand_4 g09765(new_n10142, n2515, n533);
nand_4 g09766(new_n10143, n4828, n2802);
xor_3  g09767(new_n10144, new_n10143, new_n10142);
xnor_3 g09768(new_n10145, new_n10144, new_n10141);
xnor_3 g09769(new_n10146, new_n10145, new_n10138);
nand_4 g09770(new_n10147, n7891, n5069);
not_3  g09771(new_n10148, new_n10147);
not_3  g09772(new_n10149, new_n9966);
nor_4  g09773(new_n10150, new_n9968, new_n10149);
not_3  g09774(new_n10151, new_n9965);
nor_4  g09775(new_n10152, new_n9969, new_n10151);
nor_4  g09776(new_n10153, new_n10152, new_n10150);
xnor_3 g09777(new_n10154, new_n10153, new_n10148);
xnor_3 g09778(new_n10155, new_n10154, new_n10146);
xnor_3 g09779(new_n10156, new_n10155, new_n10137);
xnor_3 g09780(new_n10157, new_n10156, new_n10134);
xnor_3 g09781(new_n10158, new_n10157, new_n10129);
xnor_3 g09782(new_n10159, new_n10158, new_n10125);
xnor_3 g09783(new_n10160, new_n10159, new_n10079);
xnor_3 g09784(new_n10161, new_n10160, new_n10075);
not_3  g09785(new_n10162, new_n9979);
nand_4 g09786(new_n10163, new_n10162, new_n9977);
nand_4 g09787(new_n10164, new_n9980, new_n9934);
nand_4 g09788(new_n10165, new_n10164, new_n10163);
nand_4 g09789(new_n10166, new_n9926, new_n9892);
nand_4 g09790(new_n10167, new_n9933, new_n9927);
nand_4 g09791(new_n10168, new_n10167, new_n10166);
nand_4 g09792(new_n10169, new_n9864, new_n9857);
not_3  g09793(new_n10170, new_n9865);
not_3  g09794(new_n10171, new_n9876);
nand_4 g09795(new_n10172, new_n10171, new_n10170);
nand_4 g09796(new_n10173, new_n10172, new_n10169);
xnor_3 g09797(new_n10174_1, new_n10173, new_n10168);
nand_4 g09798(new_n10175, new_n9880, new_n9879);
nand_4 g09799(new_n10176, new_n9882, new_n9877);
nand_4 g09800(new_n10177, new_n10176, new_n10175);
nand_4 g09801(new_n10178, n7500, n7320);
nand_4 g09802(new_n10179, n7523, n7354);
xor_3  g09803(new_n10180, new_n10179, new_n10178);
nand_4 g09804(new_n10181, n4141, n2226);
nand_4 g09805(new_n10182, n8336, n783);
not_3  g09806(new_n10183, new_n10182);
xor_3  g09807(new_n10184, new_n10183, new_n10181);
xor_3  g09808(new_n10185, new_n10184, new_n10180);
nor_4  g09809(new_n10186, new_n9868, new_n9867);
not_3  g09810(new_n10187, new_n9869);
nor_4  g09811(new_n10188, new_n9875, new_n10187);
nor_4  g09812(new_n10189, new_n10188, new_n10186);
nand_4 g09813(new_n10190, n12704, n996);
not_3  g09814(new_n10191, new_n10190);
not_3  g09815(new_n10192, new_n9871);
nor_4  g09816(new_n10193, new_n9873, new_n10192);
not_3  g09817(new_n10194, new_n9870);
nor_4  g09818(new_n10195, new_n9874, new_n10194);
nor_4  g09819(new_n10196, new_n10195, new_n10193);
nand_4 g09820(new_n10197, n6986, n4928);
nand_4 g09821(new_n10198, n10678, n1209);
xor_3  g09822(new_n10199, new_n10198, new_n10197);
nand_4 g09823(new_n10200, n10928, n8236);
nand_4 g09824(new_n10201, n5105, n1094);
xor_3  g09825(new_n10202, new_n10201, new_n10200);
xnor_3 g09826(new_n10203, new_n10202, new_n10199);
xnor_3 g09827(new_n10204, new_n10203, new_n10196);
xnor_3 g09828(new_n10205, new_n10204, new_n10191);
xnor_3 g09829(new_n10206, new_n10205, new_n10189);
xnor_3 g09830(new_n10207, new_n10206, new_n10185);
nand_4 g09831(new_n10208, new_n9903, new_n9896);
nand_4 g09832(new_n10209, new_n9916, new_n9904);
nand_4 g09833(new_n10210, new_n10209, new_n10208);
and_4  g09834(new_n10211, new_n9860, new_n9859);
not_3  g09835(new_n10212, new_n9858);
nor_4  g09836(new_n10213, new_n9862, new_n10212);
or_4   g09837(new_n10214, new_n10213, new_n10211);
xnor_3 g09838(new_n10215, new_n10214, new_n10210);
xnor_3 g09839(new_n10216, new_n10215, new_n10207);
xnor_3 g09840(new_n10217_1, new_n10216, new_n10177);
xnor_3 g09841(new_n10218, new_n10217_1, new_n10174_1);
xnor_3 g09842(new_n10219, new_n10218, new_n10165);
xnor_3 g09843(new_n10220, new_n10219, new_n10161);
nand_4 g09844(new_n10221, new_n9982, new_n9853);
nand_4 g09845(new_n10222, new_n10221, new_n9985);
xnor_3 g09846(new_n10223_1, new_n10222, new_n10220);
xnor_3 g09847(n3654, new_n10223_1, new_n10035);
xnor_3 g09848(n3661, new_n10031, new_n10030);
nor_4  g09849(new_n10226, new_n6538, new_n6537);
not_3  g09850(new_n10227, new_n10226);
nand_4 g09851(new_n10228, n1798, n1097);
nand_4 g09852(new_n10229, n12591, n5305);
nand_4 g09853(new_n10230, new_n10229, new_n10228);
not_3  g09854(new_n10231, new_n10230);
not_3  g09855(new_n10232, new_n10228);
not_3  g09856(new_n10233, new_n10229);
nand_4 g09857(new_n10234, new_n10233, new_n10232);
not_3  g09858(new_n10235, new_n10234);
nor_4  g09859(new_n10236, new_n10235, new_n10231);
nor_4  g09860(new_n10237, new_n10236, new_n10227);
nand_4 g09861(new_n10238, n7456, n5305);
nand_4 g09862(new_n10239, n5964, n3932);
not_3  g09863(new_n10240, new_n10239);
nand_4 g09864(new_n10241, new_n10240, new_n10230);
nand_4 g09865(new_n10242, new_n10241, new_n10234);
xor_3  g09866(new_n10243, new_n10242, new_n10238);
nand_4 g09867(new_n10244, n3932, n1097);
not_3  g09868(new_n10245, new_n10244);
nand_4 g09869(new_n10246, n4312, n1798);
nand_4 g09870(new_n10247, n12591, n5964);
xnor_3 g09871(new_n10248, new_n10247, new_n10246);
xor_3  g09872(new_n10249, new_n10248, new_n10245);
nor_4  g09873(new_n10250, new_n10249, new_n10243);
not_3  g09874(new_n10251, new_n10238);
xor_3  g09875(new_n10252, new_n10242, new_n10251);
xor_3  g09876(new_n10253, new_n10248, new_n10244);
nor_4  g09877(new_n10254, new_n10253, new_n10252);
nor_4  g09878(new_n10255, new_n10254, new_n10250);
nand_4 g09879(new_n10256, new_n10255, new_n10237);
nand_4 g09880(new_n10257, n11662, n5305);
nand_4 g09881(new_n10258, n7456, n5964);
nand_4 g09882(new_n10259, n4312, n3932);
nand_4 g09883(new_n10260, n12591, n1097);
nand_4 g09884(new_n10261, n12705, n1798);
xnor_3 g09885(new_n10262, new_n10261, new_n10260);
not_3  g09886(new_n10263, new_n10262);
nor_4  g09887(new_n10264, new_n10263, new_n10259);
not_3  g09888(new_n10265, new_n10259);
nor_4  g09889(new_n10266, new_n10262, new_n10265);
nor_4  g09890(new_n10267, new_n10266, new_n10264);
xnor_3 g09891(new_n10268, new_n10267, new_n10258);
and_4  g09892(new_n10269, new_n10247, new_n10246);
nor_4  g09893(new_n10270, new_n10248, new_n10245);
nor_4  g09894(new_n10271, new_n10270, new_n10269);
xnor_3 g09895(new_n10272, new_n10271, new_n10268);
not_3  g09896(new_n10273, new_n10272);
nor_4  g09897(new_n10274, new_n10273, new_n10257);
not_3  g09898(new_n10275, new_n10257);
nor_4  g09899(new_n10276, new_n10272, new_n10275);
nor_4  g09900(new_n10277, new_n10276, new_n10274);
not_3  g09901(new_n10278_1, new_n10242);
nor_4  g09902(new_n10279, new_n10278_1, new_n10238);
not_3  g09903(new_n10280, new_n10279);
nand_4 g09904(new_n10281, new_n10253, new_n10252);
nand_4 g09905(new_n10282, new_n10281, new_n10280);
xnor_3 g09906(new_n10283, new_n10282, new_n10277);
xor_3  g09907(new_n10284, new_n10283, new_n10256);
not_3  g09908(new_n10285, new_n10255);
xor_3  g09909(new_n10286, new_n10285, new_n10237);
not_3  g09910(new_n10287, new_n10286);
nand_4 g09911(new_n10288, n11023, n8759);
not_3  g09912(new_n10289, new_n10288);
nand_4 g09913(new_n10290, n8759, n3022);
nand_4 g09914(new_n10291, n12299, n6703);
nand_4 g09915(new_n10292, new_n10291, new_n10290);
nand_4 g09916(new_n10293, n9640, n6776);
not_3  g09917(new_n10294, new_n10293);
nand_4 g09918(new_n10295, new_n10294, new_n10292);
not_3  g09919(new_n10296, new_n10290);
not_3  g09920(new_n10297, new_n10291);
nand_4 g09921(new_n10298, new_n10297, new_n10296);
nand_4 g09922(new_n10299, new_n10298, new_n10295);
xor_3  g09923(new_n10300, new_n10299, new_n10289);
nand_4 g09924(new_n10301, n12299, n9640);
not_3  g09925(new_n10302, new_n10301);
nand_4 g09926(new_n10303, n6776, n3022);
not_3  g09927(new_n10304, new_n10303);
nand_4 g09928(new_n10305, n7436, n6703);
not_3  g09929(new_n10306, new_n10305);
nor_4  g09930(new_n10307, new_n10306, new_n10304);
nor_4  g09931(new_n10308, new_n10305, new_n10303);
nor_4  g09932(new_n10309, new_n10308, new_n10307);
xor_3  g09933(new_n10310, new_n10309, new_n10302);
xnor_3 g09934(new_n10311, new_n10310, new_n10300);
nor_4  g09935(new_n10312, new_n10293, new_n6530);
and_4  g09936(new_n10313, new_n10298, new_n10292);
nor_4  g09937(new_n10314, new_n10313, new_n10312);
not_3  g09938(new_n10315, new_n10314);
nor_4  g09939(new_n10316, new_n10315, new_n10293);
not_3  g09940(new_n10317, new_n10316);
xnor_3 g09941(new_n10318, new_n10317, new_n10311);
nor_4  g09942(new_n10319, new_n6556, new_n6555);
not_3  g09943(new_n10320, new_n10319);
nand_4 g09944(new_n10321, n5645, n2530);
not_3  g09945(new_n10322, new_n10321);
nand_4 g09946(new_n10323, n8665, n5331);
not_3  g09947(new_n10324, new_n10323);
nor_4  g09948(new_n10325, new_n10324, new_n10322);
nor_4  g09949(new_n10326, new_n10323, new_n10321);
nor_4  g09950(new_n10327_1, new_n10326, new_n10325);
nor_4  g09951(new_n10328, new_n10327_1, new_n10320);
not_3  g09952(new_n10329, new_n10328);
nand_4 g09953(new_n10330, n11922, n5331);
nand_4 g09954(new_n10331, n2530, n1067);
nand_4 g09955(new_n10332, n8665, n8476);
not_3  g09956(new_n10333, new_n10332);
nand_4 g09957(new_n10334, n12648, n5645);
not_3  g09958(new_n10335, new_n10334);
nor_4  g09959(new_n10336, new_n10335, new_n10333);
nor_4  g09960(new_n10337, new_n10334, new_n10332);
nor_4  g09961(new_n10338, new_n10337, new_n10336);
xnor_3 g09962(new_n10339, new_n10338, new_n10331);
not_3  g09963(new_n10340, new_n10339);
xnor_3 g09964(new_n10341, new_n10340, new_n10330);
not_3  g09965(new_n10342, new_n10325);
nand_4 g09966(new_n10343, n8476, n1067);
not_3  g09967(new_n10344, new_n10343);
nand_4 g09968(new_n10345, new_n10344, new_n10342);
not_3  g09969(new_n10346, new_n10345);
nor_4  g09970(new_n10347, new_n10346, new_n10326);
xnor_3 g09971(new_n10348, new_n10347, new_n10341);
xnor_3 g09972(new_n10349, new_n10348, new_n10329);
not_3  g09973(new_n10350, new_n10349);
nand_4 g09974(new_n10351, n7965, n2749);
nand_4 g09975(new_n10352, n7965, n3754);
nand_4 g09976(new_n10353, n11892, n11876);
nor_4  g09977(new_n10354, new_n10353, new_n10352);
not_3  g09978(new_n10355, new_n10354);
nand_4 g09979(new_n10356, new_n10353, new_n10352);
nand_4 g09980(new_n10357, n10898, n7388);
not_3  g09981(new_n10358, new_n10357);
nand_4 g09982(new_n10359, new_n10358, new_n10356);
nand_4 g09983(new_n10360, new_n10359, new_n10355);
not_3  g09984(new_n10361, new_n10360);
nor_4  g09985(new_n10362, new_n10361, new_n10351);
not_3  g09986(new_n10363, new_n10351);
nor_4  g09987(new_n10364, new_n10360, new_n10363);
nor_4  g09988(new_n10365, new_n10364, new_n10362);
nand_4 g09989(new_n10366, n11892, n10898);
nand_4 g09990(new_n10367, n7388, n3754);
nand_4 g09991(new_n10368, n11876, n2393);
xnor_3 g09992(new_n10369, new_n10368, new_n10367);
xnor_3 g09993(new_n10370, new_n10369, new_n10366);
not_3  g09994(new_n10371, new_n10370);
xnor_3 g09995(new_n10372, new_n10371, new_n10365);
not_3  g09996(new_n10373, new_n6532);
nor_4  g09997(new_n10374, new_n10357, new_n10373);
nand_4 g09998(new_n10375, new_n10356, new_n10355);
not_3  g09999(new_n10376, new_n10375);
nor_4  g10000(new_n10377, new_n10376, new_n10374);
not_3  g10001(new_n10378, new_n10377);
nor_4  g10002(new_n10379, new_n10378, new_n10357);
not_3  g10003(new_n10380, new_n10379);
xnor_3 g10004(new_n10381, new_n10380, new_n10372);
not_3  g10005(new_n10382, new_n10381);
nor_4  g10006(new_n10383, new_n10382, new_n10350);
nor_4  g10007(new_n10384, new_n10381, new_n10349);
nor_4  g10008(new_n10385, new_n10384, new_n10383);
not_3  g10009(new_n10386, new_n10385);
not_3  g10010(new_n10387, new_n6551);
nand_4 g10011(new_n10388, new_n6557, new_n6554);
nand_4 g10012(new_n10389, new_n10388, new_n10387);
nand_4 g10013(new_n10390, new_n10374, new_n10356);
nand_4 g10014(new_n10391_1, new_n10390, new_n10378);
not_3  g10015(new_n10392, new_n10391_1);
nor_4  g10016(new_n10393, new_n10392, new_n10389);
xnor_3 g10017(new_n10394, new_n10392, new_n10389);
not_3  g10018(new_n10395, new_n6531);
nor_4  g10019(new_n10396, new_n10343, new_n10395);
not_3  g10020(new_n10397, new_n10396);
nor_4  g10021(new_n10398, new_n10397, new_n10342);
not_3  g10022(new_n10399, new_n10327_1);
nor_4  g10023(new_n10400, new_n10396, new_n10399);
nor_4  g10024(new_n10401, new_n10400, new_n10398);
not_3  g10025(new_n10402, new_n10401);
nor_4  g10026(new_n10403, new_n10402, new_n10394);
nor_4  g10027(new_n10404, new_n10403, new_n10393);
xnor_3 g10028(new_n10405, new_n10404, new_n10386);
not_3  g10029(new_n10406, new_n10405);
nor_4  g10030(new_n10407, new_n10406, new_n10318);
not_3  g10031(new_n10408, new_n10318);
nor_4  g10032(new_n10409, new_n10405, new_n10408);
nor_4  g10033(new_n10410, new_n10409, new_n10407);
nand_4 g10034(new_n10411, new_n6544, new_n6541);
not_3  g10035(new_n10412, new_n10411);
nor_4  g10036(new_n10413, new_n6559, new_n10412);
not_3  g10037(new_n10414, new_n10413);
nor_4  g10038(new_n10415, new_n10295, new_n6530);
nor_4  g10039(new_n10416, new_n10415, new_n10314);
nor_4  g10040(new_n10417, new_n10416, new_n10414);
not_3  g10041(new_n10418, new_n10417);
not_3  g10042(new_n10419, new_n10394);
xor_3  g10043(new_n10420, new_n10401, new_n10419);
not_3  g10044(new_n10421, new_n10416);
nor_4  g10045(new_n10422, new_n10421, new_n10413);
nor_4  g10046(new_n10423, new_n10422, new_n10417);
nand_4 g10047(new_n10424, new_n10423, new_n10420);
nand_4 g10048(new_n10425, new_n10424, new_n10418);
xnor_3 g10049(new_n10426, new_n10425, new_n10410);
nand_4 g10050(new_n10427, new_n10426, new_n10287);
not_3  g10051(new_n10428, new_n10427);
nor_4  g10052(new_n10429, new_n10426, new_n10287);
nor_4  g10053(new_n10430, new_n10429, new_n10428);
xor_3  g10054(new_n10431, new_n10402, new_n10419);
not_3  g10055(new_n10432, new_n10423);
xnor_3 g10056(new_n10433, new_n10432, new_n10431);
not_3  g10057(new_n10434, new_n6528);
nor_4  g10058(new_n10435, new_n10239, new_n10434);
not_3  g10059(new_n10436, new_n10435);
nor_4  g10060(new_n10437, new_n10436, new_n10230);
not_3  g10061(new_n10438, new_n10236);
nor_4  g10062(new_n10439_1, new_n10435, new_n10438);
nor_4  g10063(new_n10440, new_n10439_1, new_n10437);
not_3  g10064(new_n10441, new_n10440);
nor_4  g10065(new_n10442, new_n10441, new_n10433);
nand_4 g10066(new_n10443, new_n6539, new_n6536);
nand_4 g10067(new_n10444, new_n6561, new_n6540);
nand_4 g10068(new_n10445, new_n10444, new_n10443);
xnor_3 g10069(new_n10446, new_n10441, new_n10433);
nor_4  g10070(new_n10447, new_n10446, new_n10445);
nor_4  g10071(new_n10448, new_n10447, new_n10442);
nand_4 g10072(new_n10449, new_n10448, new_n10430);
nand_4 g10073(new_n10450, new_n10449, new_n10427);
xnor_3 g10074(new_n10451_1, new_n10450, new_n10284);
nor_4  g10075(new_n10452, new_n10317, new_n10311);
nand_4 g10076(new_n10453, n10451, n8759);
nand_4 g10077(new_n10454, n11023, n6776);
not_3  g10078(new_n10455, new_n10454);
nor_4  g10079(new_n10456, new_n10308, new_n10302);
nor_4  g10080(new_n10457, new_n10456, new_n10307);
xnor_3 g10081(new_n10458, new_n10457, new_n10455);
nand_4 g10082(new_n10459, n9640, n7436);
nand_4 g10083(new_n10460, n12299, n3022);
not_3  g10084(new_n10461, new_n10460);
nand_4 g10085(new_n10462, n8276, n6703);
not_3  g10086(new_n10463, new_n10462);
nor_4  g10087(new_n10464, new_n10463, new_n10461);
not_3  g10088(new_n10465, new_n10464);
nor_4  g10089(new_n10466, new_n10462, new_n10460);
not_3  g10090(new_n10467, new_n10466);
nand_4 g10091(new_n10468, new_n10467, new_n10465);
xnor_3 g10092(new_n10469, new_n10468, new_n10459);
xnor_3 g10093(new_n10470, new_n10469, new_n10458);
nor_4  g10094(new_n10471, new_n10470, new_n10453);
not_3  g10095(new_n10472, new_n10453);
not_3  g10096(new_n10473, new_n10470);
nor_4  g10097(new_n10474, new_n10473, new_n10472);
nor_4  g10098(new_n10475, new_n10474, new_n10471);
not_3  g10099(new_n10476_1, new_n10475);
not_3  g10100(new_n10477, new_n10299);
nor_4  g10101(new_n10478, new_n10477, new_n10288);
not_3  g10102(new_n10479, new_n10478);
nand_4 g10103(new_n10480, new_n10310, new_n10300);
nand_4 g10104(new_n10481, new_n10480, new_n10479);
xnor_3 g10105(new_n10482, new_n10481, new_n10476_1);
xnor_3 g10106(new_n10483, new_n10482, new_n10452);
not_3  g10107(new_n10484, new_n10483);
nor_4  g10108(new_n10485, new_n10380, new_n10372);
nand_4 g10109(new_n10486, n7965, n159);
not_3  g10110(new_n10487, new_n10362);
nand_4 g10111(new_n10488, new_n10371, new_n10365);
nand_4 g10112(new_n10489, new_n10488, new_n10487);
not_3  g10113(new_n10490, new_n10489);
xnor_3 g10114(new_n10491, new_n10490, new_n10486);
nand_4 g10115(new_n10492, n7388, n2749);
not_3  g10116(new_n10493, new_n10492);
not_3  g10117(new_n10494, new_n10367);
not_3  g10118(new_n10495, new_n10368);
nor_4  g10119(new_n10496, new_n10495, new_n10494);
not_3  g10120(new_n10497, new_n10366);
nor_4  g10121(new_n10498, new_n10369, new_n10497);
nor_4  g10122(new_n10499, new_n10498, new_n10496);
nand_4 g10123(new_n10500, new_n10499, new_n10493);
not_3  g10124(new_n10501, new_n10500);
nor_4  g10125(new_n10502, new_n10499, new_n10493);
nor_4  g10126(new_n10503, new_n10502, new_n10501);
nand_4 g10127(new_n10504, n11892, n3754);
not_3  g10128(new_n10505, new_n10504);
nand_4 g10129(new_n10506, n11876, n5860);
nand_4 g10130(new_n10507, n10898, n2393);
xnor_3 g10131(new_n10508, new_n10507, new_n10506);
xnor_3 g10132(new_n10509, new_n10508, new_n10505);
xnor_3 g10133(new_n10510_1, new_n10509, new_n10503);
xnor_3 g10134(new_n10511, new_n10510_1, new_n10491);
xnor_3 g10135(new_n10512, new_n10511, new_n10485);
nor_4  g10136(new_n10513, new_n10348, new_n10329);
nand_4 g10137(new_n10514, n5331, n2551);
nand_4 g10138(new_n10515, n11922, n8476);
not_3  g10139(new_n10516, new_n10515);
not_3  g10140(new_n10517, new_n10331);
nor_4  g10141(new_n10518, new_n10337, new_n10517);
nor_4  g10142(new_n10519, new_n10518, new_n10336);
xnor_3 g10143(new_n10520, new_n10519, new_n10516);
nand_4 g10144(new_n10521, n12648, n1067);
not_3  g10145(new_n10522, new_n10521);
nand_4 g10146(new_n10523, n8665, n2530);
not_3  g10147(new_n10524, new_n10523);
nand_4 g10148(new_n10525, n10545, n5645);
not_3  g10149(new_n10526, new_n10525);
nor_4  g10150(new_n10527, new_n10526, new_n10524);
not_3  g10151(new_n10528, new_n10527);
nor_4  g10152(new_n10529, new_n10525, new_n10523);
not_3  g10153(new_n10530, new_n10529);
nand_4 g10154(new_n10531, new_n10530, new_n10528);
xnor_3 g10155(new_n10532, new_n10531, new_n10522);
xnor_3 g10156(new_n10533, new_n10532, new_n10520);
not_3  g10157(new_n10534, new_n10533);
nor_4  g10158(new_n10535, new_n10534, new_n10514);
not_3  g10159(new_n10536, new_n10514);
nor_4  g10160(new_n10537, new_n10533, new_n10536);
nor_4  g10161(new_n10538, new_n10537, new_n10535);
nor_4  g10162(new_n10539, new_n10340, new_n10330);
nor_4  g10163(new_n10540, new_n10347, new_n10341);
nor_4  g10164(new_n10541, new_n10540, new_n10539);
not_3  g10165(new_n10542, new_n10541);
xnor_3 g10166(new_n10543, new_n10542, new_n10538);
not_3  g10167(new_n10544, new_n10543);
nor_4  g10168(new_n10545_1, new_n10544, new_n10513);
not_3  g10169(new_n10546, new_n10513);
nor_4  g10170(new_n10547_1, new_n10543, new_n10546);
nor_4  g10171(new_n10548, new_n10547_1, new_n10545_1);
xnor_3 g10172(new_n10549, new_n10548, new_n10512);
not_3  g10173(new_n10550, new_n10549);
not_3  g10174(new_n10551, new_n10383);
not_3  g10175(new_n10552, new_n10404);
nand_4 g10176(new_n10553, new_n10552, new_n10385);
nand_4 g10177(new_n10554, new_n10553, new_n10551);
xnor_3 g10178(new_n10555, new_n10554, new_n10550);
xnor_3 g10179(new_n10556, new_n10555, new_n10484);
not_3  g10180(new_n10557, new_n10409);
nand_4 g10181(new_n10558, new_n10425, new_n10410);
nand_4 g10182(new_n10559, new_n10558, new_n10557);
xnor_3 g10183(new_n10560, new_n10559, new_n10556);
xor_3  g10184(n3677, new_n10560, new_n10451_1);
not_3  g10185(new_n10562, new_n9136);
xor_3  g10186(n3849, new_n9137_1, new_n10562);
xor_3  g10187(n4088, new_n6524, new_n6523);
xor_3  g10188(n4155, new_n1197, new_n1095);
not_3  g10189(new_n10566, new_n3091);
nand_4 g10190(new_n10567, new_n3049, new_n3048);
xnor_3 g10191(n4159, new_n10567, new_n10566);
xor_3  g10192(n4226, new_n6511, new_n6313);
nand_4 g10193(new_n10570, n12591, n4312);
not_3  g10194(new_n10571, new_n10570);
nand_4 g10195(new_n10572, new_n10261, new_n10260);
not_3  g10196(new_n10573, new_n10572);
nor_4  g10197(new_n10574, new_n10266, new_n10573);
xnor_3 g10198(new_n10575, new_n10574, new_n10571);
not_3  g10199(new_n10576, new_n10575);
nand_4 g10200(new_n10577, n12705, n3932);
nand_4 g10201(new_n10578, n12025, n1798);
not_3  g10202(new_n10579, new_n10578);
xor_3  g10203(new_n10580, new_n10579, new_n10577);
xnor_3 g10204(new_n10581, new_n10580, new_n10576);
nand_4 g10205(new_n10582, n11662, n5964);
nand_4 g10206(new_n10583, n7456, n1097);
xor_3  g10207(new_n10584, new_n10583, new_n10582);
xnor_3 g10208(new_n10585, new_n10584, new_n10581);
nor_4  g10209(new_n10586, new_n10267, new_n10258);
not_3  g10210(new_n10587, new_n10271);
nor_4  g10211(new_n10588, new_n10587, new_n10268);
nor_4  g10212(new_n10589_1, new_n10588, new_n10586);
xnor_3 g10213(new_n10590, new_n10589_1, new_n10585);
not_3  g10214(new_n10591, new_n10590);
not_3  g10215(new_n10592, new_n10274);
nand_4 g10216(new_n10593, new_n10282, new_n10277);
nand_4 g10217(new_n10594, new_n10593, new_n10592);
nand_4 g10218(new_n10595, new_n10594, new_n10591);
nor_4  g10219(new_n10596, new_n10574, new_n10571);
not_3  g10220(new_n10597, new_n10596);
nand_4 g10221(new_n10598, new_n10580, new_n10576);
nand_4 g10222(new_n10599, new_n10598, new_n10597);
nand_4 g10223(new_n10600, n10327, n5964);
nand_4 g10224(new_n10601, n11662, n1097);
nand_4 g10225(new_n10602, n9583, n5305);
not_3  g10226(new_n10603, new_n10602);
xor_3  g10227(new_n10604, new_n10603, new_n10601);
xnor_3 g10228(new_n10605, new_n10604, new_n10600);
xnor_3 g10229(new_n10606, new_n10605, new_n10599);
nor_4  g10230(new_n10607, new_n10578, new_n10577);
nand_4 g10231(new_n10608, n7456, n4312);
not_3  g10232(new_n10609, new_n10608);
xor_3  g10233(new_n10610, new_n10609, new_n10607);
not_3  g10234(new_n10611, new_n10610);
nand_4 g10235(new_n10612, n12025, n3932);
nand_4 g10236(new_n10613, n12705, n12591);
nand_4 g10237(new_n10614, n11257, n1798);
not_3  g10238(new_n10615, new_n10614);
xor_3  g10239(new_n10616, new_n10615, new_n10613);
xnor_3 g10240(new_n10617, new_n10616, new_n10612);
not_3  g10241(new_n10618, new_n10617);
nor_4  g10242(new_n10619, new_n10618, new_n10611);
nor_4  g10243(new_n10620, new_n10617, new_n10610);
nor_4  g10244(new_n10621, new_n10620, new_n10619);
xnor_3 g10245(new_n10622, new_n10621, new_n10606);
nand_4 g10246(new_n10623, new_n10584, new_n10581);
nor_4  g10247(new_n10624, new_n10583, new_n10582);
nor_4  g10248(new_n10625, new_n10589_1, new_n10585);
xnor_3 g10249(new_n10626, new_n10625, new_n10624);
nand_4 g10250(new_n10627, new_n10626, new_n10623);
xnor_3 g10251(new_n10628, new_n10627, new_n10622);
xnor_3 g10252(new_n10629, new_n10628, new_n10595);
nand_4 g10253(new_n10630, n10327, n5305);
not_3  g10254(new_n10631, new_n10630);
xnor_3 g10255(new_n10632, new_n10594, new_n10590);
nor_4  g10256(new_n10633, new_n10632, new_n10631);
nor_4  g10257(new_n10634, new_n10283, new_n10256);
xnor_3 g10258(new_n10635, new_n10632, new_n10631);
nor_4  g10259(new_n10636, new_n10635, new_n10634);
nor_4  g10260(new_n10637, new_n10636, new_n10633);
xnor_3 g10261(new_n10638, new_n10637, new_n10629);
nand_4 g10262(new_n10639, new_n10457, new_n10455);
not_3  g10263(new_n10640, new_n10458);
not_3  g10264(new_n10641, new_n10469);
nand_4 g10265(new_n10642, new_n10641, new_n10640);
nand_4 g10266(new_n10643, new_n10642, new_n10639);
nand_4 g10267(new_n10644_1, n10451, n6776);
nand_4 g10268(new_n10645, n12299, n11023);
xor_3  g10269(new_n10646, new_n10645, new_n10644_1);
xnor_3 g10270(new_n10647, new_n10646, new_n10643);
not_3  g10271(new_n10648, new_n10647);
nand_4 g10272(new_n10649, n7436, n3022);
not_3  g10273(new_n10650, new_n10649);
nand_4 g10274(new_n10651, n9640, n8276);
nand_4 g10275(new_n10652, n9241, n6703);
not_3  g10276(new_n10653, new_n10652);
xor_3  g10277(new_n10654, new_n10653, new_n10651);
xnor_3 g10278(new_n10655, new_n10654, new_n10650);
not_3  g10279(new_n10656, new_n10459);
nor_4  g10280(new_n10657, new_n10466, new_n10656);
nor_4  g10281(new_n10658, new_n10657, new_n10464);
xnor_3 g10282(new_n10659, new_n10658, new_n10655);
xnor_3 g10283(new_n10660, new_n10659, new_n10648);
not_3  g10284(new_n10661, new_n10471);
nand_4 g10285(new_n10662, new_n10481, new_n10475);
nand_4 g10286(new_n10663, new_n10662, new_n10661);
nand_4 g10287(new_n10664, new_n10663, new_n10660);
nand_4 g10288(new_n10665, new_n10654, new_n10649);
not_3  g10289(new_n10666, new_n10658);
nand_4 g10290(new_n10667, new_n10666, new_n10655);
nand_4 g10291(new_n10668, new_n10667, new_n10665);
nand_4 g10292(new_n10669, n10278, n6776);
nand_4 g10293(new_n10670, n12299, n10451);
nand_4 g10294(new_n10671, n11423, n8759);
not_3  g10295(new_n10672, new_n10671);
xor_3  g10296(new_n10673, new_n10672, new_n10670);
xnor_3 g10297(new_n10674, new_n10673, new_n10669);
not_3  g10298(new_n10675, new_n10674);
xnor_3 g10299(new_n10676, new_n10675, new_n10668);
nor_4  g10300(new_n10677, new_n10652, new_n10651);
nand_4 g10301(new_n10678_1, n11023, n7436);
not_3  g10302(new_n10679, new_n10678_1);
xor_3  g10303(new_n10680, new_n10679, new_n10677);
nand_4 g10304(new_n10681, n9640, n9241);
nand_4 g10305(new_n10682, n8276, n3022);
nand_4 g10306(new_n10683, n10510, n6703);
not_3  g10307(new_n10684, new_n10683);
xor_3  g10308(new_n10685_1, new_n10684, new_n10682);
xnor_3 g10309(new_n10686, new_n10685_1, new_n10681);
not_3  g10310(new_n10687, new_n10686);
nor_4  g10311(new_n10688, new_n10687, new_n10680);
not_3  g10312(new_n10689, new_n10680);
nor_4  g10313(new_n10690, new_n10686, new_n10689);
nor_4  g10314(new_n10691, new_n10690, new_n10688);
not_3  g10315(new_n10692, new_n10691);
xnor_3 g10316(new_n10693, new_n10692, new_n10676);
nand_4 g10317(new_n10694, new_n10646, new_n10643);
nor_4  g10318(new_n10695_1, new_n10645, new_n10644_1);
nor_4  g10319(new_n10696, new_n10659, new_n10647);
xnor_3 g10320(new_n10697, new_n10696, new_n10695_1);
nand_4 g10321(new_n10698, new_n10697, new_n10694);
xnor_3 g10322(new_n10699, new_n10698, new_n10693);
xnor_3 g10323(new_n10700, new_n10699, new_n10664);
nand_4 g10324(new_n10701, n10278, n8759);
xnor_3 g10325(new_n10702, new_n10663, new_n10660);
nor_4  g10326(new_n10703, new_n10702, new_n10701);
nand_4 g10327(new_n10704, new_n10482, new_n10452);
xnor_3 g10328(new_n10705, new_n10702, new_n10701);
nor_4  g10329(new_n10706, new_n10705, new_n10704);
nor_4  g10330(new_n10707, new_n10706, new_n10703);
xnor_3 g10331(new_n10708, new_n10707, new_n10700);
nand_4 g10332(new_n10709, n12648, n8665);
nand_4 g10333(new_n10710, n10545, n1067);
nand_4 g10334(new_n10711, n7690, n5645);
xnor_3 g10335(new_n10712, new_n10711, new_n10710);
nor_4  g10336(new_n10713, new_n10712, new_n10709);
not_3  g10337(new_n10714, new_n10709);
not_3  g10338(new_n10715, new_n10712);
nor_4  g10339(new_n10716, new_n10715, new_n10714);
nor_4  g10340(new_n10717, new_n10716, new_n10713);
nor_4  g10341(new_n10718, new_n10529, new_n10522);
nor_4  g10342(new_n10719, new_n10718, new_n10527);
xnor_3 g10343(new_n10720, new_n10719, new_n10717);
not_3  g10344(new_n10721, new_n10720);
nand_4 g10345(new_n10722, n8476, n2551);
nand_4 g10346(new_n10723, n11922, n2530);
xor_3  g10347(new_n10724, new_n10723, new_n10722);
xnor_3 g10348(new_n10725, new_n10724, new_n10721);
and_4  g10349(new_n10726, new_n10519, new_n10516);
not_3  g10350(new_n10727, new_n10532);
nor_4  g10351(new_n10728, new_n10727, new_n10520);
nor_4  g10352(new_n10729, new_n10728, new_n10726);
xnor_3 g10353(new_n10730, new_n10729, new_n10725);
not_3  g10354(new_n10731, new_n10535);
not_3  g10355(new_n10732, new_n10537);
nand_4 g10356(new_n10733, new_n10542, new_n10732);
nand_4 g10357(new_n10734, new_n10733, new_n10731);
not_3  g10358(new_n10735, new_n10734);
nor_4  g10359(new_n10736, new_n10735, new_n10730);
nor_4  g10360(new_n10737, new_n10711, new_n10710);
nand_4 g10361(new_n10738, n12648, n11922);
not_3  g10362(new_n10739, new_n10738);
xor_3  g10363(new_n10740, new_n10739, new_n10737);
nand_4 g10364(new_n10741, n7690, n1067);
not_3  g10365(new_n10742, new_n10741);
nand_4 g10366(new_n10743, n10545, n8665);
nand_4 g10367(new_n10744, n5645, n3616);
xnor_3 g10368(new_n10745, new_n10744, new_n10743);
xnor_3 g10369(new_n10746, new_n10745, new_n10742);
xnor_3 g10370(new_n10747, new_n10746, new_n10740);
not_3  g10371(new_n10748, new_n10747);
nand_4 g10372(new_n10749, new_n10719, new_n10717);
not_3  g10373(new_n10750, new_n10749);
nor_4  g10374(new_n10751, new_n10750, new_n10713);
not_3  g10375(new_n10752, new_n10751);
nand_4 g10376(new_n10753, n12826, n8476);
not_3  g10377(new_n10754, new_n10753);
nand_4 g10378(new_n10755, n2551, n2530);
nand_4 g10379(new_n10756, n5331, n4094);
xnor_3 g10380(new_n10757, new_n10756, new_n10755);
xor_3  g10381(new_n10758, new_n10757, new_n10754);
xnor_3 g10382(new_n10759, new_n10758, new_n10752);
xnor_3 g10383(new_n10760, new_n10759, new_n10748);
nand_4 g10384(new_n10761, new_n10724, new_n10721);
nor_4  g10385(new_n10762, new_n10723, new_n10722);
nor_4  g10386(new_n10763, new_n10729, new_n10725);
xnor_3 g10387(new_n10764, new_n10763, new_n10762);
nand_4 g10388(new_n10765, new_n10764, new_n10761);
xnor_3 g10389(new_n10766, new_n10765, new_n10760);
xnor_3 g10390(new_n10767, new_n10766, new_n10736);
nand_4 g10391(new_n10768, n12826, n5331);
not_3  g10392(new_n10769, new_n10768);
xnor_3 g10393(new_n10770, new_n10734, new_n10730);
nand_4 g10394(new_n10771, new_n10770, new_n10769);
not_3  g10395(new_n10772, new_n10770);
nand_4 g10396(new_n10773, new_n10772, new_n10768);
nand_4 g10397(new_n10774, new_n10773, new_n10547_1);
nand_4 g10398(new_n10775, new_n10774, new_n10771);
xnor_3 g10399(new_n10776, new_n10775, new_n10767);
not_3  g10400(new_n10777, new_n10776);
nand_4 g10401(new_n10778, n7965, n1510);
not_3  g10402(new_n10779, new_n10778);
nand_4 g10403(new_n10780, new_n10509, new_n10503);
nand_4 g10404(new_n10781, new_n10780, new_n10500);
nand_4 g10405(new_n10782, n7388, n159);
nand_4 g10406(new_n10783, n11892, n2749);
xor_3  g10407(new_n10784, new_n10783, new_n10782);
xnor_3 g10408(new_n10785, new_n10784, new_n10781);
nand_4 g10409(new_n10786, n3754, n2393);
nand_4 g10410(new_n10787, n10898, n5860);
nand_4 g10411(new_n10788, n11876, n3986);
xnor_3 g10412(new_n10789_1, new_n10788, new_n10787);
nor_4  g10413(new_n10790, new_n10789_1, new_n10786);
not_3  g10414(new_n10791, new_n10786);
not_3  g10415(new_n10792, new_n10789_1);
nor_4  g10416(new_n10793, new_n10792, new_n10791);
nor_4  g10417(new_n10794, new_n10793, new_n10790);
and_4  g10418(new_n10795, new_n10507, new_n10506);
nor_4  g10419(new_n10796, new_n10508, new_n10505);
nor_4  g10420(new_n10797, new_n10796, new_n10795);
nand_4 g10421(new_n10798, new_n10797, new_n10794);
not_3  g10422(new_n10799, new_n10798);
nor_4  g10423(new_n10800, new_n10797, new_n10794);
nor_4  g10424(new_n10801, new_n10800, new_n10799);
xnor_3 g10425(new_n10802, new_n10801, new_n10785);
nor_4  g10426(new_n10803, new_n10490, new_n10486);
nor_4  g10427(new_n10804, new_n10510_1, new_n10491);
nor_4  g10428(new_n10805, new_n10804, new_n10803);
xnor_3 g10429(new_n10806, new_n10805, new_n10802);
nand_4 g10430(new_n10807, new_n10806, new_n10779);
not_3  g10431(new_n10808, new_n10485);
nor_4  g10432(new_n10809, new_n10511, new_n10808);
xnor_3 g10433(new_n10810, new_n10806, new_n10778);
nand_4 g10434(new_n10811, new_n10810, new_n10809);
nand_4 g10435(new_n10812, new_n10811, new_n10807);
not_3  g10436(new_n10813, new_n10802);
nor_4  g10437(new_n10814, new_n10805, new_n10813);
nor_4  g10438(new_n10815, new_n10783, new_n10782);
nor_4  g10439(new_n10816, new_n10784, new_n10781);
nor_4  g10440(new_n10817, new_n10801, new_n10785);
nor_4  g10441(new_n10818, new_n10817, new_n10816);
xnor_3 g10442(new_n10819, new_n10818, new_n10815);
not_3  g10443(new_n10820, new_n10790);
nand_4 g10444(new_n10821, new_n10798, new_n10820);
nand_4 g10445(new_n10822, n7388, n1510);
not_3  g10446(new_n10823, new_n10822);
nand_4 g10447(new_n10824, n11892, n159);
not_3  g10448(new_n10825, new_n10824);
nand_4 g10449(new_n10826, n12247, n7965);
not_3  g10450(new_n10827, new_n10826);
nand_4 g10451(new_n10828, new_n10827, new_n10825);
nand_4 g10452(new_n10829, new_n10826, new_n10824);
nand_4 g10453(new_n10830, new_n10829, new_n10828);
xor_3  g10454(new_n10831, new_n10830, new_n10823);
xnor_3 g10455(new_n10832, new_n10831, new_n10821);
nor_4  g10456(new_n10833, new_n10788, new_n10787);
nand_4 g10457(new_n10834, n2749, n2393);
not_3  g10458(new_n10835, new_n10834);
xor_3  g10459(new_n10836, new_n10835, new_n10833);
not_3  g10460(new_n10837, new_n10836);
nand_4 g10461(new_n10838, n10898, n3986);
not_3  g10462(new_n10839, new_n10838);
nand_4 g10463(new_n10840, n11876, n5857);
nand_4 g10464(new_n10841, n5860, n3754);
not_3  g10465(new_n10842, new_n10841);
xor_3  g10466(new_n10843, new_n10842, new_n10840);
xnor_3 g10467(new_n10844, new_n10843, new_n10839);
xnor_3 g10468(new_n10845, new_n10844, new_n10837);
xnor_3 g10469(new_n10846, new_n10845, new_n10832);
xnor_3 g10470(new_n10847, new_n10846, new_n10819);
xnor_3 g10471(new_n10848_1, new_n10847, new_n10814);
xnor_3 g10472(new_n10849, new_n10848_1, new_n10812);
xnor_3 g10473(new_n10850, new_n10849, new_n10777);
xnor_3 g10474(new_n10851_1, new_n10810, new_n10809);
nand_4 g10475(new_n10852, new_n10773, new_n10771);
xnor_3 g10476(new_n10853, new_n10852, new_n10547_1);
not_3  g10477(new_n10854, new_n10853);
nand_4 g10478(new_n10855, new_n10854, new_n10851_1);
nor_4  g10479(new_n10856, new_n10548, new_n10512);
not_3  g10480(new_n10857, new_n10856);
nand_4 g10481(new_n10858, new_n10554, new_n10550);
nand_4 g10482(new_n10859, new_n10858, new_n10857);
xnor_3 g10483(new_n10860, new_n10853, new_n10851_1);
nand_4 g10484(new_n10861, new_n10860, new_n10859);
nand_4 g10485(new_n10862, new_n10861, new_n10855);
xnor_3 g10486(new_n10863, new_n10862, new_n10850);
xnor_3 g10487(new_n10864, new_n10863, new_n10708);
not_3  g10488(new_n10865, new_n10704);
not_3  g10489(new_n10866, new_n10705);
nor_4  g10490(new_n10867, new_n10866, new_n10865);
nor_4  g10491(new_n10868, new_n10867, new_n10706);
not_3  g10492(new_n10869, new_n10868);
not_3  g10493(new_n10870, new_n10860);
xnor_3 g10494(new_n10871, new_n10870, new_n10859);
nand_4 g10495(new_n10872, new_n10871, new_n10869);
nand_4 g10496(new_n10873, new_n10555, new_n10484);
not_3  g10497(new_n10874, new_n10873);
nor_4  g10498(new_n10875, new_n10559, new_n10556);
nor_4  g10499(new_n10876, new_n10875, new_n10874);
xnor_3 g10500(new_n10877, new_n10871, new_n10868);
nand_4 g10501(new_n10878, new_n10877, new_n10876);
nand_4 g10502(new_n10879, new_n10878, new_n10872);
xnor_3 g10503(new_n10880, new_n10879, new_n10864);
nand_4 g10504(new_n10881, new_n10880, new_n10638);
not_3  g10505(new_n10882, new_n10638);
xnor_3 g10506(new_n10883, new_n10880, new_n10882);
not_3  g10507(new_n10884, new_n10635);
xor_3  g10508(new_n10885, new_n10884, new_n10634);
not_3  g10509(new_n10886, new_n10885);
not_3  g10510(new_n10887, new_n10877);
xnor_3 g10511(new_n10888, new_n10887, new_n10876);
nand_4 g10512(new_n10889, new_n10888, new_n10886);
not_3  g10513(new_n10890, new_n10889);
nor_4  g10514(new_n10891, new_n10888, new_n10886);
nor_4  g10515(new_n10892, new_n10891, new_n10890);
not_3  g10516(new_n10893, new_n10284);
not_3  g10517(new_n10894, new_n10450);
nor_4  g10518(new_n10895, new_n10894, new_n10893);
nor_4  g10519(new_n10896, new_n10560, new_n10451_1);
nor_4  g10520(new_n10897, new_n10896, new_n10895);
nand_4 g10521(new_n10898_1, new_n10897, new_n10892);
nand_4 g10522(new_n10899, new_n10898_1, new_n10889);
nand_4 g10523(new_n10900, new_n10899, new_n10883);
nand_4 g10524(new_n10901, new_n10900, new_n10881);
nand_4 g10525(new_n10902, new_n10863, new_n10708);
not_3  g10526(new_n10903, new_n10708);
xnor_3 g10527(new_n10904, new_n10863, new_n10903);
nand_4 g10528(new_n10905, new_n10879, new_n10904);
nand_4 g10529(new_n10906, new_n10905, new_n10902);
nand_4 g10530(new_n10907, new_n10696, new_n10695_1);
nand_4 g10531(new_n10908, new_n10698, new_n10693);
nand_4 g10532(new_n10909, new_n10908, new_n10907);
and_4  g10533(new_n10910, new_n10679, new_n10677);
or_4   g10534(new_n10911, new_n10690, new_n10910);
not_3  g10535(new_n10912, new_n10670);
nor_4  g10536(new_n10913_1, new_n10672, new_n10912);
not_3  g10537(new_n10914, new_n10669);
nor_4  g10538(new_n10915, new_n10673, new_n10914);
nor_4  g10539(new_n10916, new_n10915, new_n10913_1);
nand_4 g10540(new_n10917, n12511, n7965);
xor_3  g10541(new_n10918, new_n10917, new_n10916);
nand_4 g10542(new_n10919, n8759, n2278);
nand_4 g10543(new_n10920, n10510, n9640);
xor_3  g10544(new_n10921, new_n10920, new_n10919);
xnor_3 g10545(new_n10922, new_n10921, new_n10918);
xnor_3 g10546(new_n10923, new_n10922, new_n10911);
xnor_3 g10547(new_n10924, new_n10923, new_n10909);
xnor_3 g10548(new_n10925, new_n10924, new_n10906);
nand_4 g10549(new_n10926, new_n10849, new_n10777);
not_3  g10550(new_n10927, new_n10850);
nand_4 g10551(new_n10928_1, new_n10862, new_n10927);
nand_4 g10552(new_n10929, new_n10928_1, new_n10926);
not_3  g10553(new_n10930, new_n10847);
nand_4 g10554(new_n10931, new_n10930, new_n10814);
nand_4 g10555(new_n10932, new_n10848_1, new_n10812);
nand_4 g10556(new_n10933, new_n10932, new_n10931);
nor_4  g10557(new_n10934, new_n10699, new_n10664);
nor_4  g10558(new_n10935, new_n10707, new_n10700);
nor_4  g10559(new_n10936, new_n10935, new_n10934);
nand_4 g10560(new_n10937, new_n10766, new_n10736);
not_3  g10561(new_n10938, new_n10767);
nand_4 g10562(new_n10939, new_n10775, new_n10938);
nand_4 g10563(new_n10940, new_n10939, new_n10937);
not_3  g10564(new_n10941, new_n10821);
nand_4 g10565(new_n10942, new_n10831, new_n10941);
not_3  g10566(new_n10943, new_n10845);
nand_4 g10567(new_n10944, new_n10943, new_n10832);
nand_4 g10568(new_n10945, new_n10944, new_n10942);
nand_4 g10569(new_n10946, new_n10829, new_n10823);
and_4  g10570(new_n10947, new_n10946, new_n10828);
nand_4 g10571(new_n10948, n11892, n1510);
nand_4 g10572(new_n10949_1, n2393, n159);
xor_3  g10573(new_n10950, new_n10949_1, new_n10948);
xnor_3 g10574(new_n10951, new_n10950, new_n10947);
not_3  g10575(new_n10952, new_n10840);
nor_4  g10576(new_n10953, new_n10842, new_n10952);
nor_4  g10577(new_n10954, new_n10843, new_n10839);
nor_4  g10578(new_n10955, new_n10954, new_n10953);
nand_4 g10579(new_n10956, n5860, n2749);
nand_4 g10580(new_n10957, n10685, n5331);
nand_4 g10581(new_n10958, n5645, n4499);
xor_3  g10582(new_n10959, new_n10958, new_n10957);
xnor_3 g10583(new_n10960, new_n10959, new_n10956);
xnor_3 g10584(new_n10961, new_n10960, new_n10955);
xnor_3 g10585(new_n10962, new_n10961, new_n10951);
nand_4 g10586(new_n10963, new_n10835, new_n10833);
nand_4 g10587(new_n10964, new_n10844, new_n10836);
nand_4 g10588(new_n10965_1, new_n10964, new_n10963);
nand_4 g10589(new_n10966, n12247, n7388);
not_3  g10590(new_n10967, new_n10966);
xnor_3 g10591(new_n10968, new_n10967, new_n10965_1);
xnor_3 g10592(new_n10969, new_n10968, new_n10962);
xnor_3 g10593(new_n10970, new_n10969, new_n10945);
xnor_3 g10594(new_n10971, new_n10970, new_n10940);
xnor_3 g10595(new_n10972, new_n10971, new_n10936);
xnor_3 g10596(new_n10973, new_n10972, new_n10933);
xnor_3 g10597(new_n10974, new_n10973, new_n10929);
nand_4 g10598(new_n10975, new_n10758, new_n10751);
nand_4 g10599(new_n10976, new_n10759, new_n10747);
nand_4 g10600(new_n10977, new_n10976, new_n10975);
nand_4 g10601(new_n10978, n12648, n2551);
not_3  g10602(new_n10979, new_n10978);
and_4  g10603(new_n10980, new_n10756, new_n10755);
nor_4  g10604(new_n10981, new_n10757, new_n10754);
nor_4  g10605(new_n10982, new_n10981, new_n10980);
xnor_3 g10606(new_n10983, new_n10982, new_n10979);
and_4  g10607(new_n10984, new_n10744, new_n10743);
nor_4  g10608(new_n10985, new_n10745, new_n10742);
nor_4  g10609(new_n10986, new_n10985, new_n10984);
nand_4 g10610(new_n10987, n11922, n10545);
nand_4 g10611(new_n10988, n8665, n7690);
xnor_3 g10612(new_n10989, new_n10988, new_n10987);
nand_4 g10613(new_n10990_1, n8476, n4094);
nand_4 g10614(new_n10991, n12826, n2530);
xnor_3 g10615(new_n10992, new_n10991, new_n10990_1);
xnor_3 g10616(new_n10993, new_n10992, new_n10989);
xnor_3 g10617(new_n10994, new_n10993, new_n10986);
xnor_3 g10618(new_n10995, new_n10994, new_n10983);
nand_4 g10619(new_n10996, new_n10739, new_n10737);
nand_4 g10620(new_n10997, new_n10746, new_n10740);
nand_4 g10621(new_n10998, new_n10997, new_n10996);
nand_4 g10622(new_n10999, n10547, n1798);
not_3  g10623(new_n11000, new_n10999);
xnor_3 g10624(new_n11001, new_n11000, new_n10998);
xnor_3 g10625(new_n11002, new_n11001, new_n10995);
xnor_3 g10626(new_n11003, new_n11002, new_n10977);
nand_4 g10627(new_n11004, n3616, n1067);
nand_4 g10628(new_n11005, n5305, n753);
xor_3  g10629(new_n11006, new_n11005, new_n11004);
xnor_3 g10630(new_n11007, new_n11006, new_n11003);
nand_4 g10631(new_n11008, new_n10763, new_n10762);
not_3  g10632(new_n11009, new_n10760);
nand_4 g10633(new_n11010, new_n10765, new_n11009);
nand_4 g10634(new_n11011, new_n11010, new_n11008);
xnor_3 g10635(new_n11012, new_n11011, new_n11007);
not_3  g10636(new_n11013, new_n10682);
nor_4  g10637(new_n11014, new_n10684, new_n11013);
not_3  g10638(new_n11015, new_n10681);
nor_4  g10639(new_n11016, new_n10685_1, new_n11015);
nor_4  g10640(new_n11017, new_n11016, new_n11014);
nand_4 g10641(new_n11018, n10451, n7436);
nand_4 g10642(new_n11019, n9241, n3022);
xor_3  g10643(new_n11020, new_n11019, new_n11018);
nand_4 g10644(new_n11021, n11423, n6776);
nand_4 g10645(new_n11022, n11023, n8276);
not_3  g10646(new_n11023_1, new_n11022);
xor_3  g10647(new_n11024, new_n11023_1, new_n11021);
xor_3  g10648(new_n11025, new_n11024, new_n11020);
xnor_3 g10649(new_n11026, new_n11025, new_n11017);
nand_4 g10650(new_n11027, n12299, n10278);
nand_4 g10651(new_n11028, n10644, n6703);
not_3  g10652(new_n11029, new_n11028);
xor_3  g10653(new_n11030, new_n11029, new_n11027);
xnor_3 g10654(new_n11031, new_n11030, new_n11026);
xnor_3 g10655(new_n11032, new_n11031, new_n11012);
nand_4 g10656(new_n11033, new_n10625, new_n10624);
not_3  g10657(new_n11034, new_n10622);
nand_4 g10658(new_n11035, new_n10627, new_n11034);
nand_4 g10659(new_n11036, new_n11035, new_n11033);
nand_4 g10660(new_n11037, new_n10674, new_n10668);
nand_4 g10661(new_n11038, new_n10692, new_n10676);
nand_4 g10662(new_n11039, new_n11038, new_n11037);
xnor_3 g10663(new_n11040, new_n11039, new_n11036);
xnor_3 g10664(new_n11041, new_n11040, new_n11032);
and_4  g10665(new_n11042, new_n10605, new_n10599);
not_3  g10666(new_n11043, new_n10621);
nor_4  g10667(new_n11044, new_n11043, new_n10606);
nor_4  g10668(new_n11045, new_n11044, new_n11042);
not_3  g10669(new_n11046, new_n10595);
nand_4 g10670(new_n11047, new_n10628, new_n11046);
nand_4 g10671(new_n11048, new_n10637, new_n10629);
nand_4 g10672(new_n11049, new_n11048, new_n11047);
xnor_3 g10673(new_n11050, new_n11049, new_n11045);
xnor_3 g10674(new_n11051, new_n11050, new_n11041);
nand_4 g10675(new_n11052, new_n10818, new_n10815);
not_3  g10676(new_n11053, new_n10819);
not_3  g10677(new_n11054, new_n10846);
nand_4 g10678(new_n11055, new_n11054, new_n11053);
nand_4 g10679(new_n11056, new_n11055, new_n11052);
nor_4  g10680(new_n11057, new_n10609, new_n10607);
nor_4  g10681(new_n11058, new_n10619, new_n11057);
nand_4 g10682(new_n11059, n10898, n5857);
nand_4 g10683(new_n11060, n11257, n3932);
not_3  g10684(new_n11061, new_n11060);
xor_3  g10685(new_n11062, new_n11061, new_n11059);
xor_3  g10686(new_n11063, new_n11062, new_n11058);
nand_4 g10687(new_n11064, n11876, n45);
nand_4 g10688(new_n11065, n3986, n3754);
not_3  g10689(new_n11066, new_n11065);
xor_3  g10690(new_n11067, new_n11066, new_n11064);
nand_4 g10691(new_n11068, n10327, n1097);
nand_4 g10692(new_n11069, n12705, n7456);
xor_3  g10693(new_n11070, new_n11069, new_n11068);
nand_4 g10694(new_n11071, n12591, n12025);
nand_4 g10695(new_n11072, n9583, n5964);
nand_4 g10696(new_n11073, n11662, n4312);
xor_3  g10697(new_n11074, new_n11073, new_n11072);
xor_3  g10698(new_n11075, new_n11074, new_n11071);
xnor_3 g10699(new_n11076, new_n11075, new_n11070);
not_3  g10700(new_n11077, new_n10601);
nor_4  g10701(new_n11078, new_n10603, new_n11077);
not_3  g10702(new_n11079, new_n10600);
nor_4  g10703(new_n11080, new_n10604, new_n11079);
nor_4  g10704(new_n11081, new_n11080, new_n11078);
not_3  g10705(new_n11082, new_n10613);
nor_4  g10706(new_n11083, new_n10615, new_n11082);
not_3  g10707(new_n11084, new_n10612);
nor_4  g10708(new_n11085, new_n10616, new_n11084);
nor_4  g10709(new_n11086, new_n11085, new_n11083);
xnor_3 g10710(new_n11087, new_n11086, new_n11081);
xnor_3 g10711(new_n11088, new_n11087, new_n11076);
xnor_3 g10712(new_n11089, new_n11088, new_n11067);
xnor_3 g10713(new_n11090, new_n11089, new_n11063);
xnor_3 g10714(new_n11091, new_n11090, new_n11056);
xnor_3 g10715(new_n11092, new_n11091, new_n11051);
xnor_3 g10716(new_n11093, new_n11092, new_n10974);
xnor_3 g10717(new_n11094, new_n11093, new_n10925);
xnor_3 g10718(n4230, new_n11094, new_n10901);
not_3  g10719(new_n11096, new_n6285);
xor_3  g10720(n4300, new_n11096, new_n6284);
not_3  g10721(new_n11098, new_n3830);
xor_3  g10722(n4326, new_n11098, new_n3829);
not_3  g10723(new_n11100, new_n1324);
nor_4  g10724(new_n11101, new_n11100, new_n1317);
not_3  g10725(new_n11102, new_n11101);
nand_4 g10726(new_n11103, n6687, n5320);
not_3  g10727(new_n11104, new_n1300);
nand_4 g10728(new_n11105, new_n1309, new_n11104);
not_3  g10729(new_n11106, new_n11105);
nor_4  g10730(new_n11107, new_n1316, new_n1310);
nor_4  g10731(new_n11108, new_n11107, new_n11106);
xnor_3 g10732(new_n11109, new_n11108, new_n11103);
nand_4 g10733(new_n11110, n4370, n2564);
not_3  g10734(new_n11111, new_n11110);
and_4  g10735(new_n11112, new_n1314, new_n1313);
nor_4  g10736(new_n11113, new_n1315, new_n1312);
nor_4  g10737(new_n11114, new_n11113, new_n11112);
nand_4 g10738(new_n11115, new_n11114, new_n11111);
not_3  g10739(new_n11116, new_n11115);
nor_4  g10740(new_n11117, new_n11114, new_n11111);
nor_4  g10741(new_n11118, new_n11117, new_n11116);
nand_4 g10742(new_n11119, n6770, n5212);
nand_4 g10743(new_n11120, n11877, n4189);
nand_4 g10744(new_n11121, n11407, n9920);
xnor_3 g10745(new_n11122, new_n11121, new_n11120);
xor_3  g10746(new_n11123, new_n11122, new_n11119);
nand_4 g10747(new_n11124, new_n11123, new_n11118);
not_3  g10748(new_n11125, new_n11124);
nor_4  g10749(new_n11126, new_n11123, new_n11118);
nor_4  g10750(new_n11127, new_n11126, new_n11125);
not_3  g10751(new_n11128, new_n11127);
xnor_3 g10752(new_n11129, new_n11128, new_n11109);
not_3  g10753(new_n11130, new_n11129);
xor_3  g10754(new_n11131, new_n11130, new_n11102);
not_3  g10755(new_n11132, new_n1444);
nor_4  g10756(new_n11133, new_n11132, new_n1443);
nand_4 g10757(new_n11134, n8336, n2433);
nand_4 g10758(new_n11135, n10928, n8819);
not_3  g10759(new_n11136, new_n11135);
not_3  g10760(new_n11137, new_n1434);
not_3  g10761(new_n11138, new_n1435);
nor_4  g10762(new_n11139, new_n11138, new_n11137);
nor_4  g10763(new_n11140, new_n1435, new_n1434);
nor_4  g10764(new_n11141, new_n11140, new_n1433);
nor_4  g10765(new_n11142, new_n11141, new_n11139);
xnor_3 g10766(new_n11143, new_n11142, new_n11136);
nand_4 g10767(new_n11144, n11728, n2226);
not_3  g10768(new_n11145, new_n11144);
nand_4 g10769(new_n11146, n6986, n6429);
not_3  g10770(new_n11147, new_n11146);
nand_4 g10771(new_n11148, n12709, n1094);
not_3  g10772(new_n11149, new_n11148);
nor_4  g10773(new_n11150, new_n11149, new_n11147);
nor_4  g10774(new_n11151, new_n11148, new_n11146);
nor_4  g10775(new_n11152, new_n11151, new_n11150);
xnor_3 g10776(new_n11153_1, new_n11152, new_n11145);
xnor_3 g10777(new_n11154, new_n11153_1, new_n11143);
nor_4  g10778(new_n11155, new_n11154, new_n11134);
not_3  g10779(new_n11156, new_n11134);
not_3  g10780(new_n11157, new_n11154);
nor_4  g10781(new_n11158, new_n11157, new_n11156);
nor_4  g10782(new_n11159, new_n11158, new_n11155);
nor_4  g10783(new_n11160, new_n1438, new_n1431);
not_3  g10784(new_n11161, new_n11160);
nand_4 g10785(new_n11162, new_n1442, new_n1439);
nand_4 g10786(new_n11163, new_n11162, new_n11161);
xnor_3 g10787(new_n11164, new_n11163, new_n11159);
xnor_3 g10788(new_n11165, new_n11164, new_n11133);
nand_4 g10789(new_n11166, new_n1491, new_n1445);
nand_4 g10790(new_n11167, new_n1496, new_n1499);
nand_4 g10791(new_n11168, new_n11167, new_n11166);
nand_4 g10792(new_n11169, new_n11168, new_n11165);
not_3  g10793(new_n11170, new_n11165);
not_3  g10794(new_n11171, new_n11166);
nor_4  g10795(new_n11172, new_n1498, new_n11171);
nand_4 g10796(new_n11173, new_n11172, new_n11170);
nand_4 g10797(new_n11174, new_n11173, new_n11169);
nand_4 g10798(new_n11175, n12069, n11967);
nand_4 g10799(new_n11176, n12391, n6254);
not_3  g10800(new_n11177, new_n11176);
not_3  g10801(new_n11178, new_n1453);
nor_4  g10802(new_n11179, new_n1459, new_n11178);
nor_4  g10803(new_n11180, new_n11179, new_n1458);
xnor_3 g10804(new_n11181, new_n11180, new_n11177);
nand_4 g10805(new_n11182, n7160, n7159);
not_3  g10806(new_n11183, new_n11182);
nand_4 g10807(new_n11184, n12777, n7891);
not_3  g10808(new_n11185, new_n11184);
nand_4 g10809(new_n11186, n12489, n4828);
not_3  g10810(new_n11187, new_n11186);
nor_4  g10811(new_n11188, new_n11187, new_n11185);
nor_4  g10812(new_n11189, new_n11186, new_n11184);
nor_4  g10813(new_n11190, new_n11189, new_n11188);
xnor_3 g10814(new_n11191, new_n11190, new_n11183);
xnor_3 g10815(new_n11192, new_n11191, new_n11181);
nor_4  g10816(new_n11193, new_n11192, new_n11175);
not_3  g10817(new_n11194, new_n11175);
not_3  g10818(new_n11195, new_n11192);
nor_4  g10819(new_n11196, new_n11195, new_n11194);
nor_4  g10820(new_n11197, new_n11196, new_n11193);
nand_4 g10821(new_n11198, new_n1451, new_n1447);
nor_4  g10822(new_n11199, new_n1462, new_n1452);
not_3  g10823(new_n11200, new_n11199);
nand_4 g10824(new_n11201, new_n11200, new_n11198);
xnor_3 g10825(new_n11202, new_n11201, new_n11197);
not_3  g10826(new_n11203, new_n11202);
nor_4  g10827(new_n11204, new_n11203, new_n1466);
not_3  g10828(new_n11205, new_n1466);
nor_4  g10829(new_n11206, new_n11202, new_n11205);
nor_4  g10830(new_n11207, new_n11206, new_n11204);
not_3  g10831(new_n11208, new_n11207);
nand_4 g10832(new_n11209, n12947, n11222);
nand_4 g10833(new_n11210, n11791, n11153);
not_3  g10834(new_n11211, new_n1475);
not_3  g10835(new_n11212, new_n1476);
nor_4  g10836(new_n11213, new_n11212, new_n11211);
not_3  g10837(new_n11214, new_n1474);
nor_4  g10838(new_n11215, new_n1477, new_n11214);
nor_4  g10839(new_n11216_1, new_n11215, new_n11213);
xnor_3 g10840(new_n11217, new_n11216_1, new_n11210);
nand_4 g10841(new_n11218, n5760, n996);
nand_4 g10842(new_n11219, n5314, n1478);
nand_4 g10843(new_n11220, n10990, n5767);
nand_4 g10844(new_n11221, new_n11220, new_n11219);
not_3  g10845(new_n11222_1, new_n11221);
not_3  g10846(new_n11223, new_n11219);
not_3  g10847(new_n11224, new_n11220);
nand_4 g10848(new_n11225, new_n11224, new_n11223);
not_3  g10849(new_n11226, new_n11225);
nor_4  g10850(new_n11227, new_n11226, new_n11222_1);
xnor_3 g10851(new_n11228, new_n11227, new_n11218);
xnor_3 g10852(new_n11229, new_n11228, new_n11217);
xnor_3 g10853(new_n11230, new_n11229, new_n11209);
nor_4  g10854(new_n11231, new_n1472, new_n1470);
nor_4  g10855(new_n11232, new_n1478_1, new_n1473);
nor_4  g10856(new_n11233, new_n11232, new_n11231);
xnor_3 g10857(new_n11234, new_n11233, new_n11230);
not_3  g10858(new_n11235, new_n11234);
xor_3  g10859(new_n11236, new_n11235, new_n1482);
nor_4  g10860(new_n11237, new_n1485, new_n1469);
nor_4  g10861(new_n11238, new_n1490, new_n1486);
nor_4  g10862(new_n11239, new_n11238, new_n11237);
nand_4 g10863(new_n11240, new_n11239, new_n11236);
not_3  g10864(new_n11241, new_n1482);
xor_3  g10865(new_n11242, new_n11235, new_n11241);
not_3  g10866(new_n11243, new_n11239);
nand_4 g10867(new_n11244, new_n11243, new_n11242);
nand_4 g10868(new_n11245, new_n11244, new_n11240);
xnor_3 g10869(new_n11246, new_n11245, new_n11208);
xnor_3 g10870(new_n11247, new_n11246, new_n11174);
nor_4  g10871(new_n11248, new_n11247, new_n11131);
nand_4 g10872(new_n11249, new_n11247, new_n11131);
not_3  g10873(new_n11250, new_n11249);
nor_4  g10874(new_n11251, new_n11250, new_n11248);
not_3  g10875(new_n11252, new_n1427);
nand_4 g10876(new_n11253, new_n1501, new_n1430);
nand_4 g10877(new_n11254, new_n11253, new_n11252);
xor_3  g10878(n4333, new_n11254, new_n11251);
nand_4 g10879(new_n11256, n11877, n11757);
not_3  g10880(new_n11257_1, new_n11256);
nand_4 g10881(new_n11258, n5240, n5212);
nand_4 g10882(new_n11259, n11821, n11407);
xnor_3 g10883(new_n11260, new_n11259, new_n11258);
not_3  g10884(new_n11261, new_n11260);
nor_4  g10885(new_n11262, new_n11261, new_n11257_1);
nor_4  g10886(new_n11263, new_n11260, new_n11256);
nor_4  g10887(new_n11264, new_n11263, new_n11262);
not_3  g10888(new_n11265, new_n11264);
nand_4 g10889(new_n11266, n11407, n5240);
nand_4 g10890(new_n11267, n11877, n3172);
nand_4 g10891(new_n11268, new_n11267, new_n11266);
not_3  g10892(new_n11269, new_n11268);
nand_4 g10893(new_n11270, n11757, n5212);
not_3  g10894(new_n11271, new_n11270);
xnor_3 g10895(new_n11272, new_n11267, new_n11266);
nor_4  g10896(new_n11273, new_n11272, new_n11271);
nor_4  g10897(new_n11274, new_n11273, new_n11269);
nor_4  g10898(new_n11275, new_n11274, new_n11265);
not_3  g10899(new_n11276, new_n11274);
nor_4  g10900(new_n11277, new_n11276, new_n11264);
nor_4  g10901(new_n11278, new_n11277, new_n11275);
nand_4 g10902(new_n11279, n5320, n1333);
nand_4 g10903(new_n11280, n4370, n3172);
xor_3  g10904(new_n11281, new_n11280, new_n11279);
xnor_3 g10905(new_n11282, new_n11281, new_n11278);
nand_4 g10906(new_n11283, n4370, n1333);
not_3  g10907(new_n11284, new_n11283);
nand_4 g10908(new_n11285, n11877, n1333);
not_3  g10909(new_n11286, new_n11285);
nand_4 g10910(new_n11287, n11757, n11407);
not_3  g10911(new_n11288, new_n11287);
nor_4  g10912(new_n11289, new_n11288, new_n11286);
nand_4 g10913(new_n11290, n5212, n3172);
not_3  g10914(new_n11291, new_n11290);
xnor_3 g10915(new_n11292, new_n11287, new_n11285);
nor_4  g10916(new_n11293, new_n11292, new_n11291);
nor_4  g10917(new_n11294, new_n11293, new_n11289);
nand_4 g10918(new_n11295, new_n11294, new_n11284);
not_3  g10919(new_n11296_1, new_n11295);
nor_4  g10920(new_n11297, new_n11294, new_n11284);
nor_4  g10921(new_n11298, new_n11297, new_n11296_1);
xor_3  g10922(new_n11299, new_n11272, new_n11270);
nand_4 g10923(new_n11300, new_n11299, new_n11298);
nand_4 g10924(new_n11301, new_n11300, new_n11295);
nand_4 g10925(new_n11302, new_n11301, new_n11282);
not_3  g10926(new_n11303, new_n11302);
nor_4  g10927(new_n11304, new_n11301, new_n11282);
nor_4  g10928(new_n11305, new_n11304, new_n11303);
not_3  g10929(new_n11306, new_n11305);
nand_4 g10930(new_n11307, n7862, n5320);
xnor_3 g10931(new_n11308, new_n11299, new_n11298);
nand_4 g10932(new_n11309, new_n11308, new_n11307);
xnor_3 g10933(new_n11310, new_n11308, new_n11307);
not_3  g10934(new_n11311_1, new_n11310);
nand_4 g10935(new_n11312, n7862, n4370);
not_3  g10936(new_n11313, new_n11312);
nand_4 g10937(new_n11314, n11407, n3172);
not_3  g10938(new_n11315, new_n11314);
nand_4 g10939(new_n11316, n11877, n7862);
not_3  g10940(new_n11317, new_n11316);
nor_4  g10941(new_n11318, new_n11317, new_n11315);
nand_4 g10942(new_n11319, n11407, n7862);
nor_4  g10943(new_n11320, new_n11319, new_n11267);
nand_4 g10944(new_n11321, n5212, n1333);
not_3  g10945(new_n11322, new_n11321);
nor_4  g10946(new_n11323, new_n11322, new_n11320);
nor_4  g10947(new_n11324, new_n11323, new_n11318);
and_4  g10948(new_n11325, new_n11324, new_n11313);
not_3  g10949(new_n11326_1, new_n11325);
xor_3  g10950(new_n11327, new_n11324, new_n11312);
xor_3  g10951(new_n11328, new_n11292, new_n11291);
nor_4  g10952(new_n11329, new_n11328, new_n11327);
not_3  g10953(new_n11330, new_n11329);
nand_4 g10954(new_n11331, new_n11330, new_n11326_1);
not_3  g10955(new_n11332, new_n11331);
nand_4 g10956(new_n11333, new_n11332, new_n11311_1);
nand_4 g10957(new_n11334, new_n11333, new_n11309);
nor_4  g10958(new_n11335, new_n11334, new_n11306);
not_3  g10959(new_n11336, new_n11335);
not_3  g10960(new_n11337, new_n11278);
nand_4 g10961(new_n11338, new_n11281, new_n11337);
nor_4  g10962(new_n11339, new_n11280, new_n11279);
xnor_3 g10963(new_n11340, new_n11303, new_n11339);
nand_4 g10964(new_n11341, new_n11340, new_n11338);
nor_4  g10965(new_n11342, new_n11259, new_n11258);
nand_4 g10966(new_n11343, n11757, n4370);
not_3  g10967(new_n11344, new_n11343);
xor_3  g10968(new_n11345, new_n11344, new_n11342);
nand_4 g10969(new_n11346, n11821, n5212);
not_3  g10970(new_n11347, new_n11346);
nand_4 g10971(new_n11348, n11877, n5240);
nand_4 g10972(new_n11349, n11407, n9080);
not_3  g10973(new_n11350, new_n11349);
xor_3  g10974(new_n11351, new_n11350, new_n11348);
xnor_3 g10975(new_n11352, new_n11351, new_n11347);
xnor_3 g10976(new_n11353, new_n11352, new_n11345);
nor_4  g10977(new_n11354, new_n11275, new_n11262);
nand_4 g10978(new_n11355, n12000, n1333);
nand_4 g10979(new_n11356, n5320, n3172);
nand_4 g10980(new_n11357, n9725, n7862);
not_3  g10981(new_n11358, new_n11357);
xor_3  g10982(new_n11359, new_n11358, new_n11356);
xnor_3 g10983(new_n11360, new_n11359, new_n11355);
xnor_3 g10984(new_n11361, new_n11360, new_n11354);
xnor_3 g10985(new_n11362, new_n11361, new_n11353);
xor_3  g10986(new_n11363, new_n11362, new_n11341);
xnor_3 g10987(new_n11364, new_n11363, new_n11336);
nand_4 g10988(new_n11365, n12000, n7862);
not_3  g10989(new_n11366, new_n11365);
not_3  g10990(new_n11367, new_n11334);
nor_4  g10991(new_n11368, new_n11367, new_n11305);
nor_4  g10992(new_n11369, new_n11368, new_n11335);
nor_4  g10993(new_n11370, new_n11369, new_n11366);
nor_4  g10994(new_n11371, new_n11320, new_n11318);
nand_4 g10995(new_n11372, n11407, n1333);
nand_4 g10996(new_n11373, n7862, n5212);
nor_4  g10997(new_n11374, new_n11373, new_n11372);
not_3  g10998(new_n11375, new_n11374);
nor_4  g10999(new_n11376, new_n11375, new_n11371);
not_3  g11000(new_n11377, new_n11376);
xnor_3 g11001(new_n11378, new_n11328, new_n11327);
nor_4  g11002(new_n11379, new_n11378, new_n11377);
xor_3  g11003(new_n11380, new_n11331, new_n11311_1);
nand_4 g11004(new_n11381, new_n11380, new_n11379);
not_3  g11005(new_n11382, new_n11381);
xnor_3 g11006(new_n11383, new_n11369, new_n11366);
nor_4  g11007(new_n11384, new_n11383, new_n11382);
nor_4  g11008(new_n11385, new_n11384, new_n11370);
xnor_3 g11009(new_n11386, new_n11385, new_n11364);
nand_4 g11010(new_n11387, n11311, n6429);
nand_4 g11011(new_n11388, n12709, n4203);
nand_4 g11012(new_n11389, n11728, n4187);
xnor_3 g11013(new_n11390, new_n11389, new_n11388);
nor_4  g11014(new_n11391, new_n11390, new_n11387);
not_3  g11015(new_n11392, new_n11387);
not_3  g11016(new_n11393, new_n11390);
nor_4  g11017(new_n11394, new_n11393, new_n11392);
nor_4  g11018(new_n11395, new_n11394, new_n11391);
nand_4 g11019(new_n11396, n12709, n4187);
nand_4 g11020(new_n11397, n6429, n2464);
and_4  g11021(new_n11398, new_n11397, new_n11396);
nand_4 g11022(new_n11399, n11728, n11311);
not_3  g11023(new_n11400, new_n11399);
xnor_3 g11024(new_n11401, new_n11397, new_n11396);
nor_4  g11025(new_n11402, new_n11401, new_n11400);
nor_4  g11026(new_n11403, new_n11402, new_n11398);
xnor_3 g11027(new_n11404, new_n11403, new_n11395);
nand_4 g11028(new_n11405, n9400, n2433);
nand_4 g11029(new_n11406, n8819, n2464);
xor_3  g11030(new_n11407_1, new_n11406, new_n11405);
not_3  g11031(new_n11408, new_n11407_1);
nor_4  g11032(new_n11409, new_n11408, new_n11404);
not_3  g11033(new_n11410, new_n11404);
nor_4  g11034(new_n11411, new_n11407_1, new_n11410);
nor_4  g11035(new_n11412, new_n11411, new_n11409);
nand_4 g11036(new_n11413, n9400, n8819);
not_3  g11037(new_n11414, new_n11413);
nand_4 g11038(new_n11415, n12709, n11311);
not_3  g11039(new_n11416, new_n11415);
nand_4 g11040(new_n11417, n9400, n6429);
not_3  g11041(new_n11418, new_n11417);
nor_4  g11042(new_n11419, new_n11418, new_n11416);
nand_4 g11043(new_n11420, n11728, n2464);
not_3  g11044(new_n11421, new_n11420);
xnor_3 g11045(new_n11422, new_n11417, new_n11415);
nor_4  g11046(new_n11423_1, new_n11422, new_n11421);
nor_4  g11047(new_n11424, new_n11423_1, new_n11419);
nand_4 g11048(new_n11425, new_n11424, new_n11414);
not_3  g11049(new_n11426, new_n11425);
xnor_3 g11050(new_n11427, new_n11424, new_n11414);
xnor_3 g11051(new_n11428, new_n11401, new_n11399);
nor_4  g11052(new_n11429, new_n11428, new_n11427);
nor_4  g11053(new_n11430, new_n11429, new_n11426);
not_3  g11054(new_n11431, new_n11430);
xnor_3 g11055(new_n11432, new_n11431, new_n11412);
nand_4 g11056(new_n11433, n6877, n2433);
xnor_3 g11057(new_n11434, new_n11428, new_n11427);
nor_4  g11058(new_n11435, new_n11434, new_n11433);
not_3  g11059(new_n11436, new_n11435);
not_3  g11060(new_n11437, new_n11433);
not_3  g11061(new_n11438, new_n11434);
nor_4  g11062(new_n11439, new_n11438, new_n11437);
nor_4  g11063(new_n11440, new_n11439, new_n11435);
nand_4 g11064(new_n11441, n8819, n6877);
not_3  g11065(new_n11442, new_n11441);
nand_4 g11066(new_n11443, n12709, n2464);
not_3  g11067(new_n11444, new_n11443);
nand_4 g11068(new_n11445, n6877, n6429);
not_3  g11069(new_n11446, new_n11445);
nor_4  g11070(new_n11447, new_n11446, new_n11444);
nor_4  g11071(new_n11448, new_n11445, new_n11443);
nand_4 g11072(new_n11449, n11728, n9400);
not_3  g11073(new_n11450, new_n11449);
nor_4  g11074(new_n11451, new_n11450, new_n11448);
nor_4  g11075(new_n11452, new_n11451, new_n11447);
nand_4 g11076(new_n11453, new_n11452, new_n11442);
not_3  g11077(new_n11454, new_n11453);
xnor_3 g11078(new_n11455, new_n11452, new_n11442);
and_4  g11079(new_n11456, new_n11422, new_n11421);
nor_4  g11080(new_n11457, new_n11456, new_n11423_1);
nor_4  g11081(new_n11458, new_n11457, new_n11455);
nor_4  g11082(new_n11459, new_n11458, new_n11454);
not_3  g11083(new_n11460, new_n11459);
nand_4 g11084(new_n11461, new_n11460, new_n11440);
nand_4 g11085(new_n11462, new_n11461, new_n11436);
not_3  g11086(new_n11463, new_n11462);
nor_4  g11087(new_n11464, new_n11463, new_n11432);
not_3  g11088(new_n11465, new_n11409);
nor_4  g11089(new_n11466, new_n11406, new_n11405);
nand_4 g11090(new_n11467, new_n11431, new_n11412);
not_3  g11091(new_n11468, new_n11467);
xnor_3 g11092(new_n11469, new_n11468, new_n11466);
nand_4 g11093(new_n11470, new_n11469, new_n11465);
not_3  g11094(new_n11471, new_n11391);
nand_4 g11095(new_n11472, new_n11403, new_n11395);
nand_4 g11096(new_n11473, new_n11472, new_n11471);
nand_4 g11097(new_n11474, n9400, n8717);
not_3  g11098(new_n11475, new_n11474);
nand_4 g11099(new_n11476, n2464, n2433);
nand_4 g11100(new_n11477, n7730, n6877);
not_3  g11101(new_n11478_1, new_n11477);
xor_3  g11102(new_n11479, new_n11478_1, new_n11476);
xnor_3 g11103(new_n11480, new_n11479, new_n11475);
xnor_3 g11104(new_n11481, new_n11480, new_n11473);
nor_4  g11105(new_n11482, new_n11389, new_n11388);
not_3  g11106(new_n11483, new_n11482);
nand_4 g11107(new_n11484, n11311, n8819);
xor_3  g11108(new_n11485, new_n11484, new_n11483);
nand_4 g11109(new_n11486, n11728, n4203);
nand_4 g11110(new_n11487, n6429, n4187);
nand_4 g11111(new_n11488, n12753, n12709);
not_3  g11112(new_n11489, new_n11488);
xor_3  g11113(new_n11490, new_n11489, new_n11487);
xnor_3 g11114(new_n11491, new_n11490, new_n11486);
xnor_3 g11115(new_n11492, new_n11491, new_n11485);
xnor_3 g11116(new_n11493, new_n11492, new_n11481);
xnor_3 g11117(new_n11494, new_n11493, new_n11470);
xnor_3 g11118(new_n11495, new_n11494, new_n11464);
not_3  g11119(new_n11496, new_n11495);
nand_4 g11120(new_n11497, n8717, n6877);
not_3  g11121(new_n11498, new_n11497);
not_3  g11122(new_n11499, new_n11432);
nor_4  g11123(new_n11500, new_n11462, new_n11499);
nor_4  g11124(new_n11501, new_n11500, new_n11464);
nand_4 g11125(new_n11502, new_n11501, new_n11498);
nor_4  g11126(new_n11503, new_n11448, new_n11447);
nand_4 g11127(new_n11504, n12709, n9400);
nand_4 g11128(new_n11505, n11728, n6877);
nor_4  g11129(new_n11506, new_n11505, new_n11504);
not_3  g11130(new_n11507, new_n11506);
nor_4  g11131(new_n11508, new_n11507, new_n11503);
not_3  g11132(new_n11509, new_n11508);
xnor_3 g11133(new_n11510, new_n11457, new_n11455);
nor_4  g11134(new_n11511, new_n11510, new_n11509);
not_3  g11135(new_n11512, new_n11511);
xnor_3 g11136(new_n11513, new_n11460, new_n11440);
nor_4  g11137(new_n11514, new_n11513, new_n11512);
xnor_3 g11138(new_n11515, new_n11501, new_n11497);
nand_4 g11139(new_n11516, new_n11515, new_n11514);
nand_4 g11140(new_n11517, new_n11516, new_n11502);
xnor_3 g11141(new_n11518, new_n11517, new_n11496);
nand_4 g11142(new_n11519, n11478, n6254);
not_3  g11143(new_n11520, new_n11519);
nand_4 g11144(new_n11521, n12489, n137);
not_3  g11145(new_n11522, new_n11521);
nand_4 g11146(new_n11523, n12777, n11478);
not_3  g11147(new_n11524, new_n11523);
nor_4  g11148(new_n11525, new_n11524, new_n11522);
nand_4 g11149(new_n11526, n7159, n5283);
not_3  g11150(new_n11527, new_n11526);
xnor_3 g11151(new_n11528, new_n11523, new_n11521);
nor_4  g11152(new_n11529, new_n11528, new_n11527);
nor_4  g11153(new_n11530, new_n11529, new_n11525);
nand_4 g11154(new_n11531, new_n11530, new_n11520);
nand_4 g11155(new_n11532, n7159, n137);
not_3  g11156(new_n11533, new_n11532);
nand_4 g11157(new_n11534, n12489, n6294);
nand_4 g11158(new_n11535, n12777, n5283);
xnor_3 g11159(new_n11536_1, new_n11535, new_n11534);
xnor_3 g11160(new_n11537, new_n11536_1, new_n11533);
xnor_3 g11161(new_n11538, new_n11530, new_n11519);
nand_4 g11162(new_n11539, new_n11538, new_n11537);
nand_4 g11163(new_n11540, new_n11539, new_n11531);
nand_4 g11164(new_n11541, n11967, n11478);
nand_4 g11165(new_n11542, n6254, n5283);
nor_4  g11166(new_n11543, new_n11542, new_n11541);
and_4  g11167(new_n11544, new_n11542, new_n11541);
nor_4  g11168(new_n11545, new_n11544, new_n11543);
not_3  g11169(new_n11546, new_n11545);
xnor_3 g11170(new_n11547, new_n11546, new_n11540);
nand_4 g11171(new_n11548, n12777, n137);
nand_4 g11172(new_n11549, n7159, n6294);
nand_4 g11173(new_n11550, n12489, n6797);
xnor_3 g11174(new_n11551, new_n11550, new_n11549);
nor_4  g11175(new_n11552, new_n11551, new_n11548);
not_3  g11176(new_n11553, new_n11548);
not_3  g11177(new_n11554, new_n11551);
nor_4  g11178(new_n11555, new_n11554, new_n11553);
nor_4  g11179(new_n11556, new_n11555, new_n11552);
and_4  g11180(new_n11557, new_n11535, new_n11534);
nor_4  g11181(new_n11558, new_n11536_1, new_n11533);
nor_4  g11182(new_n11559, new_n11558, new_n11557);
nand_4 g11183(new_n11560, new_n11559, new_n11556);
not_3  g11184(new_n11561, new_n11560);
nor_4  g11185(new_n11562, new_n11559, new_n11556);
nor_4  g11186(new_n11563, new_n11562, new_n11561);
nand_4 g11187(new_n11564, new_n11563, new_n11547);
xnor_3 g11188(new_n11565, new_n11545, new_n11540);
xnor_3 g11189(new_n11566, new_n11559, new_n11556);
nand_4 g11190(new_n11567, new_n11566, new_n11565);
nand_4 g11191(new_n11568, new_n11567, new_n11564);
nand_4 g11192(new_n11569, n11967, n4805);
not_3  g11193(new_n11570, new_n11569);
nand_4 g11194(new_n11571, n6254, n4805);
not_3  g11195(new_n11572, new_n11571);
nand_4 g11196(new_n11573, n12489, n5283);
not_3  g11197(new_n11574, new_n11573);
nand_4 g11198(new_n11575, n12777, n4805);
not_3  g11199(new_n11576, new_n11575);
nor_4  g11200(new_n11577, new_n11576, new_n11574);
nor_4  g11201(new_n11578, new_n11575, new_n11573);
nand_4 g11202(new_n11579, n11478, n7159);
not_3  g11203(new_n11580, new_n11579);
nor_4  g11204(new_n11581, new_n11580, new_n11578);
nor_4  g11205(new_n11582, new_n11581, new_n11577);
nand_4 g11206(new_n11583, new_n11582, new_n11572);
not_3  g11207(new_n11584, new_n11583);
nor_4  g11208(new_n11585, new_n11582, new_n11572);
nor_4  g11209(new_n11586, new_n11585, new_n11584);
xnor_3 g11210(new_n11587, new_n11528, new_n11526);
not_3  g11211(new_n11588, new_n11587);
nand_4 g11212(new_n11589, new_n11588, new_n11586);
nand_4 g11213(new_n11590, new_n11589, new_n11583);
nor_4  g11214(new_n11591, new_n11590, new_n11570);
not_3  g11215(new_n11592, new_n11591);
not_3  g11216(new_n11593, new_n11539);
nor_4  g11217(new_n11594, new_n11538, new_n11537);
nor_4  g11218(new_n11595, new_n11594, new_n11593);
not_3  g11219(new_n11596, new_n11595);
xnor_3 g11220(new_n11597, new_n11590, new_n11569);
nand_4 g11221(new_n11598, new_n11597, new_n11596);
nand_4 g11222(new_n11599, new_n11598, new_n11592);
nor_4  g11223(new_n11600, new_n11599, new_n11568);
not_3  g11224(new_n11601, new_n11552);
nand_4 g11225(new_n11602, new_n11560, new_n11601);
nand_4 g11226(new_n11603, n11478, n447);
nand_4 g11227(new_n11604, n11967, n5283);
nand_4 g11228(new_n11605, n4805, n1353);
nand_4 g11229(new_n11606, new_n11605, new_n11604);
not_3  g11230(new_n11607, new_n11604);
not_3  g11231(new_n11608, new_n11605);
nand_4 g11232(new_n11609, new_n11608, new_n11607);
nand_4 g11233(new_n11610, new_n11609, new_n11606);
xnor_3 g11234(new_n11611, new_n11610, new_n11603);
xnor_3 g11235(new_n11612, new_n11611, new_n11602);
nor_4  g11236(new_n11613, new_n11550, new_n11549);
not_3  g11237(new_n11614, new_n11613);
nand_4 g11238(new_n11615, n6254, n137);
xor_3  g11239(new_n11616, new_n11615, new_n11614);
nand_4 g11240(new_n11617, n7159, n6797);
nand_4 g11241(new_n11618, n12777, n6294);
nand_4 g11242(new_n11619, n12489, n3146);
xnor_3 g11243(new_n11620, new_n11619, new_n11618);
xnor_3 g11244(new_n11621, new_n11620, new_n11617);
xnor_3 g11245(new_n11622, new_n11621, new_n11616);
xnor_3 g11246(new_n11623, new_n11622, new_n11612);
not_3  g11247(new_n11624, new_n11540);
nor_4  g11248(new_n11625, new_n11546, new_n11624);
not_3  g11249(new_n11626, new_n11625);
not_3  g11250(new_n11627, new_n11543);
xnor_3 g11251(new_n11628, new_n11564, new_n11627);
nand_4 g11252(new_n11629, new_n11628, new_n11626);
xnor_3 g11253(new_n11630, new_n11629, new_n11623);
xnor_3 g11254(new_n11631, new_n11630, new_n11600);
nand_4 g11255(new_n11632, n4805, n447);
not_3  g11256(new_n11633, new_n11632);
xnor_3 g11257(new_n11634, new_n11590, new_n11570);
nor_4  g11258(new_n11635, new_n11634, new_n11595);
nor_4  g11259(new_n11636, new_n11635, new_n11591);
xnor_3 g11260(new_n11637, new_n11636, new_n11568);
nand_4 g11261(new_n11638, new_n11637, new_n11633);
nor_4  g11262(new_n11639, new_n11578, new_n11577);
nand_4 g11263(new_n11640, n12489, n11478);
nand_4 g11264(new_n11641, n7159, n4805);
nor_4  g11265(new_n11642, new_n11641, new_n11640);
not_3  g11266(new_n11643, new_n11642);
nor_4  g11267(new_n11644, new_n11643, new_n11639);
not_3  g11268(new_n11645, new_n11644);
xnor_3 g11269(new_n11646, new_n11588, new_n11586);
nor_4  g11270(new_n11647, new_n11646, new_n11645);
xnor_3 g11271(new_n11648, new_n11634, new_n11595);
nand_4 g11272(new_n11649, new_n11648, new_n11647);
not_3  g11273(new_n11650, new_n11649);
xnor_3 g11274(new_n11651, new_n11637, new_n11632);
nand_4 g11275(new_n11652, new_n11651, new_n11650);
nand_4 g11276(new_n11653, new_n11652, new_n11638);
xnor_3 g11277(new_n11654, new_n11653, new_n11631);
nand_4 g11278(new_n11655, n11791, n3992);
not_3  g11279(new_n11656, new_n11655);
nand_4 g11280(new_n11657, n10990, n6358);
not_3  g11281(new_n11658, new_n11657);
nand_4 g11282(new_n11659, n3992, n1478);
not_3  g11283(new_n11660, new_n11659);
nor_4  g11284(new_n11661, new_n11660, new_n11658);
nand_4 g11285(new_n11662_1, n8384, n5760);
not_3  g11286(new_n11663, new_n11662_1);
xnor_3 g11287(new_n11664, new_n11659, new_n11657);
nor_4  g11288(new_n11665, new_n11664, new_n11663);
nor_4  g11289(new_n11666, new_n11665, new_n11661);
nand_4 g11290(new_n11667, new_n11666, new_n11656);
nand_4 g11291(new_n11668, n6358, n5760);
not_3  g11292(new_n11669, new_n11668);
nand_4 g11293(new_n11670, n10990, n5198);
nand_4 g11294(new_n11671, n8384, n1478);
xnor_3 g11295(new_n11672, new_n11671, new_n11670);
xnor_3 g11296(new_n11673, new_n11672, new_n11669);
xnor_3 g11297(new_n11674, new_n11666, new_n11655);
nand_4 g11298(new_n11675, new_n11674, new_n11673);
nand_4 g11299(new_n11676, new_n11675, new_n11667);
nand_4 g11300(new_n11677, n12947, n3992);
not_3  g11301(new_n11678, new_n11677);
nand_4 g11302(new_n11679, n11791, n8384);
not_3  g11303(new_n11680, new_n11679);
nor_4  g11304(new_n11681, new_n11680, new_n11678);
nor_4  g11305(new_n11682, new_n11679, new_n11677);
nor_4  g11306(new_n11683, new_n11682, new_n11681);
not_3  g11307(new_n11684, new_n11683);
xnor_3 g11308(new_n11685, new_n11684, new_n11676);
nand_4 g11309(new_n11686, n6358, n1478);
nand_4 g11310(new_n11687, n5760, n5198);
nand_4 g11311(new_n11688, n10990, n1471);
xnor_3 g11312(new_n11689, new_n11688, new_n11687);
nor_4  g11313(new_n11690, new_n11689, new_n11686);
not_3  g11314(new_n11691, new_n11686);
not_3  g11315(new_n11692, new_n11689);
nor_4  g11316(new_n11693, new_n11692, new_n11691);
nor_4  g11317(new_n11694, new_n11693, new_n11690);
not_3  g11318(new_n11695, new_n11694);
and_4  g11319(new_n11696, new_n11671, new_n11670);
nor_4  g11320(new_n11697, new_n11672, new_n11669);
nor_4  g11321(new_n11698, new_n11697, new_n11696);
xnor_3 g11322(new_n11699, new_n11698, new_n11695);
nand_4 g11323(new_n11700, new_n11699, new_n11685);
xnor_3 g11324(new_n11701, new_n11683, new_n11676);
xnor_3 g11325(new_n11702, new_n11698, new_n11694);
nand_4 g11326(new_n11703, new_n11702, new_n11701);
nand_4 g11327(new_n11704, new_n11703, new_n11700);
nand_4 g11328(new_n11705, n12947, n7236);
not_3  g11329(new_n11706, new_n11705);
nand_4 g11330(new_n11707_1, n11791, n7236);
not_3  g11331(new_n11708, new_n11707_1);
nand_4 g11332(new_n11709, n10990, n8384);
nand_4 g11333(new_n11710, n7236, n1478);
nand_4 g11334(new_n11711, new_n11710, new_n11709);
not_3  g11335(new_n11712, new_n11711);
nor_4  g11336(new_n11713, new_n11710, new_n11709);
nand_4 g11337(new_n11714, n5760, n3992);
not_3  g11338(new_n11715, new_n11714);
nor_4  g11339(new_n11716, new_n11715, new_n11713);
nor_4  g11340(new_n11717, new_n11716, new_n11712);
nand_4 g11341(new_n11718, new_n11717, new_n11708);
not_3  g11342(new_n11719, new_n11718);
nor_4  g11343(new_n11720, new_n11717, new_n11708);
nor_4  g11344(new_n11721, new_n11720, new_n11719);
xnor_3 g11345(new_n11722, new_n11664, new_n11662_1);
not_3  g11346(new_n11723, new_n11722);
nand_4 g11347(new_n11724, new_n11723, new_n11721);
nand_4 g11348(new_n11725, new_n11724, new_n11718);
nor_4  g11349(new_n11726, new_n11725, new_n11706);
not_3  g11350(new_n11727, new_n11726);
not_3  g11351(new_n11728_1, new_n11675);
nor_4  g11352(new_n11729, new_n11674, new_n11673);
nor_4  g11353(new_n11730, new_n11729, new_n11728_1);
not_3  g11354(new_n11731, new_n11730);
xnor_3 g11355(new_n11732, new_n11725, new_n11705);
nand_4 g11356(new_n11733, new_n11732, new_n11731);
nand_4 g11357(new_n11734, new_n11733, new_n11727);
nor_4  g11358(new_n11735, new_n11734, new_n11704);
not_3  g11359(new_n11736, new_n11690);
nand_4 g11360(new_n11737, new_n11698, new_n11694);
nand_4 g11361(new_n11738, new_n11737, new_n11736);
nand_4 g11362(new_n11739, n6441, n3992);
not_3  g11363(new_n11740, new_n11739);
nand_4 g11364(new_n11741, n12947, n8384);
nand_4 g11365(new_n11742, n11999, n7236);
xnor_3 g11366(new_n11743, new_n11742, new_n11741);
and_4  g11367(new_n11744, new_n11743, new_n11740);
nor_4  g11368(new_n11745, new_n11743, new_n11740);
nor_4  g11369(new_n11746, new_n11745, new_n11744);
xnor_3 g11370(new_n11747, new_n11746, new_n11738);
nor_4  g11371(new_n11748, new_n11688, new_n11687);
nand_4 g11372(new_n11749, n11791, n6358);
not_3  g11373(new_n11750, new_n11749);
xor_3  g11374(new_n11751, new_n11750, new_n11748);
nand_4 g11375(new_n11752, n5760, n1471);
not_3  g11376(new_n11753, new_n11752);
nand_4 g11377(new_n11754, n5198, n1478);
nand_4 g11378(new_n11755_1, n10990, n7646);
xnor_3 g11379(new_n11756, new_n11755_1, new_n11754);
and_4  g11380(new_n11757_1, new_n11756, new_n11753);
nor_4  g11381(new_n11758, new_n11756, new_n11753);
nor_4  g11382(new_n11759, new_n11758, new_n11757_1);
xnor_3 g11383(new_n11760, new_n11759, new_n11751);
xnor_3 g11384(new_n11761, new_n11760, new_n11747);
not_3  g11385(new_n11762, new_n11676);
nor_4  g11386(new_n11763, new_n11684, new_n11762);
not_3  g11387(new_n11764, new_n11763);
not_3  g11388(new_n11765, new_n11682);
xnor_3 g11389(new_n11766, new_n11700, new_n11765);
nand_4 g11390(new_n11767, new_n11766, new_n11764);
xnor_3 g11391(new_n11768, new_n11767, new_n11761);
xnor_3 g11392(new_n11769, new_n11768, new_n11735);
nand_4 g11393(new_n11770, n7236, n6441);
not_3  g11394(new_n11771, new_n11770);
xnor_3 g11395(new_n11772, new_n11725, new_n11706);
nor_4  g11396(new_n11773, new_n11772, new_n11730);
nor_4  g11397(new_n11774, new_n11773, new_n11726);
xnor_3 g11398(new_n11775, new_n11774, new_n11704);
nand_4 g11399(new_n11776, new_n11775, new_n11771);
xnor_3 g11400(new_n11777, new_n11723, new_n11721);
nand_4 g11401(new_n11778, n10990, n7236);
not_3  g11402(new_n11779, new_n11778);
nor_4  g11403(new_n11780_1, new_n11779, new_n11714);
nor_4  g11404(new_n11781, new_n11780_1, new_n11711);
nor_4  g11405(new_n11782, new_n11781, new_n11713);
nor_4  g11406(new_n11783, new_n11782, new_n11714);
not_3  g11407(new_n11784, new_n11783);
nor_4  g11408(new_n11785, new_n11784, new_n11777);
xnor_3 g11409(new_n11786, new_n11772, new_n11730);
nand_4 g11410(new_n11787, new_n11786, new_n11785);
not_3  g11411(new_n11788, new_n11787);
xnor_3 g11412(new_n11789, new_n11775, new_n11770);
nand_4 g11413(new_n11790, new_n11789, new_n11788);
nand_4 g11414(new_n11791_1, new_n11790, new_n11776);
xnor_3 g11415(new_n11792, new_n11791_1, new_n11769);
nand_4 g11416(new_n11793, new_n11792, new_n11654);
not_3  g11417(new_n11794, new_n11600);
xnor_3 g11418(new_n11795, new_n11630, new_n11794);
xnor_3 g11419(new_n11796, new_n11653, new_n11795);
not_3  g11420(new_n11797, new_n11735);
xnor_3 g11421(new_n11798, new_n11768, new_n11797);
xnor_3 g11422(new_n11799, new_n11791_1, new_n11798);
nand_4 g11423(new_n11800, new_n11799, new_n11796);
nand_4 g11424(new_n11801, new_n11800, new_n11793);
xnor_3 g11425(new_n11802, new_n11599, new_n11568);
nand_4 g11426(new_n11803, new_n11802, new_n11632);
nand_4 g11427(new_n11804, new_n11803, new_n11638);
xnor_3 g11428(new_n11805, new_n11804, new_n11650);
not_3  g11429(new_n11806, new_n11805);
xnor_3 g11430(new_n11807, new_n11648, new_n11647);
xnor_3 g11431(new_n11808, new_n11786, new_n11785);
nor_4  g11432(new_n11809, new_n11808, new_n11807);
xnor_3 g11433(new_n11810, new_n11808, new_n11807);
xnor_3 g11434(new_n11811, new_n11646, new_n11644);
xnor_3 g11435(new_n11812, new_n11783, new_n11777);
nor_4  g11436(new_n11813, new_n11812, new_n11811);
not_3  g11437(new_n11814, new_n11813);
nand_4 g11438(new_n11815, n12489, n4805);
not_3  g11439(new_n11816, new_n11815);
nand_4 g11440(new_n11817, new_n11816, new_n11779);
xnor_3 g11441(new_n11818, new_n11641, new_n11640);
nand_4 g11442(new_n11819, new_n11818, new_n11817);
not_3  g11443(new_n11820, new_n11819);
xnor_3 g11444(new_n11821_1, new_n11818, new_n11817);
nand_4 g11445(new_n11822, n10990, n3992);
nand_4 g11446(new_n11823, n7236, n5760);
not_3  g11447(new_n11824, new_n11823);
xnor_3 g11448(new_n11825, new_n11824, new_n11822);
nor_4  g11449(new_n11826, new_n11825, new_n11821_1);
nor_4  g11450(new_n11827, new_n11826, new_n11820);
nand_4 g11451(new_n11828, new_n11780_1, new_n11711);
nand_4 g11452(new_n11829, new_n11828, new_n11782);
not_3  g11453(new_n11830, new_n11829);
nor_4  g11454(new_n11831, new_n11830, new_n11827);
not_3  g11455(new_n11832, new_n11831);
xnor_3 g11456(new_n11833, new_n11829, new_n11827);
nor_4  g11457(new_n11834, new_n11816, new_n11579);
and_4  g11458(new_n11835, new_n11834, new_n11577);
not_3  g11459(new_n11836, new_n11639);
nor_4  g11460(new_n11837, new_n11834, new_n11836);
nor_4  g11461(new_n11838, new_n11837, new_n11835);
nand_4 g11462(new_n11839, new_n11838, new_n11833);
nand_4 g11463(new_n11840, new_n11839, new_n11832);
not_3  g11464(new_n11841, new_n11812);
xnor_3 g11465(new_n11842, new_n11841, new_n11811);
nand_4 g11466(new_n11843, new_n11842, new_n11840);
nand_4 g11467(new_n11844, new_n11843, new_n11814);
nor_4  g11468(new_n11845, new_n11844, new_n11810);
nor_4  g11469(new_n11846, new_n11845, new_n11809);
nand_4 g11470(new_n11847, new_n11846, new_n11806);
xnor_3 g11471(new_n11848, new_n11789, new_n11788);
xnor_3 g11472(new_n11849, new_n11846, new_n11805);
nand_4 g11473(new_n11850, new_n11849, new_n11848);
nand_4 g11474(new_n11851, new_n11850, new_n11847);
xnor_3 g11475(new_n11852, new_n11851, new_n11801);
xnor_3 g11476(new_n11853, new_n11852, new_n11518);
xnor_3 g11477(new_n11854, new_n11501, new_n11498);
xnor_3 g11478(new_n11855, new_n11854, new_n11514);
xnor_3 g11479(new_n11856, new_n11513, new_n11512);
xnor_3 g11480(new_n11857, new_n11510, new_n11509);
not_3  g11481(new_n11858, new_n11857);
xnor_3 g11482(new_n11859, new_n11842, new_n11840);
nand_4 g11483(new_n11860, new_n11859, new_n11858);
not_3  g11484(new_n11861, new_n11860);
xnor_3 g11485(new_n11862, new_n11859, new_n11858);
xnor_3 g11486(new_n11863, new_n11838, new_n11833);
nand_4 g11487(new_n11864, n12709, n6877);
not_3  g11488(new_n11865, new_n11864);
nor_4  g11489(new_n11866, new_n11865, new_n11449);
and_4  g11490(new_n11867, new_n11866, new_n11447);
not_3  g11491(new_n11868, new_n11503);
nor_4  g11492(new_n11869, new_n11866, new_n11868);
nor_4  g11493(new_n11870, new_n11869, new_n11867);
not_3  g11494(new_n11871, new_n11870);
nand_4 g11495(new_n11872, new_n11871, new_n11863);
not_3  g11496(new_n11873, new_n11872);
xnor_3 g11497(new_n11874, new_n11871, new_n11863);
xnor_3 g11498(new_n11875, new_n11825, new_n11821_1);
xor_3  g11499(new_n11876_1, new_n11505, new_n11504);
nand_4 g11500(new_n11877_1, new_n11876_1, new_n11875);
not_3  g11501(new_n11878, new_n11877_1);
xor_3  g11502(new_n11879, new_n11816, new_n11778);
nor_4  g11503(new_n11880, new_n11879, new_n11864);
not_3  g11504(new_n11881, new_n11880);
xnor_3 g11505(new_n11882, new_n11876_1, new_n11875);
nor_4  g11506(new_n11883, new_n11882, new_n11881);
nor_4  g11507(new_n11884, new_n11883, new_n11878);
nor_4  g11508(new_n11885, new_n11884, new_n11874);
nor_4  g11509(new_n11886, new_n11885, new_n11873);
nor_4  g11510(new_n11887, new_n11886, new_n11862);
nor_4  g11511(new_n11888, new_n11887, new_n11861);
nand_4 g11512(new_n11889, new_n11888, new_n11856);
not_3  g11513(new_n11890, new_n11856);
xnor_3 g11514(new_n11891, new_n11888, new_n11890);
xnor_3 g11515(new_n11892_1, new_n11844, new_n11810);
nand_4 g11516(new_n11893, new_n11892_1, new_n11891);
nand_4 g11517(new_n11894, new_n11893, new_n11889);
not_3  g11518(new_n11895, new_n11894);
nor_4  g11519(new_n11896, new_n11895, new_n11855);
not_3  g11520(new_n11897, new_n11896);
not_3  g11521(new_n11898, new_n11850);
nor_4  g11522(new_n11899, new_n11849, new_n11848);
nor_4  g11523(new_n11900, new_n11899, new_n11898);
xnor_3 g11524(new_n11901, new_n11894, new_n11855);
nand_4 g11525(new_n11902, new_n11901, new_n11900);
nand_4 g11526(new_n11903, new_n11902, new_n11897);
nand_4 g11527(new_n11904, new_n11903, new_n11853);
xnor_3 g11528(new_n11905, new_n11517, new_n11495);
xnor_3 g11529(new_n11906, new_n11852, new_n11905);
not_3  g11530(new_n11907, new_n11900);
xnor_3 g11531(new_n11908, new_n11515, new_n11514);
xnor_3 g11532(new_n11909, new_n11894, new_n11908);
nor_4  g11533(new_n11910, new_n11909, new_n11907);
nor_4  g11534(new_n11911, new_n11910, new_n11896);
nand_4 g11535(new_n11912, new_n11911, new_n11906);
nand_4 g11536(new_n11913, new_n11912, new_n11904);
not_3  g11537(new_n11914, new_n11913);
nand_4 g11538(new_n11915, new_n11914, new_n11386);
xnor_3 g11539(new_n11916, new_n11913, new_n11386);
xnor_3 g11540(new_n11917_1, new_n11383, new_n11382);
not_3  g11541(new_n11918, new_n11917_1);
xnor_3 g11542(new_n11919_1, new_n11380, new_n11379);
not_3  g11543(new_n11920, new_n11892_1);
xnor_3 g11544(new_n11921, new_n11920, new_n11891);
nand_4 g11545(new_n11922_1, new_n11921, new_n11919_1);
not_3  g11546(new_n11923, new_n11919_1);
xnor_3 g11547(new_n11924, new_n11921, new_n11923);
not_3  g11548(new_n11925, new_n11378);
xor_3  g11549(new_n11926, new_n11925, new_n11376);
xnor_3 g11550(new_n11927, new_n11886, new_n11862);
not_3  g11551(new_n11928, new_n11927);
nor_4  g11552(new_n11929, new_n11928, new_n11926);
not_3  g11553(new_n11930, new_n11929);
xnor_3 g11554(new_n11931, new_n11884, new_n11874);
not_3  g11555(new_n11932, new_n11931);
not_3  g11556(new_n11933, new_n11319);
nor_4  g11557(new_n11934, new_n11321, new_n11933);
nor_4  g11558(new_n11935, new_n11934, new_n11371);
not_3  g11559(new_n11936, new_n11934);
nor_4  g11560(new_n11937, new_n11936, new_n11318);
nor_4  g11561(new_n11938, new_n11937, new_n11935);
nor_4  g11562(new_n11939, new_n11938, new_n11932);
not_3  g11563(new_n11940, new_n11939);
not_3  g11564(new_n11941, new_n11938);
nor_4  g11565(new_n11942, new_n11941, new_n11931);
nor_4  g11566(new_n11943, new_n11942, new_n11939);
xor_3  g11567(new_n11944, new_n11815, new_n11778);
nor_4  g11568(new_n11945, new_n11944, new_n11865);
nor_4  g11569(new_n11946, new_n11945, new_n11880);
nand_4 g11570(new_n11947, new_n11946, new_n11933);
not_3  g11571(new_n11948, new_n11947);
xor_3  g11572(new_n11949, new_n11373, new_n11372);
nor_4  g11573(new_n11950, new_n11949, new_n11948);
not_3  g11574(new_n11951, new_n11950);
not_3  g11575(new_n11952, new_n11882);
xor_3  g11576(new_n11953, new_n11952, new_n11881);
xor_3  g11577(new_n11954, new_n11949, new_n11948);
nand_4 g11578(new_n11955, new_n11954, new_n11953);
nand_4 g11579(new_n11956, new_n11955, new_n11951);
nand_4 g11580(new_n11957, new_n11956, new_n11943);
nand_4 g11581(new_n11958, new_n11957, new_n11940);
not_3  g11582(new_n11959, new_n11926);
nor_4  g11583(new_n11960, new_n11927, new_n11959);
nor_4  g11584(new_n11961, new_n11960, new_n11929);
nand_4 g11585(new_n11962, new_n11961, new_n11958);
nand_4 g11586(new_n11963, new_n11962, new_n11930);
nand_4 g11587(new_n11964, new_n11963, new_n11924);
nand_4 g11588(new_n11965, new_n11964, new_n11922_1);
nand_4 g11589(new_n11966, new_n11965, new_n11918);
nor_4  g11590(new_n11967_1, new_n11901, new_n11900);
nor_4  g11591(new_n11968, new_n11967_1, new_n11910);
xnor_3 g11592(new_n11969, new_n11965, new_n11917_1);
nand_4 g11593(new_n11970, new_n11969, new_n11968);
nand_4 g11594(new_n11971, new_n11970, new_n11966);
nand_4 g11595(new_n11972, new_n11971, new_n11916);
nand_4 g11596(new_n11973, new_n11972, new_n11915);
not_3  g11597(new_n11974, new_n11852);
nor_4  g11598(new_n11975, new_n11974, new_n11518);
not_3  g11599(new_n11976, new_n11904);
nor_4  g11600(new_n11977, new_n11976, new_n11975);
xnor_3 g11601(new_n11978, new_n11977, new_n11973);
nand_4 g11602(new_n11979, new_n11768, new_n11735);
nand_4 g11603(new_n11980, new_n11791_1, new_n11798);
nand_4 g11604(new_n11981, new_n11980, new_n11979);
not_3  g11605(new_n11982, new_n11494);
nand_4 g11606(new_n11983, new_n11982, new_n11464);
nand_4 g11607(new_n11984, new_n11517, new_n11495);
nand_4 g11608(new_n11985, new_n11984, new_n11983);
xnor_3 g11609(new_n11986, new_n11985, new_n11981);
nand_4 g11610(new_n11987, new_n11363, new_n11335);
nand_4 g11611(new_n11988, new_n11385, new_n11364);
nand_4 g11612(new_n11989, new_n11988, new_n11987);
not_3  g11613(new_n11990, new_n11354);
nand_4 g11614(new_n11991, new_n11360, new_n11990);
nand_4 g11615(new_n11992, new_n11361, new_n11353);
nand_4 g11616(new_n11993, new_n11992, new_n11991);
nand_4 g11617(new_n11994, n6877, n1198);
nand_4 g11618(new_n11995, n12753, n11728);
xor_3  g11619(new_n11996, new_n11995, new_n11994);
nand_4 g11620(new_n11997, n10990, n4722);
nand_4 g11621(new_n11998, n1478, n1471);
xor_3  g11622(new_n11999_1, new_n11998, new_n11997);
xor_3  g11623(new_n12000_1, new_n11999_1, new_n11996);
xnor_3 g11624(new_n12001, new_n12000_1, new_n11993);
nand_4 g11625(new_n12002, n6429, n4203);
not_3  g11626(new_n12003, new_n12002);
nand_4 g11627(new_n12004, new_n11480, new_n11473);
not_3  g11628(new_n12005_1, new_n11481);
nand_4 g11629(new_n12006, new_n11492, new_n12005_1);
nand_4 g11630(new_n12007, new_n12006, new_n12004);
xnor_3 g11631(new_n12008, new_n12007, new_n12003);
xnor_3 g11632(new_n12009, new_n12008, new_n12001);
nand_4 g11633(new_n12010, n8819, n4187);
not_3  g11634(new_n12011, new_n11476);
nor_4  g11635(new_n12012, new_n11478_1, new_n12011);
nor_4  g11636(new_n12013, new_n11479, new_n11475);
nor_4  g11637(new_n12014_1, new_n12013, new_n12012);
xor_3  g11638(new_n12015, new_n12014_1, new_n12010);
xnor_3 g11639(new_n12016, new_n12015, new_n12009);
nand_4 g11640(new_n12017, new_n11468, new_n11466);
nand_4 g11641(new_n12018, new_n11493, new_n11470);
nand_4 g11642(new_n12019, new_n12018, new_n12017);
nor_4  g11643(new_n12020_1, new_n11344, new_n11342);
not_3  g11644(new_n12021, new_n11345);
nor_4  g11645(new_n12022, new_n11352, new_n12021);
nor_4  g11646(new_n12023, new_n12022, new_n12020_1);
nand_4 g11647(new_n12024, n9080, n5212);
xor_3  g11648(new_n12025_1, new_n12024, new_n12023);
not_3  g11649(new_n12026, new_n11356);
nor_4  g11650(new_n12027, new_n11358, new_n12026);
not_3  g11651(new_n12028, new_n11355);
nor_4  g11652(new_n12029, new_n11359, new_n12028);
nor_4  g11653(new_n12030, new_n12029, new_n12027);
nand_4 g11654(new_n12031, n12709, n10174);
not_3  g11655(new_n12032, new_n12031);
nand_4 g11656(new_n12033, n12000, n3172);
nand_4 g11657(new_n12034, n5240, n4370);
xor_3  g11658(new_n12035, new_n12034, new_n12033);
xnor_3 g11659(new_n12036, new_n12035, new_n12032);
xnor_3 g11660(new_n12037, new_n12036, new_n12030);
nand_4 g11661(new_n12038, n9725, n1333);
not_3  g11662(new_n12039, new_n12038);
nand_4 g11663(new_n12040, n11757, n5320);
nand_4 g11664(new_n12041, n11877, n11821);
xor_3  g11665(new_n12042, new_n12041, new_n12040);
xnor_3 g11666(new_n12043, new_n12042, new_n12039);
not_3  g11667(new_n12044_1, new_n11348);
nor_4  g11668(new_n12045, new_n11350, new_n12044_1);
nor_4  g11669(new_n12046, new_n11351, new_n11347);
nor_4  g11670(new_n12047, new_n12046, new_n12045);
xnor_3 g11671(new_n12048, new_n12047, new_n12043);
xnor_3 g11672(new_n12049, new_n12048, new_n12037);
nand_4 g11673(new_n12050, n7646, n5760);
nand_4 g11674(new_n12051, n10022, n7236);
not_3  g11675(new_n12052, new_n12051);
xor_3  g11676(new_n12053, new_n12052, new_n12050);
xnor_3 g11677(new_n12054, new_n12053, new_n12049);
xnor_3 g11678(new_n12055, new_n12054, new_n12025_1);
xnor_3 g11679(new_n12056, new_n12055, new_n12019);
xnor_3 g11680(new_n12057, new_n12056, new_n12016);
xnor_3 g11681(new_n12058, new_n12057, new_n11989);
xnor_3 g11682(new_n12059, new_n12058, new_n11986);
not_3  g11683(new_n12060, new_n11801);
not_3  g11684(new_n12061, new_n11851);
nand_4 g11685(new_n12062, new_n12061, new_n12060);
nand_4 g11686(new_n12063, new_n12062, new_n11793);
nor_4  g11687(new_n12064, new_n11615, new_n11614);
xor_3  g11688(new_n12065, new_n11615, new_n11613);
nor_4  g11689(new_n12066, new_n11621, new_n12065);
nor_4  g11690(new_n12067, new_n12066, new_n12064);
and_4  g11691(new_n12068, new_n11742, new_n11741);
nor_4  g11692(new_n12069_1, new_n11745, new_n12068);
nand_4 g11693(new_n12070, n4805, n4436);
not_3  g11694(new_n12071, new_n12070);
not_3  g11695(new_n12072, new_n11603);
nand_4 g11696(new_n12073, new_n11606, new_n12072);
nand_4 g11697(new_n12074, new_n12073, new_n11609);
xor_3  g11698(new_n12075, new_n12074, new_n12071);
xor_3  g11699(new_n12076_1, new_n12075, new_n12069_1);
xnor_3 g11700(new_n12077, new_n12076_1, new_n12067);
nand_4 g11701(new_n12078, new_n11750, new_n11748);
not_3  g11702(new_n12079, new_n11759);
nand_4 g11703(new_n12080, new_n12079, new_n11751);
nand_4 g11704(new_n12081, new_n12080, new_n12078);
nand_4 g11705(new_n12082, n7159, n3146);
not_3  g11706(new_n12083, new_n12082);
nand_4 g11707(new_n12084, n11967, n137);
nand_4 g11708(new_n12085, n8384, n6441);
xor_3  g11709(new_n12086, new_n12085, new_n12084);
xor_3  g11710(new_n12087, new_n12086, new_n12083);
nand_4 g11711(new_n12088, n12777, n6797);
nand_4 g11712(new_n12089, n6294, n6254);
xor_3  g11713(new_n12090, new_n12089, new_n12088);
nand_4 g11714(new_n12091, n12947, n6358);
nand_4 g11715(new_n12092, n11999, n3992);
not_3  g11716(new_n12093, new_n12092);
xor_3  g11717(new_n12094, new_n12093, new_n12091);
xor_3  g11718(new_n12095, new_n12094, new_n12090);
xnor_3 g11719(new_n12096, new_n12095, new_n12087);
xnor_3 g11720(new_n12097, new_n12096, new_n12081);
nand_4 g11721(new_n12098, n11478, n1353);
nand_4 g11722(new_n12099, n7862, n6604);
nand_4 g11723(new_n12100, n11407, n6826);
xor_3  g11724(new_n12101, new_n12100, new_n12099);
xor_3  g11725(new_n12102, new_n12101, new_n12098);
nor_4  g11726(new_n12103, new_n11619, new_n11618);
not_3  g11727(new_n12104, new_n11617);
nand_4 g11728(new_n12105, new_n11619, new_n11618);
nand_4 g11729(new_n12106, new_n12105, new_n12104);
not_3  g11730(new_n12107, new_n12106);
nor_4  g11731(new_n12108, new_n12107, new_n12103);
xnor_3 g11732(new_n12109, new_n12108, new_n12102);
xnor_3 g11733(new_n12110, new_n12109, new_n12097);
xnor_3 g11734(new_n12111_1, new_n12110, new_n12077);
not_3  g11735(new_n12112, new_n11602);
nand_4 g11736(new_n12113, new_n11611, new_n12112);
xnor_3 g11737(new_n12114, new_n11621, new_n12065);
nand_4 g11738(new_n12115, new_n12114, new_n11612);
nand_4 g11739(new_n12116, new_n12115, new_n12113);
not_3  g11740(new_n12117, new_n11746);
nor_4  g11741(new_n12118, new_n12117, new_n11738);
not_3  g11742(new_n12119, new_n11747);
nor_4  g11743(new_n12120, new_n11760, new_n12119);
nor_4  g11744(new_n12121, new_n12120, new_n12118);
xor_3  g11745(new_n12122, new_n12121, new_n12116);
xnor_3 g11746(new_n12123, new_n12122, new_n12111_1);
nand_4 g11747(new_n12124, new_n11630, new_n11600);
nand_4 g11748(new_n12125, new_n11653, new_n11795);
nand_4 g11749(new_n12126, new_n12125, new_n12124);
nor_4  g11750(new_n12127, new_n11700, new_n11765);
not_3  g11751(new_n12128, new_n11767);
nor_4  g11752(new_n12129, new_n12128, new_n11761);
nor_4  g11753(new_n12130, new_n12129, new_n12127);
xnor_3 g11754(new_n12131, new_n12130, new_n12126);
nor_4  g11755(new_n12132, new_n11564, new_n11627);
not_3  g11756(new_n12133, new_n11629);
nor_4  g11757(new_n12134, new_n12133, new_n11623);
nor_4  g11758(new_n12135, new_n12134, new_n12132);
nand_4 g11759(new_n12136, new_n11303, new_n11339);
nand_4 g11760(new_n12137, new_n11362, new_n11341);
nand_4 g11761(new_n12138, new_n12137, new_n12136);
and_4  g11762(new_n12139, new_n11755_1, new_n11754);
nor_4  g11763(new_n12140, new_n11758, new_n12139);
nand_4 g11764(new_n12141, n5283, n447);
nand_4 g11765(new_n12142, n12489, n4938);
nand_4 g11766(new_n12143, n11791, n5198);
xor_3  g11767(new_n12144, new_n12143, new_n12142);
xor_3  g11768(new_n12145_1, new_n12144, new_n12141);
xnor_3 g11769(new_n12146, new_n12145_1, new_n12140);
xnor_3 g11770(new_n12147, new_n12146, new_n12138);
nand_4 g11771(new_n12148, n8717, n2464);
not_3  g11772(new_n12149, new_n12148);
nor_4  g11773(new_n12150, new_n11484, new_n11483);
not_3  g11774(new_n12151, new_n11485);
nor_4  g11775(new_n12152, new_n11491, new_n12151);
nor_4  g11776(new_n12153, new_n12152, new_n12150);
not_3  g11777(new_n12154, new_n11487);
nor_4  g11778(new_n12155, new_n11489, new_n12154);
not_3  g11779(new_n12156, new_n11486);
nor_4  g11780(new_n12157, new_n11490, new_n12156);
nor_4  g11781(new_n12158, new_n12157, new_n12155);
nand_4 g11782(new_n12159, n11311, n2433);
nand_4 g11783(new_n12160, n9400, n7730);
not_3  g11784(new_n12161, new_n12160);
xor_3  g11785(new_n12162, new_n12161, new_n12159);
xnor_3 g11786(new_n12163, new_n12162, new_n12158);
xnor_3 g11787(new_n12164, new_n12163, new_n12153);
xnor_3 g11788(new_n12165, new_n12164, new_n12149);
xnor_3 g11789(new_n12166, new_n12165, new_n12147);
xnor_3 g11790(new_n12167, new_n12166, new_n12135);
xnor_3 g11791(new_n12168, new_n12167, new_n12131);
xnor_3 g11792(new_n12169, new_n12168, new_n12123);
xnor_3 g11793(new_n12170, new_n12169, new_n12063);
xnor_3 g11794(new_n12171, new_n12170, new_n12059);
xnor_3 g11795(n4378, new_n12171, new_n11978);
xor_3  g11796(n4397, new_n4109, new_n4021);
xor_3  g11797(n4553, new_n4453, new_n4442);
xor_3  g11798(n4686, new_n1043, new_n1033);
xnor_3 g11799(n4689, new_n10023, new_n10005);
not_3  g11800(new_n12177, new_n5277);
nand_4 g11801(new_n12178, new_n5232, new_n5231);
xnor_3 g11802(n4733, new_n12178, new_n12177);
xnor_3 g11803(n4757, new_n2184, new_n2176);
not_3  g11804(new_n12181, new_n5273);
xor_3  g11805(n4971, new_n12181, new_n5271);
xnor_3 g11806(n5030, new_n7035, new_n7034);
not_3  g11807(new_n12184, new_n3089);
xor_3  g11808(n5034, new_n12184, new_n3056);
not_3  g11809(new_n12186, new_n3073);
xor_3  g11810(n5094, new_n3082, new_n12186);
nand_4 g11811(new_n12188, new_n11124, new_n11115);
nand_4 g11812(new_n12189, n5320, n2564);
nand_4 g11813(new_n12190, n4370, n4189);
xor_3  g11814(new_n12191, new_n12190, new_n12189);
xnor_3 g11815(new_n12192, new_n12191, new_n12188);
nand_4 g11816(new_n12193, n11877, n6770);
not_3  g11817(new_n12194, new_n12193);
and_4  g11818(new_n12195, new_n11121, new_n11120);
not_3  g11819(new_n12196, new_n11119);
nor_4  g11820(new_n12197, new_n11122, new_n12196);
nor_4  g11821(new_n12198, new_n12197, new_n12195);
nand_4 g11822(new_n12199, new_n12198, new_n12194);
not_3  g11823(new_n12200, new_n12199);
nor_4  g11824(new_n12201, new_n12198, new_n12194);
nor_4  g11825(new_n12202, new_n12201, new_n12200);
nand_4 g11826(new_n12203, n9920, n5212);
nand_4 g11827(new_n12204, n11407, n3627);
xor_3  g11828(new_n12205, new_n12204, new_n12203);
xnor_3 g11829(new_n12206, new_n12205, new_n12202);
xnor_3 g11830(new_n12207, new_n12206, new_n12192);
not_3  g11831(new_n12208, new_n12207);
nor_4  g11832(new_n12209, new_n11108, new_n11103);
not_3  g11833(new_n12210, new_n12209);
not_3  g11834(new_n12211, new_n11103);
xnor_3 g11835(new_n12212, new_n11108, new_n12211);
nand_4 g11836(new_n12213, new_n11127, new_n12212);
nand_4 g11837(new_n12214, new_n12213, new_n12210);
nand_4 g11838(new_n12215, new_n12214, new_n12208);
nand_4 g11839(new_n12216, new_n12205, new_n12202);
nand_4 g11840(new_n12217, new_n12216, new_n12199);
nand_4 g11841(new_n12218, n12000, n2564);
not_3  g11842(new_n12219, new_n12218);
nand_4 g11843(new_n12220, n5320, n4189);
nand_4 g11844(new_n12221_1, n9725, n6687);
xor_3  g11845(new_n12222, new_n12221_1, new_n12220);
xnor_3 g11846(new_n12223, new_n12222, new_n12219);
xnor_3 g11847(new_n12224, new_n12223, new_n12217);
nor_4  g11848(new_n12225, new_n12204, new_n12203);
nand_4 g11849(new_n12226, n6770, n4370);
not_3  g11850(new_n12227, new_n12226);
xor_3  g11851(new_n12228, new_n12227, new_n12225);
nand_4 g11852(new_n12229, n5212, n3627);
nand_4 g11853(new_n12230, n11877, n9920);
nand_4 g11854(new_n12231, n11407, n4516);
nand_4 g11855(new_n12232, new_n12231, new_n12230);
not_3  g11856(new_n12233, new_n12230);
not_3  g11857(new_n12234, new_n12231);
nand_4 g11858(new_n12235, new_n12234, new_n12233);
nand_4 g11859(new_n12236, new_n12235, new_n12232);
xor_3  g11860(new_n12237, new_n12236, new_n12229);
xnor_3 g11861(new_n12238, new_n12237, new_n12228);
not_3  g11862(new_n12239, new_n12238);
xnor_3 g11863(new_n12240, new_n12239, new_n12224);
not_3  g11864(new_n12241, new_n12240);
not_3  g11865(new_n12242, new_n12188);
not_3  g11866(new_n12243, new_n12191);
nor_4  g11867(new_n12244, new_n12243, new_n12242);
not_3  g11868(new_n12245, new_n12244);
nor_4  g11869(new_n12246, new_n12190, new_n12189);
nor_4  g11870(new_n12247_1, new_n12206, new_n12192);
xnor_3 g11871(new_n12248, new_n12247_1, new_n12246);
nand_4 g11872(new_n12249, new_n12248, new_n12245);
nor_4  g11873(new_n12250, new_n12249, new_n12241);
nand_4 g11874(new_n12251, new_n12249, new_n12241);
not_3  g11875(new_n12252, new_n12251);
nor_4  g11876(new_n12253, new_n12252, new_n12250);
xnor_3 g11877(new_n12254, new_n12253, new_n12215);
nand_4 g11878(new_n12255, n12000, n6687);
not_3  g11879(new_n12256, new_n12255);
xnor_3 g11880(new_n12257, new_n12214, new_n12208);
not_3  g11881(new_n12258, new_n12257);
nand_4 g11882(new_n12259, new_n12258, new_n12256);
nor_4  g11883(new_n12260, new_n11129, new_n11102);
xnor_3 g11884(new_n12261, new_n12257, new_n12256);
nand_4 g11885(new_n12262, new_n12261, new_n12260);
nand_4 g11886(new_n12263, new_n12262, new_n12259);
xnor_3 g11887(new_n12264, new_n12263, new_n12254);
not_3  g11888(new_n12265, new_n12264);
nand_4 g11889(new_n12266, n8717, n8336);
nand_4 g11890(new_n12267, n6429, n2226);
nand_4 g11891(new_n12268, n11728, n1094);
nand_4 g11892(new_n12269, n12709, n10678);
xnor_3 g11893(new_n12270, new_n12269, new_n12268);
nor_4  g11894(new_n12271, new_n12270, new_n12267);
not_3  g11895(new_n12272, new_n12267);
not_3  g11896(new_n12273, new_n12270);
nor_4  g11897(new_n12274, new_n12273, new_n12272);
nor_4  g11898(new_n12275, new_n12274, new_n12271);
nor_4  g11899(new_n12276, new_n11151, new_n11145);
nor_4  g11900(new_n12277, new_n12276, new_n11150);
xnor_3 g11901(new_n12278, new_n12277, new_n12275);
nand_4 g11902(new_n12279, n10928, n2433);
nand_4 g11903(new_n12280, n8819, n6986);
xor_3  g11904(new_n12281, new_n12280, new_n12279);
xnor_3 g11905(new_n12282, new_n12281, new_n12278);
nand_4 g11906(new_n12283, new_n11142, new_n11136);
not_3  g11907(new_n12284, new_n12283);
nor_4  g11908(new_n12285, new_n11153_1, new_n11143);
nor_4  g11909(new_n12286, new_n12285, new_n12284);
not_3  g11910(new_n12287, new_n12286);
nand_4 g11911(new_n12288, new_n12287, new_n12282);
not_3  g11912(new_n12289, new_n12288);
nor_4  g11913(new_n12290, new_n12287, new_n12282);
nor_4  g11914(new_n12291, new_n12290, new_n12289);
not_3  g11915(new_n12292, new_n11155);
nand_4 g11916(new_n12293, new_n11163, new_n11159);
nand_4 g11917(new_n12294, new_n12293, new_n12292);
xnor_3 g11918(new_n12295, new_n12294, new_n12291);
nor_4  g11919(new_n12296, new_n12295, new_n12266);
not_3  g11920(new_n12297, new_n12296);
not_3  g11921(new_n12298, new_n11133);
nor_4  g11922(new_n12299_1, new_n11164, new_n12298);
not_3  g11923(new_n12300, new_n12266);
xnor_3 g11924(new_n12301, new_n12295, new_n12300);
nand_4 g11925(new_n12302, new_n12301, new_n12299_1);
nand_4 g11926(new_n12303, new_n12302, new_n12297);
nand_4 g11927(new_n12304, new_n12294, new_n12291);
not_3  g11928(new_n12305, new_n12271);
nand_4 g11929(new_n12306, new_n12277, new_n12275);
and_4  g11930(new_n12307, new_n12306, new_n12305);
nand_4 g11931(new_n12308, n10928, n8717);
not_3  g11932(new_n12309, new_n12308);
nand_4 g11933(new_n12310, n6986, n2433);
nand_4 g11934(new_n12311, n8336, n7730);
not_3  g11935(new_n12312, new_n12311);
xor_3  g11936(new_n12313, new_n12312, new_n12310);
xnor_3 g11937(new_n12314, new_n12313, new_n12309);
xnor_3 g11938(new_n12315, new_n12314, new_n12307);
nor_4  g11939(new_n12316, new_n12269, new_n12268);
not_3  g11940(new_n12317, new_n12316);
nand_4 g11941(new_n12318, n8819, n2226);
xor_3  g11942(new_n12319, new_n12318, new_n12317);
nand_4 g11943(new_n12320, n11728, n10678);
nand_4 g11944(new_n12321, n6429, n1094);
nand_4 g11945(new_n12322, n12709, n7320);
not_3  g11946(new_n12323, new_n12322);
xor_3  g11947(new_n12324, new_n12323, new_n12321);
xnor_3 g11948(new_n12325, new_n12324, new_n12320);
xnor_3 g11949(new_n12326, new_n12325, new_n12319);
xnor_3 g11950(new_n12327, new_n12326, new_n12315);
not_3  g11951(new_n12328, new_n12278);
nand_4 g11952(new_n12329, new_n12281, new_n12328);
nor_4  g11953(new_n12330, new_n12280, new_n12279);
xnor_3 g11954(new_n12331, new_n12289, new_n12330);
nand_4 g11955(new_n12332, new_n12331, new_n12329);
xnor_3 g11956(new_n12333, new_n12332, new_n12327);
xnor_3 g11957(new_n12334, new_n12333, new_n12304);
xnor_3 g11958(new_n12335, new_n12334, new_n12303);
xnor_3 g11959(new_n12336, new_n12301, new_n12299_1);
not_3  g11960(new_n12337, new_n11169);
not_3  g11961(new_n12338, new_n11173);
nor_4  g11962(new_n12339, new_n11246, new_n12338);
nor_4  g11963(new_n12340, new_n12339, new_n12337);
nor_4  g11964(new_n12341, new_n12340, new_n12336);
not_3  g11965(new_n12342, new_n12341);
nand_4 g11966(new_n12343, new_n12340, new_n12336);
nor_4  g11967(new_n12344, new_n11234, new_n11241);
not_3  g11968(new_n12345, new_n12344);
nand_4 g11969(new_n12346, n11222, n6441);
not_3  g11970(new_n12347, new_n11210);
nand_4 g11971(new_n12348, new_n11216_1, new_n12347);
nand_4 g11972(new_n12349, new_n11228, new_n11217);
nand_4 g11973(new_n12350, new_n12349, new_n12348);
nand_4 g11974(new_n12351, n12947, n11153);
nand_4 g11975(new_n12352, n11791, n5314);
xor_3  g11976(new_n12353, new_n12352, new_n12351);
xnor_3 g11977(new_n12354, new_n12353, new_n12350);
nand_4 g11978(new_n12355, n1478, n996);
nand_4 g11979(new_n12356, n10990, n5319);
nand_4 g11980(new_n12357, n5767, n5760);
xnor_3 g11981(new_n12358, new_n12357, new_n12356);
nor_4  g11982(new_n12359, new_n12358, new_n12355);
not_3  g11983(new_n12360, new_n12355);
not_3  g11984(new_n12361, new_n12358);
nor_4  g11985(new_n12362, new_n12361, new_n12360);
nor_4  g11986(new_n12363, new_n12362, new_n12359);
nand_4 g11987(new_n12364, new_n11225, new_n11218);
nand_4 g11988(new_n12365, new_n12364, new_n11221);
xor_3  g11989(new_n12366, new_n12365, new_n12363);
xnor_3 g11990(new_n12367, new_n12366, new_n12354);
nor_4  g11991(new_n12368, new_n11229, new_n11209);
nor_4  g11992(new_n12369, new_n11233, new_n11230);
nor_4  g11993(new_n12370, new_n12369, new_n12368);
nor_4  g11994(new_n12371, new_n12370, new_n12367);
not_3  g11995(new_n12372, new_n12367);
not_3  g11996(new_n12373, new_n12370);
nor_4  g11997(new_n12374, new_n12373, new_n12372);
nor_4  g11998(new_n12375, new_n12374, new_n12371);
xnor_3 g11999(new_n12376, new_n12375, new_n12346);
xnor_3 g12000(new_n12377, new_n12376, new_n12345);
not_3  g12001(new_n12378, new_n11206);
nand_4 g12002(new_n12379, n12069, n447);
nand_4 g12003(new_n12380, n12777, n7160);
nand_4 g12004(new_n12381, n7159, n4828);
nand_4 g12005(new_n12382, n12489, n2515);
xnor_3 g12006(new_n12383, new_n12382, new_n12381);
nor_4  g12007(new_n12384, new_n12383, new_n12380);
not_3  g12008(new_n12385, new_n12380);
not_3  g12009(new_n12386, new_n12383);
nor_4  g12010(new_n12387, new_n12386, new_n12385);
nor_4  g12011(new_n12388, new_n12387, new_n12384);
nor_4  g12012(new_n12389, new_n11189, new_n11183);
nor_4  g12013(new_n12390, new_n12389, new_n11188);
xnor_3 g12014(new_n12391_1, new_n12390, new_n12388);
nand_4 g12015(new_n12392, n12391, n11967);
nand_4 g12016(new_n12393, n7891, n6254);
not_3  g12017(new_n12394, new_n12393);
xor_3  g12018(new_n12395, new_n12394, new_n12392);
xnor_3 g12019(new_n12396, new_n12395, new_n12391_1);
and_4  g12020(new_n12397, new_n11180, new_n11177);
nor_4  g12021(new_n12398, new_n11191, new_n11181);
nor_4  g12022(new_n12399, new_n12398, new_n12397);
not_3  g12023(new_n12400, new_n12399);
xnor_3 g12024(new_n12401, new_n12400, new_n12396);
not_3  g12025(new_n12402, new_n11193);
nand_4 g12026(new_n12403, new_n11201, new_n11197);
nand_4 g12027(new_n12404, new_n12403, new_n12402);
xnor_3 g12028(new_n12405, new_n12404, new_n12401);
xnor_3 g12029(new_n12406, new_n12405, new_n12379);
not_3  g12030(new_n12407, new_n12406);
nor_4  g12031(new_n12408, new_n12407, new_n12378);
nor_4  g12032(new_n12409, new_n12406, new_n11206);
nor_4  g12033(new_n12410, new_n12409, new_n12408);
not_3  g12034(new_n12411, new_n12410);
nand_4 g12035(new_n12412, new_n11244, new_n11207);
nand_4 g12036(new_n12413, new_n12412, new_n11240);
xnor_3 g12037(new_n12414, new_n12413, new_n12411);
xnor_3 g12038(new_n12415, new_n12414, new_n12377);
nand_4 g12039(new_n12416, new_n12415, new_n12343);
nand_4 g12040(new_n12417, new_n12416, new_n12342);
xnor_3 g12041(new_n12418, new_n12417, new_n12335);
not_3  g12042(new_n12419, new_n12363);
nor_4  g12043(new_n12420, new_n12365, new_n12419);
nor_4  g12044(new_n12421, new_n12420, new_n12359);
not_3  g12045(new_n12422, new_n12421);
nand_4 g12046(new_n12423, n11153, n6441);
nand_4 g12047(new_n12424, n12947, n5314);
nand_4 g12048(new_n12425, n11999, n11222);
not_3  g12049(new_n12426, new_n12425);
xor_3  g12050(new_n12427, new_n12426, new_n12424);
xnor_3 g12051(new_n12428, new_n12427, new_n12423);
xnor_3 g12052(new_n12429, new_n12428, new_n12422);
nor_4  g12053(new_n12430, new_n12357, new_n12356);
nand_4 g12054(new_n12431, n11791, n996);
xor_3  g12055(new_n12432, new_n12431, new_n12430);
nand_4 g12056(new_n12433, n5760, n5319);
nand_4 g12057(new_n12434, n5767, n1478);
nand_4 g12058(new_n12435, n10990, n9457);
not_3  g12059(new_n12436, new_n12435);
xor_3  g12060(new_n12437, new_n12436, new_n12434);
xnor_3 g12061(new_n12438, new_n12437, new_n12433);
xnor_3 g12062(new_n12439, new_n12438, new_n12432);
not_3  g12063(new_n12440, new_n12439);
xnor_3 g12064(new_n12441, new_n12440, new_n12429);
nand_4 g12065(new_n12442, new_n12353, new_n12350);
nor_4  g12066(new_n12443, new_n12352, new_n12351);
nor_4  g12067(new_n12444_1, new_n12366, new_n12354);
xnor_3 g12068(new_n12445, new_n12444_1, new_n12443);
nand_4 g12069(new_n12446, new_n12445, new_n12442);
xnor_3 g12070(new_n12447, new_n12446, new_n12441);
xnor_3 g12071(new_n12448, new_n12447, new_n12371);
not_3  g12072(new_n12449, new_n12346);
nand_4 g12073(new_n12450, new_n12375, new_n12449);
nand_4 g12074(new_n12451, new_n12376, new_n12344);
nand_4 g12075(new_n12452, new_n12451, new_n12450);
xnor_3 g12076(new_n12453, new_n12452, new_n12448);
not_3  g12077(new_n12454, new_n12401);
not_3  g12078(new_n12455, new_n12404);
nor_4  g12079(new_n12456, new_n12455, new_n12454);
not_3  g12080(new_n12457, new_n12456);
nand_4 g12081(new_n12458, new_n12390, new_n12388);
not_3  g12082(new_n12459, new_n12458);
nor_4  g12083(new_n12460, new_n12459, new_n12384);
not_3  g12084(new_n12461, new_n12460);
nand_4 g12085(new_n12462, n12391, n447);
not_3  g12086(new_n12463, new_n12462);
nand_4 g12087(new_n12464, n11967, n7891);
nand_4 g12088(new_n12465, n12069, n1353);
nand_4 g12089(new_n12466, new_n12465, new_n12464);
not_3  g12090(new_n12467, new_n12464);
not_3  g12091(new_n12468, new_n12465);
nand_4 g12092(new_n12469, new_n12468, new_n12467);
nand_4 g12093(new_n12470, new_n12469, new_n12466);
xor_3  g12094(new_n12471, new_n12470, new_n12463);
xnor_3 g12095(new_n12472, new_n12471, new_n12461);
nor_4  g12096(new_n12473, new_n12382, new_n12381);
nand_4 g12097(new_n12474, n7160, n6254);
xor_3  g12098(new_n12475, new_n12474, new_n12473);
nand_4 g12099(new_n12476, n7159, n2515);
not_3  g12100(new_n12477, new_n12476);
nand_4 g12101(new_n12478, n12777, n4828);
nand_4 g12102(new_n12479, n12489, n1199);
nand_4 g12103(new_n12480, new_n12479, new_n12478);
not_3  g12104(new_n12481, new_n12478);
not_3  g12105(new_n12482, new_n12479);
nand_4 g12106(new_n12483, new_n12482, new_n12481);
nand_4 g12107(new_n12484, new_n12483, new_n12480);
xor_3  g12108(new_n12485, new_n12484, new_n12477);
xnor_3 g12109(new_n12486, new_n12485, new_n12475);
not_3  g12110(new_n12487, new_n12486);
xnor_3 g12111(new_n12488, new_n12487, new_n12472);
nor_4  g12112(new_n12489_1, new_n12395, new_n12391_1);
not_3  g12113(new_n12490, new_n12489_1);
nor_4  g12114(new_n12491, new_n12393, new_n12392);
nor_4  g12115(new_n12492, new_n12399, new_n12396);
xnor_3 g12116(new_n12493, new_n12492, new_n12491);
nand_4 g12117(new_n12494, new_n12493, new_n12490);
xnor_3 g12118(new_n12495, new_n12494, new_n12488);
xnor_3 g12119(new_n12496, new_n12495, new_n12457);
not_3  g12120(new_n12497, new_n12379);
not_3  g12121(new_n12498, new_n12405);
nor_4  g12122(new_n12499, new_n12498, new_n12497);
nor_4  g12123(new_n12500, new_n12409, new_n12499);
xnor_3 g12124(new_n12501, new_n12500, new_n12496);
xnor_3 g12125(new_n12502, new_n12501, new_n12453);
nand_4 g12126(new_n12503, new_n12413, new_n12411);
xnor_3 g12127(new_n12504, new_n12413, new_n12410);
nand_4 g12128(new_n12505, new_n12504, new_n12377);
nand_4 g12129(new_n12506, new_n12505, new_n12503);
xnor_3 g12130(new_n12507, new_n12506, new_n12502);
not_3  g12131(new_n12508, new_n12507);
xnor_3 g12132(new_n12509, new_n12508, new_n12418);
not_3  g12133(new_n12510, new_n12509);
nand_4 g12134(new_n12511_1, new_n12510, new_n12265);
nand_4 g12135(new_n12512, new_n12509, new_n12264);
nand_4 g12136(new_n12513, new_n12512, new_n12511_1);
not_3  g12137(new_n12514, new_n12262);
nor_4  g12138(new_n12515, new_n12261, new_n12260);
nor_4  g12139(new_n12516, new_n12515, new_n12514);
nor_4  g12140(new_n12517, new_n11254, new_n11248);
nor_4  g12141(new_n12518, new_n12517, new_n11250);
nor_4  g12142(new_n12519, new_n12518, new_n12516);
xnor_3 g12143(new_n12520, new_n12518, new_n12516);
xnor_3 g12144(new_n12521, new_n12504, new_n12377);
not_3  g12145(new_n12522, new_n12336);
xnor_3 g12146(new_n12523, new_n11245, new_n11207);
nand_4 g12147(new_n12524, new_n12523, new_n11173);
nand_4 g12148(new_n12525, new_n12524, new_n11169);
nor_4  g12149(new_n12526, new_n12525, new_n12522);
nor_4  g12150(new_n12527, new_n12526, new_n12341);
xnor_3 g12151(new_n12528, new_n12527, new_n12521);
nor_4  g12152(new_n12529, new_n12528, new_n12520);
nor_4  g12153(new_n12530, new_n12529, new_n12519);
xnor_3 g12154(n5132, new_n12530, new_n12513);
xor_3  g12155(n5191, new_n11946, new_n11933);
nor_4  g12156(new_n12533, new_n3991, new_n3845);
nor_4  g12157(new_n12534, new_n12533, new_n3848);
nor_4  g12158(new_n12535, new_n3977, new_n3940);
nor_4  g12159(new_n12536, new_n3982, new_n3978);
nor_4  g12160(new_n12537, new_n12536, new_n12535);
not_3  g12161(new_n12538, new_n12537);
not_3  g12162(new_n12539, new_n3352);
nand_4 g12163(new_n12540, new_n3384, new_n12539);
nand_4 g12164(new_n12541, new_n3407, new_n3385);
nand_4 g12165(new_n12542, new_n12541, new_n12540);
nor_4  g12166(new_n12543, new_n3906, new_n3903);
nor_4  g12167(new_n12544, new_n3921, new_n3907);
nor_4  g12168(new_n12545, new_n12544, new_n12543);
xnor_3 g12169(new_n12546, new_n12545, new_n12542);
nand_4 g12170(new_n12547, n1835, n1333);
nand_4 g12171(new_n12548, n9637, n3172);
xor_3  g12172(new_n12549, new_n12548, new_n12547);
nand_4 g12173(new_n12550, n9080, n4921);
nand_4 g12174(new_n12551, n11917, n11821);
xor_3  g12175(new_n12552, new_n12551, new_n12550);
xor_3  g12176(new_n12553, new_n12552, new_n12549);
xnor_3 g12177(new_n12554, new_n12553, new_n12546);
xnor_3 g12178(new_n12555, new_n12554, new_n12538);
nor_4  g12179(new_n12556, new_n3887, new_n3851);
nor_4  g12180(new_n12557, new_n3501, new_n3466);
nor_4  g12181(new_n12558, new_n3890, new_n12557);
nand_4 g12182(new_n12559, new_n12558, new_n3465);
nand_4 g12183(new_n12560, new_n12559, new_n3889);
nor_4  g12184(new_n12561, new_n12560, new_n3888);
nor_4  g12185(new_n12562, new_n12561, new_n12556);
nand_4 g12186(new_n12563, new_n3970, new_n3969);
not_3  g12187(new_n12564, new_n3967);
nand_4 g12188(new_n12565, new_n3972, new_n12564);
nand_4 g12189(new_n12566, new_n12565, new_n12563);
nand_4 g12190(new_n12567, n10174, n3719);
nand_4 g12191(new_n12568, n6877, n4190);
nand_4 g12192(new_n12569, n12753, n3602);
xor_3  g12193(new_n12570, new_n12569, new_n12568);
nand_4 g12194(new_n12571, n4086, n1471);
nand_4 g12195(new_n12572, n8065, n2464);
nand_4 g12196(new_n12573, n11311, n10439);
xor_3  g12197(new_n12574, new_n12573, new_n12572);
xnor_3 g12198(new_n12575, new_n12574, new_n12571);
nand_4 g12199(new_n12576, n7236, n1357);
nand_4 g12200(new_n12577, n7646, n405);
xnor_3 g12201(new_n12578, new_n12577, new_n12576);
nand_4 g12202(new_n12579, n6126, n4203);
nand_4 g12203(new_n12580, n10391, n9400);
xnor_3 g12204(new_n12581, new_n12580, new_n12579);
xnor_3 g12205(new_n12582, new_n12581, new_n12578);
nor_4  g12206(new_n12583, new_n3858, new_n3857);
nand_4 g12207(new_n12584, new_n3858, new_n3857);
nand_4 g12208(new_n12585, new_n12584, new_n3856);
not_3  g12209(new_n12586, new_n12585);
nor_4  g12210(new_n12587, new_n12586, new_n12583);
xnor_3 g12211(new_n12588, new_n12587, new_n12582);
xnor_3 g12212(new_n12589, new_n12588, new_n12575);
xnor_3 g12213(new_n12590, new_n12589, new_n12570);
nand_4 g12214(new_n12591_1, n5240, n3842);
not_3  g12215(new_n12592, new_n12591_1);
nand_4 g12216(new_n12593, n8595, n4187);
nand_4 g12217(new_n12594, n8433, n4722);
xor_3  g12218(new_n12595, new_n12594, new_n12593);
xnor_3 g12219(new_n12596, new_n12595, new_n12592);
nand_4 g12220(new_n12597, new_n3865_1, new_n3863);
nand_4 g12221(new_n12598, new_n3872, new_n3866);
nand_4 g12222(new_n12599, new_n12598, new_n12597);
and_4  g12223(new_n12600, new_n3870, new_n3869);
nor_4  g12224(new_n12601, new_n3871, new_n3868);
nor_4  g12225(new_n12602, new_n12601, new_n12600);
xnor_3 g12226(new_n12603, new_n12602, new_n12599);
xnor_3 g12227(new_n12604, new_n12603, new_n12596);
xnor_3 g12228(new_n12605, new_n12604, new_n12590);
not_3  g12229(new_n12606, new_n3854);
nand_4 g12230(new_n12607, new_n3860, new_n12606);
nand_4 g12231(new_n12608, new_n3873, new_n3861);
nand_4 g12232(new_n12609, new_n12608, new_n12607);
nor_4  g12233(new_n12610, new_n3359, new_n3358);
nand_4 g12234(new_n12611, new_n3359, new_n3358);
nand_4 g12235(new_n12612, new_n12611, new_n3357);
not_3  g12236(new_n12613, new_n12612);
nor_4  g12237(new_n12614, new_n12613, new_n12610);
xnor_3 g12238(new_n12615, new_n12614, new_n12609);
xnor_3 g12239(new_n12616, new_n12615, new_n12605);
xnor_3 g12240(new_n12617, new_n12616, new_n12567);
xnor_3 g12241(new_n12618, new_n12617, new_n12566);
nor_4  g12242(new_n12619, new_n3886, new_n3875);
nor_4  g12243(new_n12620, new_n12619, new_n3882);
not_3  g12244(new_n12621, new_n3355);
nand_4 g12245(new_n12622, new_n3361, new_n12621);
not_3  g12246(new_n12623, new_n3377);
nand_4 g12247(new_n12624, new_n12623, new_n3362);
nand_4 g12248(new_n12625, new_n12624, new_n12622);
nor_4  g12249(new_n12626, new_n3365, new_n3364);
nor_4  g12250(new_n12627, new_n3376, new_n12626);
not_3  g12251(new_n12628, new_n3368);
nor_4  g12252(new_n12629, new_n3370, new_n12628);
not_3  g12253(new_n12630, new_n3367);
nor_4  g12254(new_n12631, new_n3371, new_n12630);
nor_4  g12255(new_n12632, new_n12631, new_n12629);
nand_4 g12256(new_n12633, n11757, n2577);
not_3  g12257(new_n12634, new_n12633);
xnor_3 g12258(new_n12635, new_n12634, new_n12632);
xnor_3 g12259(new_n12636, new_n12635, new_n12627);
xnor_3 g12260(new_n12637, new_n12636, new_n12625);
xnor_3 g12261(new_n12638, new_n12637, new_n12620);
xnor_3 g12262(new_n12639, new_n12638, new_n12618);
xnor_3 g12263(new_n12640, new_n12639, new_n12562);
nand_4 g12264(new_n12641, new_n3973, new_n3943);
not_3  g12265(new_n12642, new_n3974);
not_3  g12266(new_n12643, new_n3976);
nand_4 g12267(new_n12644, new_n12643, new_n12642);
nand_4 g12268(new_n12645, new_n12644, new_n12641);
or_4   g12269(new_n12646, new_n3917, new_n3912);
not_3  g12270(new_n12647, new_n12646);
nor_4  g12271(new_n12648_1, new_n12647, new_n3918);
xnor_3 g12272(new_n12649, new_n12648_1, new_n12645);
xnor_3 g12273(new_n12650, new_n12649, new_n12640);
xnor_3 g12274(new_n12651, new_n12650, new_n12555);
not_3  g12275(new_n12652, new_n3893);
nand_4 g12276(new_n12653, new_n3983, new_n12652);
nand_4 g12277(new_n12654, new_n3990, new_n3984);
nand_4 g12278(new_n12655, new_n12654, new_n12653);
nor_4  g12279(new_n12656, new_n3930, new_n3896);
nor_4  g12280(new_n12657, new_n3939, new_n3931);
nor_4  g12281(new_n12658, new_n12657, new_n12656);
not_3  g12282(new_n12659, new_n3949);
nor_4  g12283(new_n12660, new_n3954, new_n12659);
not_3  g12284(new_n12661, new_n3955);
nor_4  g12285(new_n12662, new_n3966, new_n12661);
nor_4  g12286(new_n12663, new_n12662, new_n12660);
nand_4 g12287(new_n12664, new_n3381, new_n3380);
not_3  g12288(new_n12665, new_n3378);
nand_4 g12289(new_n12666, new_n3383, new_n12665);
nand_4 g12290(new_n12667, new_n12666, new_n12664);
nand_4 g12291(new_n12668, new_n3927, new_n3925);
nand_4 g12292(new_n12669, new_n3929, new_n3922);
nand_4 g12293(new_n12670, new_n12669, new_n12668);
nand_4 g12294(new_n12671, new_n3910, new_n3908);
not_3  g12295(new_n12672, new_n3920);
nand_4 g12296(new_n12673, new_n12672, new_n3911);
nand_4 g12297(new_n12674, new_n12673, new_n12671);
nand_4 g12298(new_n12675, n5283, n503);
not_3  g12299(new_n12676, new_n12675);
not_3  g12300(new_n12677, new_n3899);
nor_4  g12301(new_n12678, new_n3901, new_n12677);
nor_4  g12302(new_n12679, new_n3902, new_n3898);
nor_4  g12303(new_n12680, new_n12679, new_n12678);
xnor_3 g12304(new_n12681, new_n12680, new_n12676);
xnor_3 g12305(new_n12682, new_n12681, new_n12674);
nor_4  g12306(new_n12683, new_n3958, new_n3957);
not_3  g12307(new_n12684, new_n3959);
nor_4  g12308(new_n12685, new_n3965, new_n12684);
nor_4  g12309(new_n12686, new_n12685, new_n12683);
not_3  g12310(new_n12687, new_n3945);
nor_4  g12311(new_n12688, new_n3947, new_n12687);
not_3  g12312(new_n12689, new_n3944);
nor_4  g12313(new_n12690, new_n3948, new_n12689);
nor_4  g12314(new_n12691, new_n12690, new_n12688);
nand_4 g12315(new_n12692, n5198, n217);
not_3  g12316(new_n12693, new_n12692);
nand_4 g12317(new_n12694, n11296, n3992);
nand_4 g12318(new_n12695, n6611, n6358);
xor_3  g12319(new_n12696, new_n12695, new_n12694);
xnor_3 g12320(new_n12697, new_n12696, new_n12693);
xnor_3 g12321(new_n12698, new_n12697, new_n12691);
xnor_3 g12322(new_n12699, new_n12698, new_n12686);
nand_4 g12323(new_n12700, n4970, n137);
nand_4 g12324(new_n12701, n6797, n4826);
nand_4 g12325(new_n12702, n7610, n6294);
xor_3  g12326(new_n12703, new_n12702, new_n12701);
xnor_3 g12327(new_n12704_1, new_n12703, new_n12700);
nor_4  g12328(new_n12705_1, new_n3963, new_n3962);
nand_4 g12329(new_n12706_1, new_n3963, new_n3962);
nand_4 g12330(new_n12707, new_n12706_1, new_n3961);
not_3  g12331(new_n12708, new_n12707);
nor_4  g12332(new_n12709_1, new_n12708, new_n12705_1);
xnor_3 g12333(new_n12710, new_n12709_1, new_n12704_1);
nand_4 g12334(new_n12711, n11478, n10965);
not_3  g12335(new_n12712, new_n12711);
nand_4 g12336(new_n12713, n11536, n7862);
nand_4 g12337(new_n12714, n9956, n6826);
xor_3  g12338(new_n12715, new_n12714, new_n12713);
xnor_3 g12339(new_n12716, new_n12715, new_n12712);
nand_4 g12340(new_n12717, n8384, n6359);
nand_4 g12341(new_n12718, n7733, n3146);
xor_3  g12342(new_n12719, new_n12718, new_n12717);
nand_4 g12343(new_n12720_1, n12925, n4938);
nand_4 g12344(new_n12721, n7546, n4805);
xor_3  g12345(new_n12722, new_n12721, new_n12720_1);
xnor_3 g12346(new_n12723, new_n12722, new_n12719);
xnor_3 g12347(new_n12724, new_n12723, new_n12716);
xnor_3 g12348(new_n12725, new_n12724, new_n12710);
xnor_3 g12349(new_n12726, new_n12725, new_n12699);
xnor_3 g12350(new_n12727, new_n12726, new_n12682);
xnor_3 g12351(new_n12728, new_n12727, new_n12670);
xnor_3 g12352(new_n12729, new_n12728, new_n12667);
xnor_3 g12353(new_n12730, new_n12729, new_n12663);
xnor_3 g12354(new_n12731, new_n12730, new_n12658);
not_3  g12355(new_n12732, new_n12731);
xnor_3 g12356(new_n12733, new_n12732, new_n12655);
nand_4 g12357(new_n12734, new_n12733, new_n12651);
xnor_3 g12358(new_n12735, new_n12554, new_n12537);
xnor_3 g12359(new_n12736, new_n12650, new_n12735);
xnor_3 g12360(new_n12737, new_n12731, new_n12655);
nand_4 g12361(new_n12738, new_n12737, new_n12736);
nand_4 g12362(new_n12739, new_n12738, new_n12734);
xnor_3 g12363(n5257, new_n12739, new_n12534);
not_3  g12364(new_n12741, new_n11956);
xor_3  g12365(n5411, new_n12741, new_n11943);
xor_3  g12366(n5435, new_n3832, new_n3823);
xor_3  g12367(n5641, new_n6535, new_n6528);
not_3  g12368(new_n12745, new_n9129);
xor_3  g12369(n5670, new_n9139, new_n12745);
not_3  g12370(new_n12747, new_n5275);
xor_3  g12371(n5693, new_n12747, new_n5240_1);
not_3  g12372(new_n12749, new_n1411);
xor_3  g12373(n5934, new_n1424, new_n12749);
not_3  g12374(new_n12751, new_n11958);
xor_3  g12375(n6089, new_n11961, new_n12751);
not_3  g12376(new_n12753_1, new_n8290);
nand_4 g12377(new_n12754, new_n8292, new_n12753_1);
nor_4  g12378(new_n12755, new_n8271, new_n8267);
not_3  g12379(new_n12756, new_n12755);
nand_4 g12380(new_n12757, new_n8278, new_n8272);
nand_4 g12381(new_n12758, new_n12757, new_n12756);
nand_4 g12382(new_n12759, n2564, n2253);
nand_4 g12383(new_n12760, n9195, n4189);
nand_4 g12384(new_n12761, n6687, n3865);
nand_4 g12385(new_n12762, new_n12761, new_n12760);
not_3  g12386(new_n12763, new_n12760);
not_3  g12387(new_n12764, new_n12761);
nand_4 g12388(new_n12765, new_n12764, new_n12763);
nand_4 g12389(new_n12766, new_n12765, new_n12762);
xnor_3 g12390(new_n12767, new_n12766, new_n12759);
xnor_3 g12391(new_n12768, new_n12767, new_n12758);
not_3  g12392(new_n12769, new_n12768);
nor_4  g12393(new_n12770, new_n8270, new_n8269);
nand_4 g12394(new_n12771, n6770, n4634);
xor_3  g12395(new_n12772, new_n12771, new_n12770);
nand_4 g12396(new_n12773, n3627, n2879);
not_3  g12397(new_n12774, new_n12773);
nand_4 g12398(new_n12775, n10223, n9920);
nand_4 g12399(new_n12776, n7265, n4516);
xnor_3 g12400(new_n12777_1, new_n12776, new_n12775);
xnor_3 g12401(new_n12778, new_n12777_1, new_n12774);
not_3  g12402(new_n12779, new_n12778);
xnor_3 g12403(new_n12780, new_n12779, new_n12772);
not_3  g12404(new_n12781, new_n12780);
xor_3  g12405(new_n12782, new_n12781, new_n12769);
nand_4 g12406(new_n12783, new_n8283, new_n8280);
nor_4  g12407(new_n12784, new_n8282, new_n8281);
nor_4  g12408(new_n12785, new_n8289, new_n8285);
xnor_3 g12409(new_n12786, new_n12785, new_n12784);
nand_4 g12410(new_n12787, new_n12786, new_n12783);
xnor_3 g12411(new_n12788, new_n12787, new_n12782);
xnor_3 g12412(new_n12789, new_n12788, new_n12754);
nor_4  g12413(new_n12790, new_n8293, new_n8266);
nor_4  g12414(new_n12791, new_n8294, new_n8264);
nor_4  g12415(new_n12792, new_n12791, new_n12790);
xnor_3 g12416(new_n12793, new_n12792, new_n12789);
nand_4 g12417(new_n12794, new_n8337, new_n8303_1);
xnor_3 g12418(new_n12795, new_n8337, new_n8302);
nand_4 g12419(new_n12796, new_n12795, new_n8301);
nand_4 g12420(new_n12797, new_n12796, new_n12794);
not_3  g12421(new_n12798, new_n8308);
nand_4 g12422(new_n12799, new_n8317, new_n8312);
nand_4 g12423(new_n12800, new_n12799, new_n12798);
nand_4 g12424(new_n12801, n12221, n10928);
nand_4 g12425(new_n12802, n12145, n6986);
nand_4 g12426(new_n12803, n10217, n8336);
xnor_3 g12427(new_n12804, new_n12803, new_n12802);
xnor_3 g12428(new_n12805, new_n12804, new_n12801);
xnor_3 g12429(new_n12806, new_n12805, new_n12800);
nor_4  g12430(new_n12807_1, new_n8306, new_n8305);
nand_4 g12431(new_n12808, n2522, n2226);
xor_3  g12432(new_n12809, new_n12808, new_n12807_1);
nand_4 g12433(new_n12810, n10678, n2024);
not_3  g12434(new_n12811, new_n12810);
nand_4 g12435(new_n12812, n9189, n1094);
nand_4 g12436(new_n12813, n7946, n7320);
xnor_3 g12437(new_n12814, new_n12813, new_n12812);
and_4  g12438(new_n12815, new_n12814, new_n12811);
nor_4  g12439(new_n12816, new_n12814, new_n12811);
nor_4  g12440(new_n12817, new_n12816, new_n12815);
xnor_3 g12441(new_n12818, new_n12817, new_n12809);
not_3  g12442(new_n12819, new_n12818);
xor_3  g12443(new_n12820, new_n12819, new_n12806);
not_3  g12444(new_n12821, new_n12820);
nand_4 g12445(new_n12822, new_n8322, new_n8319);
nor_4  g12446(new_n12823, new_n8321, new_n8320);
nor_4  g12447(new_n12824, new_n8328, new_n8324);
xnor_3 g12448(new_n12825, new_n12824, new_n12823);
nand_4 g12449(new_n12826_1, new_n12825, new_n12822);
xnor_3 g12450(new_n12827, new_n12826_1, new_n12821);
xnor_3 g12451(new_n12828, new_n12827, new_n8334);
xnor_3 g12452(new_n12829, new_n12828, new_n12797);
nor_4  g12453(new_n12830, new_n8372, new_n8369);
nor_4  g12454(new_n12831, new_n8358, new_n8357);
nand_4 g12455(new_n12832, n7160, n521);
not_3  g12456(new_n12833, new_n12832);
xor_3  g12457(new_n12834, new_n12833, new_n12831);
nand_4 g12458(new_n12835, n2515, n2498);
nand_4 g12459(new_n12836, n2558, n1199);
nand_4 g12460(new_n12837, n5579, n4828);
not_3  g12461(new_n12838, new_n12837);
xor_3  g12462(new_n12839, new_n12838, new_n12836);
xnor_3 g12463(new_n12840, new_n12839, new_n12835);
not_3  g12464(new_n12841, new_n12840);
nand_4 g12465(new_n12842, new_n12841, new_n12834);
not_3  g12466(new_n12843, new_n12842);
nor_4  g12467(new_n12844, new_n12841, new_n12834);
nor_4  g12468(new_n12845, new_n12844, new_n12843);
not_3  g12469(new_n12846, new_n8355);
nand_4 g12470(new_n12847, new_n8359, new_n8356);
nand_4 g12471(new_n12848, new_n12847, new_n12846);
nand_4 g12472(new_n12849, n12391, n5798);
nand_4 g12473(new_n12850, n7891, n6016);
nand_4 g12474(new_n12851, n12069, n2347);
not_3  g12475(new_n12852, new_n12851);
xor_3  g12476(new_n12853, new_n12852, new_n12850);
xnor_3 g12477(new_n12854, new_n12853, new_n12849);
xnor_3 g12478(new_n12855, new_n12854, new_n12848);
xnor_3 g12479(new_n12856, new_n12855, new_n12845);
not_3  g12480(new_n12857, new_n8360);
not_3  g12481(new_n12858, new_n8364);
nand_4 g12482(new_n12859, new_n12858, new_n12857);
nor_4  g12483(new_n12860, new_n8362, new_n8361);
nor_4  g12484(new_n12861, new_n8368, new_n8365);
xnor_3 g12485(new_n12862, new_n12861, new_n12860);
nand_4 g12486(new_n12863, new_n12862, new_n12859);
xnor_3 g12487(new_n12864, new_n12863, new_n12856);
xnor_3 g12488(new_n12865, new_n12864, new_n12830);
nor_4  g12489(new_n12866, new_n8373, new_n8349);
nor_4  g12490(new_n12867, new_n8374, new_n8348);
nor_4  g12491(new_n12868, new_n12867, new_n12866);
xnor_3 g12492(new_n12869, new_n12868, new_n12865);
nor_4  g12493(new_n12870, new_n8402, new_n8398_1);
not_3  g12494(new_n12871, new_n12870);
nand_4 g12495(new_n12872, new_n8388, new_n8386);
not_3  g12496(new_n12873, new_n12872);
nor_4  g12497(new_n12874, new_n12873, new_n8382);
not_3  g12498(new_n12875, new_n12874);
nand_4 g12499(new_n12876, n11153, n5153);
nand_4 g12500(new_n12877, n7270, n5314);
nand_4 g12501(new_n12878, n11222, n2507);
not_3  g12502(new_n12879, new_n12878);
xor_3  g12503(new_n12880, new_n12879, new_n12877);
xnor_3 g12504(new_n12881, new_n12880, new_n12876);
xnor_3 g12505(new_n12882, new_n12881, new_n12875);
nor_4  g12506(new_n12883, new_n8380, new_n8379);
not_3  g12507(new_n12884, new_n12883);
nand_4 g12508(new_n12885, n996, n806);
xor_3  g12509(new_n12886, new_n12885, new_n12884);
nand_4 g12510(new_n12887, n9111, n5319);
nand_4 g12511(new_n12888, n5767, n3342);
nand_4 g12512(new_n12889, n9763, n9457);
not_3  g12513(new_n12890, new_n12889);
xor_3  g12514(new_n12891, new_n12890, new_n12888);
xnor_3 g12515(new_n12892, new_n12891, new_n12887);
xnor_3 g12516(new_n12893, new_n12892, new_n12886);
xnor_3 g12517(new_n12894, new_n12893, new_n12882);
nand_4 g12518(new_n12895, new_n8393, new_n8390);
nor_4  g12519(new_n12896, new_n8392, new_n8391);
nor_4  g12520(new_n12897, new_n8397, new_n8394);
xnor_3 g12521(new_n12898, new_n12897, new_n12896);
nand_4 g12522(new_n12899, new_n12898, new_n12895);
xnor_3 g12523(new_n12900, new_n12899, new_n12894);
xnor_3 g12524(new_n12901, new_n12900, new_n12871);
not_3  g12525(new_n12902, new_n8377);
not_3  g12526(new_n12903, new_n8403);
nor_4  g12527(new_n12904, new_n12903, new_n12902);
nor_4  g12528(new_n12905, new_n8407, new_n12904);
xnor_3 g12529(new_n12906, new_n12905, new_n12901);
xnor_3 g12530(new_n12907, new_n12906, new_n12869);
nand_4 g12531(new_n12908, new_n8416, new_n8409);
nand_4 g12532(new_n12909, new_n12908, new_n8412);
xnor_3 g12533(new_n12910, new_n12909, new_n12907);
xnor_3 g12534(new_n12911, new_n12910, new_n12829);
nand_4 g12535(new_n12912, new_n8344, new_n8339);
nor_4  g12536(new_n12913, new_n8344, new_n8339);
not_3  g12537(new_n12914, new_n12912);
nor_4  g12538(new_n12915, new_n12914, new_n12913);
nand_4 g12539(new_n12916, new_n8417, new_n12915);
nand_4 g12540(new_n12917, new_n12916, new_n12912);
xnor_3 g12541(new_n12918, new_n12917, new_n12911);
not_3  g12542(new_n12919, new_n12918);
nand_4 g12543(new_n12920, new_n12919, new_n12793);
not_3  g12544(new_n12921, new_n12793);
nand_4 g12545(new_n12922, new_n12918, new_n12921);
nor_4  g12546(new_n12923, new_n8299, new_n8295);
nor_4  g12547(new_n12924, new_n8420, new_n12923);
nand_4 g12548(new_n12925_1, new_n12924, new_n12922);
nand_4 g12549(new_n12926, new_n12925_1, new_n12920);
nor_4  g12550(new_n12927, new_n12910, new_n12829);
nor_4  g12551(new_n12928, new_n12917, new_n12911);
nor_4  g12552(new_n12929, new_n12928, new_n12927);
not_3  g12553(new_n12930, new_n12869);
not_3  g12554(new_n12931, new_n12906);
nand_4 g12555(new_n12932, new_n12931, new_n12930);
nand_4 g12556(new_n12933, new_n12906, new_n12869);
nand_4 g12557(new_n12934, new_n12909, new_n12933);
nand_4 g12558(new_n12935, new_n12934, new_n12932);
nand_4 g12559(new_n12936, new_n12861, new_n12860);
not_3  g12560(new_n12937, new_n12856);
nand_4 g12561(new_n12938, new_n12863, new_n12937);
nand_4 g12562(new_n12939, new_n12938, new_n12936);
nand_4 g12563(new_n12940, new_n12785, new_n12784);
not_3  g12564(new_n12941, new_n12782);
nand_4 g12565(new_n12942, new_n12787, new_n12941);
nand_4 g12566(new_n12943, new_n12942, new_n12940);
nand_4 g12567(new_n12944, n5579, n2515);
nand_4 g12568(new_n12945, n4828, n521);
not_3  g12569(new_n12946, new_n12945);
xor_3  g12570(new_n12947_1, new_n12946, new_n12944);
nor_4  g12571(new_n12948, new_n12837, new_n12836);
not_3  g12572(new_n12949, new_n12835);
nand_4 g12573(new_n12950, new_n12837, new_n12836);
nand_4 g12574(new_n12951, new_n12950, new_n12949);
not_3  g12575(new_n12952, new_n12951);
nor_4  g12576(new_n12953, new_n12952, new_n12948);
nand_4 g12577(new_n12954, n7891, n5798);
nand_4 g12578(new_n12955, n12391, n2347);
xor_3  g12579(new_n12956, new_n12955, new_n12954);
nand_4 g12580(new_n12957, n6687, n2512);
nand_4 g12581(new_n12958, n7265, n2087);
xor_3  g12582(new_n12959, new_n12958, new_n12957);
xnor_3 g12583(new_n12960, new_n12959, new_n12956);
xnor_3 g12584(new_n12961, new_n12960, new_n12953);
xnor_3 g12585(new_n12962, new_n12961, new_n12947_1);
nand_4 g12586(new_n12963, n2498, n1199);
nand_4 g12587(new_n12964, new_n12833, new_n12831);
nand_4 g12588(new_n12965, new_n12842, new_n12964);
xor_3  g12589(new_n12966, new_n12965, new_n12963);
xnor_3 g12590(new_n12967, new_n12966, new_n12962);
xnor_3 g12591(new_n12968, new_n12967, new_n12943);
xnor_3 g12592(new_n12969, new_n12968, new_n12939);
xnor_3 g12593(new_n12970, new_n12969, new_n12935);
nand_4 g12594(new_n12971, new_n12864, new_n12830);
nor_4  g12595(new_n12972, new_n12868, new_n12865);
not_3  g12596(new_n12973, new_n12972);
nand_4 g12597(new_n12974, new_n12973, new_n12971);
nand_4 g12598(new_n12975, new_n12900, new_n12870);
nand_4 g12599(new_n12976, new_n12905, new_n12901);
nand_4 g12600(new_n12977, new_n12976, new_n12975);
nand_4 g12601(new_n12978, new_n12897, new_n12896);
not_3  g12602(new_n12979, new_n12894);
nand_4 g12603(new_n12980, new_n12899, new_n12979);
nand_4 g12604(new_n12981, new_n12980, new_n12978);
not_3  g12605(new_n12982, new_n12807_1);
nand_4 g12606(new_n12983, new_n12808, new_n12982);
not_3  g12607(new_n12984, new_n12809);
nand_4 g12608(new_n12985, new_n12817, new_n12984);
nand_4 g12609(new_n12986, new_n12985, new_n12983);
nand_4 g12610(new_n12987, n9457, n9111);
nand_4 g12611(new_n12988, n10678, n9189);
nand_4 g12612(new_n12989, n11222, n6431);
xor_3  g12613(new_n12990, new_n12989, new_n12988);
xnor_3 g12614(new_n12991, new_n12990, new_n12987);
xnor_3 g12615(new_n12992, new_n12991, new_n12986);
nand_4 g12616(new_n12993, n12145, n2226);
nand_4 g12617(new_n12994, n9763, n4817);
nand_4 g12618(new_n12995, n5319, n3342);
xor_3  g12619(new_n12996, new_n12995, new_n12994);
nand_4 g12620(new_n12997, n12221, n6986);
nand_4 g12621(new_n12998, n2522, n1094);
xor_3  g12622(new_n12999, new_n12998, new_n12997);
xnor_3 g12623(new_n13000, new_n12999, new_n12996);
xnor_3 g12624(new_n13001, new_n13000, new_n12993);
nand_4 g12625(new_n13002, n10928, n10217);
not_3  g12626(new_n13003, new_n12812);
not_3  g12627(new_n13004, new_n12813);
nor_4  g12628(new_n13005, new_n13004, new_n13003);
nor_4  g12629(new_n13006, new_n12816, new_n13005);
xor_3  g12630(new_n13007, new_n13006, new_n13002);
xnor_3 g12631(new_n13008, new_n13007, new_n13001);
xnor_3 g12632(new_n13009, new_n13008, new_n12992);
xnor_3 g12633(new_n13010, new_n13009, new_n12981);
nor_4  g12634(new_n13011, new_n12885, new_n12884);
not_3  g12635(new_n13012, new_n12886);
nor_4  g12636(new_n13013, new_n12892, new_n13012);
nor_4  g12637(new_n13014, new_n13013, new_n13011);
not_3  g12638(new_n13015, new_n12888);
nor_4  g12639(new_n13016, new_n12890, new_n13015);
not_3  g12640(new_n13017, new_n12887);
nor_4  g12641(new_n13018, new_n12891, new_n13017);
nor_4  g12642(new_n13019, new_n13018, new_n13016);
nand_4 g12643(new_n13020, n11153, n2507);
nand_4 g12644(new_n13021, n5314, n5153);
not_3  g12645(new_n13022, new_n13021);
xor_3  g12646(new_n13023, new_n13022, new_n13020);
xnor_3 g12647(new_n13024, new_n13023, new_n13019);
xnor_3 g12648(new_n13025, new_n13024, new_n13014);
nand_4 g12649(new_n13026, n7946, n7523);
nand_4 g12650(new_n13027, n9920, n4634);
xor_3  g12651(new_n13028, new_n13027, new_n13026);
nand_4 g12652(new_n13029, n8336, n7823);
nand_4 g12653(new_n13030, n7320, n2024);
xor_3  g12654(new_n13031, new_n13030, new_n13029);
xnor_3 g12655(new_n13032, new_n13031, new_n13028);
not_3  g12656(new_n13033, new_n12759);
nand_4 g12657(new_n13034, new_n12762, new_n13033);
and_4  g12658(new_n13035, new_n13034, new_n12765);
nand_4 g12659(new_n13036, n10223, n3627);
nand_4 g12660(new_n13037, n4516, n2879);
xor_3  g12661(new_n13038, new_n13037, new_n13036);
xnor_3 g12662(new_n13039, new_n13038, new_n13035);
xnor_3 g12663(new_n13040, new_n13039, new_n13032);
xnor_3 g12664(new_n13041, new_n13040, new_n13025);
not_3  g12665(new_n13042, new_n12758);
nand_4 g12666(new_n13043, new_n12767, new_n13042);
nand_4 g12667(new_n13044, new_n12780, new_n12768);
nand_4 g12668(new_n13045, new_n13044, new_n13043);
not_3  g12669(new_n13046, new_n12771);
nor_4  g12670(new_n13047, new_n13046, new_n12770);
nor_4  g12671(new_n13048, new_n12778, new_n12772);
nor_4  g12672(new_n13049, new_n13048, new_n13047);
nand_4 g12673(new_n13050, n6578, n2558);
and_4  g12674(new_n13051, new_n12776, new_n12775);
nor_4  g12675(new_n13052, new_n12777_1, new_n12774);
nor_4  g12676(new_n13053, new_n13052, new_n13051);
nand_4 g12677(new_n13054, n9195, n6770);
nand_4 g12678(new_n13055, n4189, n2253);
nand_4 g12679(new_n13056, n3865, n2564);
xnor_3 g12680(new_n13057, new_n13056, new_n13055);
xnor_3 g12681(new_n13058, new_n13057, new_n13054);
xnor_3 g12682(new_n13059, new_n13058, new_n13053);
xnor_3 g12683(new_n13060, new_n13059, new_n13050);
xnor_3 g12684(new_n13061, new_n13060, new_n13049);
xnor_3 g12685(new_n13062, new_n13061, new_n13045);
not_3  g12686(new_n13063, new_n12800);
nand_4 g12687(new_n13064, new_n12805, new_n13063);
nand_4 g12688(new_n13065, new_n12818, new_n12806);
nand_4 g12689(new_n13066, new_n13065, new_n13064);
nor_4  g12690(new_n13067, new_n12803, new_n12802);
not_3  g12691(new_n13068, new_n12801);
nand_4 g12692(new_n13069, new_n12803, new_n12802);
nand_4 g12693(new_n13070, new_n13069, new_n13068);
not_3  g12694(new_n13071, new_n13070);
nor_4  g12695(new_n13072, new_n13071, new_n13067);
xnor_3 g12696(new_n13073, new_n13072, new_n13066);
xnor_3 g12697(new_n13074, new_n13073, new_n13062);
xnor_3 g12698(new_n13075, new_n13074, new_n13041);
xnor_3 g12699(new_n13076, new_n13075, new_n13010);
xnor_3 g12700(new_n13077, new_n13076, new_n12977);
xnor_3 g12701(new_n13078, new_n13077, new_n12974);
not_3  g12702(new_n13079, new_n12754);
nand_4 g12703(new_n13080, new_n12788, new_n13079);
nand_4 g12704(new_n13081, new_n12792, new_n12789);
nand_4 g12705(new_n13082, new_n13081, new_n13080);
nand_4 g12706(new_n13083, new_n12824, new_n12823);
nand_4 g12707(new_n13084, new_n12826_1, new_n12820);
nand_4 g12708(new_n13085, new_n13084, new_n13083);
nand_4 g12709(new_n13086, new_n12881, new_n12874);
not_3  g12710(new_n13087, new_n12893);
nand_4 g12711(new_n13088, new_n13087, new_n12882);
nand_4 g12712(new_n13089, new_n13088, new_n13086);
not_3  g12713(new_n13090, new_n12877);
nor_4  g12714(new_n13091, new_n12879, new_n13090);
not_3  g12715(new_n13092, new_n12876);
nor_4  g12716(new_n13093, new_n12880, new_n13092);
nor_4  g12717(new_n13094, new_n13093, new_n13091);
nand_4 g12718(new_n13095, n12069, n1576);
nand_4 g12719(new_n13096, n7270, n996);
nand_4 g12720(new_n13097, n5767, n806);
xor_3  g12721(new_n13098, new_n13097, new_n13096);
xor_3  g12722(new_n13099, new_n13098, new_n13095);
xnor_3 g12723(new_n13100, new_n13099, new_n13094);
xnor_3 g12724(new_n13101, new_n13100, new_n13089);
xnor_3 g12725(new_n13102, new_n13101, new_n13085);
xnor_3 g12726(new_n13103, new_n13102, new_n13082);
xnor_3 g12727(new_n13104, new_n13103, new_n13078);
xnor_3 g12728(new_n13105, new_n13104, new_n12970);
nand_4 g12729(new_n13106, new_n12827, new_n8334);
not_3  g12730(new_n13107, new_n12828);
nand_4 g12731(new_n13108, new_n13107, new_n12797);
nand_4 g12732(new_n13109, new_n13108, new_n13106);
not_3  g12733(new_n13110, new_n12848);
nand_4 g12734(new_n13111, new_n12854, new_n13110);
not_3  g12735(new_n13112, new_n12845);
nand_4 g12736(new_n13113, new_n12855, new_n13112);
nand_4 g12737(new_n13114, new_n13113, new_n13111);
nand_4 g12738(new_n13115, n7160, n6016);
not_3  g12739(new_n13116, new_n12850);
nor_4  g12740(new_n13117, new_n12852, new_n13116);
not_3  g12741(new_n13118, new_n12849);
nor_4  g12742(new_n13119, new_n12853, new_n13118);
nor_4  g12743(new_n13120, new_n13119, new_n13117);
xor_3  g12744(new_n13121, new_n13120, new_n13115);
xor_3  g12745(new_n13122, new_n13121, new_n13114);
xnor_3 g12746(new_n13123, new_n13122, new_n13109);
xnor_3 g12747(new_n13124, new_n13123, new_n13105);
xnor_3 g12748(new_n13125, new_n13124, new_n12929);
xnor_3 g12749(n6192, new_n13125, new_n12926);
xor_3  g12750(n6273, new_n1060, new_n1024);
xnor_3 g12751(n6445, new_n8246, new_n8245);
nand_4 g12752(new_n13129, new_n9999, new_n9998);
xnor_3 g12753(n6645, new_n13129, new_n10025);
not_3  g12754(new_n13131, new_n8472);
xor_3  g12755(n6689, new_n8475, new_n13131);
xor_3  g12756(n6742, new_n1412, new_n1320);
not_3  g12757(new_n13134, new_n2154);
xnor_3 g12758(n6809, new_n2195, new_n13134);
not_3  g12759(new_n13136, new_n7257);
xor_3  g12760(n6822, new_n7259, new_n13136);
not_3  g12761(new_n13138, new_n11954);
xor_3  g12762(n6860, new_n13138, new_n11953);
not_3  g12763(new_n13140, new_n10013);
xor_3  g12764(n7193, new_n10021, new_n13140);
nand_4 g12765(new_n13142, new_n8237, new_n8236_1);
xnor_3 g12766(n7568, new_n13142, new_n8248);
not_3  g12767(new_n13144, new_n1422);
xor_3  g12768(n7676, new_n13144, new_n1421);
nand_4 g12769(new_n13146, new_n471, new_n464);
not_3  g12770(new_n13147, new_n483);
nand_4 g12771(new_n13148, new_n13147, new_n472);
nand_4 g12772(new_n13149, new_n13148, new_n13146);
nand_4 g12773(new_n13150, n10644, n7354);
xor_3  g12774(new_n13151, new_n13150, new_n13149);
nand_4 g12775(new_n13152, new_n969, new_n959);
nand_4 g12776(new_n13153, new_n982, new_n970);
nand_4 g12777(new_n13154, new_n13153, new_n13152);
not_3  g12778(new_n13155, new_n977);
nor_4  g12779(new_n13156, new_n979, new_n13155);
nor_4  g12780(new_n13157, new_n980, new_n976);
nor_4  g12781(new_n13158, new_n13157, new_n13156);
xnor_3 g12782(new_n13159, new_n13158, new_n13154);
xnor_3 g12783(new_n13160, new_n13159, new_n13151);
nor_4  g12784(new_n13161, new_n475, new_n474);
not_3  g12785(new_n13162, new_n476);
nor_4  g12786(new_n13163, new_n482, new_n13162);
nor_4  g12787(new_n13164, new_n13163, new_n13161);
nand_4 g12788(new_n13165, n3986, n1980);
not_3  g12789(new_n13166, new_n13165);
nor_4  g12790(new_n13167, new_n480, new_n479);
nand_4 g12791(new_n13168, new_n480, new_n479);
nand_4 g12792(new_n13169, new_n13168, new_n478);
not_3  g12793(new_n13170, new_n13169);
nor_4  g12794(new_n13171, new_n13170, new_n13167);
nand_4 g12795(new_n13172, n7436, n4141);
nand_4 g12796(new_n13173, n9241, n1209);
not_3  g12797(new_n13174, new_n13173);
xor_3  g12798(new_n13175, new_n13174, new_n13172);
nand_4 g12799(new_n13176, n8276, n5105);
nand_4 g12800(new_n13177, n8236, n6776);
xor_3  g12801(new_n13178, new_n13177, new_n13176);
xor_3  g12802(new_n13179, new_n13178, new_n13175);
xnor_3 g12803(new_n13180, new_n13179, new_n13171);
xnor_3 g12804(new_n13181, new_n13180, new_n13166);
xnor_3 g12805(new_n13182, new_n13181, new_n13164);
or_4   g12806(new_n13183, new_n489, new_n488);
not_3  g12807(new_n13184, new_n484);
nand_4 g12808(new_n13185, new_n491, new_n13184);
nand_4 g12809(new_n13186, new_n13185, new_n13183);
xnor_3 g12810(new_n13187, new_n13186, new_n13182);
xnor_3 g12811(new_n13188, new_n13187, new_n13160);
nand_4 g12812(new_n13189, new_n620, new_n586);
not_3  g12813(new_n13190, new_n642);
nand_4 g12814(new_n13191, new_n13190, new_n621);
nand_4 g12815(new_n13192, new_n13191, new_n13189);
nand_4 g12816(new_n13193, new_n751, new_n719);
not_3  g12817(new_n13194, new_n752);
nand_4 g12818(new_n13195, new_n773, new_n13194);
nand_4 g12819(new_n13196, new_n13195, new_n13193);
nand_4 g12820(new_n13197, n12706, n5964);
nand_4 g12821(new_n13198, n4005, n1097);
xor_3  g12822(new_n13199, new_n13198, new_n13197);
nand_4 g12823(new_n13200, n12720, n12025);
nand_4 g12824(new_n13201, n11257, n2509);
xor_3  g12825(new_n13202, new_n13201, new_n13200);
xor_3  g12826(new_n13203, new_n13202, new_n13199);
nand_4 g12827(new_n13204, n12705, n2508);
not_3  g12828(new_n13205, new_n961);
nand_4 g12829(new_n13206, new_n964, new_n13205);
and_4  g12830(new_n13207, new_n13206, new_n967);
xor_3  g12831(new_n13208, new_n13207, new_n13204);
xnor_3 g12832(new_n13209, new_n13208, new_n13203);
xnor_3 g12833(new_n13210, new_n13209, new_n13196);
xnor_3 g12834(new_n13211, new_n13210, new_n13192);
nand_4 g12835(new_n13212, new_n617, new_n615_1);
not_3  g12836(new_n13213, new_n612);
nand_4 g12837(new_n13214, new_n619, new_n13213);
nand_4 g12838(new_n13215, new_n13214, new_n13212);
not_3  g12839(new_n13216, new_n985);
nor_4  g12840(new_n13217, new_n986, new_n13216);
nor_4  g12841(new_n13218, new_n988, new_n984);
nor_4  g12842(new_n13219, new_n13218, new_n13217);
xnor_3 g12843(new_n13220, new_n13219, new_n13215);
nand_4 g12844(new_n13221, n12704, n2393);
not_3  g12845(new_n13222, new_n732);
nor_4  g12846(new_n13223, new_n743, new_n13222);
nor_4  g12847(new_n13224, new_n13223, new_n731);
not_3  g12848(new_n13225, new_n724);
nor_4  g12849(new_n13226, new_n726, new_n13225);
not_3  g12850(new_n13227, new_n723);
nor_4  g12851(new_n13228, new_n727, new_n13227);
nor_4  g12852(new_n13229, new_n13228, new_n13226);
nand_4 g12853(new_n13230, n4499, n1564);
nand_4 g12854(new_n13231, n12648, n6806);
xor_3  g12855(new_n13232, new_n13231, new_n13230);
nand_4 g12856(new_n13233, n10547, n6038);
nand_4 g12857(new_n13234, n5069, n2530);
xor_3  g12858(new_n13235, new_n13234, new_n13233);
xnor_3 g12859(new_n13236, new_n13235, new_n13232);
xnor_3 g12860(new_n13237, new_n13236, new_n13229);
nand_4 g12861(new_n13238, n5694, n5331);
nand_4 g12862(new_n13239, n7388, n4903);
not_3  g12863(new_n13240, new_n13239);
xor_3  g12864(new_n13241, new_n13240, new_n13238);
xnor_3 g12865(new_n13242, new_n13241, new_n13237);
nor_4  g12866(new_n13243, new_n735, new_n734);
not_3  g12867(new_n13244, new_n736);
nor_4  g12868(new_n13245, new_n742, new_n13244);
nor_4  g12869(new_n13246, new_n13245, new_n13243);
not_3  g12870(new_n13247, new_n738);
nor_4  g12871(new_n13248, new_n740, new_n13247);
not_3  g12872(new_n13249, new_n737);
nor_4  g12873(new_n13250, new_n741, new_n13249);
nor_4  g12874(new_n13251, new_n13250, new_n13248);
nand_4 g12875(new_n13252, n7294, n5860);
nand_4 g12876(new_n13253, n11892, n5814);
xor_3  g12877(new_n13254, new_n13253, new_n13252);
xnor_3 g12878(new_n13255, new_n13254, new_n13251);
xnor_3 g12879(new_n13256, new_n13255, new_n13246);
xnor_3 g12880(new_n13257, new_n13256, new_n13242);
xnor_3 g12881(new_n13258, new_n13257, new_n13224);
xnor_3 g12882(new_n13259, new_n13258, new_n13221);
and_4  g12883(new_n13260, new_n748, new_n747);
not_3  g12884(new_n13261, new_n750);
nor_4  g12885(new_n13262, new_n13261, new_n744);
nor_4  g12886(new_n13263, new_n13262, new_n13260);
nand_4 g12887(new_n13264, new_n597, new_n590);
not_3  g12888(new_n13265, new_n611);
nand_4 g12889(new_n13266, new_n13265, new_n598);
nand_4 g12890(new_n13267, new_n13266, new_n13264);
not_3  g12891(new_n13268, new_n593);
nor_4  g12892(new_n13269, new_n595, new_n13268);
not_3  g12893(new_n13270, new_n592);
nor_4  g12894(new_n13271, new_n596, new_n13270);
nor_4  g12895(new_n13272, new_n13271, new_n13269);
not_3  g12896(new_n13273, new_n606);
nor_4  g12897(new_n13274, new_n608, new_n13273);
nor_4  g12898(new_n13275, new_n609, new_n605);
nor_4  g12899(new_n13276, new_n13275, new_n13274);
xnor_3 g12900(new_n13277, new_n13276, new_n13272);
nand_4 g12901(new_n13278, n10545, n2802);
nand_4 g12902(new_n13279, n12044, n8476);
xor_3  g12903(new_n13280, new_n13279, new_n13278);
nand_4 g12904(new_n13281, n7690, n533);
nand_4 g12905(new_n13282, n3616, n1512);
xor_3  g12906(new_n13283, new_n13282, new_n13281);
xnor_3 g12907(new_n13284, new_n13283, new_n13280);
xnor_3 g12908(new_n13285, new_n13284, new_n13277);
nand_4 g12909(new_n13286, n5305, n615);
not_3  g12910(new_n13287, new_n13286);
nand_4 g12911(new_n13288, new_n601, new_n599);
nand_4 g12912(new_n13289, new_n610, new_n602);
nand_4 g12913(new_n13290, new_n13289, new_n13288);
xnor_3 g12914(new_n13291, new_n13290, new_n13287);
xnor_3 g12915(new_n13292, new_n13291, new_n13285);
xnor_3 g12916(new_n13293, new_n13292, new_n13267);
nand_4 g12917(new_n13294, n10848, n5857);
nand_4 g12918(new_n13295, n7965, n1906);
not_3  g12919(new_n13296, new_n13295);
xor_3  g12920(new_n13297, new_n13296, new_n13294);
not_3  g12921(new_n13298, new_n467);
nor_4  g12922(new_n13299, new_n469, new_n13298);
not_3  g12923(new_n13300, new_n466);
nor_4  g12924(new_n13301, new_n470, new_n13300);
nor_4  g12925(new_n13302, new_n13301, new_n13299);
nand_4 g12926(new_n13303, n8028, n45);
nand_4 g12927(new_n13304, n12299, n4928);
xor_3  g12928(new_n13305, new_n13304, new_n13303);
xnor_3 g12929(new_n13306, new_n13305, new_n13302);
xnor_3 g12930(new_n13307, new_n13306, new_n13297);
nand_4 g12931(new_n13308, new_n973, new_n971);
nand_4 g12932(new_n13309, new_n981, new_n974);
nand_4 g12933(new_n13310, new_n13309, new_n13308);
nand_4 g12934(new_n13311, n8759, n783);
nand_4 g12935(new_n13312, n10510, n7500);
xor_3  g12936(new_n13313, new_n13312, new_n13311);
xnor_3 g12937(new_n13314, new_n13313, new_n13310);
xnor_3 g12938(new_n13315, new_n13314, new_n13307);
xnor_3 g12939(new_n13316, new_n13315, new_n13293);
xnor_3 g12940(new_n13317, new_n13316, new_n13263);
xnor_3 g12941(new_n13318, new_n13317, new_n13259);
xnor_3 g12942(new_n13319, new_n13318, new_n13220);
xnor_3 g12943(new_n13320, new_n13319, new_n13211);
xnor_3 g12944(new_n13321, new_n13320, new_n13188);
nor_4  g12945(new_n13322, new_n989, new_n955);
not_3  g12946(new_n13323, new_n1010);
nor_4  g12947(new_n13324, new_n13323, new_n990);
nor_4  g12948(new_n13325, new_n13324, new_n13322);
nor_4  g12949(new_n13326, new_n774, new_n643);
nor_4  g12950(new_n13327, new_n826, new_n775);
nor_4  g12951(new_n13328, new_n13327, new_n13326);
xnor_3 g12952(new_n13329, new_n13328, new_n13325);
xnor_3 g12953(new_n13330, new_n13329, new_n13321);
not_3  g12954(new_n13331, new_n513);
nand_4 g12955(new_n13332, new_n827, new_n13331);
nand_4 g12956(new_n13333, new_n878, new_n828);
nand_4 g12957(new_n13334, new_n13333, new_n13332);
not_3  g12958(new_n13335, new_n461);
nand_4 g12959(new_n13336, new_n492, new_n13335);
nand_4 g12960(new_n13337, new_n512, new_n493);
nand_4 g12961(new_n13338, new_n13337, new_n13336);
nand_4 g12962(new_n13339, n4312, n2585);
xor_3  g12963(new_n13340, new_n13339, new_n13338);
xnor_3 g12964(new_n13341, new_n13340, new_n13334);
not_3  g12965(new_n13342, new_n1065);
nand_4 g12966(new_n13343, new_n1066, new_n879);
nand_4 g12967(new_n13344, new_n13343, new_n13342);
xnor_3 g12968(new_n13345, new_n13344, new_n13341);
xnor_3 g12969(n7966, new_n13345, new_n13330);
not_3  g12970(new_n13347, new_n12924);
nand_4 g12971(new_n13348, new_n12922, new_n12920);
xnor_3 g12972(n7981, new_n13348, new_n13347);
nand_4 g12973(new_n13350, new_n12530, new_n12512);
nand_4 g12974(new_n13351, new_n13350, new_n12511_1);
nor_4  g12975(new_n13352, new_n12521, new_n12526);
nor_4  g12976(new_n13353, new_n13352, new_n12341);
nor_4  g12977(new_n13354, new_n13353, new_n12335);
xnor_3 g12978(new_n13355, new_n13353, new_n12335);
nor_4  g12979(new_n13356, new_n12507, new_n13355);
nor_4  g12980(new_n13357, new_n13356, new_n13354);
not_3  g12981(new_n13358, new_n12215);
nand_4 g12982(new_n13359, new_n12253, new_n13358);
nand_4 g12983(new_n13360, new_n12263, new_n12254);
nand_4 g12984(new_n13361, new_n13360, new_n13359);
nand_4 g12985(new_n13362, new_n12247_1, new_n12246);
nand_4 g12986(new_n13363, new_n12251, new_n13362);
nand_4 g12987(new_n13364, n12391, n1353);
not_3  g12988(new_n13365, new_n13364);
nand_4 g12989(new_n13366, new_n12471, new_n12460);
nand_4 g12990(new_n13367, new_n12486, new_n12472);
nand_4 g12991(new_n13368, new_n13367, new_n13366);
not_3  g12992(new_n13369, new_n12473);
nor_4  g12993(new_n13370, new_n12474, new_n13369);
nor_4  g12994(new_n13371, new_n12485, new_n12475);
nor_4  g12995(new_n13372, new_n13371, new_n13370);
nand_4 g12996(new_n13373, n7891, n447);
nand_4 g12997(new_n13374, new_n12466, new_n12463);
nand_4 g12998(new_n13375, new_n13374, new_n12469);
xor_3  g12999(new_n13376, new_n13375, new_n13373);
nand_4 g13000(new_n13377, new_n12480, new_n12477);
and_4  g13001(new_n13378, new_n13377, new_n12483);
nand_4 g13002(new_n13379, n11407, n2087);
nand_4 g13003(new_n13380, n6687, n6604);
xor_3  g13004(new_n13381, new_n13380, new_n13379);
xnor_3 g13005(new_n13382, new_n13381, new_n13378);
xnor_3 g13006(new_n13383, new_n13382, new_n13376);
xnor_3 g13007(new_n13384, new_n13383, new_n13372);
xnor_3 g13008(new_n13385, new_n13384, new_n13368);
nand_4 g13009(new_n13386, new_n12428, new_n12421);
nand_4 g13010(new_n13387, new_n12439, new_n12429);
nand_4 g13011(new_n13388, new_n13387, new_n13386);
not_3  g13012(new_n13389, new_n12424);
nor_4  g13013(new_n13390, new_n12426, new_n13389);
not_3  g13014(new_n13391, new_n12423);
nor_4  g13015(new_n13392, new_n12427, new_n13391);
nor_4  g13016(new_n13393, new_n13392, new_n13390);
xnor_3 g13017(new_n13394, new_n13393, new_n13388);
xnor_3 g13018(new_n13395, new_n13394, new_n13385);
xnor_3 g13019(new_n13396, new_n13395, new_n13365);
not_3  g13020(new_n13397, new_n12431);
nand_4 g13021(new_n13398, new_n13397, new_n12430);
not_3  g13022(new_n13399, new_n12432);
not_3  g13023(new_n13400, new_n12438);
nand_4 g13024(new_n13401, new_n13400, new_n13399);
nand_4 g13025(new_n13402, new_n13401, new_n13398);
nand_4 g13026(new_n13403, n12709, n7523);
nand_4 g13027(new_n13404, n12777, n2515);
xor_3  g13028(new_n13405, new_n13404, new_n13403);
xor_3  g13029(new_n13406, new_n13405, new_n13402);
nand_4 g13030(new_n13407, n7159, n1199);
nand_4 g13031(new_n13408, n6441, n5314);
xor_3  g13032(new_n13409, new_n13408, new_n13407);
nand_4 g13033(new_n13410, n11791, n5767);
nand_4 g13034(new_n13411, n6254, n4828);
xor_3  g13035(new_n13412, new_n13411, new_n13410);
xnor_3 g13036(new_n13413, new_n13412, new_n13409);
nand_4 g13037(new_n13414, n12069, n4436);
nand_4 g13038(new_n13415, n11999, n11153);
xor_3  g13039(new_n13416, new_n13415, new_n13414);
nand_4 g13040(new_n13417, n12489, n6578);
nand_4 g13041(new_n13418, n12947, n996);
xor_3  g13042(new_n13419, new_n13418, new_n13417);
xnor_3 g13043(new_n13420, new_n13419, new_n13416);
xnor_3 g13044(new_n13421, new_n13420, new_n13413);
nand_4 g13045(new_n13422, n11967, n7160);
not_3  g13046(new_n13423, new_n13422);
not_3  g13047(new_n13424, new_n12434);
nor_4  g13048(new_n13425, new_n12436, new_n13424);
not_3  g13049(new_n13426, new_n12433);
nor_4  g13050(new_n13427, new_n12437, new_n13426);
nor_4  g13051(new_n13428, new_n13427, new_n13425);
xnor_3 g13052(new_n13429, new_n13428, new_n13423);
xnor_3 g13053(new_n13430, new_n13429, new_n13421);
xnor_3 g13054(new_n13431, new_n13430, new_n13406);
xnor_3 g13055(new_n13432, new_n13431, new_n13396);
xnor_3 g13056(new_n13433, new_n13432, new_n13363);
xnor_3 g13057(new_n13434, new_n13433, new_n13361);
not_3  g13058(new_n13435, new_n12304);
nand_4 g13059(new_n13436, new_n12333, new_n13435);
nand_4 g13060(new_n13437, new_n12334, new_n12303);
nand_4 g13061(new_n13438, new_n13437, new_n13436);
nor_4  g13062(new_n13439, new_n12221_1, new_n12220);
and_4  g13063(new_n13440, new_n12221_1, new_n12220);
or_4   g13064(new_n13441, new_n13440, new_n12218);
not_3  g13065(new_n13442, new_n13441);
nor_4  g13066(new_n13443, new_n13442, new_n13439);
nand_4 g13067(new_n13444, n11877, n3627);
nand_4 g13068(new_n13445, n8336, n1198);
nand_4 g13069(new_n13446, n6770, n5320);
xor_3  g13070(new_n13447, new_n13446, new_n13445);
xor_3  g13071(new_n13448, new_n13447, new_n13444);
xnor_3 g13072(new_n13449, new_n13448, new_n13443);
xnor_3 g13073(new_n13450, new_n13449, new_n13438);
and_4  g13074(new_n13451, new_n12492, new_n12491);
not_3  g13075(new_n13452, new_n12494);
nor_4  g13076(new_n13453, new_n13452, new_n12488);
nor_4  g13077(new_n13454, new_n13453, new_n13451);
nand_4 g13078(new_n13455, new_n12495, new_n12456);
nand_4 g13079(new_n13456, new_n12500, new_n12496);
nand_4 g13080(new_n13457, new_n13456, new_n13455);
xnor_3 g13081(new_n13458, new_n13457, new_n13454);
xnor_3 g13082(new_n13459, new_n13458, new_n13450);
xnor_3 g13083(new_n13460, new_n13459, new_n13434);
not_3  g13084(new_n13461, new_n12501);
nand_4 g13085(new_n13462, new_n13461, new_n12453);
nand_4 g13086(new_n13463, new_n12506, new_n12502);
nand_4 g13087(new_n13464, new_n13463, new_n13462);
nand_4 g13088(new_n13465, new_n12447, new_n12371);
not_3  g13089(new_n13466, new_n12448);
nand_4 g13090(new_n13467, new_n12452, new_n13466);
nand_4 g13091(new_n13468, new_n13467, new_n13465);
nor_4  g13092(new_n13469, new_n12318, new_n12317);
not_3  g13093(new_n13470, new_n12319);
nor_4  g13094(new_n13471, new_n12325, new_n13470);
nor_4  g13095(new_n13472, new_n13471, new_n13469);
nand_4 g13096(new_n13473, n5319, n1478);
not_3  g13097(new_n13474, new_n13473);
nand_4 g13098(new_n13475, n11728, n7320);
nand_4 g13099(new_n13476, n10990, n4817);
xor_3  g13100(new_n13477, new_n13476, new_n13475);
xnor_3 g13101(new_n13478, new_n13477, new_n13474);
not_3  g13102(new_n13479, new_n12310);
nor_4  g13103(new_n13480, new_n12312, new_n13479);
nor_4  g13104(new_n13481, new_n12313, new_n12309);
nor_4  g13105(new_n13482, new_n13481, new_n13480);
xnor_3 g13106(new_n13483, new_n13482, new_n13478);
nand_4 g13107(new_n13484, n5212, n4516);
nand_4 g13108(new_n13485, n12000, n4189);
nand_4 g13109(new_n13486, n9725, n2564);
xor_3  g13110(new_n13487, new_n13486, new_n13485);
xnor_3 g13111(new_n13488, new_n13487, new_n13484);
nand_4 g13112(new_n13489, n8819, n1094);
nand_4 g13113(new_n13490, n8717, n6986);
xor_3  g13114(new_n13491, new_n13490, new_n13489);
xnor_3 g13115(new_n13492, new_n13491, new_n13488);
xnor_3 g13116(new_n13493, new_n13492, new_n13483);
xnor_3 g13117(new_n13494, new_n13493, new_n13472);
nand_4 g13118(new_n13495, n2433, n2226);
nand_4 g13119(new_n13496, n10678, n6429);
xor_3  g13120(new_n13497, new_n13496, new_n13495);
not_3  g13121(new_n13498, new_n12321);
nor_4  g13122(new_n13499, new_n12323, new_n13498);
not_3  g13123(new_n13500, new_n12320);
nor_4  g13124(new_n13501, new_n12324, new_n13500);
nor_4  g13125(new_n13502, new_n13501, new_n13499);
nand_4 g13126(new_n13503, n10928, n7730);
xnor_3 g13127(new_n13504, new_n13503, new_n13502);
xnor_3 g13128(new_n13505, new_n13504, new_n13497);
nand_4 g13129(new_n13506, new_n12227, new_n12225);
nand_4 g13130(new_n13507, new_n12237, new_n12228);
nand_4 g13131(new_n13508, new_n13507, new_n13506);
nand_4 g13132(new_n13509, n9457, n5760);
nand_4 g13133(new_n13510, n11222, n10022);
xor_3  g13134(new_n13511, new_n13510, new_n13509);
xnor_3 g13135(new_n13512, new_n13511, new_n13508);
xnor_3 g13136(new_n13513, new_n13512, new_n13505);
not_3  g13137(new_n13514, new_n12307);
nor_4  g13138(new_n13515, new_n12314, new_n13514);
not_3  g13139(new_n13516, new_n12315);
nor_4  g13140(new_n13517, new_n12326, new_n13516);
nor_4  g13141(new_n13518, new_n13517, new_n13515);
xnor_3 g13142(new_n13519, new_n13518, new_n13513);
xnor_3 g13143(new_n13520, new_n13519, new_n13494);
nand_4 g13144(new_n13521, new_n12444_1, new_n12443);
not_3  g13145(new_n13522, new_n12441);
nand_4 g13146(new_n13523, new_n12446, new_n13522);
nand_4 g13147(new_n13524, new_n13523, new_n13521);
nand_4 g13148(new_n13525, new_n12289, new_n12330);
not_3  g13149(new_n13526, new_n12327);
nand_4 g13150(new_n13527, new_n12332, new_n13526);
nand_4 g13151(new_n13528, new_n13527, new_n13525);
not_3  g13152(new_n13529, new_n12217);
nand_4 g13153(new_n13530, new_n12223, new_n13529);
nand_4 g13154(new_n13531, new_n12238, new_n12224);
nand_4 g13155(new_n13532, new_n13531, new_n13530);
nand_4 g13156(new_n13533, n9920, n4370);
not_3  g13157(new_n13534, new_n12229);
nand_4 g13158(new_n13535, new_n12232, new_n13534);
nand_4 g13159(new_n13536, new_n13535, new_n12235);
xor_3  g13160(new_n13537, new_n13536, new_n13533);
xnor_3 g13161(new_n13538, new_n13537, new_n13532);
xnor_3 g13162(new_n13539, new_n13538, new_n13528);
xnor_3 g13163(new_n13540, new_n13539, new_n13524);
xnor_3 g13164(new_n13541, new_n13540, new_n13520);
xnor_3 g13165(new_n13542, new_n13541, new_n13468);
xnor_3 g13166(new_n13543, new_n13542, new_n13464);
xnor_3 g13167(new_n13544, new_n13543, new_n13460);
xnor_3 g13168(new_n13545, new_n13544, new_n13357);
xnor_3 g13169(n8100, new_n13545, new_n13351);
not_3  g13170(new_n13547, new_n10018);
xor_3  g13171(n8138, new_n10019, new_n13547);
not_3  g13172(new_n13549, new_n6278);
xor_3  g13173(n8202, new_n6280, new_n13549);
xor_3  g13174(n8303, new_n3825, new_n3812);
not_3  g13175(new_n13552, new_n3079);
xor_3  g13176(n8398, new_n3080, new_n13552);
not_3  g13177(new_n13554, new_n4460);
xor_3  g13178(n9137, new_n4461, new_n13554);
not_3  g13179(new_n13556, new_n7375);
xor_3  g13180(n9387, new_n13556, new_n7374);
not_3  g13181(new_n13558, new_n11969);
xor_3  g13182(n9571, new_n13558, new_n11968);
nor_4  g13183(new_n13560, new_n1018, new_n1015);
xor_3  g13184(n9578, new_n13560, new_n1062);
xor_3  g13185(n9706, new_n1212, new_n1209_1);
not_3  g13186(new_n13563, new_n4450);
xor_3  g13187(n9756, new_n4463, new_n13563);
nand_4 g13188(new_n13565, new_n7039, new_n7015);
nand_4 g13189(new_n13566, new_n13565, new_n7018);
not_3  g13190(new_n13567, new_n6988);
nand_4 g13191(new_n13568, new_n13567, new_n6768);
nand_4 g13192(new_n13569, new_n7013, new_n6989);
nand_4 g13193(new_n13570, new_n13569, new_n13568);
not_3  g13194(new_n13571, new_n6614);
nand_4 g13195(new_n13572, new_n6648, new_n13571);
nand_4 g13196(new_n13573, new_n6665, new_n6649);
nand_4 g13197(new_n13574, new_n13573, new_n13572);
nor_4  g13198(new_n13575, new_n6830, new_n6829);
not_3  g13199(new_n13576, new_n6831);
nor_4  g13200(new_n13577, new_n6837, new_n13576);
nor_4  g13201(new_n13578, new_n13577, new_n13575);
xnor_3 g13202(new_n13579, new_n13578, new_n13574);
not_3  g13203(new_n13580, new_n6947);
nand_4 g13204(new_n13581, new_n13580, new_n6912);
nand_4 g13205(new_n13582, new_n6962, new_n6948);
nand_4 g13206(new_n13583, new_n13582, new_n13581);
nor_4  g13207(new_n13584, new_n6733, new_n6732);
nor_4  g13208(new_n13585, new_n6741, new_n6735);
nor_4  g13209(new_n13586, new_n13585, new_n13584);
not_3  g13210(new_n13587, new_n6737);
nor_4  g13211(new_n13588, new_n6739, new_n13587);
not_3  g13212(new_n13589, new_n6736);
nor_4  g13213(new_n13590, new_n6740, new_n13589);
nor_4  g13214(new_n13591, new_n13590, new_n13588);
nand_4 g13215(new_n13592, n10451, n2226);
xnor_3 g13216(new_n13593, new_n13592, new_n13591);
xnor_3 g13217(new_n13594, new_n13593, new_n13586);
nand_4 g13218(new_n13595, n10278, n6986);
nand_4 g13219(new_n13596, n11423, n10928);
xor_3  g13220(new_n13597, new_n13596, new_n13595);
not_3  g13221(new_n13598, new_n6725);
nor_4  g13222(new_n13599, new_n6727, new_n13598);
not_3  g13223(new_n13600, new_n6724);
nor_4  g13224(new_n13601, new_n6728, new_n13600);
nor_4  g13225(new_n13602, new_n13601, new_n13599);
nand_4 g13226(new_n13603, n10678, n3022);
xnor_3 g13227(new_n13604, new_n13603, new_n13602);
xnor_3 g13228(new_n13605, new_n13604, new_n13597);
xnor_3 g13229(new_n13606, new_n13605, new_n13594);
nand_4 g13230(new_n13607, n10327, n4189);
nand_4 g13231(new_n13608, new_n6629, new_n6627);
nand_4 g13232(new_n13609, new_n6639, new_n6630);
nand_4 g13233(new_n13610, new_n13609, new_n13608);
nand_4 g13234(new_n13611, n9583, n2564);
not_3  g13235(new_n13612, new_n13611);
xnor_3 g13236(new_n13613, new_n13612, new_n13610);
xnor_3 g13237(new_n13614, new_n13613, new_n13607);
xnor_3 g13238(new_n13615, new_n13614, new_n13606);
nand_4 g13239(new_n13616, new_n6729, new_n6722);
nand_4 g13240(new_n13617, new_n6742_1, new_n6730);
nand_4 g13241(new_n13618, new_n13617, new_n13616);
nand_4 g13242(new_n13619, n11023, n1094);
nand_4 g13243(new_n13620, n9920, n7456);
not_3  g13244(new_n13621, new_n6631);
nand_4 g13245(new_n13622, new_n6634, new_n13621);
nand_4 g13246(new_n13623, new_n13622, new_n6637);
xor_3  g13247(new_n13624, new_n13623, new_n13620);
xor_3  g13248(new_n13625, new_n13624, new_n13619);
xnor_3 g13249(new_n13626, new_n13625, new_n13618);
xnor_3 g13250(new_n13627, new_n13626, new_n13615);
xnor_3 g13251(new_n13628, new_n13627, new_n13583);
xnor_3 g13252(new_n13629, new_n13628, new_n13579);
not_3  g13253(new_n13630, new_n6719);
nand_4 g13254(new_n13631, new_n6752, new_n13630);
nand_4 g13255(new_n13632, new_n6766, new_n6753);
nand_4 g13256(new_n13633, new_n13632, new_n13631);
nand_4 g13257(new_n13634, n11662, n6770);
nand_4 g13258(new_n13635, new_n6645_1, new_n6644);
not_3  g13259(new_n13636, new_n6642);
nand_4 g13260(new_n13637, new_n6647, new_n13636);
nand_4 g13261(new_n13638, new_n13637, new_n13635);
xnor_3 g13262(new_n13639, new_n13638, new_n13634);
nand_4 g13263(new_n13640, new_n6625, new_n6618);
nand_4 g13264(new_n13641, new_n6640, new_n6626);
nand_4 g13265(new_n13642, new_n13641, new_n13640);
not_3  g13266(new_n13643, new_n6621);
nor_4  g13267(new_n13644, new_n6623, new_n13643);
not_3  g13268(new_n13645, new_n6620);
nor_4  g13269(new_n13646, new_n6624, new_n13645);
nor_4  g13270(new_n13647, new_n13646, new_n13644);
nand_4 g13271(new_n13648, n9640, n7320);
not_3  g13272(new_n13649, new_n13648);
nand_4 g13273(new_n13650, n8336, n2278);
nand_4 g13274(new_n13651, n7523, n6703);
xor_3  g13275(new_n13652, new_n13651, new_n13650);
nand_4 g13276(new_n13653, n12591, n3627);
nand_4 g13277(new_n13654, n4516, n3932);
xor_3  g13278(new_n13655, new_n13654, new_n13653);
xnor_3 g13279(new_n13656, new_n13655, new_n13652);
xnor_3 g13280(new_n13657, new_n13656, new_n13649);
xnor_3 g13281(new_n13658, new_n13657, new_n13647);
xnor_3 g13282(new_n13659, new_n13658, new_n13642);
nand_4 g13283(new_n13660, n12247, n11153);
not_3  g13284(new_n13661, new_n13660);
nor_4  g13285(new_n13662, new_n6835, new_n6834);
nand_4 g13286(new_n13663, new_n6835, new_n6834);
nand_4 g13287(new_n13664, new_n13663, new_n6833);
not_3  g13288(new_n13665, new_n13664);
nor_4  g13289(new_n13666, new_n13665, new_n13662);
nand_4 g13290(new_n13667, n6687, n753);
nand_4 g13291(new_n13668, n2087, n1798);
xor_3  g13292(new_n13669, new_n13668, new_n13667);
nand_4 g13293(new_n13670, n12826, n7891);
nand_4 g13294(new_n13671, n12391, n4094);
xor_3  g13295(new_n13672, new_n13671, new_n13670);
xnor_3 g13296(new_n13673, new_n13672, new_n13669);
xnor_3 g13297(new_n13674, new_n13673, new_n13666);
xnor_3 g13298(new_n13675, new_n13674, new_n13661);
xnor_3 g13299(new_n13676, new_n13675, new_n13659);
nand_4 g13300(new_n13677, new_n6749, new_n6747);
nand_4 g13301(new_n13678, new_n6751, new_n6743);
nand_4 g13302(new_n13679, new_n13678, new_n13677);
nand_4 g13303(new_n13680, new_n6929, new_n6922);
nand_4 g13304(new_n13681, new_n6944, new_n6931);
nand_4 g13305(new_n13682, new_n13681, new_n13680);
xnor_3 g13306(new_n13683, new_n13682, new_n13679);
xnor_3 g13307(new_n13684, new_n13683, new_n13676);
xnor_3 g13308(new_n13685, new_n13684, new_n13639);
xnor_3 g13309(new_n13686, new_n13685, new_n13633);
xnor_3 g13310(new_n13687, new_n13686, new_n13629);
nand_4 g13311(new_n13688, new_n6986_1, new_n6963);
nor_4  g13312(new_n13689, new_n6984, new_n6966);
xnor_3 g13313(new_n13690, new_n13689, new_n6963);
nand_4 g13314(new_n13691, new_n13690, new_n6863);
nand_4 g13315(new_n13692, new_n13691, new_n13688);
nand_4 g13316(new_n13693, new_n6847, new_n6815);
nand_4 g13317(new_n13694, new_n6862, new_n6848);
nand_4 g13318(new_n13695, new_n13694, new_n13693);
nand_4 g13319(new_n13696, new_n6934, new_n6932);
nand_4 g13320(new_n13697, new_n6943, new_n6935);
nand_4 g13321(new_n13698, new_n13697, new_n13696);
not_3  g13322(new_n13699, new_n6822_1);
nor_4  g13323(new_n13700, new_n6824, new_n13699);
not_3  g13324(new_n13701, new_n6821);
nor_4  g13325(new_n13702, new_n6825, new_n13701);
nor_4  g13326(new_n13703, new_n13702, new_n13700);
xnor_3 g13327(new_n13704, new_n13703, new_n13698);
nand_4 g13328(new_n13705, n10898, n9457);
nand_4 g13329(new_n13706, n12511, n11222);
not_3  g13330(new_n13707, new_n13706);
xor_3  g13331(new_n13708, new_n13707, new_n13705);
nand_4 g13332(new_n13709, n11876, n4817);
nand_4 g13333(new_n13710, n5319, n3754);
xor_3  g13334(new_n13711, new_n13710, new_n13709);
xor_3  g13335(new_n13712, new_n13711, new_n13708);
xnor_3 g13336(new_n13713, new_n13712, new_n13704);
nand_4 g13337(new_n13714, n12069, n10685);
not_3  g13338(new_n13715, new_n13714);
not_3  g13339(new_n13716, new_n6925);
nor_4  g13340(new_n13717, new_n6927, new_n13716);
nor_4  g13341(new_n13718, new_n6928, new_n6924);
nor_4  g13342(new_n13719, new_n13718, new_n13717);
nand_4 g13343(new_n13720, n6578, n5645);
not_3  g13344(new_n13721, new_n13720);
xnor_3 g13345(new_n13722, new_n13721, new_n13719);
nand_4 g13346(new_n13723, n11922, n4828);
nand_4 g13347(new_n13724, n8665, n2515);
not_3  g13348(new_n13725, new_n13724);
xor_3  g13349(new_n13726, new_n13725, new_n13723);
xnor_3 g13350(new_n13727, new_n13726, new_n13722);
xnor_3 g13351(new_n13728, new_n13727, new_n13715);
xnor_3 g13352(new_n13729, new_n13728, new_n13713);
nand_4 g13353(new_n13730, new_n6826_1, new_n6819);
not_3  g13354(new_n13731, new_n6838);
nand_4 g13355(new_n13732, new_n13731, new_n6827);
nand_4 g13356(new_n13733, new_n13732, new_n13730);
nand_4 g13357(new_n13734, n996, n159);
nand_4 g13358(new_n13735, n5767, n2749);
xor_3  g13359(new_n13736, new_n13735, new_n13734);
nand_4 g13360(new_n13737, n1199, n1067);
nand_4 g13361(new_n13738, n5314, n1510);
xor_3  g13362(new_n13739, new_n13738, new_n13737);
xor_3  g13363(new_n13740, new_n13739, new_n13736);
nand_4 g13364(new_n13741, n7160, n2551);
not_3  g13365(new_n13742, new_n6939);
nor_4  g13366(new_n13743, new_n6941, new_n13742);
nor_4  g13367(new_n13744, new_n6942, new_n6938);
nor_4  g13368(new_n13745, new_n13744, new_n13743);
xnor_3 g13369(new_n13746, new_n13745, new_n13741);
xnor_3 g13370(new_n13747, new_n13746, new_n13740);
xnor_3 g13371(new_n13748, new_n13747, new_n13733);
xnor_3 g13372(new_n13749, new_n13748, new_n13729);
nand_4 g13373(new_n13750, new_n6917, new_n6916);
nand_4 g13374(new_n13751, new_n6946, new_n6919);
nand_4 g13375(new_n13752, new_n13751, new_n13750);
nand_4 g13376(new_n13753, new_n6844, new_n6843);
not_3  g13377(new_n13754, new_n6839);
nand_4 g13378(new_n13755, new_n6846, new_n13754);
nand_4 g13379(new_n13756, new_n13755, new_n13753);
xnor_3 g13380(new_n13757, new_n13756, new_n13752);
xnor_3 g13381(new_n13758, new_n13757, new_n13749);
xnor_3 g13382(new_n13759, new_n13758, new_n13695);
xnor_3 g13383(new_n13760, new_n13759, new_n13692);
xnor_3 g13384(new_n13761, new_n13760, new_n13687);
xnor_3 g13385(new_n13762, new_n13761, new_n13570);
xnor_3 g13386(n9767, new_n13762, new_n13566);
not_3  g13387(new_n13764, new_n2180);
xor_3  g13388(n9820, new_n2182, new_n13764);
nand_4 g13389(new_n13766, new_n9990, new_n9989);
xnor_3 g13390(n9938, new_n13766, new_n10033);
xor_3  g13391(n10476, new_n1058, new_n1055);
xor_3  g13392(n10589, new_n1052, new_n1041);
not_3  g13393(new_n13770, new_n1205);
xor_3  g13394(n10695, new_n1207, new_n13770);
not_3  g13395(new_n13772, new_n3842_1);
nor_4  g13396(new_n13773, new_n3794, new_n3793);
xnor_3 g13397(n10789, new_n13773, new_n13772);
xor_3  g13398(n10851, new_n3074, new_n3064);
not_3  g13399(new_n13776, new_n5260);
xor_3  g13400(n10913, new_n5269, new_n13776);
xnor_3 g13401(n10949, new_n7512, new_n7379);
xnor_3 g13402(n11216, new_n11971, new_n11916);
xor_3  g13403(n11326, new_n5261, new_n5251);
not_3  g13404(new_n13781, new_n5571);
not_3  g13405(new_n13782, new_n5806);
nor_4  g13406(new_n13783, new_n13782, new_n13781);
nor_4  g13407(new_n13784, new_n5806, new_n5571);
nor_4  g13408(new_n13785, new_n5942, new_n13784);
nor_4  g13409(new_n13786, new_n13785, new_n13783);
nand_4 g13410(new_n13787, new_n5883, new_n5853);
not_3  g13411(new_n13788, new_n5884);
nand_4 g13412(new_n13789, new_n5887, new_n13788);
nand_4 g13413(new_n13790, new_n13789, new_n13787);
nand_4 g13414(new_n13791, n9763, n45);
nand_4 g13415(new_n13792, new_n5553, new_n5552);
not_3  g13416(new_n13793, new_n5550);
nand_4 g13417(new_n13794, new_n5555, new_n13793);
nand_4 g13418(new_n13795, new_n13794, new_n13792);
xnor_3 g13419(new_n13796, new_n13795, new_n13791);
xnor_3 g13420(new_n13797, new_n13796, new_n13790);
not_3  g13421(new_n13798, new_n5528);
nand_4 g13422(new_n13799, new_n5556, new_n13798);
nand_4 g13423(new_n13800, new_n5570, new_n5557);
nand_4 g13424(new_n13801, new_n13800, new_n13799);
nand_4 g13425(new_n13802, new_n5843, new_n5811);
nand_4 g13426(new_n13803, new_n5844, new_n5810);
nand_4 g13427(new_n13804, new_n13803, new_n13802);
xnor_3 g13428(new_n13805, new_n13804, new_n13801);
xnor_3 g13429(new_n13806, new_n13805, new_n13797);
nand_4 g13430(new_n13807, new_n5924, new_n5892);
nand_4 g13431(new_n13808, new_n5926, new_n5925);
nand_4 g13432(new_n13809, new_n13808, new_n13807);
nor_4  g13433(new_n13810, new_n5541, new_n5540);
not_3  g13434(new_n13811, new_n5542);
nor_4  g13435(new_n13812, new_n5548, new_n13811);
nor_4  g13436(new_n13813, new_n13812, new_n13810);
xnor_3 g13437(new_n13814, new_n13813, new_n13809);
not_3  g13438(new_n13815, new_n5814_1);
nand_4 g13439(new_n13816, new_n5820, new_n13815);
nand_4 g13440(new_n13817, new_n5835, new_n5821);
nand_4 g13441(new_n13818, new_n13817, new_n13816);
nand_4 g13442(new_n13819, n2253, n1097);
not_3  g13443(new_n13820, new_n5816);
nor_4  g13444(new_n13821, new_n5818, new_n13820);
not_3  g13445(new_n13822, new_n5815);
nor_4  g13446(new_n13823, new_n5819, new_n13822);
nor_4  g13447(new_n13824, new_n13823, new_n13821);
xnor_3 g13448(new_n13825, new_n13824, new_n13819);
not_3  g13449(new_n13826, new_n5826);
nand_4 g13450(new_n13827, new_n5829, new_n13826);
and_4  g13451(new_n13828, new_n13827, new_n5832);
nand_4 g13452(new_n13829, n12299, n12221);
nand_4 g13453(new_n13830, n9241, n9189);
xor_3  g13454(new_n13831, new_n13830, new_n13829);
xnor_3 g13455(new_n13832, new_n13831, new_n13828);
xnor_3 g13456(new_n13833, new_n13832, new_n13825);
nand_4 g13457(new_n13834, n12145, n7436);
not_3  g13458(new_n13835, new_n13834);
nand_4 g13459(new_n13836, n10217, n6776);
nand_4 g13460(new_n13837, n8276, n2522);
xor_3  g13461(new_n13838, new_n13837, new_n13836);
xnor_3 g13462(new_n13839, new_n13838, new_n13835);
nand_4 g13463(new_n13840, new_n5824, new_n5822);
nand_4 g13464(new_n13841, new_n5834, new_n5825);
nand_4 g13465(new_n13842, new_n13841, new_n13840);
xnor_3 g13466(new_n13843, new_n13842, new_n13839);
xnor_3 g13467(new_n13844, new_n13843, new_n13833);
xnor_3 g13468(new_n13845, new_n13844, new_n13818);
nand_4 g13469(new_n13846, new_n5921, new_n5919);
nand_4 g13470(new_n13847, new_n5923, new_n5915);
nand_4 g13471(new_n13848, new_n13847, new_n13846);
not_3  g13472(new_n13849, new_n5544);
nor_4  g13473(new_n13850, new_n5546, new_n13849);
not_3  g13474(new_n13851, new_n5543);
nor_4  g13475(new_n13852, new_n5547, new_n13851);
nor_4  g13476(new_n13853, new_n13852, new_n13850);
nand_4 g13477(new_n13854, n5964, n3865);
nand_4 g13478(new_n13855, n12705, n4634);
xor_3  g13479(new_n13856, new_n13855, new_n13854);
xor_3  g13480(new_n13857, new_n13856, new_n13853);
xnor_3 g13481(new_n13858, new_n13857, new_n13848);
xnor_3 g13482(new_n13859, new_n13858, new_n13845);
not_3  g13483(new_n13860, new_n5896);
nand_4 g13484(new_n13861, new_n5901, new_n13860);
nand_4 g13485(new_n13862, new_n5913, new_n5902);
nand_4 g13486(new_n13863, new_n13862, new_n13861);
not_3  g13487(new_n13864, new_n5904);
nand_4 g13488(new_n13865, new_n13864, new_n5903);
nand_4 g13489(new_n13866, new_n5911, new_n5905);
nand_4 g13490(new_n13867, new_n13866, new_n13865);
nand_4 g13491(new_n13868, n3616, n2498);
not_3  g13492(new_n13869, new_n13868);
nand_4 g13493(new_n13870, n10545, n521);
nand_4 g13494(new_n13871, n7690, n5579);
xnor_3 g13495(new_n13872, new_n13871, new_n13870);
xnor_3 g13496(new_n13873, new_n13872, new_n13869);
xnor_3 g13497(new_n13874, new_n13873, new_n13867);
and_4  g13498(new_n13875, new_n5899, new_n5898);
not_3  g13499(new_n13876, new_n5897);
nor_4  g13500(new_n13877, new_n5900, new_n13876);
nor_4  g13501(new_n13878, new_n13877, new_n13875);
nand_4 g13502(new_n13879, n5860, n806);
nand_4 g13503(new_n13880, n4499, n2558);
nand_4 g13504(new_n13881, n7270, n2393);
xnor_3 g13505(new_n13882, new_n13881, new_n13880);
nand_4 g13506(new_n13883, n5331, n1576);
nand_4 g13507(new_n13884, n7388, n2507);
xnor_3 g13508(new_n13885, new_n13884, new_n13883);
xnor_3 g13509(new_n13886, new_n13885, new_n13882);
xnor_3 g13510(new_n13887, new_n13886, new_n13879);
xnor_3 g13511(new_n13888, new_n13887, new_n13878);
xnor_3 g13512(new_n13889, new_n13888, new_n13874);
xnor_3 g13513(new_n13890, new_n13889, new_n13863);
not_3  g13514(new_n13891, new_n5856);
nand_4 g13515(new_n13892, new_n5861, new_n13891);
nand_4 g13516(new_n13893, new_n5873, new_n5862);
nand_4 g13517(new_n13894, new_n13893, new_n13892);
not_3  g13518(new_n13895, new_n5864);
nand_4 g13519(new_n13896, new_n13895, new_n5863);
nand_4 g13520(new_n13897, new_n5871, new_n5865);
nand_4 g13521(new_n13898, new_n13897, new_n13896);
and_4  g13522(new_n13899, new_n5869, new_n5868);
nor_4  g13523(new_n13900, new_n5870, new_n5867);
nor_4  g13524(new_n13901, new_n13900, new_n13899);
xnor_3 g13525(new_n13902, new_n13901, new_n13898);
nand_4 g13526(new_n13903, n5305, n2512);
nand_4 g13527(new_n13904, n12648, n6016);
nand_4 g13528(new_n13905, n11892, n5153);
xnor_3 g13529(new_n13906, new_n13905, new_n13904);
xnor_3 g13530(new_n13907, new_n13906, new_n13903);
nor_4  g13531(new_n13908, new_n5859, new_n5858);
not_3  g13532(new_n13909, new_n5857_1);
nand_4 g13533(new_n13910, new_n5859, new_n5858);
nand_4 g13534(new_n13911, new_n13910, new_n13909);
not_3  g13535(new_n13912, new_n13911);
nor_4  g13536(new_n13913, new_n13912, new_n13908);
nand_4 g13537(new_n13914, n5798, n2530);
nand_4 g13538(new_n13915, n10547, n7265);
nand_4 g13539(new_n13916, n8476, n2347);
xnor_3 g13540(new_n13917, new_n13916, new_n13915);
xnor_3 g13541(new_n13918, new_n13917, new_n13914);
xnor_3 g13542(new_n13919, new_n13918, new_n13913);
xnor_3 g13543(new_n13920, new_n13919, new_n13907);
xnor_3 g13544(new_n13921, new_n13920, new_n13902);
xnor_3 g13545(new_n13922, new_n13921, new_n13894);
xnor_3 g13546(new_n13923, new_n13922, new_n13890);
nand_4 g13547(new_n13924, n3986, n3342);
nand_4 g13548(new_n13925, n11257, n2879);
nand_4 g13549(new_n13926, n8759, n7823);
xor_3  g13550(new_n13927, new_n13926, new_n13925);
xor_3  g13551(new_n13928, new_n13927, new_n13924);
xnor_3 g13552(new_n13929, new_n13928, new_n13923);
and_4  g13553(new_n13930, new_n5909, new_n5908);
nor_4  g13554(new_n13931, new_n5910, new_n5907);
nor_4  g13555(new_n13932, new_n13931, new_n13930);
nand_4 g13556(new_n13933, new_n5880, new_n5878);
nand_4 g13557(new_n13934, new_n5882, new_n5874);
nand_4 g13558(new_n13935, new_n13934, new_n13933);
xnor_3 g13559(new_n13936, new_n13935, new_n13932);
xnor_3 g13560(new_n13937, new_n13936, new_n13929);
nand_4 g13561(new_n13938, new_n5839, new_n5838);
nand_4 g13562(new_n13939, new_n5841, new_n5836);
nand_4 g13563(new_n13940, new_n13939, new_n13938);
not_3  g13564(new_n13941, new_n5531);
nand_4 g13565(new_n13942, new_n5537, new_n13941);
not_3  g13566(new_n13943, new_n5549);
nand_4 g13567(new_n13944, new_n13943, new_n5538);
nand_4 g13568(new_n13945, new_n13944, new_n13942);
not_3  g13569(new_n13946, new_n5533);
nor_4  g13570(new_n13947, new_n5535, new_n13946);
not_3  g13571(new_n13948, new_n5532);
nor_4  g13572(new_n13949, new_n5536, new_n13948);
nor_4  g13573(new_n13950, new_n13949, new_n13947);
nand_4 g13574(new_n13951, n9195, n4312);
nand_4 g13575(new_n13952, n12025, n10223);
xor_3  g13576(new_n13953, new_n13952, new_n13951);
nand_4 g13577(new_n13954, n10510, n2024);
nand_4 g13578(new_n13955, n10644, n7946);
xor_3  g13579(new_n13956, new_n13955, new_n13954);
xnor_3 g13580(new_n13957, new_n13956, new_n13953);
xnor_3 g13581(new_n13958, new_n13957, new_n13950);
xnor_3 g13582(new_n13959, new_n13958, new_n13945);
xnor_3 g13583(new_n13960, new_n13959, new_n13940);
xnor_3 g13584(new_n13961, new_n13960, new_n13937);
xnor_3 g13585(new_n13962, new_n13961, new_n13859);
xnor_3 g13586(new_n13963, new_n13962, new_n13814);
xnor_3 g13587(new_n13964, new_n13963, new_n13806);
nand_4 g13588(new_n13965, n9111, n5857);
nand_4 g13589(new_n13966, n7965, n6431);
xor_3  g13590(new_n13967, new_n13966, new_n13965);
not_3  g13591(new_n13968, new_n13967);
xnor_3 g13592(new_n13969, new_n13968, new_n13964);
not_3  g13593(new_n13970, new_n5845);
nand_4 g13594(new_n13971, new_n5849, new_n13970);
not_3  g13595(new_n13972, new_n5941);
nand_4 g13596(new_n13973, new_n13972, new_n5850);
nand_4 g13597(new_n13974, new_n13973, new_n13971);
not_3  g13598(new_n13975, new_n5931);
not_3  g13599(new_n13976, new_n5938);
nand_4 g13600(new_n13977, new_n13976, new_n13975);
xnor_3 g13601(new_n13978, new_n13977, new_n13974);
xnor_3 g13602(new_n13979, new_n13978, new_n13969);
xnor_3 g13603(n11707, new_n13979, new_n13786);
not_3  g13604(new_n13981, new_n6521);
xor_3  g13605(n11755, new_n13981, new_n6520);
xor_3  g13606(n11780, new_n3838, new_n3834);
not_3  g13607(new_n13984, new_n10445);
xor_3  g13608(n11919, new_n10446, new_n13984);
xor_3  g13609(n12005, new_n10448, new_n10430);
xnor_3 g13610(n12014, new_n10897, new_n10892);
not_3  g13611(new_n13988, new_n9143);
xnor_3 g13612(n12020, new_n13988, new_n9100);
not_3  g13613(new_n13990, new_n11924);
xor_3  g13614(n12076, new_n11963, new_n13990);
xnor_3 g13615(n12111, new_n12528, new_n12520);
xnor_3 g13616(n12444, new_n10899, new_n10883);
nor_4  g13617(new_n13994, new_n5790, new_n5788);
xnor_3 g13618(n12807, new_n13994, new_n5804);
endmodule


