// Benchmark "top_810222779_843330999_776144567_776418743_1234615" written by ABC on Fri Jun 14 22:41:39 2024

module top_810222779_843330999_776144567_776418743_1234615 ( 
    n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82, n86,
    n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200, n219,
    n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273, n284,
    n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341, n344,
    n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420, n430,
    n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560, n561,
    n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609, n626,
    n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729, n734,
    n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831, n832,
    n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961, n969,
    n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061, n1071,
    n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164, n1172,
    n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246, n1250,
    n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305, n1345,
    n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411, n1415,
    n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470, n1474,
    n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536, n1566,
    n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627, n1644,
    n1647, n1656, n1750, n1753,
    n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181,
    n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362,
    n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501,
    n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669,
    n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918,
    n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063,
    n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285,
    n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368,
    n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588,
    n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752  );
  input  n11, n21, n29, n40, n45, n50, n52, n54, n56, n58, n71, n77, n82,
    n86, n87, n94, n107, n117, n138, n143, n153, n155, n156, n159, n200,
    n219, n220, n222, n223, n243, n244, n246, n251, n254, n262, n268, n273,
    n284, n288, n293, n299, n300, n307, n310, n312, n314, n315, n318, n341,
    n344, n346, n374, n376, n380, n391, n392, n399, n408, n409, n416, n420,
    n430, n477, n478, n487, n489, n502, n506, n507, n510, n545, n559, n560,
    n561, n567, n574, n581, n582, n589, n593, n598, n600, n607, n608, n609,
    n626, n641, n645, n663, n671, n676, n690, n695, n701, n710, n727, n729,
    n734, n742, n743, n755, n769, n775, n778, n779, n787, n790, n823, n831,
    n832, n839, n849, n879, n882, n885, n905, n920, n936, n947, n953, n961,
    n969, n980, n984, n986, n992, n997, n1023, n1040, n1044, n1054, n1061,
    n1071, n1095, n1103, n1114, n1121, n1138, n1152, n1154, n1156, n1164,
    n1172, n1175, n1187, n1191, n1193, n1205, n1225, n1227, n1239, n1246,
    n1250, n1263, n1278, n1281, n1283, n1286, n1289, n1299, n1301, n1305,
    n1345, n1346, n1350, n1361, n1386, n1387, n1389, n1393, n1401, n1411,
    n1415, n1418, n1428, n1435, n1438, n1443, n1446, n1448, n1463, n1470,
    n1474, n1476, n1500, n1502, n1506, n1516, n1520, n1521, n1523, n1536,
    n1566, n1569, n1576, n1586, n1592, n1609, n1613, n1616, n1626, n1627,
    n1644, n1647, n1656, n1750, n1753;
  output n22, n23, n27, n30, n85, n112, n126, n130, n161, n164, n173, n181,
    n184, n216, n230, n233, n247, n275, n292, n301, n304, n337, n352, n362,
    n364, n370, n378, n396, n417, n428, n453, n457, n460, n497, n498, n501,
    n509, n516, n517, n534, n553, n585, n595, n597, n625, n638, n640, n669,
    n693, n714, n719, n726, n773, n782, n794, n821, n842, n894, n916, n918,
    n952, n990, n1006, n1017, n1042, n1050, n1051, n1058, n1060, n1063,
    n1065, n1177, n1186, n1195, n1209, n1211, n1231, n1234, n1253, n1285,
    n1288, n1292, n1296, n1302, n1306, n1320, n1322, n1337, n1359, n1368,
    n1375, n1391, n1420, n1421, n1427, n1527, n1534, n1547, n1548, n1588,
    n1594, n1632, n1639, n1645, n1687, n1729, n1738, n1752;
  wire new_n316, new_n317, new_n318_1, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n334, new_n335,
    new_n336, new_n337_1, new_n338, new_n339, new_n340, new_n341_1,
    new_n342, new_n343, new_n344_1, new_n345, new_n346_1, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352_1, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362_1, new_n363, new_n364_1, new_n365, new_n366, new_n367,
    new_n368, new_n369, new_n370_1, new_n371, new_n372, new_n373,
    new_n374_1, new_n375, new_n376_1, new_n377, new_n378_1, new_n379,
    new_n380_1, new_n381, new_n382, new_n383, new_n384, new_n385, new_n386,
    new_n387, new_n388, new_n389, new_n390, new_n391_1, new_n392_1,
    new_n393, new_n394, new_n395, new_n396_1, new_n397, new_n398,
    new_n399_1, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408_1, new_n409_1, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416_1, new_n417_1,
    new_n418, new_n419, new_n420_1, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428_1, new_n429, new_n430_1,
    new_n431, new_n432, new_n433, new_n434, new_n435, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n443, new_n444,
    new_n445, new_n446, new_n447, new_n448, new_n449, new_n450, new_n451,
    new_n452, new_n453_1, new_n454, new_n455, new_n456, new_n457_1,
    new_n458, new_n459, new_n460_1, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477_1,
    new_n478_1, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487_1, new_n488, new_n489_1, new_n490,
    new_n491, new_n492, new_n493, new_n494, new_n495, new_n496, new_n497_1,
    new_n498_1, new_n499, new_n500, new_n501_1, new_n502_1, new_n503,
    new_n504, new_n505, new_n506_1, new_n507_1, new_n508, new_n509_1,
    new_n510_1, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516_1, new_n517_1, new_n518, new_n519, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534_1, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545_1, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553_1, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559_1, new_n560_1, new_n561_1, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567_1, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574_1, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581_1, new_n582_1,
    new_n583, new_n584, new_n585_1, new_n586, new_n587, new_n588,
    new_n589_1, new_n590, new_n591, new_n592, new_n593_1, new_n594,
    new_n595_1, new_n596, new_n597_1, new_n598_1, new_n599, new_n600_1,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607_1,
    new_n608_1, new_n609_1, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625_1, new_n626_1,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638_1, new_n639,
    new_n640_1, new_n641_1, new_n642, new_n643, new_n644, new_n645_1,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n660, new_n661, new_n663_1,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669_1, new_n670,
    new_n671_1, new_n672, new_n673, new_n674, new_n675, new_n676_1,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690_1,
    new_n691, new_n692, new_n693_1, new_n694, new_n695_1, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701_1, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710_1,
    new_n711, new_n712, new_n713, new_n714_1, new_n715, new_n716, new_n717,
    new_n718, new_n719_1, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726_1, new_n727_1, new_n728, new_n729_1, new_n730,
    new_n731, new_n732, new_n733, new_n734_1, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742_1, new_n743_1,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755_1, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769_1, new_n770, new_n771,
    new_n772, new_n773_1, new_n774, new_n775_1, new_n776, new_n777,
    new_n778_1, new_n779_1, new_n780, new_n781, new_n782_1, new_n783,
    new_n784, new_n785, new_n786, new_n787_1, new_n788, new_n789,
    new_n790_1, new_n791, new_n792, new_n793, new_n794_1, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821_1, new_n822,
    new_n823_1, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831_1, new_n832_1, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839_1, new_n840, new_n841,
    new_n842_1, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849_1, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879_1, new_n880, new_n881, new_n882_1,
    new_n883, new_n884, new_n885_1, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894_1, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905_1, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916_1, new_n917,
    new_n918_1, new_n919, new_n920_1, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936_1, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947_1, new_n948, new_n949, new_n950, new_n951,
    new_n952_1, new_n953_1, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961_1, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969_1, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980_1, new_n981, new_n982, new_n983, new_n984_1,
    new_n985, new_n986_1, new_n987, new_n988, new_n989, new_n990_1,
    new_n991, new_n992_1, new_n993, new_n994, new_n995, new_n996,
    new_n997_1, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006_1, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017_1, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023_1, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040_1, new_n1041, new_n1042_1, new_n1043, new_n1044_1, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050_1, new_n1051_1,
    new_n1052, new_n1053, new_n1054_1, new_n1055, new_n1056, new_n1057,
    new_n1058_1, new_n1059, new_n1060_1, new_n1061_1, new_n1062,
    new_n1063_1, new_n1064, new_n1065_1, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071_1, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095_1,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103_1, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114_1,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121_1, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138_1,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152_1, new_n1153, new_n1154_1, new_n1155, new_n1156_1,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164_1, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1172_1, new_n1173, new_n1174, new_n1175_1,
    new_n1176, new_n1177_1, new_n1178, new_n1179, new_n1182, new_n1184,
    new_n1185, new_n1186_1, new_n1187_1, new_n1189, new_n1191_1, new_n1192,
    new_n1193_1, new_n1194, new_n1195_1, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205_1, new_n1206, new_n1207, new_n1208, new_n1209_1, new_n1210,
    new_n1211_1, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225_1, new_n1226, new_n1227_1, new_n1228,
    new_n1229, new_n1230, new_n1231_1, new_n1232, new_n1233, new_n1234_1,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239_1, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246_1,
    new_n1247, new_n1248, new_n1249, new_n1250_1, new_n1251, new_n1252,
    new_n1253_1, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263_1, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278_1, new_n1279, new_n1280, new_n1281_1, new_n1282,
    new_n1283_1, new_n1284, new_n1285_1, new_n1286_1, new_n1287, new_n1290,
    new_n1291, new_n1292_1, new_n1293, new_n1294, new_n1295, new_n1296_1,
    new_n1297, new_n1298, new_n1299_1, new_n1300, new_n1301_1, new_n1303,
    new_n1305_1, new_n1306_1, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1318,
    new_n1319, new_n1320_1, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1328, new_n1329, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1335, new_n1336, new_n1337_1, new_n1338,
    new_n1339, new_n1340, new_n1341, new_n1342, new_n1343, new_n1344,
    new_n1345_1, new_n1346_1, new_n1347, new_n1348, new_n1349, new_n1350_1,
    new_n1351, new_n1352, new_n1353, new_n1354, new_n1355, new_n1356,
    new_n1357, new_n1358, new_n1359_1, new_n1360, new_n1361_1, new_n1362,
    new_n1363, new_n1364, new_n1366, new_n1367, new_n1368_1, new_n1373,
    new_n1374, new_n1375_1, new_n1376, new_n1377, new_n1379, new_n1380,
    new_n1382, new_n1384, new_n1385, new_n1386_1, new_n1387_1, new_n1388,
    new_n1389_1, new_n1390, new_n1391_1, new_n1392, new_n1393_1, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401_1, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411_1, new_n1412,
    new_n1413, new_n1414, new_n1415_1, new_n1416, new_n1417, new_n1418_1,
    new_n1419, new_n1420_1, new_n1421_1, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427_1, new_n1428_1, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435_1, new_n1436,
    new_n1437, new_n1438_1, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443_1, new_n1444, new_n1445, new_n1446_1, new_n1447, new_n1448_1,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1453, new_n1454,
    new_n1455, new_n1457, new_n1458, new_n1459, new_n1460, new_n1461,
    new_n1462, new_n1463_1, new_n1464, new_n1465, new_n1466, new_n1467,
    new_n1468, new_n1469, new_n1470_1, new_n1471, new_n1472, new_n1473,
    new_n1474_1, new_n1475, new_n1476_1, new_n1477, new_n1478, new_n1479,
    new_n1480, new_n1481, new_n1482, new_n1483, new_n1484, new_n1485,
    new_n1486, new_n1487, new_n1488, new_n1489, new_n1490, new_n1491,
    new_n1492, new_n1493, new_n1494, new_n1495, new_n1496, new_n1497,
    new_n1498, new_n1499, new_n1500_1, new_n1501, new_n1502_1, new_n1503,
    new_n1504, new_n1505, new_n1506_1, new_n1507, new_n1508, new_n1509,
    new_n1510, new_n1511, new_n1512, new_n1513, new_n1514, new_n1515,
    new_n1516_1, new_n1517, new_n1518, new_n1519, new_n1520_1, new_n1522,
    new_n1523_1, new_n1524, new_n1525, new_n1526, new_n1527_1, new_n1528,
    new_n1529, new_n1530, new_n1531, new_n1532, new_n1533, new_n1534_1,
    new_n1535, new_n1536_1, new_n1537, new_n1538, new_n1539, new_n1540,
    new_n1541, new_n1542, new_n1543, new_n1544, new_n1545, new_n1546,
    new_n1547_1, new_n1548_1, new_n1549, new_n1550, new_n1551, new_n1552,
    new_n1553, new_n1554, new_n1555, new_n1556, new_n1557, new_n1558,
    new_n1559, new_n1560, new_n1561, new_n1562, new_n1563, new_n1564,
    new_n1565, new_n1566_1, new_n1567, new_n1568, new_n1569_1, new_n1570,
    new_n1571, new_n1572, new_n1573, new_n1574, new_n1575, new_n1576_1,
    new_n1577, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1584, new_n1586_1, new_n1587, new_n1588_1, new_n1589,
    new_n1590, new_n1591, new_n1592_1, new_n1593, new_n1594_1, new_n1595,
    new_n1598, new_n1599, new_n1600, new_n1603, new_n1604, new_n1606,
    new_n1607, new_n1608, new_n1609_1, new_n1610, new_n1612, new_n1613_1,
    new_n1615, new_n1618, new_n1619, new_n1620, new_n1621, new_n1622,
    new_n1623, new_n1624, new_n1625, new_n1626_1, new_n1627_1, new_n1628,
    new_n1629, new_n1630, new_n1631, new_n1632_1, new_n1633, new_n1634,
    new_n1635, new_n1636, new_n1637, new_n1638, new_n1639_1, new_n1640,
    new_n1641, new_n1642, new_n1643, new_n1644_1, new_n1645_1, new_n1646,
    new_n1647_1, new_n1648, new_n1649, new_n1650, new_n1651, new_n1652,
    new_n1653, new_n1654, new_n1655, new_n1656_1, new_n1657, new_n1658,
    new_n1659, new_n1660, new_n1661, new_n1662, new_n1663, new_n1664,
    new_n1665, new_n1666, new_n1667, new_n1668, new_n1671, new_n1675,
    new_n1676, new_n1677, new_n1681, new_n1683, new_n1684;
not_3  g0000(new_n316, n1263);
nand_4 g0001(new_n317, n984, n11);
not_3  g0002(new_n318_1, new_n317);
not_3  g0003(new_n319, n1239);
nor_4  g0004(new_n320, new_n319, n220);
nor_4  g0005(new_n321, new_n320, new_n318_1);
nand_4 g0006(new_n322, new_n321, new_n316);
not_3  g0007(new_n323, new_n321);
nand_4 g0008(new_n324, new_n323, n1263);
nand_4 g0009(new_n325, new_n324, new_n322);
nor_4  g0010(new_n326, new_n319, n391);
nor_4  g0011(new_n327, new_n326, new_n318_1);
not_3  g0012(new_n328, new_n327);
nor_4  g0013(new_n329, new_n328, n346);
not_3  g0014(new_n330, n346);
nor_4  g0015(new_n331, new_n327, new_n330);
nor_4  g0016(new_n332, new_n319, n905);
nor_4  g0017(new_n333, new_n332, new_n318_1);
not_3  g0018(new_n334, new_n333);
nor_4  g0019(new_n335, new_n334, n399);
not_3  g0020(new_n336, n399);
nor_4  g0021(new_n337_1, new_n333, new_n336);
nor_4  g0022(new_n338, n1278, new_n319);
nor_4  g0023(new_n339, new_n338, new_n318_1);
not_3  g0024(new_n340, new_n339);
nor_4  g0025(new_n341_1, new_n340, n980);
not_3  g0026(new_n342, new_n341_1);
nor_4  g0027(new_n343, new_n342, new_n337_1);
nor_4  g0028(new_n344_1, new_n343, new_n335);
nor_4  g0029(new_n345, new_n344_1, new_n331);
nor_4  g0030(new_n346_1, new_n345, new_n329);
not_3  g0031(new_n347, new_n346_1);
not_3  g0032(new_n348, n318);
nor_4  g0033(new_n349, n1435, new_n319);
nor_4  g0034(new_n350, new_n349, new_n318_1);
or_4   g0035(new_n351, new_n350, new_n348);
nand_4 g0036(new_n352_1, new_n350, new_n348);
nand_4 g0037(new_n353, n1415, n1239);
not_3  g0038(new_n354, new_n353);
not_3  g0039(new_n355, n1246);
nor_4  g0040(new_n356, new_n355, n1239);
nor_4  g0041(new_n357, new_n356, new_n354);
nor_4  g0042(new_n358, new_n357, n1345);
not_3  g0043(new_n359, n1345);
not_3  g0044(new_n360, new_n357);
nor_4  g0045(new_n361, new_n360, new_n359);
nor_4  g0046(new_n362_1, new_n361, new_n358);
not_3  g0047(new_n363, new_n362_1);
nand_4 g0048(new_n364_1, n1239, n58);
not_3  g0049(new_n365, new_n364_1);
not_3  g0050(new_n366, n1443);
nor_4  g0051(new_n367, new_n366, n1239);
nor_4  g0052(new_n368, new_n367, new_n365);
xor_3  g0053(new_n369, new_n368, n1616);
not_3  g0054(new_n370_1, new_n369);
not_3  g0055(new_n371, n1446);
nand_4 g0056(new_n372, n1239, n598);
not_3  g0057(new_n373, new_n372);
not_3  g0058(new_n374_1, n1647);
nor_4  g0059(new_n375, new_n374_1, n1239);
nor_4  g0060(new_n376_1, new_n375, new_n373);
not_3  g0061(new_n377, new_n376_1);
nor_4  g0062(new_n378_1, new_n377, new_n371);
nor_4  g0063(new_n379, new_n376_1, n1446);
nor_4  g0064(new_n380_1, new_n379, new_n378_1);
not_3  g0065(new_n381, new_n380_1);
nor_4  g0066(new_n382, new_n381, new_n370_1);
not_3  g0067(new_n383, new_n382);
nor_4  g0068(new_n384, new_n383, new_n363);
not_3  g0069(new_n385, new_n384);
nand_4 g0070(new_n386, n1474, n1239);
not_3  g0071(new_n387, new_n386);
not_3  g0072(new_n388, n1506);
nor_4  g0073(new_n389, new_n388, n1239);
nor_4  g0074(new_n390, new_n389, new_n387);
and_4  g0075(new_n391_1, new_n390, n1592);
nor_4  g0076(new_n392_1, new_n390, n1592);
nor_4  g0077(new_n393, new_n392_1, new_n391_1);
not_3  g0078(new_n394, new_n393);
nor_4  g0079(new_n395, new_n394, new_n385);
not_3  g0080(new_n396_1, new_n395);
nand_4 g0081(new_n397, n1350, n1239);
not_3  g0082(new_n398, new_n397);
not_3  g0083(new_n399_1, n262);
nor_4  g0084(new_n400, n1239, new_n399_1);
nor_4  g0085(new_n401, new_n400, new_n398);
nor_4  g0086(new_n402, new_n401, n1301);
not_3  g0087(new_n403, n1301);
not_3  g0088(new_n404, new_n401);
nor_4  g0089(new_n405, new_n404, new_n403);
nand_4 g0090(new_n406, n1239, n676);
not_3  g0091(new_n407, new_n406);
not_3  g0092(new_n408_1, n1154);
nor_4  g0093(new_n409_1, n1239, new_n408_1);
nor_4  g0094(new_n410, new_n409_1, new_n407);
nor_4  g0095(new_n411, new_n410, n1566);
not_3  g0096(new_n412, n1566);
not_3  g0097(new_n413, new_n410);
nor_4  g0098(new_n414, new_n413, new_n412);
nand_4 g0099(new_n415, n1289, n1239);
not_3  g0100(new_n416_1, new_n415);
not_3  g0101(new_n417_1, n1193);
nor_4  g0102(new_n418, n1239, new_n417_1);
nor_4  g0103(new_n419, new_n418, new_n416_1);
and_4  g0104(new_n420_1, new_n419, n920);
nand_4 g0105(new_n421, n1239, n244);
not_3  g0106(new_n422, new_n421);
not_3  g0107(new_n423, n641);
nor_4  g0108(new_n424, n1239, new_n423);
nor_4  g0109(new_n425, new_n424, new_n422);
nor_4  g0110(new_n426, new_n425, n293);
nor_4  g0111(new_n427, new_n419, n920);
nor_4  g0112(new_n428_1, new_n427, new_n426);
nor_4  g0113(new_n429, new_n428_1, new_n420_1);
not_3  g0114(new_n430_1, new_n429);
nor_4  g0115(new_n431, new_n430_1, new_n414);
nor_4  g0116(new_n432, new_n431, new_n411);
nor_4  g0117(new_n433, new_n432, new_n405);
nor_4  g0118(new_n434, new_n433, new_n402);
not_3  g0119(new_n435, new_n434);
not_3  g0120(new_n436, n293);
not_3  g0121(new_n437, new_n425);
nor_4  g0122(new_n438, new_n437, new_n436);
nor_4  g0123(new_n439, new_n438, new_n426);
nand_4 g0124(new_n440, n1239, n251);
not_3  g0125(new_n441, new_n440);
not_3  g0126(new_n442, n1172);
nor_4  g0127(new_n443, n1239, new_n442);
nor_4  g0128(new_n444, new_n443, new_n441);
and_4  g0129(new_n445, new_n444, n408);
nor_4  g0130(new_n446, new_n444, n408);
not_3  g0131(new_n447, n1476);
nand_4 g0132(new_n448, n1516, n1239);
not_3  g0133(new_n449, new_n448);
not_3  g0134(new_n450, n710);
nor_4  g0135(new_n451, n1239, new_n450);
nor_4  g0136(new_n452, new_n451, new_n449);
not_3  g0137(new_n453_1, new_n452);
nor_4  g0138(new_n454, new_n453_1, new_n447);
nand_4 g0139(new_n455, n1239, n82);
not_3  g0140(new_n456, new_n455);
not_3  g0141(new_n457_1, n1061);
nor_4  g0142(new_n458, n1239, new_n457_1);
nor_4  g0143(new_n459, new_n458, new_n456);
nor_4  g0144(new_n460_1, new_n459, n1401);
not_3  g0145(new_n461, n1401);
not_3  g0146(new_n462, new_n459);
nor_4  g0147(new_n463, new_n462, new_n461);
nor_4  g0148(new_n464, new_n463, new_n460_1);
not_3  g0149(new_n465, new_n464);
nand_4 g0150(new_n466, n1239, n790);
not_3  g0151(new_n467, new_n466);
not_3  g0152(new_n468, n1521);
nor_4  g0153(new_n469, new_n468, n1239);
nor_4  g0154(new_n470, new_n469, new_n467);
and_4  g0155(new_n471, new_n470, n823);
nor_4  g0156(new_n472, new_n470, n823);
nor_4  g0157(new_n473, new_n472, new_n471);
not_3  g0158(new_n474, new_n473);
nand_4 g0159(new_n475, n1576, n1239);
not_3  g0160(new_n476, new_n475);
not_3  g0161(new_n477_1, n1283);
nor_4  g0162(new_n478_1, new_n477_1, n1239);
nor_4  g0163(new_n479, new_n478_1, new_n476);
and_4  g0164(new_n480, new_n479, n153);
nor_4  g0165(new_n481, new_n479, n153);
nor_4  g0166(new_n482, new_n481, new_n480);
not_3  g0167(new_n483, new_n482);
nor_4  g0168(new_n484, new_n483, new_n474);
not_3  g0169(new_n485, new_n484);
nor_4  g0170(new_n486, new_n485, new_n465);
not_3  g0171(new_n487_1, new_n486);
nor_4  g0172(new_n488, new_n487_1, new_n454);
not_3  g0173(new_n489_1, n374);
nand_4 g0174(new_n490, n1239, n645);
not_3  g0175(new_n491, new_n490);
not_3  g0176(new_n492, n87);
nor_4  g0177(new_n493, n1239, new_n492);
nor_4  g0178(new_n494, new_n493, new_n491);
not_3  g0179(new_n495, new_n494);
nor_4  g0180(new_n496, new_n495, new_n489_1);
nand_4 g0181(new_n497_1, new_n495, new_n489_1);
not_3  g0182(new_n498_1, n567);
nand_4 g0183(new_n499, n1239, n268);
not_3  g0184(new_n500, new_n499);
not_3  g0185(new_n501_1, n600);
nor_4  g0186(new_n502_1, n1239, new_n501_1);
nor_4  g0187(new_n503, new_n502_1, new_n500);
not_3  g0188(new_n504, new_n503);
nor_4  g0189(new_n505, new_n504, new_n498_1);
not_3  g0190(new_n506_1, new_n505);
nor_4  g0191(new_n507_1, new_n503, n567);
not_3  g0192(new_n508, new_n507_1);
nand_4 g0193(new_n509_1, n1393, n1239);
not_3  g0194(new_n510_1, new_n509_1);
not_3  g0195(new_n511, n254);
nor_4  g0196(new_n512, n1239, new_n511);
nor_4  g0197(new_n513, new_n512, new_n510_1);
nor_4  g0198(new_n514, new_n513, n1463);
not_3  g0199(new_n515, n1463);
not_3  g0200(new_n516_1, new_n513);
nor_4  g0201(new_n517_1, new_n516_1, new_n515);
nor_4  g0202(new_n518, new_n517_1, new_n514);
nand_4 g0203(new_n519, n1239, n312);
not_3  g0204(new_n520, new_n519);
not_3  g0205(new_n521, n307);
nor_4  g0206(new_n522, n1239, new_n521);
nor_4  g0207(new_n523, new_n522, new_n520);
nor_4  g0208(new_n524, new_n523, n222);
not_3  g0209(new_n525, n222);
not_3  g0210(new_n526, new_n523);
nor_4  g0211(new_n527, new_n526, new_n525);
nor_4  g0212(new_n528, new_n527, new_n524);
nand_4 g0213(new_n529, new_n528, new_n518);
not_3  g0214(new_n530, n608);
nand_4 g0215(new_n531, n1609, n1239);
not_3  g0216(new_n532, new_n531);
not_3  g0217(new_n533, n54);
nor_4  g0218(new_n534_1, n1239, new_n533);
nor_4  g0219(new_n535, new_n534_1, new_n532);
not_3  g0220(new_n536, new_n535);
nor_4  g0221(new_n537, new_n536, new_n530);
not_3  g0222(new_n538, new_n537);
nor_4  g0223(new_n539, new_n535, n608);
not_3  g0224(new_n540, new_n539);
nand_4 g0225(new_n541, n1239, n310);
not_3  g0226(new_n542, new_n541);
not_3  g0227(new_n543, n1175);
nor_4  g0228(new_n544, n1239, new_n543);
nor_4  g0229(new_n545_1, new_n544, new_n542);
nor_4  g0230(new_n546, new_n545_1, n1071);
not_3  g0231(new_n547, new_n546);
not_3  g0232(new_n548, n1071);
not_3  g0233(new_n549, new_n545_1);
nor_4  g0234(new_n550, new_n549, new_n548);
not_3  g0235(new_n551, new_n550);
nand_4 g0236(new_n552, n1239, n219);
not_3  g0237(new_n553_1, new_n552);
not_3  g0238(new_n554, n409);
nor_4  g0239(new_n555, n1239, new_n554);
nor_4  g0240(new_n556, new_n555, new_n553_1);
nor_4  g0241(new_n557, new_n556, n45);
not_3  g0242(new_n558, new_n557);
nand_4 g0243(new_n559_1, new_n556, n45);
not_3  g0244(new_n560_1, n695);
nand_4 g0245(new_n561_1, n1569, n1239);
not_3  g0246(new_n562, n1250);
nor_4  g0247(new_n563, new_n562, n1239);
not_3  g0248(new_n564, new_n563);
nand_4 g0249(new_n565, new_n564, new_n561_1);
nand_4 g0250(new_n566, new_n565, new_n560_1);
not_3  g0251(new_n567_1, new_n561_1);
nor_4  g0252(new_n568, new_n563, new_n567_1);
nand_4 g0253(new_n569, new_n568, n695);
nand_4 g0254(new_n570, new_n319, n510);
nor_4  g0255(new_n571, new_n570, n1205);
nand_4 g0256(new_n572, new_n571, new_n569);
nand_4 g0257(new_n573, new_n572, new_n566);
nand_4 g0258(new_n574_1, new_n573, new_n559_1);
nand_4 g0259(new_n575, new_n574_1, new_n558);
nand_4 g0260(new_n576, new_n575, new_n551);
nand_4 g0261(new_n577, new_n576, new_n547);
not_3  g0262(new_n578, new_n559_1);
nor_4  g0263(new_n579, new_n578, new_n557);
not_3  g0264(new_n580, new_n566);
not_3  g0265(new_n581_1, new_n569);
nor_4  g0266(new_n582_1, new_n581_1, new_n580);
nand_4 g0267(new_n583, new_n582_1, new_n579);
not_3  g0268(new_n584, n545);
not_3  g0269(new_n585_1, new_n571);
nor_4  g0270(new_n586, n1239, n510);
nand_4 g0271(new_n587, new_n586, n1205);
nand_4 g0272(new_n588, new_n587, new_n585_1);
nor_4  g0273(new_n589_1, new_n588, new_n584);
nor_4  g0274(new_n590, new_n550, new_n546);
nand_4 g0275(new_n591, new_n590, new_n589_1);
nor_4  g0276(new_n592, new_n591, new_n583);
nor_4  g0277(new_n593_1, new_n592, new_n577);
nand_4 g0278(new_n594, new_n593_1, new_n540);
nand_4 g0279(new_n595_1, new_n594, new_n538);
nor_4  g0280(new_n596, new_n595_1, new_n529);
not_3  g0281(new_n597_1, new_n524);
nor_4  g0282(new_n598_1, new_n597_1, new_n517_1);
nor_4  g0283(new_n599, new_n598_1, new_n514);
not_3  g0284(new_n600_1, new_n599);
nor_4  g0285(new_n601, new_n600_1, new_n596);
nand_4 g0286(new_n602, new_n601, new_n508);
nand_4 g0287(new_n603, new_n602, new_n506_1);
nand_4 g0288(new_n604, new_n603, new_n497_1);
not_3  g0289(new_n605, new_n604);
nor_4  g0290(new_n606, new_n605, new_n496);
nand_4 g0291(new_n607_1, new_n606, new_n488);
nor_4  g0292(new_n608_1, new_n452, n1476);
not_3  g0293(new_n609_1, new_n460_1);
nor_4  g0294(new_n610, new_n480, new_n609_1);
nor_4  g0295(new_n611, new_n481, new_n472);
not_3  g0296(new_n612, new_n611);
nor_4  g0297(new_n613, new_n612, new_n610);
nor_4  g0298(new_n614, new_n613, new_n471);
nor_4  g0299(new_n615, new_n614, new_n608_1);
nor_4  g0300(new_n616, new_n615, new_n454);
not_3  g0301(new_n617, new_n616);
nand_4 g0302(new_n618, new_n617, new_n607_1);
nor_4  g0303(new_n619, new_n618, new_n446);
nor_4  g0304(new_n620, new_n619, new_n445);
nand_4 g0305(new_n621, new_n620, new_n439);
nor_4  g0306(new_n622, new_n427, new_n420_1);
not_3  g0307(new_n623, new_n622);
nor_4  g0308(new_n624, new_n405, new_n402);
nor_4  g0309(new_n625_1, new_n414, new_n411);
and_4  g0310(new_n626_1, new_n625_1, new_n624);
not_3  g0311(new_n627, new_n626_1);
nor_4  g0312(new_n628, new_n627, new_n623);
not_3  g0313(new_n629, new_n628);
nor_4  g0314(new_n630, new_n629, new_n621);
nor_4  g0315(new_n631, new_n630, new_n435);
nor_4  g0316(new_n632, new_n631, new_n396_1);
not_3  g0317(new_n633, n1616);
not_3  g0318(new_n634, new_n368);
nand_4 g0319(new_n635, new_n634, new_n633);
nor_4  g0320(new_n636, new_n379, new_n358);
not_3  g0321(new_n637, new_n636);
nor_4  g0322(new_n638_1, new_n634, new_n633);
nor_4  g0323(new_n639, new_n378_1, new_n638_1);
nand_4 g0324(new_n640_1, new_n639, new_n637);
nand_4 g0325(new_n641_1, new_n640_1, new_n635);
nor_4  g0326(new_n642, new_n641_1, new_n392_1);
nor_4  g0327(new_n643, new_n642, new_n391_1);
nor_4  g0328(new_n644, new_n643, new_n632);
nand_4 g0329(new_n645_1, new_n644, new_n352_1);
nand_4 g0330(new_n646, new_n645_1, new_n351);
nor_4  g0331(new_n647, new_n331, new_n329);
nor_4  g0332(new_n648, new_n337_1, new_n335);
not_3  g0333(new_n649, new_n648);
xor_3  g0334(new_n650, new_n340, n980);
not_3  g0335(new_n651, new_n650);
nor_4  g0336(new_n652, new_n651, new_n649);
nand_4 g0337(new_n653, new_n652, new_n647);
nor_4  g0338(new_n654, new_n653, new_n646);
nor_4  g0339(new_n655, new_n654, new_n347);
xor_3  g0340(n22, new_n655, new_n325);
not_3  g0341(new_n657, n1361);
nand_4 g0342(n30, n1387, new_n657);
xor_3  g0343(n112, new_n620, new_n439);
nand_4 g0344(new_n660, n1613, n1520);
nand_4 g0345(new_n661, n574, n284);
or_4   g0346(n126, new_n661, new_n660);
nor_4  g0347(new_n663_1, new_n319, n223);
nor_4  g0348(new_n664, new_n663_1, new_n318_1);
not_3  g0349(new_n665, n300);
nor_4  g0350(new_n666, n1239, new_n665);
nor_4  g0351(new_n667, n1470, new_n319);
nor_4  g0352(new_n668, new_n667, new_n666);
not_3  g0353(new_n669_1, new_n668);
nor_4  g0354(new_n670, new_n669_1, new_n664);
nor_4  g0355(new_n671_1, new_n319, n86);
nor_4  g0356(new_n672, new_n671_1, new_n318_1);
not_3  g0357(new_n673, n561);
nor_4  g0358(new_n674, n1239, new_n673);
nor_4  g0359(new_n675, new_n319, n138);
or_4   g0360(new_n676_1, new_n675, new_n674);
nor_4  g0361(new_n677, new_n676_1, new_n672);
nor_4  g0362(new_n678, new_n677, new_n670);
not_3  g0363(new_n679, new_n678);
nand_4 g0364(new_n680, new_n676_1, new_n672);
nor_4  g0365(new_n681, n1299, new_n319);
nor_4  g0366(new_n682, new_n681, new_n318_1);
not_3  g0367(new_n683, n879);
nor_4  g0368(new_n684, n1239, new_n683);
nor_4  g0369(new_n685, new_n319, n769);
nor_4  g0370(new_n686, new_n685, new_n684);
not_3  g0371(new_n687, new_n686);
nand_4 g0372(new_n688, new_n687, new_n682);
nand_4 g0373(new_n689, new_n688, new_n680);
nor_4  g0374(new_n690_1, n1502, new_n319);
nor_4  g0375(new_n691, new_n690_1, new_n318_1);
not_3  g0376(new_n692, n143);
nor_4  g0377(new_n693_1, n1239, new_n692);
nor_4  g0378(new_n694, new_n319, n626);
nor_4  g0379(new_n695_1, new_n694, new_n693_1);
not_3  g0380(new_n696, new_n695_1);
nor_4  g0381(new_n697, new_n696, new_n691);
nor_4  g0382(new_n698, new_n687, new_n682);
nor_4  g0383(new_n699, new_n698, new_n697);
not_3  g0384(new_n700, new_n699);
not_3  g0385(new_n701_1, n663);
nor_4  g0386(new_n702, n1239, new_n701_1);
nor_4  g0387(new_n703, n1656, new_n319);
nor_4  g0388(new_n704, new_n703, new_n702);
nor_4  g0389(new_n705, new_n704, new_n318_1);
not_3  g0390(new_n706, new_n691);
nor_4  g0391(new_n707, new_n695_1, new_n706);
nor_4  g0392(new_n708, new_n707, new_n705);
nor_4  g0393(new_n709, new_n708, new_n700);
nor_4  g0394(new_n710_1, new_n709, new_n689);
nor_4  g0395(new_n711, new_n710_1, new_n679);
nor_4  g0396(new_n712, new_n319, n787);
nor_4  g0397(new_n713, new_n712, new_n318_1);
not_3  g0398(new_n714_1, n1164);
nor_4  g0399(new_n715, n1239, new_n714_1);
nor_4  g0400(new_n716, new_n319, n399);
nor_4  g0401(new_n717, new_n716, new_n715);
not_3  g0402(new_n718, new_n717);
nor_4  g0403(new_n719_1, new_n718, new_n713);
nor_4  g0404(new_n720, new_n319, n727);
nor_4  g0405(new_n721, new_n720, new_n318_1);
not_3  g0406(new_n722, n40);
nor_4  g0407(new_n723, n1239, new_n722);
nor_4  g0408(new_n724, n1263, new_n319);
nor_4  g0409(new_n725, new_n724, new_n723);
not_3  g0410(new_n726_1, new_n725);
nor_4  g0411(new_n727_1, new_n726_1, new_n721);
nor_4  g0412(new_n728, new_n319, n94);
nor_4  g0413(new_n729_1, new_n728, new_n318_1);
not_3  g0414(new_n730, n489);
nor_4  g0415(new_n731, n1239, new_n730);
nor_4  g0416(new_n732, new_n319, n346);
nor_4  g0417(new_n733, new_n732, new_n731);
not_3  g0418(new_n734_1, new_n733);
nor_4  g0419(new_n735, new_n734_1, new_n729_1);
nor_4  g0420(new_n736, new_n735, new_n727_1);
not_3  g0421(new_n737, new_n736);
nor_4  g0422(new_n738, new_n737, new_n719_1);
not_3  g0423(new_n739, new_n738);
not_3  g0424(new_n740, new_n713);
nor_4  g0425(new_n741, new_n717, new_n740);
nor_4  g0426(new_n742_1, new_n319, n609);
nor_4  g0427(new_n743_1, new_n742_1, new_n318_1);
not_3  g0428(new_n744, new_n743_1);
not_3  g0429(new_n745, n71);
nor_4  g0430(new_n746, n1239, new_n745);
nor_4  g0431(new_n747, new_n319, n980);
nor_4  g0432(new_n748, new_n747, new_n746);
nor_4  g0433(new_n749, new_n748, new_n744);
nor_4  g0434(new_n750, new_n749, new_n741);
nor_4  g0435(new_n751, new_n750, new_n739);
not_3  g0436(new_n752, new_n721);
nor_4  g0437(new_n753, new_n725, new_n752);
not_3  g0438(new_n754, new_n729_1);
nor_4  g0439(new_n755_1, new_n733, new_n754);
nor_4  g0440(new_n756, new_n755_1, new_n753);
nor_4  g0441(new_n757, new_n756, new_n727_1);
nor_4  g0442(new_n758, new_n757, new_n751);
nor_4  g0443(new_n759, new_n319, n839);
nor_4  g0444(new_n760, new_n759, new_n318_1);
not_3  g0445(new_n761, new_n760);
not_3  g0446(new_n762, n1523);
nor_4  g0447(new_n763, new_n762, n1239);
nor_4  g0448(new_n764, new_n319, n318);
nor_4  g0449(new_n765, new_n764, new_n763);
nand_4 g0450(new_n766, new_n765, new_n761);
not_3  g0451(new_n767, new_n750);
not_3  g0452(new_n768, new_n748);
nor_4  g0453(new_n769_1, new_n768, new_n743_1);
nor_4  g0454(new_n770, new_n769_1, new_n767);
nand_4 g0455(new_n771, new_n770, new_n738);
nor_4  g0456(new_n772, new_n765, new_n761);
nand_4 g0457(new_n773_1, n1239, n953);
not_3  g0458(new_n774, new_n773_1);
nor_4  g0459(new_n775_1, new_n774, new_n389);
not_3  g0460(new_n776, n1305);
nor_4  g0461(new_n777, new_n776, n1239);
nor_4  g0462(new_n778_1, n1592, new_n319);
nor_4  g0463(new_n779_1, new_n778_1, new_n777);
nor_4  g0464(new_n780, new_n779_1, new_n775_1);
nor_4  g0465(new_n781, new_n780, new_n772);
and_4  g0466(new_n782_1, new_n779_1, new_n775_1);
nand_4 g0467(new_n783, n1239, n52);
not_3  g0468(new_n784, new_n783);
nor_4  g0469(new_n785, new_n784, new_n367);
not_3  g0470(new_n786, n1418);
nor_4  g0471(new_n787_1, new_n786, n1239);
nor_4  g0472(new_n788, n1616, new_n319);
nor_4  g0473(new_n789, new_n788, new_n787_1);
nor_4  g0474(new_n790_1, new_n789, new_n785);
not_3  g0475(new_n791, new_n785);
not_3  g0476(new_n792, new_n789);
nor_4  g0477(new_n793, new_n792, new_n791);
nand_4 g0478(new_n794_1, n1428, n1239);
not_3  g0479(new_n795, new_n794_1);
nor_4  g0480(new_n796, new_n795, new_n375);
not_3  g0481(new_n797, new_n796);
not_3  g0482(new_n798, n1156);
nor_4  g0483(new_n799, n1239, new_n798);
nor_4  g0484(new_n800, n1446, new_n319);
nor_4  g0485(new_n801, new_n800, new_n799);
not_3  g0486(new_n802, new_n801);
nor_4  g0487(new_n803, new_n802, new_n797);
nor_4  g0488(new_n804, new_n803, new_n793);
nor_4  g0489(new_n805, new_n801, new_n796);
nand_4 g0490(new_n806, n1239, n607);
not_3  g0491(new_n807, new_n806);
nor_4  g0492(new_n808, new_n807, new_n356);
not_3  g0493(new_n809, n969);
nor_4  g0494(new_n810, n1239, new_n809);
nor_4  g0495(new_n811, n1345, new_n319);
nor_4  g0496(new_n812, new_n811, new_n810);
nor_4  g0497(new_n813, new_n812, new_n808);
nor_4  g0498(new_n814, new_n813, new_n805);
not_3  g0499(new_n815, new_n814);
and_4  g0500(new_n816, new_n815, new_n804);
nor_4  g0501(new_n817, new_n816, new_n790_1);
or_4   g0502(new_n818, new_n817, new_n782_1);
nand_4 g0503(new_n819, new_n818, new_n781);
nand_4 g0504(new_n820, n1239, n376);
not_3  g0505(new_n821_1, new_n820);
nor_4  g0506(new_n822, new_n821_1, new_n400);
not_3  g0507(new_n823_1, new_n822);
not_3  g0508(new_n824, n779);
nor_4  g0509(new_n825, n1239, new_n824);
nor_4  g0510(new_n826, n1301, new_n319);
nor_4  g0511(new_n827, new_n826, new_n825);
not_3  g0512(new_n828, new_n827);
nor_4  g0513(new_n829, new_n828, new_n823_1);
not_3  g0514(new_n830, new_n829);
nor_4  g0515(new_n831_1, new_n827, new_n822);
nand_4 g0516(new_n832_1, n1239, n273);
not_3  g0517(new_n833, new_n832_1);
nor_4  g0518(new_n834, new_n833, new_n409_1);
not_3  g0519(new_n835, n507);
nor_4  g0520(new_n836, n1239, new_n835);
nor_4  g0521(new_n837, n1566, new_n319);
nor_4  g0522(new_n838, new_n837, new_n836);
nor_4  g0523(new_n839_1, new_n838, new_n834);
nor_4  g0524(new_n840, new_n839_1, new_n831_1);
and_4  g0525(new_n841, new_n838, new_n834);
nand_4 g0526(new_n842_1, n1239, n885);
not_3  g0527(new_n843, new_n842_1);
nor_4  g0528(new_n844, new_n843, new_n418);
not_3  g0529(new_n845, n107);
nor_4  g0530(new_n846, n1239, new_n845);
nor_4  g0531(new_n847, new_n319, n920);
nor_4  g0532(new_n848, new_n847, new_n846);
and_4  g0533(new_n849_1, new_n848, new_n844);
nor_4  g0534(new_n850, new_n849_1, new_n841);
nor_4  g0535(new_n851, new_n848, new_n844);
nand_4 g0536(new_n852, n1239, n50);
not_3  g0537(new_n853, new_n852);
nor_4  g0538(new_n854, new_n853, new_n424);
not_3  g0539(new_n855, n1448);
nor_4  g0540(new_n856, new_n855, n1239);
nor_4  g0541(new_n857, new_n319, n293);
nor_4  g0542(new_n858, new_n857, new_n856);
nor_4  g0543(new_n859, new_n858, new_n854);
nor_4  g0544(new_n860, new_n859, new_n851);
nand_4 g0545(new_n861, n1239, n734);
not_3  g0546(new_n862, new_n861);
nor_4  g0547(new_n863, new_n862, new_n443);
not_3  g0548(new_n864, new_n863);
not_3  g0549(new_n865, n1152);
nor_4  g0550(new_n866, n1239, new_n865);
nor_4  g0551(new_n867, new_n319, n408);
nor_4  g0552(new_n868, new_n867, new_n866);
not_3  g0553(new_n869, new_n868);
nor_4  g0554(new_n870, new_n869, new_n864);
and_4  g0555(new_n871, new_n858, new_n854);
nor_4  g0556(new_n872, new_n871, new_n870);
nand_4 g0557(new_n873, n1586, n1239);
not_3  g0558(new_n874, new_n873);
nor_4  g0559(new_n875, new_n874, new_n451);
not_3  g0560(new_n876, n1386);
nor_4  g0561(new_n877, new_n876, n1239);
nor_4  g0562(new_n878, n1476, new_n319);
nor_4  g0563(new_n879_1, new_n878, new_n877);
nor_4  g0564(new_n880, new_n879_1, new_n875);
not_3  g0565(new_n881, new_n880);
nor_4  g0566(new_n882_1, new_n868, new_n863);
nand_4 g0567(new_n883, n1239, n1114);
not_3  g0568(new_n884, new_n883);
nor_4  g0569(new_n885_1, new_n884, new_n478_1);
not_3  g0570(new_n886, n1627);
nor_4  g0571(new_n887, new_n886, n1239);
nor_4  g0572(new_n888, new_n319, n153);
nor_4  g0573(new_n889, new_n888, new_n887);
nor_4  g0574(new_n890, new_n889, new_n885_1);
nand_4 g0575(new_n891, n1239, n77);
not_3  g0576(new_n892, new_n891);
nor_4  g0577(new_n893, new_n892, new_n469);
not_3  g0578(new_n894_1, n882);
nor_4  g0579(new_n895, n1239, new_n894_1);
nor_4  g0580(new_n896, new_n319, n823);
nor_4  g0581(new_n897, new_n896, new_n895);
nor_4  g0582(new_n898, new_n897, new_n893);
nor_4  g0583(new_n899, new_n898, new_n890);
not_3  g0584(new_n900, new_n899);
nand_4 g0585(new_n901, n1239, n344);
not_3  g0586(new_n902, new_n901);
nor_4  g0587(new_n903, new_n902, new_n458);
not_3  g0588(new_n904, n1227);
nor_4  g0589(new_n905_1, n1239, new_n904);
nor_4  g0590(new_n906, n1401, new_n319);
nor_4  g0591(new_n907, new_n906, new_n905_1);
or_4   g0592(new_n908, new_n907, new_n903);
not_3  g0593(new_n909, new_n885_1);
not_3  g0594(new_n910, new_n889);
nor_4  g0595(new_n911, new_n910, new_n909);
nor_4  g0596(new_n912, new_n911, new_n908);
nor_4  g0597(new_n913, new_n912, new_n900);
and_4  g0598(new_n914, new_n897, new_n893);
and_4  g0599(new_n915, new_n879_1, new_n875);
or_4   g0600(new_n916_1, new_n915, new_n914);
nor_4  g0601(new_n917, new_n916_1, new_n913);
nor_4  g0602(new_n918_1, new_n917, new_n882_1);
nand_4 g0603(new_n919, new_n918_1, new_n881);
nand_4 g0604(new_n920_1, new_n919, new_n872);
nand_4 g0605(new_n921, new_n920_1, new_n860);
nand_4 g0606(new_n922, new_n921, new_n850);
nand_4 g0607(new_n923, new_n922, new_n840);
nand_4 g0608(new_n924, new_n923, new_n830);
nand_4 g0609(new_n925, n1239, n288);
not_3  g0610(new_n926, new_n925);
nor_4  g0611(new_n927, new_n926, new_n502_1);
not_3  g0612(new_n928, new_n927);
not_3  g0613(new_n929, n936);
nor_4  g0614(new_n930, n1239, new_n929);
nor_4  g0615(new_n931, new_n319, n567);
nor_4  g0616(new_n932, new_n931, new_n930);
not_3  g0617(new_n933, new_n932);
nand_4 g0618(new_n934, new_n933, new_n928);
nor_4  g0619(new_n935, new_n933, new_n928);
nand_4 g0620(new_n936_1, n1239, n416);
not_3  g0621(new_n937, new_n936_1);
nor_4  g0622(new_n938, new_n937, new_n512);
not_3  g0623(new_n939, n159);
nor_4  g0624(new_n940, n1239, new_n939);
nor_4  g0625(new_n941, n1463, new_n319);
nor_4  g0626(new_n942, new_n941, new_n940);
or_4   g0627(new_n943, new_n942, new_n938);
nand_4 g0628(new_n944, n1239, n506);
not_3  g0629(new_n945, new_n944);
nor_4  g0630(new_n946, new_n945, new_n522);
not_3  g0631(new_n947_1, n243);
nor_4  g0632(new_n948, n1239, new_n947_1);
nor_4  g0633(new_n949, new_n319, n222);
nor_4  g0634(new_n950, new_n949, new_n948);
nand_4 g0635(new_n951, new_n950, new_n946);
or_4   g0636(new_n952_1, new_n950, new_n946);
nand_4 g0637(new_n953_1, n1239, n671);
not_3  g0638(new_n954, new_n953_1);
nor_4  g0639(new_n955, new_n954, new_n544);
not_3  g0640(new_n956, n341);
nor_4  g0641(new_n957, n1239, new_n956);
nor_4  g0642(new_n958, new_n319, n1071);
nor_4  g0643(new_n959, new_n958, new_n957);
or_4   g0644(new_n960, new_n959, new_n955);
nand_4 g0645(new_n961_1, n1239, n392);
not_3  g0646(new_n962, new_n961_1);
nor_4  g0647(new_n963, new_n962, new_n534_1);
not_3  g0648(new_n964, n742);
nor_4  g0649(new_n965, n1239, new_n964);
nor_4  g0650(new_n966, new_n319, n608);
nor_4  g0651(new_n967, new_n966, new_n965);
nor_4  g0652(new_n968, new_n967, new_n963);
nand_4 g0653(new_n969_1, n1239, n29);
not_3  g0654(new_n970, new_n969_1);
nor_4  g0655(new_n971, new_n970, new_n555);
not_3  g0656(new_n972, new_n971);
not_3  g0657(new_n973, n849);
nor_4  g0658(new_n974, n1239, new_n973);
nor_4  g0659(new_n975, new_n319, n45);
nor_4  g0660(new_n976, new_n975, new_n974);
not_3  g0661(new_n977, new_n976);
nor_4  g0662(new_n978, new_n977, new_n972);
nand_4 g0663(new_n979, n1239, n778);
not_3  g0664(new_n980_1, new_n979);
nor_4  g0665(new_n981, new_n980_1, new_n563);
not_3  g0666(new_n982, n502);
nor_4  g0667(new_n983, n1239, new_n982);
nor_4  g0668(new_n984_1, new_n319, n695);
nor_4  g0669(new_n985, new_n984_1, new_n983);
nand_4 g0670(new_n986_1, new_n985, new_n981);
not_3  g0671(new_n987, n690);
nor_4  g0672(new_n988, n1239, n729);
or_4   g0673(new_n989, new_n988, new_n987);
not_3  g0674(new_n990_1, new_n570);
or_4   g0675(new_n991, n729, n690);
nand_4 g0676(new_n992_1, new_n991, new_n990_1);
nand_4 g0677(new_n993, new_n992_1, new_n989);
nand_4 g0678(new_n994, new_n993, new_n986_1);
nor_4  g0679(new_n995, new_n976, new_n971);
nor_4  g0680(new_n996, new_n985, new_n981);
nor_4  g0681(new_n997_1, new_n996, new_n995);
nand_4 g0682(new_n998, new_n997_1, new_n994);
nand_4 g0683(new_n999, new_n959, new_n955);
nand_4 g0684(new_n1000, new_n999, new_n998);
nor_4  g0685(new_n1001, new_n1000, new_n978);
nor_4  g0686(new_n1002, new_n1001, new_n968);
nand_4 g0687(new_n1003, new_n1002, new_n960);
nand_4 g0688(new_n1004, new_n967, new_n963);
nand_4 g0689(new_n1005, new_n1004, new_n1003);
nand_4 g0690(new_n1006_1, new_n1005, new_n952_1);
nand_4 g0691(new_n1007, new_n1006_1, new_n951);
nand_4 g0692(new_n1008, new_n1007, new_n943);
nand_4 g0693(new_n1009, new_n942, new_n938);
nand_4 g0694(new_n1010, new_n1009, new_n1008);
nor_4  g0695(new_n1011, new_n1010, new_n935);
nand_4 g0696(new_n1012, n1753, n1239);
not_3  g0697(new_n1013, new_n1012);
nor_4  g0698(new_n1014, new_n1013, new_n493);
not_3  g0699(new_n1015, n755);
nor_4  g0700(new_n1016, n1239, new_n1015);
nor_4  g0701(new_n1017_1, new_n319, n374);
nor_4  g0702(new_n1018, new_n1017_1, new_n1016);
nor_4  g0703(new_n1019, new_n1018, new_n1014);
nor_4  g0704(new_n1020, new_n1019, new_n1011);
nand_4 g0705(new_n1021, new_n1020, new_n934);
nand_4 g0706(new_n1022, new_n1018, new_n1014);
nor_4  g0707(new_n1023_1, new_n911, new_n882_1);
nand_4 g0708(new_n1024, new_n1023_1, new_n1022);
nand_4 g0709(new_n1025, new_n872, new_n860);
nor_4  g0710(new_n1026, new_n1025, new_n916_1);
nor_4  g0711(new_n1027, new_n880, new_n829);
nand_4 g0712(new_n1028, new_n1027, new_n840);
and_4  g0713(new_n1029, new_n899, new_n850);
xor_3  g0714(new_n1030, new_n907, new_n903);
nand_4 g0715(new_n1031, new_n1030, new_n1029);
nor_4  g0716(new_n1032, new_n1031, new_n1028);
nand_4 g0717(new_n1033, new_n1032, new_n1026);
nor_4  g0718(new_n1034, new_n1033, new_n1024);
nand_4 g0719(new_n1035, new_n1034, new_n1021);
nand_4 g0720(n1306, new_n1035, new_n924);
nand_4 g0721(new_n1037, new_n812, new_n808);
and_4  g0722(new_n1038, new_n814, new_n781);
nand_4 g0723(new_n1039, new_n1038, new_n1037);
nor_4  g0724(new_n1040_1, new_n790_1, new_n782_1);
nand_4 g0725(new_n1041, new_n1040_1, new_n804);
nor_4  g0726(new_n1042_1, new_n1041, new_n1039);
nand_4 g0727(new_n1043, new_n1042_1, n1306);
not_3  g0728(new_n1044_1, new_n1043);
nor_4  g0729(new_n1045, new_n1044_1, new_n819);
nor_4  g0730(new_n1046, new_n1045, new_n771);
nand_4 g0731(new_n1047, new_n1046, new_n766);
nand_4 g0732(new_n1048, new_n1047, new_n758);
nand_4 g0733(new_n1049, new_n704, new_n318_1);
nand_4 g0734(new_n1050_1, new_n1049, new_n708);
not_3  g0735(new_n1051_1, new_n664);
nor_4  g0736(new_n1052, new_n668, new_n1051_1);
or_4   g0737(new_n1053, new_n1052, new_n700);
nor_4  g0738(new_n1054_1, new_n1053, new_n689);
nand_4 g0739(new_n1055, new_n1054_1, new_n678);
nor_4  g0740(new_n1056, new_n1055, new_n1050_1);
nand_4 g0741(new_n1057, new_n1056, new_n1048);
not_3  g0742(new_n1058_1, n986);
nor_4  g0743(new_n1059, n589, n559);
and_4  g0744(new_n1060_1, new_n1059, n156);
or_4   g0745(new_n1061_1, new_n1060_1, new_n1058_1);
not_3  g0746(new_n1062, new_n1061_1);
nor_4  g0747(new_n1063_1, new_n1062, new_n1052);
nand_4 g0748(new_n1064, new_n1063_1, new_n1057);
nor_4  g0749(new_n1065_1, new_n1064, new_n711);
nand_4 g0750(new_n1066, n589, n559);
nand_4 g0751(new_n1067, new_n1066, n156);
nor_4  g0752(new_n1068, new_n1067, n986);
nor_4  g0753(n161, new_n1068, new_n1065_1);
xor_3  g0754(new_n1070, new_n350, new_n348);
not_3  g0755(new_n1071_1, new_n1070);
xor_3  g0756(n164, new_n1071_1, new_n644);
xor_3  g0757(n181, new_n651, new_n646);
nor_4  g0758(new_n1074, new_n319, n477);
nor_4  g0759(new_n1075, new_n1074, new_n318_1);
not_3  g0760(new_n1076, new_n1075);
nor_4  g0761(new_n1077, new_n1076, n769);
not_3  g0762(new_n1078, n769);
nor_4  g0763(new_n1079, new_n1075, new_n1078);
nor_4  g0764(new_n1080, new_n1079, new_n1077);
not_3  g0765(new_n1081, n626);
nor_4  g0766(new_n1082, new_n319, n1191);
nor_4  g0767(new_n1083, new_n1082, new_n318_1);
nand_4 g0768(new_n1084, new_n1083, new_n1081);
not_3  g0769(new_n1085, new_n1084);
nor_4  g0770(new_n1086, new_n319, n430);
nor_4  g0771(new_n1087, new_n1086, new_n318_1);
not_3  g0772(new_n1088, new_n1087);
nor_4  g0773(new_n1089, new_n1088, n1656);
nor_4  g0774(new_n1090, new_n1089, new_n1085);
nand_4 g0775(new_n1091, new_n655, new_n322);
nand_4 g0776(new_n1092, new_n1091, new_n324);
nand_4 g0777(new_n1093, new_n1092, new_n1090);
nor_4  g0778(new_n1094, new_n1083, new_n1081);
not_3  g0779(new_n1095_1, n1656);
nor_4  g0780(new_n1096, new_n1087, new_n1095_1);
nor_4  g0781(new_n1097, new_n1096, new_n1094);
nor_4  g0782(new_n1098, new_n1097, new_n1085);
not_3  g0783(new_n1099, new_n1098);
nand_4 g0784(new_n1100, new_n1099, new_n1093);
xnor_3 g0785(n216, new_n1100, new_n1080);
not_3  g0786(new_n1102, new_n574_1);
nor_4  g0787(new_n1103_1, new_n573, new_n557);
nor_4  g0788(new_n1104, new_n1103_1, new_n1102);
not_3  g0789(new_n1105, new_n590);
nor_4  g0790(new_n1106, new_n539, new_n537);
xor_3  g0791(new_n1107, new_n1106, new_n1105);
not_3  g0792(new_n1108, new_n1107);
xor_3  g0793(new_n1109, new_n1108, new_n588);
nor_4  g0794(new_n1110, new_n1109, new_n571);
nor_4  g0795(new_n1111, new_n1108, new_n585_1);
nor_4  g0796(new_n1112, new_n1111, new_n1110);
xor_3  g0797(new_n1113, new_n1112, new_n1104);
not_3  g0798(new_n1114_1, new_n577);
xor_3  g0799(new_n1115, new_n582_1, new_n579);
xor_3  g0800(new_n1116, new_n1115, new_n1114_1);
nor_4  g0801(new_n1117, new_n1116, new_n1113);
nand_4 g0802(new_n1118, new_n1116, new_n1113);
nand_4 g0803(new_n1119, new_n1118, new_n584);
nor_4  g0804(new_n1120, new_n1119, new_n1117);
nor_4  g0805(new_n1121_1, new_n587, new_n580);
nor_4  g0806(new_n1122, new_n1121_1, new_n581_1);
xor_3  g0807(new_n1123, new_n1122, new_n1115);
not_3  g0808(new_n1124, new_n587);
nand_4 g0809(new_n1125, new_n1124, new_n575);
not_3  g0810(new_n1126, new_n575);
nor_4  g0811(new_n1127, new_n588, new_n583);
nor_4  g0812(new_n1128, new_n1127, new_n1124);
nand_4 g0813(new_n1129, new_n1128, new_n1126);
nand_4 g0814(new_n1130, new_n1129, new_n1125);
xor_3  g0815(new_n1131, new_n1130, new_n1123);
not_3  g0816(new_n1132, new_n1109);
not_3  g0817(new_n1133, new_n1127);
nor_4  g0818(new_n1134, new_n1133, new_n550);
nor_4  g0819(new_n1135, new_n1134, new_n577);
xor_3  g0820(new_n1136, new_n1135, new_n1132);
nor_4  g0821(new_n1137, new_n1136, new_n1131);
nand_4 g0822(new_n1138_1, new_n1136, new_n1131);
nand_4 g0823(new_n1139, new_n1138_1, n545);
nor_4  g0824(new_n1140, new_n1139, new_n1137);
nor_4  g0825(new_n1141, new_n1140, new_n1120);
nor_4  g0826(new_n1142, new_n599, new_n507_1);
nor_4  g0827(new_n1143, new_n1142, new_n505);
not_3  g0828(new_n1144, new_n529);
not_3  g0829(new_n1145, new_n527);
nor_4  g0830(new_n1146, new_n1145, new_n517_1);
nor_4  g0831(new_n1147, new_n527, new_n514);
nor_4  g0832(new_n1148, new_n1147, new_n1146);
nor_4  g0833(new_n1149, new_n1148, new_n1144);
xor_3  g0834(new_n1150, new_n494, n374);
not_3  g0835(new_n1151, new_n1150);
xor_3  g0836(new_n1152_1, new_n1151, new_n1149);
xor_3  g0837(new_n1153, new_n1152_1, new_n1143);
nand_4 g0838(new_n1154_1, new_n1153, new_n595_1);
not_3  g0839(new_n1155, new_n595_1);
nor_4  g0840(new_n1156_1, new_n600_1, new_n1144);
nor_4  g0841(new_n1157, new_n1156_1, new_n505);
and_4  g0842(new_n1158, new_n1156_1, new_n508);
nor_4  g0843(new_n1159, new_n1158, new_n1157);
nor_4  g0844(new_n1160, new_n524, new_n518);
not_3  g0845(new_n1161, new_n598_1);
nor_4  g0846(new_n1162, new_n1161, new_n514);
nor_4  g0847(new_n1163, new_n1162, new_n1160);
nor_4  g0848(new_n1164_1, new_n507_1, new_n505);
not_3  g0849(new_n1165, new_n1164_1);
xor_3  g0850(new_n1166, new_n1165, new_n1151);
xor_3  g0851(new_n1167, new_n1166, new_n1163);
xor_3  g0852(new_n1168, new_n1167, new_n1159);
nand_4 g0853(new_n1169, new_n1168, new_n1155);
nand_4 g0854(new_n1170, new_n1169, new_n1154_1);
xnor_3 g0855(n233, new_n1170, new_n1141);
xor_3  g0856(new_n1172_1, new_n452, new_n447);
not_3  g0857(new_n1173, new_n606);
nor_4  g0858(new_n1174, new_n1173, new_n465);
nor_4  g0859(new_n1175_1, new_n1174, new_n460_1);
nor_4  g0860(new_n1176, new_n1175_1, new_n483);
nor_4  g0861(new_n1177_1, new_n1176, new_n481);
nor_4  g0862(new_n1178, new_n1177_1, new_n474);
nor_4  g0863(new_n1179, new_n1178, new_n472);
xor_3  g0864(n247, new_n1179, new_n1172_1);
not_3  g0865(n275, n992);
nand_4 g0866(new_n1182, n832, n420);
not_3  g0867(n304, new_n1182);
nor_4  g0868(new_n1184, new_n651, new_n646);
nor_4  g0869(new_n1185, new_n1184, new_n341_1);
nor_4  g0870(new_n1186_1, new_n1185, new_n649);
nor_4  g0871(new_n1187_1, new_n1186_1, new_n335);
xnor_3 g0872(n364, new_n1187_1, new_n647);
nor_4  g0873(new_n1189, new_n446, new_n445);
xor_3  g0874(n370, new_n1189, new_n618);
not_3  g0875(new_n1191_1, new_n1092);
not_3  g0876(new_n1192, n138);
nor_4  g0877(new_n1193_1, n1500, new_n319);
nor_4  g0878(new_n1194, new_n1193_1, new_n318_1);
nor_4  g0879(new_n1195_1, new_n1194, new_n1192);
nor_4  g0880(new_n1196, new_n1084, new_n1079);
nor_4  g0881(new_n1197, new_n1196, new_n1077);
not_3  g0882(new_n1198, new_n1197);
nor_4  g0883(new_n1199, new_n1198, new_n1089);
not_3  g0884(new_n1200, new_n1080);
nor_4  g0885(new_n1201, new_n1094, new_n1085);
not_3  g0886(new_n1202, new_n1201);
nor_4  g0887(new_n1203, new_n1202, new_n1200);
nor_4  g0888(new_n1204, new_n1203, new_n1198);
nor_4  g0889(new_n1205_1, new_n1204, new_n1199);
not_3  g0890(new_n1206, new_n1194);
nor_4  g0891(new_n1207, new_n1206, n138);
nor_4  g0892(new_n1208, new_n1207, new_n1205_1);
nor_4  g0893(new_n1209_1, new_n1208, new_n1195_1);
not_3  g0894(new_n1210, new_n1209_1);
nor_4  g0895(new_n1211_1, new_n1207, new_n1195_1);
nor_4  g0896(new_n1212, new_n319, n582);
nor_4  g0897(new_n1213, new_n1212, new_n318_1);
not_3  g0898(new_n1214, new_n1213);
nor_4  g0899(new_n1215, new_n1214, n1470);
not_3  g0900(new_n1216, n1470);
nor_4  g0901(new_n1217, new_n1213, new_n1216);
nor_4  g0902(new_n1218, new_n1217, new_n1215);
xor_3  g0903(new_n1219, new_n1218, new_n1211_1);
nor_4  g0904(new_n1220, new_n1094, new_n1090);
xor_3  g0905(new_n1221, new_n1220, new_n1219);
xor_3  g0906(new_n1222, new_n1221, new_n1210);
not_3  g0907(new_n1223, new_n1205_1);
not_3  g0908(new_n1224, new_n1211_1);
not_3  g0909(new_n1225_1, new_n1218);
nor_4  g0910(new_n1226, new_n1225_1, new_n1224);
not_3  g0911(new_n1227_1, new_n1226);
nor_4  g0912(new_n1228, new_n1227_1, new_n1223);
not_3  g0913(new_n1229, new_n1207);
nor_4  g0914(new_n1230, new_n1217, new_n1229);
nor_4  g0915(new_n1231_1, new_n1230, new_n1215);
not_3  g0916(new_n1232, new_n1231_1);
nor_4  g0917(new_n1233, new_n1232, new_n1228);
nand_4 g0918(new_n1234_1, n487, n156);
nand_4 g0919(new_n1235, n200, n156);
not_3  g0920(new_n1236, new_n1235);
nor_4  g0921(new_n1237, new_n1236, n986);
xor_3  g0922(new_n1238, new_n1237, new_n1234_1);
and_4  g0923(new_n1239_1, new_n1238, new_n1233);
not_3  g0924(new_n1240, new_n1234_1);
nor_4  g0925(new_n1241, new_n1240, n986);
nor_4  g0926(new_n1242, new_n1235, new_n1058_1);
and_4  g0927(new_n1243, new_n1242, n487);
nor_4  g0928(new_n1244, new_n1243, new_n1241);
not_3  g0929(new_n1245, new_n1244);
nor_4  g0930(new_n1246_1, new_n1236, new_n1240);
nor_4  g0931(new_n1247, new_n1246_1, new_n1245);
not_3  g0932(new_n1248, new_n1247);
nor_4  g0933(new_n1249, new_n1248, new_n1233);
nor_4  g0934(new_n1250_1, new_n1249, new_n1239_1);
xnor_3 g0935(new_n1251, new_n1250_1, new_n1222);
xor_3  g0936(new_n1252, new_n1201, new_n1200);
nor_4  g0937(new_n1253_1, new_n1096, new_n1089);
not_3  g0938(new_n1254, new_n1089);
nor_4  g0939(new_n1255, new_n1204, new_n1254);
nor_4  g0940(new_n1256, new_n1255, new_n1199);
nor_4  g0941(new_n1257, new_n1256, new_n1253_1);
not_3  g0942(new_n1258, new_n1253_1);
nor_4  g0943(new_n1259, new_n1258, new_n1197);
nor_4  g0944(new_n1260, new_n1259, new_n1257);
xor_3  g0945(new_n1261, new_n1260, new_n1252);
xnor_3 g0946(new_n1262, new_n1261, new_n1251);
nor_4  g0947(new_n1263_1, new_n1262, new_n1191_1);
not_3  g0948(new_n1264, new_n1233);
not_3  g0949(new_n1265, new_n1203);
nor_4  g0950(new_n1266, new_n1258, new_n1265);
not_3  g0951(new_n1267, new_n1266);
nor_4  g0952(new_n1268, new_n1267, new_n1224);
not_3  g0953(new_n1269, new_n1268);
nor_4  g0954(new_n1270, new_n1269, new_n1225_1);
nor_4  g0955(new_n1271, new_n1270, new_n1264);
and_4  g0956(new_n1272, new_n1271, new_n1238);
nor_4  g0957(new_n1273, new_n1271, new_n1248);
or_4   g0958(new_n1274, new_n1273, new_n1272);
and_4  g0959(new_n1275, new_n1256, new_n1252);
not_3  g0960(new_n1276, new_n1256);
nand_4 g0961(new_n1277, new_n1267, new_n1252);
and_4  g0962(new_n1278_1, new_n1277, new_n1276);
nor_4  g0963(new_n1279, new_n1278_1, new_n1275);
xor_3  g0964(new_n1280, new_n1279, new_n1219);
nor_4  g0965(new_n1281_1, new_n1210, new_n1099);
nor_4  g0966(new_n1282, new_n1268, new_n1098);
and_4  g0967(new_n1283_1, new_n1282, new_n1210);
nor_4  g0968(new_n1284, new_n1283_1, new_n1281_1);
xnor_3 g0969(new_n1285_1, new_n1284, new_n1280);
xnor_3 g0970(new_n1286_1, new_n1285_1, new_n1274);
nor_4  g0971(new_n1287, new_n1286_1, new_n1092);
nor_4  g0972(n378, new_n1287, new_n1263_1);
xor_3  g0973(n396, new_n1185, new_n649);
nor_4  g0974(new_n1290, new_n1258, new_n1092);
nand_4 g0975(new_n1291, new_n1290, new_n1203);
nand_4 g0976(new_n1292_1, new_n1291, new_n1223);
nand_4 g0977(new_n1293, new_n1292_1, new_n1226);
nand_4 g0978(new_n1294, new_n1293, new_n1231_1);
nand_4 g0979(new_n1295, new_n1294, new_n1238);
nand_4 g0980(new_n1296_1, new_n1253_1, new_n1191_1);
nor_4  g0981(new_n1297, new_n1296_1, new_n1265);
nor_4  g0982(new_n1298, new_n1297, new_n1205_1);
nor_4  g0983(new_n1299_1, new_n1298, new_n1227_1);
nor_4  g0984(new_n1300, new_n1299_1, new_n1232);
nand_4 g0985(new_n1301_1, new_n1300, new_n1248);
nand_4 g0986(n428, new_n1301_1, new_n1295);
nor_4  g0987(new_n1303, new_n1242, new_n1237);
xnor_3 g0988(n453, new_n1303, new_n1294);
or_4   g0989(new_n1305_1, new_n429, new_n411);
nor_4  g0990(new_n1306_1, new_n1305_1, new_n620);
not_3  g0991(new_n1307, new_n432);
not_3  g0992(new_n1308, new_n439);
nor_4  g0993(new_n1309, new_n1308, new_n414);
and_4  g0994(new_n1310, new_n1309, new_n622);
nor_4  g0995(new_n1311, new_n1310, new_n1307);
nor_4  g0996(new_n1312, new_n1311, new_n1306_1);
xor_3  g0997(n517, new_n1312, new_n624);
nor_4  g0998(new_n1314, new_n631, new_n363);
nor_4  g0999(new_n1315, new_n1314, new_n637);
nor_4  g1000(new_n1316, new_n1315, new_n378_1);
xor_3  g1001(n534, new_n1316, new_n369);
nor_4  g1002(new_n1318, new_n1294, new_n1244);
or_4   g1003(new_n1319, new_n1246_1, n986);
not_3  g1004(new_n1320_1, new_n1319);
nor_4  g1005(n553, new_n1320_1, new_n1318);
xor_3  g1006(n597, new_n588, new_n584);
nor_4  g1007(new_n1323, new_n481, new_n460_1);
nor_4  g1008(new_n1324, new_n1323, new_n610);
xor_3  g1009(new_n1325, new_n1324, new_n614);
xor_3  g1010(new_n1326, new_n482, new_n474);
xor_3  g1011(new_n1327, new_n1189, new_n1172_1);
xor_3  g1012(new_n1328, new_n1327, new_n1326);
xor_3  g1013(new_n1329, new_n617, new_n464);
not_3  g1014(new_n1330, new_n1329);
xnor_3 g1015(new_n1331, new_n1330, new_n1328);
xnor_3 g1016(new_n1332, new_n1331, new_n1325);
nand_4 g1017(new_n1333, new_n1332, new_n1173);
nor_4  g1018(new_n1334, new_n1329, new_n488);
xor_3  g1019(new_n1335, new_n614, new_n463);
nor_4  g1020(new_n1336, new_n1335, new_n486);
not_3  g1021(new_n1337_1, new_n463);
nor_4  g1022(new_n1338, new_n481, new_n1337_1);
nor_4  g1023(new_n1339, new_n1338, new_n480);
xnor_3 g1024(new_n1340, new_n1339, new_n1328);
xnor_3 g1025(new_n1341, new_n1340, new_n1336);
xnor_3 g1026(new_n1342, new_n1341, new_n1334);
nand_4 g1027(new_n1343, new_n1342, new_n606);
nand_4 g1028(new_n1344, new_n1343, new_n1333);
xor_3  g1029(new_n1345_1, new_n625_1, new_n624);
not_3  g1030(new_n1346_1, new_n428_1);
not_3  g1031(new_n1347, new_n438);
nor_4  g1032(new_n1348, new_n1347, new_n420_1);
nor_4  g1033(new_n1349, new_n1348, new_n1346_1);
not_3  g1034(new_n1350_1, new_n426);
not_3  g1035(new_n1351, new_n427);
nor_4  g1036(new_n1352, new_n1351, new_n1350_1);
nor_4  g1037(new_n1353, new_n1352, new_n1349);
xor_3  g1038(new_n1354, new_n1353, new_n1345_1);
xor_3  g1039(new_n1355, new_n1354, new_n1311);
nand_4 g1040(new_n1356, new_n1355, new_n620);
not_3  g1041(new_n1357, new_n620);
xor_3  g1042(new_n1358, new_n623, new_n438);
not_3  g1043(new_n1359_1, new_n431);
nand_4 g1044(new_n1360, new_n1305_1, new_n1359_1);
xnor_3 g1045(new_n1361_1, new_n1360, new_n1345_1);
xor_3  g1046(new_n1362, new_n1361_1, new_n1358);
nand_4 g1047(new_n1363, new_n1362, new_n1357);
nand_4 g1048(new_n1364, new_n1363, new_n1356);
xnor_3 g1049(n625, new_n1364, new_n1344);
nand_4 g1050(new_n1366, n1536, n1438);
nand_4 g1051(new_n1367, n997, n315);
nor_4  g1052(new_n1368_1, new_n1367, new_n1366);
not_3  g1053(n669, new_n1368_1);
xor_3  g1054(n693, new_n1175_1, new_n483);
xor_3  g1055(n714, new_n1151, new_n603);
or_4   g1056(n719, n1361, n1225);
not_3  g1057(new_n1373, new_n579);
not_3  g1058(new_n1374, new_n582_1);
nor_4  g1059(new_n1375_1, new_n589_1, new_n571);
nor_4  g1060(new_n1376, new_n1375_1, new_n1374);
nor_4  g1061(new_n1377, new_n1376, new_n580);
xor_3  g1062(n794, new_n1377, new_n1373);
nand_4 g1063(new_n1379, new_n1316, new_n369);
nand_4 g1064(new_n1380, new_n1379, new_n635);
xor_3  g1065(n894, new_n1380, new_n393);
nor_4  g1066(new_n1382, new_n1253_1, new_n1191_1);
nor_4  g1067(n916, new_n1382, new_n1290);
nand_4 g1068(new_n1384, n1411, n1239);
nand_4 g1069(new_n1385, new_n1384, new_n570);
xor_3  g1070(new_n1386_1, new_n1385, new_n981);
xor_3  g1071(new_n1387_1, new_n971, new_n938);
xor_3  g1072(new_n1388, new_n1387_1, new_n1386_1);
xor_3  g1073(new_n1389_1, new_n1388, new_n963);
xor_3  g1074(new_n1390, new_n955, new_n946);
not_3  g1075(new_n1391_1, n299);
nor_4  g1076(new_n1392, n1239, new_n1391_1);
nand_4 g1077(new_n1393_1, n1239, n1044);
not_3  g1078(new_n1394, new_n1393_1);
nor_4  g1079(new_n1395, new_n1394, new_n1392);
xor_3  g1080(new_n1396, new_n1014, new_n927);
xor_3  g1081(new_n1397, new_n1396, new_n1395);
xor_3  g1082(new_n1398, new_n1397, new_n1390);
nor_4  g1083(new_n1399, new_n1398, new_n1389_1);
and_4  g1084(new_n1400, new_n1398, new_n1389_1);
nor_4  g1085(new_n1401_1, new_n1400, new_n1399);
nor_4  g1086(new_n1402, new_n318_1, new_n319);
not_3  g1087(new_n1403, n56);
xor_3  g1088(new_n1404, n1389, n246);
xor_3  g1089(new_n1405, new_n1404, new_n1403);
and_4  g1090(new_n1406, new_n1405, new_n1402);
and_4  g1091(new_n1407, new_n690_1, new_n682);
not_3  g1092(new_n1408, new_n681);
nor_4  g1093(new_n1409, new_n706, new_n1408);
nor_4  g1094(new_n1410, new_n1409, new_n1407);
not_3  g1095(new_n1411_1, new_n671_1);
nor_4  g1096(new_n1412, new_n1411_1, new_n1051_1);
and_4  g1097(new_n1413, new_n672, new_n663_1);
nor_4  g1098(new_n1414, new_n1413, new_n1412);
xor_3  g1099(new_n1415_1, new_n1414, new_n1410);
xor_3  g1100(new_n1416, new_n1415_1, new_n1406);
nor_4  g1101(new_n1417, new_n1416, new_n1401_1);
not_3  g1102(new_n1418_1, new_n712);
nor_4  g1103(new_n1419, new_n744, new_n1418_1);
not_3  g1104(new_n1420_1, new_n742_1);
nor_4  g1105(new_n1421_1, new_n1420_1, new_n740);
nor_4  g1106(new_n1422, new_n1421_1, new_n1419);
not_3  g1107(new_n1423, n1103);
nor_4  g1108(new_n1424, n1239, new_n1423);
nand_4 g1109(new_n1425, n1239, n1023);
not_3  g1110(new_n1426, new_n1425);
nor_4  g1111(new_n1427_1, new_n1426, new_n1424);
xor_3  g1112(new_n1428_1, new_n1427_1, new_n808);
xor_3  g1113(new_n1429, new_n1428_1, new_n1422);
xor_3  g1114(new_n1430, new_n797, new_n785);
not_3  g1115(new_n1431, new_n728);
nor_4  g1116(new_n1432, new_n1431, new_n752);
not_3  g1117(new_n1433, new_n720);
nor_4  g1118(new_n1434, new_n754, new_n1433);
nor_4  g1119(new_n1435_1, new_n1434, new_n1432);
xor_3  g1120(new_n1436, new_n775_1, new_n760);
xor_3  g1121(new_n1437, new_n1436, new_n1435_1);
xor_3  g1122(new_n1438_1, new_n1437, new_n1430);
xnor_3 g1123(new_n1439, new_n1438_1, new_n1429);
xor_3  g1124(new_n1440, new_n854, new_n834);
not_3  g1125(new_n1441, n1121);
nor_4  g1126(new_n1442, n1239, new_n1441);
nand_4 g1127(new_n1443_1, n1239, n560);
not_3  g1128(new_n1444, new_n1443_1);
nor_4  g1129(new_n1445, new_n1444, new_n1442);
xor_3  g1130(new_n1446_1, new_n1445, new_n909);
xor_3  g1131(new_n1447, new_n1446_1, new_n1440);
xor_3  g1132(new_n1448_1, new_n903, new_n864);
xor_3  g1133(new_n1449, new_n1448_1, new_n1447);
not_3  g1134(new_n1450, new_n893);
xor_3  g1135(new_n1451, new_n1450, new_n844);
xor_3  g1136(new_n1452, new_n1451, new_n875);
xor_3  g1137(new_n1453, new_n1452, new_n823_1);
xnor_3 g1138(new_n1454, new_n1453, new_n1449);
nor_4  g1139(new_n1455, new_n1454, new_n1439);
nand_4 g1140(n1375, new_n1455, new_n1417);
xor_3  g1141(new_n1457, new_n479, new_n459);
xor_3  g1142(new_n1458, new_n444, new_n413);
xor_3  g1143(new_n1459, new_n1458, new_n1457);
xor_3  g1144(new_n1460, new_n1459, new_n419);
xor_3  g1145(new_n1461, new_n452, new_n401);
nand_4 g1146(new_n1462, n1239, n314);
not_3  g1147(new_n1463_1, new_n1462);
nor_4  g1148(new_n1464, new_n1463_1, new_n1442);
xor_3  g1149(new_n1465, new_n470, new_n437);
xor_3  g1150(new_n1466, new_n1465, new_n1464);
xor_3  g1151(new_n1467, new_n1466, new_n1461);
xnor_3 g1152(new_n1468, new_n1467, new_n1460);
xor_3  g1153(new_n1469, new_n503, new_n495);
xor_3  g1154(new_n1470_1, new_n523, new_n513);
xor_3  g1155(new_n1471, new_n1470_1, new_n1469);
nand_4 g1156(new_n1472, n1281, n1239);
not_3  g1157(new_n1473, new_n1472);
nor_4  g1158(new_n1474_1, new_n1473, new_n1392);
nand_4 g1159(new_n1475, n1239, n961);
not_3  g1160(new_n1476_1, new_n1475);
nor_4  g1161(new_n1477, new_n1476_1, new_n990_1);
xor_3  g1162(new_n1478, new_n1477, new_n1474_1);
xor_3  g1163(new_n1479, new_n556, new_n549);
xor_3  g1164(new_n1480, new_n1479, new_n1478);
xor_3  g1165(new_n1481, new_n568, new_n535);
xor_3  g1166(new_n1482, new_n1481, new_n1480);
xnor_3 g1167(new_n1483, new_n1482, new_n1471);
nor_4  g1168(new_n1484, new_n1483, new_n1468);
not_3  g1169(new_n1485, new_n320);
nor_4  g1170(new_n1486, new_n328, new_n1485);
not_3  g1171(new_n1487, new_n326);
nor_4  g1172(new_n1488, new_n1487, new_n323);
nor_4  g1173(new_n1489, new_n1488, new_n1486);
xor_3  g1174(new_n1490, new_n634, new_n350);
xor_3  g1175(new_n1491, new_n1490, new_n1489);
xor_3  g1176(new_n1492, new_n390, new_n376_1);
not_3  g1177(new_n1493, new_n332);
nor_4  g1178(new_n1494, new_n340, new_n1493);
not_3  g1179(new_n1495, new_n338);
nor_4  g1180(new_n1496, new_n1495, new_n334);
nor_4  g1181(new_n1497, new_n1496, new_n1494);
nand_4 g1182(new_n1498, n1239, n117);
not_3  g1183(new_n1499, new_n1498);
nor_4  g1184(new_n1500_1, new_n1499, new_n1424);
xor_3  g1185(new_n1501, new_n1500_1, new_n357);
xor_3  g1186(new_n1502_1, new_n1501, new_n1497);
xor_3  g1187(new_n1503, new_n1502_1, new_n1492);
xnor_3 g1188(new_n1504, new_n1503, new_n1491);
not_3  g1189(new_n1505, n430);
xor_3  g1190(new_n1506_1, n1626, n775);
xor_3  g1191(new_n1507, new_n1506_1, new_n1505);
and_4  g1192(new_n1508, new_n1507, new_n1402);
not_3  g1193(new_n1509, new_n1212);
nor_4  g1194(new_n1510, new_n1509, new_n1206);
not_3  g1195(new_n1511, new_n1193_1);
nor_4  g1196(new_n1512, new_n1214, new_n1511);
nor_4  g1197(new_n1513, new_n1512, new_n1510);
and_4  g1198(new_n1514, new_n1083, new_n1074);
not_3  g1199(new_n1515, new_n1082);
nor_4  g1200(new_n1516_1, new_n1515, new_n1076);
nor_4  g1201(new_n1517, new_n1516_1, new_n1514);
xor_3  g1202(new_n1518, new_n1517, new_n1513);
xor_3  g1203(new_n1519, new_n1518, new_n1508);
nor_4  g1204(new_n1520_1, new_n1519, new_n1504);
nand_4 g1205(n1288, new_n1520_1, new_n1484);
nor_4  g1206(new_n1522, n1288, n1375);
not_3  g1207(new_n1523_1, n1346);
nor_4  g1208(new_n1524, new_n1523_1, n1239);
nor_4  g1209(new_n1525, new_n319, n831);
nor_4  g1210(new_n1526, new_n1525, new_n1524);
xor_3  g1211(new_n1527_1, new_n695_1, new_n686);
xor_3  g1212(new_n1528, new_n1527_1, new_n1526);
not_3  g1213(new_n1529, new_n1066);
nor_4  g1214(new_n1530, new_n1529, new_n1059);
nor_4  g1215(new_n1531, new_n1530, n1239);
xor_3  g1216(new_n1532, n487, n200);
nor_4  g1217(new_n1533, new_n1532, new_n319);
or_4   g1218(new_n1534_1, new_n1533, new_n1531);
not_3  g1219(new_n1535, new_n1534_1);
xor_3  g1220(new_n1536_1, new_n676_1, new_n668);
xor_3  g1221(new_n1537, new_n1536_1, new_n704);
xnor_3 g1222(new_n1538, new_n1537, new_n1535);
xnor_3 g1223(new_n1539, new_n1538, new_n1528);
nand_4 g1224(new_n1540, n1239, n21);
not_3  g1225(new_n1541, new_n1540);
nor_4  g1226(new_n1542, n1644, n1239);
nor_4  g1227(new_n1543, new_n1542, new_n1541);
xor_3  g1228(new_n1544, new_n1543, new_n779_1);
xor_3  g1229(new_n1545, new_n765, new_n734_1);
xor_3  g1230(new_n1546, new_n1545, new_n1544);
xor_3  g1231(new_n1547_1, new_n792, new_n717);
xor_3  g1232(new_n1548_1, new_n812, new_n801);
xor_3  g1233(new_n1549, new_n1548_1, new_n1547_1);
xor_3  g1234(new_n1550, new_n748, new_n726_1);
xor_3  g1235(new_n1551, new_n1550, new_n1549);
xnor_3 g1236(new_n1552, new_n1551, new_n1546);
nor_4  g1237(new_n1553, new_n1552, new_n1539);
nand_4 g1238(new_n1554, n1239, n947);
not_3  g1239(new_n1555, new_n1554);
nor_4  g1240(new_n1556, n1750, n1239);
nor_4  g1241(new_n1557, new_n1556, new_n1555);
xor_3  g1242(new_n1558, new_n1557, new_n879_1);
xor_3  g1243(new_n1559, new_n897, new_n869);
xor_3  g1244(new_n1560, new_n858, new_n838);
xor_3  g1245(new_n1561, new_n1560, new_n1559);
xor_3  g1246(new_n1562, new_n907, new_n910);
xor_3  g1247(new_n1563, new_n848, new_n827);
xor_3  g1248(new_n1564, new_n1563, new_n1562);
xnor_3 g1249(new_n1565, new_n1564, new_n1561);
xnor_3 g1250(new_n1566_1, new_n1565, new_n1558);
nand_4 g1251(new_n1567, n1239, n1205);
not_3  g1252(new_n1568, new_n1567);
nor_4  g1253(new_n1569_1, new_n1568, new_n988);
xor_3  g1254(new_n1570, new_n1569_1, new_n1018);
not_3  g1255(new_n1571, new_n942);
nand_4 g1256(new_n1572, n1239, n1138);
not_3  g1257(new_n1573, new_n1572);
nor_4  g1258(new_n1574, n1239, n155);
nor_4  g1259(new_n1575, new_n1574, new_n1573);
xor_3  g1260(new_n1576_1, new_n1575, new_n1571);
xor_3  g1261(new_n1577, new_n1576_1, new_n1570);
xor_3  g1262(new_n1578, new_n985, new_n977);
xor_3  g1263(new_n1579, new_n967, new_n959);
xor_3  g1264(new_n1580, new_n1579, new_n1578);
xor_3  g1265(new_n1581, new_n950, new_n932);
xor_3  g1266(new_n1582, new_n1581, new_n1580);
xnor_3 g1267(new_n1583, new_n1582, new_n1577);
nor_4  g1268(new_n1584, new_n1583, new_n1566_1);
nand_4 g1269(n1322, new_n1584, new_n1553);
nand_4 g1270(new_n1586_1, n1095, n743);
nand_4 g1271(new_n1587, n581, n478);
nor_4  g1272(new_n1588_1, new_n1587, new_n1586_1);
nand_4 g1273(new_n1589, n1286, n1054);
nand_4 g1274(new_n1590, n1040, n593);
nor_4  g1275(new_n1591, new_n1590, new_n1589);
nand_4 g1276(new_n1592_1, new_n1591, new_n1368_1);
nor_4  g1277(new_n1593, new_n1592_1, n126);
nand_4 g1278(new_n1594_1, new_n1593, new_n1588_1);
nor_4  g1279(new_n1595, new_n1594_1, n1322);
nand_4 g1280(n918, new_n1595, new_n1522);
xor_3  g1281(n952, new_n1177_1, new_n474);
not_3  g1282(new_n1598, new_n1195_1);
nand_4 g1283(new_n1599, new_n1291, new_n1208);
nand_4 g1284(new_n1600, new_n1599, new_n1598);
xnor_3 g1285(n990, new_n1600, new_n1218);
xor_3  g1286(n1006, new_n1155, new_n528);
not_3  g1287(new_n1603, n380);
nor_4  g1288(new_n1604, n1361, new_n1603);
nand_4 g1289(n1050, new_n1604, n701);
not_3  g1290(new_n1606, new_n378_1);
nand_4 g1291(new_n1607, new_n1315, new_n1606);
nor_4  g1292(new_n1608, new_n1314, new_n358);
nor_4  g1293(new_n1609_1, new_n1608, new_n380_1);
not_3  g1294(new_n1610, new_n1609_1);
nand_4 g1295(n1051, new_n1610, new_n1607);
nor_4  g1296(new_n1612, new_n1377, new_n1373);
nor_4  g1297(new_n1613_1, new_n1612, new_n557);
xor_3  g1298(n1058, new_n1613_1, new_n1105);
nand_4 g1299(new_n1615, new_n621, new_n1350_1);
xor_3  g1300(n1060, new_n1615, new_n622);
xor_3  g1301(n1063, new_n606, new_n464);
not_3  g1302(new_n1618, new_n631);
xor_3  g1303(new_n1619, new_n380_1, new_n370_1);
xor_3  g1304(new_n1620, new_n1071_1, new_n393);
xor_3  g1305(new_n1621, new_n1620, new_n1619);
not_3  g1306(new_n1622, new_n1621);
not_3  g1307(new_n1623, new_n358);
nor_4  g1308(new_n1624, new_n378_1, new_n1623);
nor_4  g1309(new_n1625, new_n1624, new_n636);
xor_3  g1310(new_n1626_1, new_n1625, new_n641_1);
xor_3  g1311(new_n1627_1, new_n1626_1, new_n1622);
xor_3  g1312(new_n1628, new_n643, new_n363);
xor_3  g1313(new_n1629, new_n1628, new_n1627_1);
nor_4  g1314(new_n1630, new_n1629, new_n1618);
xor_3  g1315(new_n1631, new_n641_1, new_n361);
nor_4  g1316(new_n1632_1, new_n1631, new_n384);
nand_4 g1317(new_n1633, new_n1632_1, new_n1628);
not_3  g1318(new_n1634, new_n1628);
nor_4  g1319(new_n1635, new_n1632_1, new_n395);
nand_4 g1320(new_n1636, new_n1635, new_n1634);
nand_4 g1321(new_n1637, new_n1636, new_n1633);
not_3  g1322(new_n1638, new_n361);
nor_4  g1323(new_n1639_1, new_n379, new_n1638);
nor_4  g1324(new_n1640, new_n1639_1, new_n378_1);
xor_3  g1325(new_n1641, new_n1640, new_n1622);
xor_3  g1326(new_n1642, new_n1641, new_n1637);
nor_4  g1327(new_n1643, new_n1642, new_n631);
nor_4  g1328(new_n1644_1, new_n1643, new_n1630);
not_3  g1329(new_n1645_1, new_n335);
nor_4  g1330(new_n1646, new_n650, new_n1645_1);
not_3  g1331(new_n1647_1, new_n344_1);
nor_4  g1332(new_n1648, new_n652, new_n1647_1);
not_3  g1333(new_n1649, new_n1648);
and_4  g1334(new_n1650, new_n651, new_n337_1);
nor_4  g1335(new_n1651, new_n1650, new_n1649);
nor_4  g1336(new_n1652, new_n1651, new_n1646);
xor_3  g1337(new_n1653, new_n647, new_n325);
xor_3  g1338(new_n1654, new_n1653, new_n342);
not_3  g1339(new_n1655, new_n1654);
xor_3  g1340(new_n1656_1, new_n1655, new_n1652);
xor_3  g1341(new_n1657, new_n1656_1, new_n347);
nand_4 g1342(new_n1658, new_n1657, new_n646);
not_3  g1343(new_n1659, new_n329);
nor_4  g1344(new_n1660, new_n1649, new_n1659);
not_3  g1345(new_n1661, new_n331);
nor_4  g1346(new_n1662, new_n1648, new_n1661);
nor_4  g1347(new_n1663, new_n1662, new_n1660);
xor_3  g1348(new_n1664, new_n1663, new_n1655);
xor_3  g1349(new_n1665, new_n1664, new_n648);
nor_4  g1350(new_n1666, new_n1665, new_n646);
not_3  g1351(new_n1667, new_n1666);
nand_4 g1352(new_n1668, new_n1667, new_n1658);
xnor_3 g1353(n1065, new_n1668, new_n1644_1);
xor_3  g1354(n1195, new_n1165, new_n601);
nor_4  g1355(new_n1671, new_n1290, new_n1089);
xnor_3 g1356(n1302, new_n1671, new_n1201);
xnor_3 g1357(n1391, new_n1292_1, new_n1224);
xor_3  g1358(n1420, new_n1375_1, new_n1374);
nand_4 g1359(new_n1675, new_n1155, new_n528);
and_4  g1360(new_n1676, new_n1675, new_n1160);
or_4   g1361(new_n1677, new_n1676, new_n596);
nor_4  g1362(n1427, new_n1677, new_n1162);
xor_3  g1363(n1527, new_n631, new_n363);
not_3  g1364(n1594, new_n1591);
not_3  g1365(new_n1681, new_n593_1);
xor_3  g1366(n1639, new_n1106, new_n1681);
nor_4  g1367(new_n1683, new_n1615, new_n623);
nor_4  g1368(new_n1684, new_n1683, new_n420_1);
xor_3  g1369(n1687, new_n1684, new_n625_1);
not_3  g1370(n1752, new_n1588_1);
buf_2  g1371(n23, n346);
buf_2  g1372(n27, n947);
buf_2  g1373(n85, n153);
buf_2  g1374(n130, n1592);
buf_2  g1375(n173, n823);
buf_2  g1376(n184, n420);
buf_2  g1377(n230, n831);
buf_2  g1378(n292, n408);
buf_2  g1379(n301, n318);
buf_2  g1380(n337, n626);
buf_2  g1381(n352, n1463);
nand_4 g1382(n362, n1387, new_n657);
buf_2  g1383(n417, n399);
nor_4  g1384(n457, new_n1068, new_n1065_1);
buf_2  g1385(n460, n21);
buf_2  g1386(n497, n1656);
buf_2  g1387(n498, n293);
buf_2  g1388(n501, n200);
buf_2  g1389(n509, n769);
buf_2  g1390(n516, n1187);
nor_4  g1391(n585, new_n1320_1, new_n1318);
buf_2  g1392(n595, n1301);
buf_2  g1393(n638, n420);
buf_2  g1394(n640, n1345);
not_3  g1395(n726, n992);
buf_2  g1396(n773, n980);
buf_2  g1397(n782, n222);
buf_2  g1398(n821, n374);
buf_2  g1399(n842, n1205);
buf_2  g1400(n1017, n1476);
buf_2  g1401(n1042, n1566);
buf_2  g1402(n1177, n487);
nor_4  g1403(n1186, new_n1320_1, new_n1318);
buf_2  g1404(n1209, n1071);
nor_4  g1405(n1211, new_n1068, new_n1065_1);
buf_2  g1406(n1231, n1470);
buf_2  g1407(n1234, n608);
nand_4 g1408(n1253, new_n1604, n701);
buf_2  g1409(n1285, n1401);
buf_2  g1410(n1292, n1616);
not_3  g1411(n1296, n992);
buf_2  g1412(n1320, n1263);
buf_2  g1413(n1337, n1138);
xnor_3 g1414(n1359, new_n1303, new_n1294);
buf_2  g1415(n1368, n420);
buf_2  g1416(n1421, n695);
buf_2  g1417(n1534, n920);
buf_2  g1418(n1547, n420);
buf_2  g1419(n1548, n567);
nand_4 g1420(n1588, new_n1301_1, new_n1295);
nor_4  g1421(n1632, new_n1320_1, new_n1318);
buf_2  g1422(n1645, n1446);
buf_2  g1423(n1729, n138);
buf_2  g1424(n1738, n45);
endmodule


