
module top_810026173_826291639_946996917_1246901 (n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213, n223, n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414, n424, n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649, n653, n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788, n801, n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968, n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332, n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530, n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747, n1757, n1763, n1764, n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156, n174, n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299, n317, n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457, n460, n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547, n549, n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648, n665, n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773, n790, n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888, n891, n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989, n991, n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103, n1113, n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183, n1191, n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255, n1260, n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347, n1348, n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426, n1440, n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502, n1507, n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633, n1635, n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690, n1721, n1727, n1729, n1731, n1737, n1746);
input n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213, n223, n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414, n424, n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649, n653, n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788, n801, n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968, n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332, n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530, n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747, n1757, n1763, n1764;
output n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156, n174, n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299, n317, n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457, n460, n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547, n549, n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648, n665, n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773, n790, n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888, n891, n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989, n991, n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103, n1113, n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183, n1191, n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255, n1260, n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347, n1348, n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426, n1440, n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502, n1507, n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633, n1635, n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690, n1721, n1727, n1729, n1731, n1737, n1746;
wire n0, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n16, n18, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n34, n35, n37, n38, n39, n40, n41, n42, n43, n45, n47, n48, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61, n62, n63, n64, n65, n68, n70, n71, n72, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n127, n128, n129, n130, n131, n132, n133, n134, n136, n137, n138, n139, n140, n141, n142, n143, n144, n146, n147, n148, n149, n150, n151, n152, n153, n154, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n172, n173, n175, n176, n177, n178, n179, n180, n182, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n209, n210, n211, n212, n214, n215, n217, n219, n220, n221, n222, n224, n225, n226, n227, n228, n229, n230, n232, n233, n234, n235, n236, n237, n239, n240, n241, n242, n243, n244, n245, n246, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268, n269, n271, n272, n273, n274, n275, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n291, n293, n294, n295, n296, n297, n298, n300, n301, n302, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n348, n349, n350, n351, n352, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n373, n374, n375, n376, n377, n380, n381, n382, n383, n384, n385, n386, n388, n389, n390, n392, n393, n394, n395, n396, n397, n398, n399, n400, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n415, n417, n418, n419, n420, n421, n422, n425, n427, n428, n430, n431, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n445, n446, n447, n448, n449, n450, n451, n453, n454, n455, n456, n458, n459, n461, n462, n463, n464, n465, n466, n467, n468, n470, n471, n473, n474, n475, n477, n478, n479, n480, n481, n483, n484, n485, n486, n487, n489, n490, n491, n492, n494, n495, n496, n497, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n511, n512, n513, n514, n515, n516, n518, n519, n520, n521, n523, n524, n525, n526, n527, n528, n529, n530, n531, n533, n535, n536, n537, n538, n539, n540, n542, n543, n544, n545, n546, n548, n550, n551, n552, n553, n554, n556, n558, n560, n561, n562, n563, n564, n565, n566, n567, n568, n570, n571, n572, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n586, n587, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n601, n602, n603, n604, n605, n606, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n639, n640, n641, n642, n644, n645, n650, n651, n652, n654, n656, n657, n658, n659, n660, n661, n662, n663, n664, n666, n667, n668, n669, n670, n671, n672, n673, n674, n676, n677, n678, n679, n680, n681, n685, n686, n687, n688, n689, n690, n691, n692, n694, n696, n697, n698, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n713, n714, n716, n717, n718, n719, n720, n721, n722, n723, n726, n727, n728, n730, n732, n733, n734, n735, n736, n737, n739, n740, n741, n742, n743, n744, n745, n746, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n760, n762, n763, n764, n765, n766, n767, n768, n769, n771, n772, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n789, n791, n793, n794, n795, n796, n797, n798, n799, n800, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n814, n815, n816, n817, n818, n819, n820, n821, n822, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n837, n838, n840, n841, n842, n843, n844, n845, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n859, n860, n861, n863, n864, n866, n868, n869, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n884, n885, n886, n887, n889, n890, n893, n894, n895, n896, n897, n898, n899, n900, n901, n903, n904, n907, n908, n909, n910, n911, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n928, n929, n930, n932, n933, n934, n936, n937, n938, n939, n940, n941, n943, n945, n946, n947, n948, n949, n950, n951, n954, n955, n956, n957, n958, n959, n960, n962, n963, n964, n965, n966, n967, n969, n970, n971, n972, n973, n975, n976, n977, n978, n981, n982, n983, n984, n985, n986, n987, n988, n990, n992, n993, n994, n995, n996, n997, n998, n999, n1001, n1002, n1003, n1004, n1006, n1007, n1008, n1009, n1010, n1011, n1013, n1014, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1026, n1027, n1028, n1029, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1063, n1064, n1065, n1066, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1114, n1115, n1116, n1117, n1118, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1136, n1137, n1139, n1141, n1143, n1144, n1146, n1147, n1148, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1173, n1174, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1192, n1193, n1195, n1196, n1197, n1198, n1200, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1236, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1250, n1251, n1252, n1253, n1254, n1256, n1257, n1258, n1259, n1261, n1262, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1279, n1280, n1281, n1282, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1316, n1317, n1318, n1319, n1320, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1331, n1333, n1334, n1335, n1336, n1337, n1339, n1342, n1343, n1344, n1345, n1346, n1350, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1364, n1365, n1366, n1367, n1368, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1382, n1384, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1394, n1395, n1396, n1397, n1398, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1423, n1424, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1436, n1437, n1438, n1439, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1454, n1455, n1456, n1458, n1459, n1462, n1464, n1465, n1466, n1467, n1468, n1469, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1496, n1497, n1499, n1500, n1503, n1504, n1505, n1506, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1526, n1528, n1529, n1531, n1532, n1533, n1534, n1536, n1538, n1539, n1540, n1541, n1542, n1543, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1596, n1598, n1599, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1623, n1624, n1625, n1626, n1627, n1628, n1630, n1631, n1632, n1634, n1636, n1637, n1638, n1639, n1640, n1641, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1655, n1656, n1658, n1659, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1676, n1679, n1680, n1681, n1682, n1684, n1685, n1687, n1689, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1722, n1723, n1724, n1725, n1726, n1728, n1730, n1732, n1733, n1734, n1735, n1736, n1738, n1739, n1740, n1741, n1742, n1744, n1745, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1758, n1759, n1760, n1761, n1762, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773;
assign n1251 = n235 | n1266;
assign n1565 = ~n527;
assign n1312 = ~n1653;
assign n1414 = n1090 | n673;
assign n1352 = ~(n298 ^ n1568);
assign n599 = ~(n416 ^ n1403);
assign n1037 = n188 | n554;
assign n540 = ~(n654 | n986);
assign n1181 = n1582 | n72;
assign n473 = n562 | n1653;
assign n1146 = ~n911;
assign n1432 = ~(n265 ^ n953);
assign n188 = n952 & n329;
assign n229 = ~(n283 ^ n557);
assign n13 = n1085 & n1290;
assign n1272 = n1312 & n214;
assign n1716 = ~n390;
assign n361 = n1429 & n1126;
assign n1523 = ~(n1390 ^ n1645);
assign n702 = n1750 & n582;
assign n1368 = ~(n1343 | n816);
assign n662 = ~(n1371 | n1169);
assign n1015 = ~(n960 ^ n458);
assign n1156 = n874 | n193;
assign n696 = n1263 | n1444;
assign n1596 = n1316 | n316;
assign n827 = n1255 & n1155;
assign n1079 = n441 | n264;
assign n1502 = ~(n255 ^ n727);
assign n1725 = n898 & n1171;
assign n1318 = n1692 & n589;
assign n1384 = ~(n1174 | n48);
assign n744 = ~(n257 | n552);
assign n1697 = n101 & n283;
assign n308 = n1170 | n392;
assign n78 = n326 | n1680;
assign n1634 = ~n1282;
assign n1391 = ~(n128 ^ n92);
assign n1003 = ~(n1607 ^ n1764);
assign n20 = ~(n1671 ^ n305);
assign n1664 = n473 & n1404;
assign n1410 = ~n722;
assign n1155 = ~(n962 ^ n259);
assign n88 = n1527 | n46;
assign n228 = n1409 & n1099;
assign n458 = n96 | n698;
assign n1499 = n1642 | n1232;
assign n1234 = ~(n1458 ^ n569);
assign n35 = n543 | n706;
assign n726 = ~(n816 ^ n1579);
assign n819 = n1622 & n1346;
assign n12 = n922 & n1508;
assign n485 = n1057 | n463;
assign n704 = ~n1037;
assign n1770 = ~n1104;
assign n434 = n202 & n1276;
assign n63 = n503 & n1547;
assign n846 = ~(n604 ^ n286);
assign n1602 = n227 & n367;
assign n580 = n1727 & n1663;
assign n1046 = ~(n1643 ^ n1707);
assign n1773 = ~n1007;
assign n1722 = ~(n164 | n347);
assign n1702 = n1461 & n1381;
assign n665 = ~(n831 ^ n1698);
assign n1756 = n1734 | n1639;
assign n1174 = ~n123;
assign n843 = ~n133;
assign n529 = ~n119;
assign n398 = ~n936;
assign n902 = ~(n1099 ^ n1359);
assign n925 = ~(n1768 | n1167);
assign n1005 = ~(n125 ^ n103);
assign n1647 = ~n331;
assign n146 = n1381 | n1116;
assign n1715 = ~(n555 | n1014);
assign n125 = ~n550;
assign n1609 = ~(n1254 ^ n243);
assign n192 = n1329 | n266;
assign n1398 = ~(n5 ^ n260);
assign n428 = ~(n16 ^ n254);
assign n1730 = ~(n815 ^ n1357);
assign n1284 = ~(n1204 ^ n112);
assign n1322 = ~n203;
assign n584 = ~n362;
assign n1614 = n1337 & n131;
assign n1739 = n1658 & n179;
assign n371 = ~n682;
assign n42 = ~(n1442 | n994);
assign n1366 = ~n1363;
assign n947 = ~(n195 | n565);
assign n367 = n1381 | n601;
assign n73 = ~n1578;
assign n1243 = n1511 & n1767;
assign n1173 = n1473 & n1769;
assign n387 = ~(n1271 ^ n1425);
assign n834 = n789 | n249;
assign n474 = ~n954;
assign n1018 = ~n111;
assign n1456 = n382 & n474;
assign n443 = ~(n46 | n805);
assign n1327 = n1381 | n309;
assign n1762 = ~(n1146 ^ n497);
assign n639 = n1566 & n1771;
assign n1090 = ~(n1442 | n1335);
assign n590 = ~(n1643 | n1709);
assign n157 = ~n953;
assign n1106 = ~(n268 ^ n486);
assign n901 = n1626 | n1164;
assign n1688 = ~(n1168 ^ n898);
assign n470 = n605 | n548;
assign n1147 = n568 & n1076;
assign n177 = ~n379;
assign n535 = n472 & n99;
assign n921 = n332 & n1055;
assign n258 = n1543 | n233;
assign n77 = ~(n1469 | n558);
assign n338 = n1100 & n826;
assign n1317 = n1219 | n312;
assign n312 = ~n1280;
assign n767 = n820 | n1167;
assign n924 = n895 | n596;
assign n911 = n1323 | n640;
assign n158 = n1532 | n1472;
assign n857 = ~(n99 ^ n1743);
assign n108 = n1684 & n39;
assign n539 = n1112 & n1048;
assign n715 = ~n1408;
assign n368 = ~(n1443 ^ n213);
assign n55 = ~(n626 ^ n898);
assign n408 = ~n275;
assign n1211 = n40 | n75;
assign n1388 = ~(n1259 | n593);
assign n1486 = n1678 & n1381;
assign n971 = ~(n1065 | n1598);
assign n1268 = ~n1420;
assign n536 = ~n810;
assign n1606 = n57 | n1685;
assign n708 = ~n449;
assign n582 = ~(n1709 ^ n1474);
assign n1259 = n1310 | n1590;
assign n1517 = n102 | n191;
assign n129 = n562 | n73;
assign n370 = n1121 & n1367;
assign n160 = ~(n952 | n197);
assign n1353 = ~(n275 ^ n600);
assign n1210 = n1261 & n611;
assign n212 = n175 | n1374;
assign n278 = n947 | n1567;
assign n1719 = n827 & n1244;
assign n1621 = ~(n876 | n570);
assign n676 = ~n495;
assign n1242 = n1497 | n1061;
assign n749 = n391 & n536;
assign n1245 = ~(n1642 | n1617);
assign n1367 = n10 | n12;
assign n1407 = ~(n673 ^ n1733);
assign n1302 = ~(n1057 ^ n1169);
assign n1320 = ~n753;
assign n90 = n295 & n1215;
assign n1700 = ~n1592;
assign n809 = ~n839;
assign n669 = ~n70;
assign n1586 = n226 & n386;
assign n946 = n1532 | n296;
assign n1082 = ~n1115;
assign n849 = ~(n633 ^ n303);
assign n1119 = ~n471;
assign n1449 = n1435 & n1532;
assign n735 = ~n1448;
assign n820 = ~n247;
assign n1316 = ~n1381;
assign n570 = n667 | n166;
assign n938 = n1435 & n1167;
assign n1641 = n1274 ^ n247;
assign n376 = ~(n1512 ^ n1581);
assign n863 = n164 | n1381;
assign n710 = ~n1571;
assign n1550 = n657 & n308;
assign n807 = n94 | n1405;
assign n1324 = n926 & n211;
assign n1749 = ~n288;
assign n170 = ~(n1606 ^ n1222);
assign n1323 = n1381 & n1101;
assign n1054 = n1063 & n1414;
assign n374 = n1084 & n244;
assign n70 = n301 | n1506;
assign n45 = n978 & n924;
assign n237 = ~(n353 | n655);
assign n534 = ~(n923 | n660);
assign n68 = ~(n397 | n769);
assign n714 = n1044 & n995;
assign n1563 = n166 | n1353;
assign n1639 = ~(n1120 ^ n437);
assign n169 = n360 & n998;
assign n124 = n262 | n361;
assign n1365 = n23 | n996;
assign n654 = ~n737;
assign n915 = ~n1456;
assign n648 = ~(n511 ^ n1352);
assign n53 = n869 & n350;
assign n1637 = ~n1062;
assign n366 = ~n16;
assign n687 = ~(n1607 ^ n1062);
assign n1463 = ~(n28 ^ n139);
assign n1455 = n738 & n1485;
assign n246 = n366 | n137;
assign n932 = n579 | n354;
assign n76 = ~(n1673 ^ n133);
assign n148 = ~(n863 | n1611);
assign n235 = ~n1527;
assign n1292 = ~(n1469 | n1111);
assign n541 = n829 | n527;
assign n22 = n413 & n764;
assign n122 = n1416 & n701;
assign n1539 = n720 & n185;
assign n873 = n711 | n908;
assign n487 = n343 | n1606;
assign n121 = ~(n223 | n1584);
assign n71 = ~n1224;
assign n1084 = n1287 | n1528;
assign n826 = n110 | n1594;
assign n442 = ~(n1217 | n679);
assign n325 = n1082 | n1639;
assign n1349 = ~(n1239 ^ n1373);
assign n1385 = ~n614;
assign n659 = ~n787;
assign n1053 = ~(n253 | n1042);
assign n1280 = ~(n326 ^ n93);
assign n522 = ~(n323 ^ n352);
assign n1149 = ~(n652 ^ n851);
assign n322 = ~n1480;
assign n561 = ~n112;
assign n1112 = n1568 | n298;
assign n1065 = ~(n780 ^ n277);
assign n422 = n79 | n1627;
assign n96 = ~n1601;
assign n1182 = n1544 & n749;
assign n1477 = n806 & n1117;
assign n903 = ~(n952 | n265);
assign n477 = ~(n1597 | n266);
assign n1304 = ~(n1300 ^ n271);
assign n742 = ~n1636;
assign n996 = n219 & n395;
assign n642 = n825 | n832;
assign n586 = n1316 | n269;
assign n1121 = n291 | n1089;
assign n382 = ~n1185;
assign n754 = n1604 | n234;
assign n1040 = n1422 | n696;
assign n764 = ~n1762;
assign n462 = ~(n952 ^ n653);
assign n234 = ~(n507 ^ n796);
assign n777 = ~n763;
assign n1676 = ~(n1266 ^ n4);
assign n525 = n1386 & n631;
assign n825 = ~n1115;
assign n840 = n533 | n1662;
assign n1213 = ~(n1154 ^ n862);
assign n1286 = n1344 | n704;
assign n810 = n1328 | n453;
assign n1685 = ~n1154;
assign n271 = ~n75;
assign n1279 = n1585 | n279;
assign n948 = ~(n1604 ^ n1169);
assign n943 = n1694 & n1638;
assign n1342 = ~n797;
assign n748 = ~(n1203 ^ n242);
assign n1503 = ~n246;
assign n1769 = ~n1519;
assign n890 = ~(n1576 ^ n46);
assign n1511 = n490 | n281;
assign n1068 = ~(n1391 ^ n1755);
assign n664 = n322 | n407;
assign n306 = ~(n1575 ^ n736);
assign n1165 = ~(n1602 ^ n390);
assign n759 = ~(n30 ^ n1766);
assign n1475 = ~(n73 ^ n200);
assign n1138 = ~n284;
assign n851 = ~n78;
assign n1201 = ~(n1331 ^ n1714);
assign n951 = ~(n1365 ^ n693);
assign n190 = n141 & n1038;
assign n869 = ~n721;
assign n47 = ~(n1643 | n36);
assign n1199 = ~(n644 ^ n215);
assign n51 = ~(n1190 ^ n1708);
assign n611 = n853 | n1054;
assign n260 = ~(n1618 ^ n1763);
assign n448 = ~n411;
assign n595 = n1652 & n60;
assign n889 = ~n856;
assign n1126 = n1510 | n415;
assign n200 = ~n1225;
assign n84 = n1316 | n618;
assign n481 = n272 | n1102;
assign n321 = ~(n447 | n516);
assign n305 = ~(n1034 ^ n1643);
assign n1023 = ~(n555 ^ n1172);
assign n597 = n164 | n574;
assign n514 = ~(n654 | n692);
assign n98 = n80 | n551;
assign n551 = ~(n563 | n1306);
assign n454 = n1479 | n576;
assign n208 = ~(n994 ^ n117);
assign n1081 = ~(n39 ^ n1684);
assign n1684 = ~(n27 ^ n738);
assign n888 = ~(n1567 ^ n1552);
assign n144 = n1073 & n934;
assign n44 = ~(n1731 ^ n87);
assign n484 = ~(n1371 | n1555);
assign n1333 = n1259 & n436;
assign n173 = n1666 | n1710;
assign n916 = ~n819;
assign n65 = ~(n1014 ^ n555);
assign n113 = n1532 | n1593;
assign n1184 = ~n1483;
assign n1558 = ~n1501;
assign n1665 = ~n718;
assign n0 = ~n1763;
assign n1588 = ~(n722 | n1717);
assign n1001 = n1394 & n1141;
assign n41 = n1195 | n75;
assign n1047 = ~(n1473 | n1769);
assign n1509 = ~(n1275 | n1751);
assign n976 = ~(n199 | n1531);
assign n546 = n1588 | n190;
assign n345 = n794 | n758;
assign n1030 = ~(n1180 ^ n1326);
assign n900 = ~(n1207 ^ n31);
assign n1216 = n578 & n1156;
assign n1560 = ~(n720 ^ n1370);
assign n1459 = n1146 | n1004;
assign n1418 = n535 | n68;
assign n1070 = ~n489;
assign n523 = ~n1014;
assign n1694 = n509 | n1505;
assign n1582 = ~(n1240 ^ n1332);
assign n50 = n969 & n1184;
assign n1289 = n222 & n1008;
assign n572 = ~(n203 ^ n1579);
assign n731 = ~(n63 ^ n1676);
assign n400 = ~(n969 ^ n1483);
assign n1295 = ~(n584 | n1354);
assign n617 = ~(n620 ^ n803);
assign n1116 = n206 & n597;
assign n456 = n1139 | n832;
assign n1029 = ~n1748;
assign n482 = ~(n13 ^ n194);
assign n352 = ~(n879 ^ n268);
assign n1620 = n171 & n1499;
assign n39 = ~n861;
assign n393 = n1000 | n1040;
assign n1729 = ~(n998 ^ n1049);
assign n1230 = ~(n1564 ^ n1544);
assign n497 = n1250 & n1534;
assign n395 = ~n1618;
assign n604 = n1400 & n267;
assign n1592 = n1034 & n1129;
assign n1064 = ~(n24 ^ n781);
assign n449 = ~(n412 ^ n1661);
assign n409 = ~(n555 ^ n1140);
assign n1425 = ~(n1673 ^ n1108);
assign n254 = n528 & n1433;
assign n1050 = n232 | n894;
assign n268 = ~n1284;
assign n980 = ~(n1084 | n1272);
assign n1690 = ~(n118 ^ n610);
assign n1133 = n886 | n1137;
assign n1546 = n1317 & n431;
assign n9 = ~n832;
assign n1220 = ~(n741 | n1158);
assign n627 = n824 & n1271;
assign n349 = ~(n1208 | n104);
assign n1129 = ~n637;
assign n351 = ~n658;
assign n496 = ~(n121 | n1216);
assign n32 = ~n501;
assign n493 = ~n1078;
assign n241 = ~n393;
assign n1319 = n1124 & n1650;
assign n1013 = ~n994;
assign n1031 = ~(n454 ^ n1432);
assign n1457 = ~n1609;
assign n1595 = ~(n990 ^ n1348);
assign n524 = ~(n1513 | n402);
assign n1467 = ~(n478 | n475);
assign n973 = n1533 & n412;
assign n1346 = ~n987;
assign n1135 = ~(n35 ^ n1333);
assign n33 = ~(n639 ^ n273);
assign n1451 = ~(n1082 ^ n351);
assign n1667 = ~n698;
assign n1576 = ~n163;
assign n802 = ~n695;
assign n153 = n34 & n1728;
assign n287 = ~(n855 | n1671);
assign n883 = ~(n1165 ^ n1074);
assign n1099 = ~n1353;
assign n1334 = n1741 & n774;
assign n814 = n682 & n1371;
assign n618 = ~(n1620 | n283);
assign n1239 = n456 & n808;
assign n1115 = ~n123;
assign n830 = n1381 | n615;
assign n339 = ~n838;
assign n928 = n1568 & n298;
assign n1657 = ~(n2 ^ n1138);
assign n530 = ~n607;
assign n452 = ~(n1273 ^ n1523);
assign n479 = ~(n555 | n1172);
assign n717 = ~(n852 | n1052);
assign n249 = n957 & n1679;
assign n222 = n1723 | n1505;
assign n112 = n972 | n1018;
assign n641 = ~n54;
assign n786 = ~(n353 ^ n655);
assign n1376 = n906 & n819;
assign n858 = ~(n1491 ^ n500);
assign n1492 = ~n1444;
assign n1430 = ~(n98 ^ n353);
assign n750 = ~(n1324 | n616);
assign n1130 = ~(n101 | n402);
assign n1100 = n359 | n1374;
assign n1669 = ~(n1322 | n228);
assign n189 = n101 | n335;
assign n1476 = ~(n1265 | n795);
assign n307 = ~(n797 ^ n433);
assign n1720 = n1300 & n1581;
assign n1369 = n864 | n1333;
assign n1594 = n955 & n1454;
assign n1087 = n737 | n302;
assign n1552 = ~(n435 ^ n195);
assign n1372 = ~(n1217 ^ n379);
assign n316 = n723 & n1232;
assign n811 = ~(n585 | n402);
assign n1161 = ~(n1141 ^ n828);
assign n451 = n505 & n933;
assign n528 = n1691 | n477;
assign n727 = ~(n104 ^ n1480);
assign n1711 = n543 & n1224;
assign n1542 = ~n464;
assign n1077 = ~(n197 ^ n472);
assign n204 = n1152 | n1327;
assign n293 = ~n696;
assign n1420 = n1051 | n775;
assign n1699 = ~(n66 | n1442);
assign n1528 = n91 & n144;
assign n1257 = ~n1190;
assign n871 = ~n1617;
assign n1378 = n240 | n620;
assign n824 = n1093 & n1724;
assign n511 = ~n122;
assign n194 = ~(n825 ^ n48);
assign n1659 = n177 & n88;
assign n917 = ~n396;
assign n1445 = ~n1105;
assign n1091 = ~(n667 | n266);
assign n1608 = n223 & n1584;
assign n217 = ~n1474;
assign n1249 = ~n711;
assign n1011 = n1177 & n1110;
assign n673 = n833 & n1096;
assign n1709 = n1486 | n384;
assign n1580 = n177 | n879;
assign n818 = ~(n1450 ^ n587);
assign n762 = n659 | n312;
assign n1331 = n1231 & n251;
assign n56 = ~(n1143 ^ n172);
assign n1437 = n1607 | n440;
assign n1488 = ~(n1217 | n1280);
assign n757 = n1375 & n331;
assign n680 = ~(n338 ^ n65);
assign n1589 = ~(n257 | n1725);
assign n743 = ~(n1461 | n402);
assign n1512 = ~n489;
assign n1765 = n486 | n268;
assign n1753 = n1695 | n209;
assign n100 = n1708 & n1257;
assign n678 = n1580 & n1738;
assign n83 = ~n849;
assign n1741 = n1415 | n658;
assign n1308 = ~(n624 | n1147);
assign n202 = n1300 | n72;
assign n1401 = n675 & n1214;
assign n432 = ~(n233 ^ n773);
assign n711 = ~(n1307 ^ n1397);
assign n336 = n413 | n764;
assign n131 = n1699 | n21;
assign n1471 = ~(n543 | n1224);
assign n209 = n1269 & n118;
assign n1673 = ~n1093;
assign n815 = ~(n361 ^ n1021);
assign n460 = ~(n1605 ^ n728);
assign n573 = ~(n1625 ^ n948);
assign n1613 = n591 | n1658;
assign n274 = ~(n447 ^ n1084);
assign n30 = n336 & n765;
assign n583 = ~(n1768 | n402);
assign n500 = ~(n1581 ^ n1265);
assign n829 = n1721 & n406;
assign n300 = ~(n447 | n1312);
assign n548 = n860 & n1605;
assign n1473 = ~(n1437 ^ n462);
assign n1496 = n504 | n676;
assign n1759 = ~(n953 | n265);
assign n227 = n1316 | n229;
assign n1223 = ~n960;
assign n1392 = ~(n1371 | n1645);
assign n291 = ~n555;
assign n935 = ~(n1149 ^ n162);
assign n165 = ~n252;
assign n995 = n1043 | n1075;
assign n733 = ~n1499;
assign n616 = n164 | n355;
assign n1556 = ~(n1426 ^ n96);
assign n800 = ~(n1217 | n268);
assign n1364 = ~(n678 ^ n1166);
assign n273 = ~(n509 ^ n1357);
assign n346 = n326 | n64;
assign n118 = n1148 | n1293;
assign n1058 = n1060 ^ n171;
assign n1026 = n1213 | n1581;
assign n1055 = n1000 | n619;
assign n907 = n1259 & n593;
assign n886 = ~(n805 | n1320);
assign n1491 = n1644 & n752;
assign n518 = ~n480;
assign n993 = ~(n50 ^ n1192);
assign n1150 = n149 | n1053;
assign n10 = ~(n555 | n927);
assign n756 = n155 & n1000;
assign n1300 = ~n1070;
assign n304 = ~n896;
assign n861 = ~(n1636 ^ n1039);
assign n558 = n581 & n529;
assign n48 = ~n1639;
assign n808 = n920 | n1319;
assign n436 = n845 & n545;
assign n1137 = n41 & n844;
assign n619 = ~(n508 ^ n379);
assign n1632 = n1643 & n761;
assign n1073 = ~(n1307 ^ n480);
assign n1469 = ~n730;
assign n1615 = ~n162;
assign n720 = ~n1307;
assign n499 = ~n1187;
assign n21 = ~n691;
assign n461 = ~(n266 | n184);
assign n1340 = ~(n745 ^ n1752);
assign n1696 = ~n1539;
assign n876 = ~n968;
assign n1148 = n1065 & n1598;
assign n578 = n1713 | n1443;
assign n1760 = ~(n952 ^ n329);
assign n43 = n143 | n413;
assign n1056 = ~(n634 | n1357);
assign n111 = n1029 & n868;
assign n1404 = n300 | n28;
assign n1360 = ~n977;
assign n15 = ~(n1763 | n395);
assign n219 = ~n422;
assign n835 = ~(n410 | n1578);
assign n95 = n1149 & n1615;
assign n28 = n129 & n11;
assign n1736 = ~(n1139 ^ n9);
assign n734 = n455 & n467;
assign n1124 = n815 | n281;
assign n1383 = n1388 | n907;
assign n1555 = ~n234;
assign n1014 = n1041 | n661;
assign n1110 = n337 | n30;
assign n564 = ~n542;
assign n383 = n687 & n83;
assign n404 = n926 | n1492;
assign n1744 = ~n1159;
assign n1297 = n652 | n78;
assign n792 = ~(n153 ^ n1032);
assign n929 = n417 & n1019;
assign n1127 = n682 | n1371;
assign n406 = ~n1739;
assign n1113 = ~(n849 ^ n898);
assign n899 = ~(n787 | n1280);
assign n465 = ~(n921 | n1549);
assign n1644 = n1750 | n582;
assign n1247 = ~n788;
assign n193 = ~n1418;
assign n1640 = ~(n562 | n993);
assign n770 = n35 & n1333;
assign n594 = ~n1003;
assign n1326 = ~(n386 ^ n226);
assign n568 = n291 | n939;
assign n236 = ~n498;
assign n638 = ~(n470 ^ n721);
assign n1180 = ~n1356;
assign n1122 = ~(n410 | n1560);
assign n806 = n1195 | n1581;
assign n437 = ~n1559;
assign n643 = n128 & n538;
assign n1177 = n1266 | n1612;
assign n985 = n926 | n562;
assign n1403 = ~n1658;
assign n1144 = ~(n562 ^ n923);
assign n668 = n682 | n1000;
assign n1604 = ~n1045;
assign n965 = ~(n607 | n1678);
assign n358 = ~n801;
assign n1169 = ~(n1034 ^ n637);
assign n966 = ~(n353 ^ n498);
assign n369 = ~n171;
assign n1212 = ~n173;
assign n136 = n1381 | n89;
assign n716 = ~n818;
assign n964 = ~n1505;
assign n1431 = n1532 | n1163;
assign n1572 = ~n1610;
assign n1359 = ~n1409;
assign n571 = n1527 | n61;
assign n257 = ~n1033;
assign n732 = ~n1073;
assign n186 = ~n841;
assign n1021 = ~(n353 ^ n695);
assign n301 = n1157 & n1190;
assign n1141 = n1640 | n451;
assign n1004 = ~n497;
assign n334 = ~(n1082 ^ n37);
assign n29 = n1410 | n1612;
assign n1754 = n1123 | n249;
assign n290 = ~(n1171 ^ n594);
assign n1290 = n1585 | n42;
assign n1444 = n379 | n709;
assign n216 = ~(n894 ^ n1128);
assign n1132 = n556 | n1745;
assign n856 = ~n1655;
assign n954 = n757 | n348;
assign n1771 = n744 | n1031;
assign n1311 = n369 | n1167;
assign n1400 = n1266 | n407;
assign n844 = n1294 | n525;
assign n1107 = n1607 | n1536;
assign n565 = ~n435;
assign n979 = ~(n1646 ^ n755);
assign n57 = ~n862;
assign n1203 = ~n714;
assign n1723 = ~(n191 ^ n966);
assign n552 = ~n1591;
assign n75 = ~(n528 ^ n1592);
assign n531 = n1674 & n420;
assign n988 = n1476 | n1491;
assign n1224 = n1263 | n1548;
assign n180 = n115 & n356;
assign n318 = n1146 | n1496;
assign n1409 = ~(n1607 ^ n183);
assign n1629 = ~(n383 ^ n1325);
assign n99 = ~n249;
assign n1266 = ~n1740;
assign n5 = n220 | n398;
assign n838 = n158 & n1406;
assign n1660 = ~(n1391 ^ n793);
assign n1628 = ~n684;
assign n897 = n1758 | n1243;
assign n1693 = n166 | n1168;
assign n501 = n973 | n915;
assign n884 = n1597 & n1512;
assign n201 = ~n1274;
assign n874 = ~(n444 | n977);
assign n1638 = n697 | n1331;
assign n1088 = n1532 | n189;
assign n357 = ~(n1678 | n402);
assign n513 = ~(n693 | n1365);
assign n354 = n754 & n1557;
assign n1208 = ~n1104;
assign n1085 = n509 | n1013;
assign n127 = ~n17;
assign n1645 = ~n582;
assign n93 = n1744 & n1361;
assign n556 = ~(n555 | n788);
assign n605 = ~(n629 | n713);
assign n1513 = ~n26;
assign n958 = n310 | n1551;
assign n1233 = n1246 | n678;
assign n1406 = n1000 | n1131;
assign n280 = n1626 & n1164;
assign n603 = n257 & n1725;
assign n1571 = n105 | n881;
assign n1607 = ~n1145;
assign n1195 = ~n1070;
assign n576 = ~n633;
assign n384 = ~(n1196 | n1236);
assign n480 = n666 & n1749;
assign n1658 = n1237 & n1609;
assign n143 = ~n46;
assign n1545 = n650 | n134;
assign n242 = ~(n104 ^ n1770);
assign n1745 = n1080 & n1286;
assign n238 = ~(n1019 ^ n645);
assign n864 = ~(n1259 | n436);
assign n1450 = n956 & n1445;
assign n1521 = ~(n879 ^ n679);
assign n314 = ~(n1341 | n1014);
assign n1691 = n607 & n266;
assign n1191 = ~(n1664 ^ n58);
assign n1748 = ~(n16 ^ n324);
assign n1439 = n885 | n539;
assign n288 = n742 | n1002;
assign n142 = ~n1221;
assign n79 = n870 & n1000;
assign n1692 = n359 | n636;
assign n1265 = ~n1213;
assign n1315 = ~(n1727 ^ n1619);
assign n495 = n399 | n1205;
assign n2 = n614 | n364;
assign n1299 = ~(n413 ^ n1320);
assign n677 = ~(n1584 ^ n223);
assign n1283 = ~(n1725 ^ n1494);
assign n549 = ~(n821 | n53);
assign n505 = n362 | n663;
assign n918 = ~(n1160 | n1532);
assign n543 = ~n1422;
assign n1167 = ~n266;
assign n162 = n1083 | n87;
assign n455 = n1225 | n1578;
assign n1742 = ~n692;
assign n905 = ~(n1054 ^ n334);
assign n1387 = ~n628;
assign n405 = ~(n1576 ^ n435);
assign n850 = ~(n1173 | n791);
assign n3 = n1597 | n1512;
assign n983 = ~n1288;
assign n364 = ~n580;
assign n488 = ~(n166 ^ n347);
assign n184 = n1583 & n61;
assign n593 = n845 & n1421;
assign n647 = n962 & n1703;
assign n1231 = n1229 | n1563;
assign n289 = ~n414;
assign n1508 = n237 | n710;
assign n1206 = n562 | n713;
assign n385 = n1122 | n625;
assign n244 = n1670 | n1336;
assign n787 = ~(n1732 ^ n839);
assign n1274 = n1513 | n1313;
assign n37 = ~n1164;
assign n1727 = ~(n504 ^ n495);
assign n389 = ~n144;
assign n671 = ~n1022;
assign n1458 = n617 | n1719;
assign n658 = ~(n1448 ^ n411);
assign n637 = n735 | n448;
assign n596 = n999 & n1517;
assign n1309 = ~(n703 | n604);
assign n1083 = ~n1731;
assign n1186 = ~n1111;
assign n1581 = ~(n504 ^ n1228);
assign n763 = n1431 & n176;
assign n836 = ~(n552 ^ n694);
assign n1250 = ~n504;
assign n423 = ~(n1007 ^ n751);
assign n1142 = ~(n1221 ^ n660);
assign n1017 = ~n1496;
assign n506 = n1123 | n1134;
assign n728 = ~(n713 ^ n629);
assign n168 = n486 & n268;
assign n1443 = ~n977;
assign n712 = ~(n1519 ^ n919);
assign n624 = ~(n1643 | n1707);
assign n81 = ~(n952 | n653);
assign n1278 = n1413 & n793;
assign n634 = ~n1109;
assign n774 = n577 | n1289;
assign n609 = n43 & n1772;
assign n1577 = ~n1172;
assign n25 = n962 | n160;
assign n1766 = ~(n1208 ^ n1612);
assign n123 = ~(n1745 ^ n785);
assign n419 = ~(n816 ^ n968);
assign n206 = n820 | n402;
assign n187 = n205 & n225;
assign n1269 = n252 | n400;
assign n417 = n613 | n679;
assign n719 = n730 | n1186;
assign n85 = n1711 | n566;
assign n765 = n22 | n1477;
assign n520 = ~(n1371 | n716);
assign n698 = ~(n1545 ^ n779);
assign n1232 = ~n544;
assign n491 = ~(n1709 ^ n1643);
assign n1686 = ~(n869 ^ n1681);
assign n1028 = n1636 | n1209;
assign n1134 = ~n729;
assign n8 = n1542 | n1773;
assign n1683 = ~n617;
assign n224 = ~n1623;
assign n1294 = ~(n1512 | n271);
assign n411 = n1603 | n1291;
assign n821 = n1673 | n843;
assign n1498 = ~(n1289 ^ n1395);
assign n1006 = ~(n1264 | n524);
assign n537 = ~n1433;
assign n134 = ~(n1066 | n1614);
assign n978 = n291 | n1366;
assign n1045 = ~n900;
assign n467 = n168 | n311;
assign n1330 = ~(n1396 ^ n686);
assign n956 = n1751 | n1226;
assign n666 = ~n1575;
assign n310 = ~(n1263 | n483);
assign n489 = ~(n173 ^ n1501);
assign n58 = ~(n362 ^ n374);
assign n919 = ~(n1473 ^ n791);
assign n1514 = ~(n257 | n261);
assign n355 = ~(n926 | n211);
assign n569 = ~n20;
assign n1506 = ~n50;
assign n340 = n1151 | n671;
assign n67 = ~(n1653 ^ n214);
assign n1549 = n531 & n1446;
assign n365 = ~n1490;
assign n877 = n730 | n373;
assign n333 = n212 & n1587;
assign n633 = n1702 | n445;
assign n755 = ~(n1300 ^ n298);
assign n243 = ~(n265 ^ n952);
assign n937 = ~n1434;
assign n997 = n1520 & n1016;
assign n1202 = ~(n647 ^ n646);
assign n476 = ~(n1071 ^ n1069);
assign n674 = ~n265;
assign n1235 = ~(n1364 ^ n719);
assign n779 = ~(n1371 ^ n682);
assign n297 = ~n600;
assign n172 = ~(n1230 ^ n602);
assign n1625 = n1464 & n1200;
assign n793 = n567 | n1074;
assign n1178 = ~(n353 | n1351);
assign n950 = ~(n1612 ^ n722);
assign n1252 = n1607 | n893;
assign n1196 = ~(n164 | n682);
assign n547 = ~(n691 ^ n1718);
assign n372 = ~(n83 ^ n1189);
assign n1687 = ~n1450;
assign n1569 = n740 | n1389;
assign n799 = ~n656;
assign n1470 = n77 | n1421;
assign n156 = ~(n1602 ^ n342);
assign n279 = ~(n464 | n1007);
assign n137 = ~n254;
assign n776 = n899 | n550;
assign n1656 = ~n539;
assign n430 = n869 & n470;
assign n566 = n266 | n1471;
assign n606 = n86 & n592;
assign n341 = n226 | n386;
assign n1248 = ~n346;
assign n986 = n1223 & n553;
assign n270 = ~(n1364 ^ n877);
assign n502 = n1114 | n705;
assign n1325 = ~(n1253 ^ n1031);
assign n483 = ~n1548;
assign n1022 = n1687 & n1424;
assign n893 = ~n931;
assign n1405 = ~(n1456 ^ n783);
assign n775 = ~n996;
assign n805 = ~n163;
assign n1772 = n443 | n880;
assign n736 = n742 & n1503;
assign n399 = ~(n1275 | n18);
assign n1194 = ~(n1118 ^ n1087);
assign n24 = ~n1405;
assign n1386 = n1390 | n463;
assign n1357 = ~n281;
assign n74 = ~(n983 ^ n1630);
assign n631 = n662 | n1625;
assign n1636 = n767 & n345;
assign n377 = ~n1678;
assign n120 = ~(n241 | n100);
assign n1276 = n1350 | n1303;
assign n1185 = ~(n331 ^ n606);
assign n626 = ~(n936 ^ n1530);
assign n718 = n1426 | n96;
assign n853 = ~(n1174 | n37);
assign n429 = ~(n873 ^ n493);
assign n1733 = ~(n490 ^ n1335);
assign n746 = ~(n132 | n383);
assign n1553 = ~(n1575 ^ n1490);
assign n1677 = ~(n570 ^ n419);
assign n1214 = n1537 & n896;
assign n1601 = ~(n1614 ^ n521);
assign n721 = ~(n441 ^ n1539);
assign n1706 = ~n940;
assign n199 = ~(n164 | n968);
assign n164 = ~n402;
assign n550 = n29 & n546;
assign n969 = ~(n1623 ^ n799);
assign n267 = n349 | n714;
assign n396 = n449 & n32;
assign n1354 = ~n400;
assign n89 = ~(n583 | n1092);
assign n1731 = ~(n326 ^ n1227);
assign n1237 = ~(n633 ^ n1145);
assign n181 = ~(n960 ^ n1541);
assign n828 = ~(n562 ^ n1221);
assign n1111 = n581 & n804;
assign n507 = n766 & n1559;
assign n645 = ~(n679 ^ n613);
assign n790 = ~(n525 ^ n1304);
assign n1345 = n1301 | n609;
assign n441 = ~n1427;
assign n650 = n1435 & n1174;
assign n154 = ~(n213 | n1360);
assign n1570 = ~(n1626 ^ n37);
assign n1454 = n1254 | n903;
assign n1561 = n359 | n977;
assign n343 = ~n1222;
assign n486 = ~(n519 ^ n649);
assign n694 = ~(n1229 ^ n1031);
assign n1460 = ~(n261 ^ n670);
assign n1103 = n715 ^ n1565;
assign n933 = n1295 | n169;
assign n1270 = ~n228;
assign n1567 = n1181 & n1436;
assign n1012 = ~(n1599 ^ n575);
assign n1192 = ~n301;
assign n970 = n834 & n481;
assign n282 = n1489 & n167;
assign n313 = n1026 & n988;
assign n533 = n1734 & n1639;
assign n1310 = ~n35;
assign n1618 = n918 | n1241;
assign n1541 = n718 | n698;
assign n1060 = n1768 | n871;
assign n221 = n471 | n152;
assign n1735 = n101 | n1167;
assign n1209 = ~n1002;
assign n1162 = n540 | n804;
assign n581 = ~n1118;
assign n1429 = n1123 | n1153;
assign n207 = ~(n1480 | n104);
assign n1548 = n379 | n571;
assign n1044 = n413 | n1405;
assign n1655 = ~n1401;
assign n681 = n1747 & n1455;
assign n245 = n291 | n1247;
assign n1654 = ~(n1477 ^ n319);
assign n656 = n1238 & n872;
assign n1067 = ~(n502 ^ n1106);
assign n119 = n737 | n1742;
assign n521 = ~(n1174 ^ n1435);
assign n130 = ~n88;
assign n688 = n1253 | n1;
assign n1710 = ~(n47 | n1207);
assign n875 = ~(n1643 | n424);
assign n1288 = n1756 & n840;
assign n1016 = ~n1244;
assign n344 = ~(n1643 ^ n469);
assign n1154 = n1632 | n984;
assign n630 = ~(n1300 ^ n967);
assign n1380 = n1059 & n818;
assign n1500 = n1381 & n1697;
assign n225 = n1669 | n1579;
assign n478 = ~(n562 | n1664);
assign n16 = n913 | n461;
assign n117 = ~(n490 ^ n1585);
assign n1519 = n1003 & n1171;
assign n1651 = n1027 & n1482;
assign n1008 = n161 | n187;
assign n772 = n1381 | n743;
assign n1157 = n838 | n1187;
assign n589 = n1178 | n320;
assign n1066 = ~(n1435 | n1174);
assign n1703 = n1145 | n275;
assign n1102 = ~(n1743 | n197);
assign n1348 = ~(n128 ^ n538);
assign n1379 = n815 & n281;
assign n1761 = ~(n170 | n1762);
assign n1377 = ~(n69 | n98);
assign n356 = n479 | n375;
assign n1516 = ~(n555 ^ n1363);
assign n1484 = n1341 & n1014;
assign n1104 = ~n1740;
assign n1187 = n656 & n224;
assign n723 = n820 | n1402;
assign n620 = n1561 & n1569;
assign n1218 = n1684 | n39;
assign n957 = n1160 | n1167;
assign n450 = ~(n369 | n402);
assign n62 = n1390 | n582;
assign n182 = n1497 & n1061;
assign n107 = ~(n90 | n513);
assign n1048 = n928 | n122;
assign n1559 = n909 | n107;
assign n151 = n442 | n1550;
assign n1305 = ~(n35 ^ n907);
assign n796 = ~n757;
assign n601 = ~(n1130 | n1220);
assign n852 = n177 & n571;
assign n284 = ~(n318 ^ n1159);
assign n1438 = n1461 & n1000;
assign n1397 = n666 | n1193;
assign n741 = n543 & n159;
assign n1260 = ~(n76 ^ n430);
assign n152 = n428 | n258;
assign n967 = ~n72;
assign n1452 = n291 | n735;
assign n519 = ~n1182;
assign n504 = n1524 & n204;
assign n97 = ~n1151;
assign n6 = ~(n257 | n1382);
assign n1337 = n1329 | n490;
assign n833 = n1229 | n1693;
assign n1554 = n359 | n802;
assign n1433 = n1509 | n287;
assign n1143 = n285 & n278;
assign n1061 = ~(n1418 ^ n1010);
assign n360 = n410 | n400;
assign n211 = n379 | n88;
assign n1675 = ~(n228 ^ n572);
assign n753 = ~(n16 ^ n114);
assign n1415 = ~(n596 ^ n1516);
assign n447 = ~n889;
assign n1671 = n1452 & n1378;
assign n166 = ~n438;
assign n608 = ~n91;
assign n975 = n1266 | n602;
assign n54 = n1631 & n668;
assign n1002 = n16 | n1462;
assign n804 = ~n1087;
assign n23 = n422 & n1618;
assign n1507 = ~(n1319 ^ n1736);
assign n999 = n359 | n236;
assign n832 = ~(n333 ^ n1668);
assign n685 = n1380 | n425;
assign n991 = ~(n933 ^ n1098);
assign n1442 = ~n1109;
assign n1226 = n735 & n977;
assign n1650 = n1379 | n651;
assign n868 = ~n340;
assign n1681 = n1206 & n385;
assign n1109 = ~n612;
assign n86 = n965 | n946;
assign n962 = n1607 | n408;
assign n72 = ~(n1022 ^ n97);
assign n239 = ~(n952 ^ n729);
assign n803 = ~(n1448 ^ n555);
assign n215 = ~(n1371 ^ n1555);
assign n538 = n1602 | n1297;
assign n1382 = ~n1563;
assign n1168 = ~(n275 ^ n801);
assign n1585 = ~(n90 ^ n951);
assign n1489 = n157 | n674;
assign n1339 = ~n195;
assign n632 = n1123 | n289;
assign n1497 = ~(n320 ^ n248);
assign n185 = ~n1370;
assign n373 = ~n558;
assign n1139 = ~(n375 ^ n1023);
assign n1543 = ~(n1468 ^ n537);
assign n1591 = n166 | n849;
assign n1536 = ~n183;
assign n1534 = ~n1228;
assign n895 = ~(n555 | n1363);
assign n1728 = n800 | n323;
assign n859 = n1195 | n298;
assign n1052 = n266 | n784;
assign n1095 = n720 & n178;
assign n457 = n514 | n529;
assign n1515 = n562 | n386;
assign n1505 = ~(n970 ^ n368);
assign n984 = ~(n1682 | n180);
assign n679 = ~n1553;
assign n1605 = n854 | n929;
assign n1373 = ~(n1750 ^ n1645);
assign n255 = ~n847;
assign n1436 = n1362 | n831;
assign n1240 = n198 | n1308;
assign n1538 = ~(n1266 ^ n39);
assign n1575 = n925 | n717;
assign n1653 = ~(n389 ^ n608);
assign n1518 = n82 | n1334;
assign n912 = ~(n1118 ^ n119);
assign n657 = n1266 | n861;
assign n1680 = ~n1227;
assign n386 = ~(n652 ^ n346);
assign n294 = n814 | n1562;
assign n683 = ~(n1150 ^ n1081);
assign n1419 = n1218 & n1150;
assign n544 = n820 & n1402;
assign n1573 = ~(n1643 ^ n424);
assign n210 = n150 | n1441;
assign n1635 = n1649 | n250;
assign n265 = n492 | n976;
assign n1672 = ~(n396 ^ n1434);
assign n1007 = n1047 | n850;
assign n1256 = ~n156;
assign n706 = n985 & n1233;
assign n771 = ~(n764 ^ n170);
assign n990 = n1256 | n1487;
assign n1648 = ~(n926 | n1548);
assign n1423 = ~n870;
assign n1599 = ~n1011;
assign n163 = ~n307;
assign n1198 = n325 & n380;
assign n865 = ~n306;
assign n1416 = n1282 | n234;
assign n872 = n1000 | n388;
assign n1713 = ~n444;
assign n1176 = ~(n555 ^ n927);
assign n1131 = ~(n293 ^ n1422);
assign n816 = ~n515;
assign n615 = ~(n155 | n402);
assign n1344 = ~(n353 | n747);
assign n87 = n284 | n2;
assign n1689 = ~(n379 | n1217);
assign n977 = n109 & n192;
assign n410 = ~n889;
assign n1447 = n1285 | n371;
assign n940 = n1597 | n682;
assign n453 = ~n1240;
assign n1329 = ~n66;
assign n1170 = ~(n1208 | n39);
assign n335 = n369 | n1060;
assign n1408 = ~(n1651 ^ n491);
assign n690 = ~(n1706 ^ n46);
assign n1704 = ~(n1466 | n745);
assign n760 = ~n1549;
assign n1101 = ~(n26 ^ n607);
assign n139 = ~(n562 ^ n1312);
assign n1246 = ~(n1263 | n447);
assign n1287 = n1673 & n1079;
assign n1411 = ~n49;
assign n232 = n40 & n75;
assign n1171 = ~n626;
assign n660 = n663 & n1753;
assign n1468 = ~n528;
assign n955 = n1123 | n674;
assign n1424 = n1608 | n496;
assign n401 = ~(n190 ^ n950);
assign n992 = n280 | n817;
assign n560 = ~n747;
assign n691 = n1621 | n1368;
assign n378 = ~(n1662 ^ n328);
assign n38 = ~n1204;
assign n892 = n1413 & n1755;
assign n1009 = n143 & n1285;
assign n471 = ~(n1636 ^ n246);
assign n1587 = n1377 | n282;
assign n418 = ~(n952 | n329);
assign n286 = ~(n1672 ^ n1217);
assign n914 = ~(n1428 ^ n239);
assign n848 = ~(n353 ^ n747);
assign n1057 = ~(n45 ^ n1573);
assign n1767 = n1056 | n639;
assign n1529 = ~(n1643 | n469);
assign n831 = n1465 & n685;
assign n1020 = n207 | n847;
assign n784 = ~(n177 | n571);
assign n327 = ~n655;
assign n782 = ~n1616;
assign n426 = ~(n1243 ^ n1701);
assign n251 = n6 | n1579;
assign n930 = ~(n952 ^ n1296);
assign n114 = ~n466;
assign n446 = n1219 | n1553;
assign n559 = ~(n434 ^ n405);
assign n1480 = ~(n916 ^ n906);
assign n644 = ~n1198;
assign n1758 = ~(n1174 | n9);
assign n256 = n413 | n753;
assign n179 = ~(n1594 ^ n1430);
assign n459 = n884 | n421;
assign n1328 = ~n1332;
assign n115 = n291 | n1577;
assign n579 = n1195 & n298;
assign n1074 = n1515 & n1522;
assign n1395 = ~(n1415 ^ n351);
assign n942 = ~(n152 ^ n1119);
assign n1175 = ~(n221 ^ n865);
assign n296 = ~n1313;
assign n1531 = n1381 | n811;
assign n1 = ~n383;
assign n1394 = n362 | n142;
assign n1336 = ~n1528;
assign n1136 = ~n972;
assign n1205 = ~(n590 | n1651);
assign n1350 = ~(n1512 | n967);
assign n1532 = ~n1000;
assign n463 = ~n1169;
assign n1737 = ~(n76 ^ n53);
assign n320 = n506 & n1036;
assign n1590 = ~(n1422 | n230);
assign n1282 = ~(n370 ^ n344);
assign n262 = ~(n353 | n695);
assign n1027 = n291 | n523;
assign n1434 = n465 | n224;
assign n981 = ~(n1497 ^ n1335);
assign n567 = ~n1165;
assign n1163 = n866 | n201;
assign n598 = n1392 | n1273;
assign n468 = ~(n1059 ^ n716);
assign n910 = n235 | n143;
assign n699 = ~(n1188 ^ n1144);
assign n1117 = n1720 | n635;
assign n1600 = ~(n943 ^ n1451);
assign n92 = n1602 | n1716;
assign n1682 = ~(n1643 | n761);
assign n218 = ~(n187 ^ n381);
assign n350 = ~n1681;
assign n440 = ~n1764;
assign n1041 = n155 & n1381;
assign n1708 = n1088 & n393;
assign n1652 = n914 | n798;
assign n841 = n606 & n1647;
assign n1698 = ~(n1582 ^ n967);
assign n1630 = ~(n1555 ^ n1634);
assign n1128 = ~(n40 ^ n271);
assign n794 = ~(n1527 | n1009);
assign n309 = ~(n607 | n402);
assign n105 = n952 & n653;
assign n233 = n20 | n1458;
assign n403 = ~(n584 ^ n1560);
assign n1448 = n1540 | n938;
assign n972 = n1028 & n288;
assign n909 = n693 & n1365;
assign n1229 = ~n515;
assign n1623 = n778 | n760;
assign n526 = n1586 | n1356;
assign n879 = ~n1712;
assign n1189 = ~n687;
assign n517 = ~(n1550 ^ n1521);
assign n686 = ~(n1672 ^ n1065);
assign n1495 = ~(n595 ^ n981);
assign n381 = ~(n1723 ^ n964);
assign n1356 = n762 & n776;
assign n752 = n702 | n1239;
assign n1718 = ~(n490 ^ n66);
assign n1428 = n1607 | n1628;
assign n1105 = n1751 & n1226;
assign n317 = ~(n313 ^ n771);
assign n427 = ~(n1529 | n370);
assign n494 = ~n1095;
assign n503 = n413 | n435;
assign n281 = ~(n282 ^ n1267);
assign n778 = ~n921;
assign n397 = n358 | n408;
assign n272 = n297 | n408;
assign n1241 = ~(n876 | n1000);
assign n701 = n116 | n1288;
assign n191 = n632 & n945;
assign n109 = n1423 | n1167;
assign n636 = ~n1351;
assign n1485 = n961 & n1387;
assign n31 = ~(n1643 ^ n36);
assign n34 = n1219 | n1284;
assign n614 = ~(n911 ^ n1017);
assign n302 = ~n986;
assign n1487 = ~n95;
assign n591 = n1183 & n1457;
assign n661 = ~(n1417 | n830);
assign n766 = ~n1120;
assign n231 = ~(n467 ^ n1475);
assign n1093 = n1355 & n71;
assign n1051 = n756 | n1449;
assign n934 = n38 & n561;
assign n1275 = ~n1643;
assign n259 = ~(n99 ^ n952);
assign n150 = n1643 & n424;
assign n553 = ~n458;
assign n923 = n120 | n669;
assign n1510 = n1607 | n1637;
assign n908 = n306 | n221;
assign n1738 = n1689 | n542;
assign n1755 = n567 | n707;
assign n348 = ~n507;
assign n1562 = n1127 & n1545;
assign n421 = n3 & n294;
assign n1631 = n1532 | n1678;
assign n1303 = n512 & n1412;
assign n707 = n341 & n526;
assign n881 = ~(n1437 | n81);
assign n1402 = n1513 & n530;
assign n439 = ~(n628 ^ n961);
assign n1108 = ~n1724;
assign n1396 = n664 & n1020;
assign n789 = ~n1743;
assign n960 = ~(n294 ^ n941);
assign n904 = ~(n439 ^ n753);
assign n751 = ~(n1585 ^ n1542);
assign n175 = ~n69;
assign n621 = ~(n450 | n750);
assign n791 = ~n1398;
assign n1152 = ~(n164 | n1597);
assign n1307 = n1311 & n958;
assign n1158 = n164 | n768;
assign n141 = n330 | n764;
assign n1446 = ~n412;
assign n1624 = ~n159;
assign n713 = ~n1560;
assign n887 = n1527 & n1009;
assign n1335 = ~n1061;
assign n1679 = n876 | n266;
assign n725 = n997 | n1719;
assign n982 = ~(n667 | n1000);
assign n1244 = ~(n1389 ^ n812);
assign n298 = ~(n1185 ^ n954);
assign n128 = n148 | n1500;
assign n1123 = ~n952;
assign n1200 = n1358 | n943;
assign n610 = ~(n1354 ^ n165);
assign n1238 = n1532 | n1058;
assign n1159 = n1596 & n146;
assign n1227 = n1744 & n394;
assign n651 = n688 & n1097;
assign n867 = ~(n392 ^ n1538);
assign n161 = n1723 & n1505;
assign n994 = n603 | n59;
assign n823 = ~(n651 ^ n1730);
assign n1421 = ~n877;
assign n822 = ~(n952 | n414);
assign n769 = ~(n472 | n197);
assign n739 = ~(n200 | n73);
assign n240 = ~(n555 | n1448);
assign n331 = n641 | n1420;
assign n101 = ~n557;
assign n1221 = ~(n70 ^ n51);
assign n1086 = ~n609;
assign n878 = ~(n562 | n1221);
assign n1522 = n321 | n1546;
assign n1390 = ~n1045;
assign n1207 = n245 & n1132;
assign n1301 = ~(n1527 | n1208);
assign n697 = ~(n634 | n964);
assign n4 = ~n602;
assign n388 = n404 & n696;
assign n252 = n277 & n1376;
assign n1441 = ~(n875 | n45);
assign n1049 = ~(n362 ^ n400);
assign n508 = ~n709;
assign n435 = ~(n1748 ^ n340);
assign n299 = ~(n821 | n430);
assign n1494 = ~(n257 ^ n1398);
assign n91 = ~(n441 ^ n264);
assign n1633 = ~(n1467 ^ n274);
assign n1253 = ~(n1510 ^ n930);
assign n1096 = n1514 | n138;
assign n1740 = ~(n304 ^ n1537);
assign n178 = ~n1397;
assign n1375 = n54 | n1268;
assign n1273 = n642 & n897;
assign n1649 = ~(n1665 | n1667);
assign n1039 = n366 | n466;
assign n59 = ~(n1589 | n791);
assign n896 = n433 & n1342;
assign n936 = n1438 | n982;
assign n623 = ~(n314 | n333);
assign n1298 = ~n210;
assign n1306 = n1381 | n1035;
assign n1701 = ~(n825 ^ n9);
assign n588 = ~(n625 ^ n403);
assign n1188 = n878 | n1001;
assign n625 = n446 & n151;
assign n167 = n454 | n1759;
assign n328 = ~(n1734 ^ n48);
assign n1619 = n1408 | n527;
assign n276 = ~(n1210 ^ n689);
assign n1166 = ~(n562 ^ n1263);
assign n332 = n1245 | n113;
assign n574 = n910 & n88;
assign n140 = ~(n1601 | n1667);
assign n1557 = n484 | n1198;
assign n920 = n1139 & n832;
assign n1125 = ~(n952 | n729);
assign n1493 = ~n1455;
assign n1746 = ~(n635 ^ n376);
assign n812 = ~(n1443 ^ n353);
assign n842 = ~(n1770 ^ n1527);
assign n253 = ~(n439 | n1320);
assign n159 = n1263 | n211;
assign n703 = n879 & n1672;
assign n959 = ~n1214;
assign n1343 = n876 & n570;
assign n1338 = ~(n1303 ^ n630);
assign n1751 = n1478 & n963;
assign n1490 = n742 & n1726;
assign n1464 = n1082 | n658;
assign n527 = n680 & n1739;
assign n1076 = n1705 | n1318;
assign n1025 = ~(n374 ^ n1272);
assign n285 = n1339 | n435;
assign n783 = ~n973;
assign n509 = ~n612;
assign n1285 = ~n1597;
assign n1481 = ~(n1353 ^ n898);
assign n1264 = ~(n164 | n46);
assign n1071 = ~n1168;
assign n1374 = ~n98;
assign n1271 = n1078 | n873;
assign n1190 = n339 | n499;
assign n315 = ~n652;
assign n1626 = ~(n1318 ^ n409);
assign n261 = ~n1693;
assign n652 = n84 & n672;
assign n475 = ~(n374 | n1179);
assign n324 = n1468 & n1105;
assign n1610 = n1258 | n427;
assign n622 = ~(n1643 ^ n761);
assign n464 = ~(n1571 ^ n786);
assign n490 = ~n612;
assign n197 = ~n249;
assign n1043 = ~(n805 | n24);
assign n532 = n1292 | n545;
assign n337 = n1266 & n1612;
assign n1466 = ~n914;
assign n1399 = ~(n1382 ^ n726);
assign n138 = ~(n397 ^ n1077);
assign n1603 = n213 & n1360;
assign n562 = ~n856;
assign n1075 = n859 & n932;
assign n894 = n485 & n1518;
assign n837 = ~(n1230 | n4);
assign n1228 = n18 | n217;
assign n1568 = ~(n1610 ^ n49);
assign n880 = ~n459;
assign n1462 = ~n324;
assign n1078 = ~(n441 ^ n1095);
assign n1267 = ~(n98 ^ n69);
assign n1258 = n1643 & n469;
assign n939 = ~n1140;
assign n1705 = ~(n555 | n1140);
assign n19 = ~(n196 ^ n1262);
assign n275 = n147 | n1091;
assign n1033 = ~(n1252 ^ n1760);
assign n1236 = n1381 | n357;
assign n1504 = ~(n1576 | n565);
assign n1646 = ~n354;
assign n1314 = ~(n959 ^ n675);
assign n737 = ~(n459 ^ n890);
assign n795 = ~n1581;
assign n380 = n1384 | n13;
assign n1535 = ~(n817 ^ n1570);
assign n1668 = ~(n1014 ^ n1341);
assign n1042 = n1211 & n1050;
assign n492 = ~(n1160 | n1316);
assign n1080 = n359 | n560;
assign n941 = ~(n1512 ^ n1597);
assign n1721 = ~n680;
assign n27 = ~n1485;
assign n722 = ~(n487 ^ n1757);
assign n133 = n1427 | n1696;
assign n1474 = n1484 | n623;
assign n1024 = n235 | n782;
assign n94 = ~n781;
assign n1662 = n8 & n1279;
assign n1526 = n379 & n130;
assign n1371 = ~n900;
assign n813 = ~(n1334 ^ n1302);
assign n1574 = n52 | n63;
assign n577 = n1415 & n658;
assign n116 = ~(n1634 | n1555);
assign n1059 = ~(n1147 ^ n1046);
assign n855 = ~(n1643 | n1034);
assign n592 = n1000 | n1094;
assign n1670 = ~n1287;
assign n135 = ~(n425 ^ n468);
assign n359 = ~n353;
assign n1666 = n1643 & n36;
assign n1197 = n164 | n1526;
assign n392 = n256 & n1133;
assign n1215 = n5 | n15;
assign n60 = n1704 | n138;
assign n1277 = ~(n908 ^ n1249);
assign n1164 = ~(n1216 ^ n677);
assign n1413 = n128 & n92;
assign n330 = ~n170;
assign n545 = ~n719;
assign n1219 = ~n1712;
assign n885 = ~(n781 | n24);
assign n563 = ~(n164 | n66);
assign n220 = ~n1530;
assign n195 = ~(n810 ^ n391);
assign n1179 = n584 & n1664;
assign n1417 = ~(n164 | n1435);
assign n1724 = n1427 | n494;
assign n1118 = ~(n1086 ^ n842);
assign n612 = ~(n1037 ^ n848);
assign n1063 = n490 | n1061;
assign n1524 = n1316 | n607;
assign n1098 = ~(n410 ^ n663);
assign n1482 = n1715 | n338;
assign n390 = n315 & n1248;
assign n781 = ~(n987 ^ n1622);
assign n323 = n975 & n1574;
assign n198 = n1643 & n1707;
assign n1281 = n1024 & n709;
assign n740 = ~(n353 | n1360);
assign n1768 = ~n1642;
assign n7 = n182 | n595;
assign n963 = n371 | n266;
assign n1611 = n1422 | n159;
assign n18 = ~n1709;
assign n1714 = ~(n509 ^ n964);
assign n1069 = ~n949;
assign n104 = ~n407;
assign n817 = n1242 & n7;
assign n1479 = ~n303;
assign n724 = ~(n258 ^ n145);
assign n730 = ~(n564 ^ n1372);
assign n987 = n1411 | n1572;
assign n445 = ~(n1722 | n772);
assign n1347 = ~(n993 ^ n1753);
assign n945 = n1107 | n822;
assign n326 = n586 & n136;
assign n375 = n1554 & n124;
assign n1750 = ~(n180 ^ n622);
assign n1010 = ~(n1443 ^ n444);
assign n542 = n1251 & n1345;
assign n295 = n0 | n1618;
assign n646 = ~n1155;
assign n438 = ~(n1607 ^ n931);
assign n1089 = ~n927;
assign n780 = ~n1376;
assign n203 = ~(n1107 ^ n700);
assign n1193 = ~n736;
assign n80 = ~(n1423 | n1316);
assign n1593 = ~n1060;
assign n1453 = n140 | n553;
assign n214 = n739 | n734;
assign n640 = ~(n1381 | n1006);
assign n250 = ~n1541;
assign n1072 = ~n1757;
assign n283 = n369 & n733;
assign n82 = n1057 & n463;
assign n1566 = n1229 | n1591;
assign n1540 = n155 & n266;
assign n1361 = ~n1459;
assign n407 = ~(n501 ^ n708);
assign n515 = ~n1033;
assign n1120 = ~(n996 ^ n1051);
assign n1291 = ~(n154 | n970);
assign n745 = n949 & n1071;
assign n1255 = ~n647;
assign n1092 = ~(n1659 | n1197);
assign n1389 = n1754 & n25;
assign n1578 = ~(n934 ^ n732);
assign n989 = ~(n1137 ^ n1299);
assign n1225 = n649 & n1182;
assign n1726 = ~n1039;
assign n758 = n266 | n887;
assign n554 = ~(n1252 | n418);
assign n342 = ~n1297;
assign n628 = n127 | n1298;
assign n319 = ~(n805 ^ n764);
assign n149 = n439 & n1320;
assign n61 = ~n1009;
assign n1254 = n1607 | n576;
assign n944 = ~(n1042 ^ n904);
assign n1533 = n763 | n841;
assign n1584 = ~(n1448 ^ n1360);
assign n1094 = n1447 & n940;
assign n1097 = n746 | n1031;
assign n1520 = ~n827;
assign n147 = n1461 & n266;
assign n425 = n901 & n992;
assign n1426 = ~n547;
assign n1293 = ~(n971 | n1396);
assign n1151 = ~(n1468 ^ n1445);
assign n263 = ~(n584 ^ n516);
assign n102 = ~(n353 | n498);
assign n587 = ~n1424;
assign n1483 = n937 | n917;
assign n798 = ~n745;
assign n11 = n835 | n153;
assign n230 = ~n706;
assign n1663 = ~n1619;
assign n1616 = n46 | n940;
assign n672 = n1381 | n621;
assign n248 = ~(n353 ^ n1351);
assign n412 = n777 | n186;
assign n700 = ~(n952 ^ n414);
assign n1034 = ~n1751;
assign n1370 = n666 | n365;
assign n1114 = n1230 & n4;
assign n1734 = ~(n12 ^ n1176);
assign n1362 = n1582 & n72;
assign n667 = ~n347;
assign n226 = n809 | n1732;
assign n1183 = ~n1237;
assign n1261 = n825 | n1164;
assign n1661 = ~n531;
assign n1674 = n1532 | n1641;
assign n866 = ~(n26 | n296);
assign n413 = ~n307;
assign n768 = n1422 & n1624;
assign n431 = n1488 | n1011;
assign n394 = ~n318;
assign n926 = ~n1263;
assign n785 = ~(n555 ^ n788);
assign n1732 = n1072 | n487;
assign n629 = ~n681;
assign n1440 = n643 & n990;
assign n512 = n1604 | n818;
assign n466 = n1468 | n1700;
assign n847 = n807 & n1439;
assign n362 = ~n1655;
assign n510 = ~(n1546 ^ n263);
assign n269 = ~(n544 ^ n1642);
assign n416 = ~n179;
assign n1695 = ~(n165 | n1354);
assign n1035 = ~(n870 | n402);
assign n705 = ~(n837 | n1143);
assign n1579 = ~(n272 ^ n857);
assign n689 = ~(n1604 ^ n716);
assign n264 = n720 | n518;
assign n1617 = n247 & n201;
assign n205 = n203 | n1270;
assign n891 = ~(n1165 ^ n707);
assign n1583 = n143 | n1285;
assign n103 = ~(n1280 ^ n787);
assign n363 = ~(n1219 | n1672);
assign n52 = ~(n1770 | n4);
assign n1627 = ~(n1329 | n1000);
assign n797 = n1558 | n1212;
assign n998 = n363 | n1309;
assign n635 = n62 & n598;
assign n106 = n156 ^ n95;
assign n1598 = ~n1672;
assign n773 = ~n1543;
assign n709 = n1527 | n1616;
assign n575 = ~(n1280 ^ n1217);
assign n311 = n1765 & n502;
assign n1393 = ~(n1656 ^ n1064);
assign n1472 = n335 ^ n557;
assign n1038 = n1761 | n313;
assign n854 = n613 & n679;
assign n415 = ~(n952 | n1296);
assign n1355 = ~(n1422 | n266);
assign n1019 = n108 | n1419;
assign n1547 = n1504 | n434;
assign n1032 = ~(n562 ^ n1578);
assign n602 = ~(n111 ^ n1136);
assign n126 = n580 ^ n1385;
assign n176 = n1000 | n690;
assign n1427 = n1735 & n85;
assign n613 = ~(n1493 ^ n1747);
assign n913 = ~(n1513 | n1167);
assign n1564 = ~n749;
assign n663 = ~n993;
assign n949 = ~(n1607 ^ n684);
assign n692 = n1223 & n250;
assign n1465 = n1059 | n818;
assign n1262 = ~(n1576 ^ n24);
assign n1358 = ~(n1174 | n351);
assign n1036 = n1428 | n1125;
assign n845 = ~n1364;
assign n1612 = ~n1717;
assign n922 = n359 | n327;
assign n1412 = n520 | n1210;
assign n1551 = n266 | n1648;
assign n132 = ~n1253;
assign n64 = ~n93;
assign n860 = n681 | n1560;
assign n1313 = n530 | n377;
assign n974 = n35 & n907;
assign n1752 = ~(n914 ^ n138);
assign n1525 = ~(n1719 ^ n1683);
assign n1153 = ~n1296;
assign n1160 = ~n585;
assign n196 = ~n1075;
assign n1204 = ~(n666 ^ n288);
assign n40 = ~(n210 ^ n17);
assign n670 = ~(n816 ^ n138);
assign n420 = n1000 | n1281;
assign n1717 = ~(n1744 ^ n1459);
assign n516 = ~n386;
assign n1478 = n377 | n1167;
assign n110 = ~(n353 | n98);
assign n145 = ~n428;
endmodule
