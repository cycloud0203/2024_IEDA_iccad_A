
module top_810026173_843396535_809698999_829556405_809567927 (n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089, n27104, n27120, n27134, n27188, n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298, n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548, n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819, n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984, n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196, n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518, n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703, n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891, n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105, n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374, n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555, n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703, n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929, n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125, n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332, n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555, n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755, n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932, n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103, n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173, n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340, n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552, n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770, n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952, n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120, n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325, n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564, n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742, n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911, n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084, n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271, n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407, n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558, n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655, n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802, n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983, n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236, n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349, n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558, n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643, n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834, n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031, n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149, n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339, n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519, n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744, n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911, n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129, n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308, n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451, n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633, n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767, n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919, n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101, n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295, n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387, n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525, n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653, n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851, n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078, n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138, n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326, n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398, n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515, n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710, n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843, n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157, n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304, n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397, n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540, n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665, n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783, n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904, n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043, n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168, n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407, n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501, n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754, n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059, n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190, n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342, n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475, n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763, n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944, n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052, n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180, n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353, n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470, n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573, n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793, n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889, n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062, n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215, n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350, n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433, n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527, n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656, n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841, n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075, n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202, n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344, n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450, n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592, n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855, n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976, n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152, n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310, n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414, n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515, n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679, n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830, n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919, n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141, n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233, n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385, n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523, n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749, n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923, n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086, n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330, n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441, n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602, n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691, n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761, n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936, n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154, n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238, n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404, n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665, n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874, n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076, n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157, n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484, n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714, n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903, n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014, n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289, n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433, n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619, n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719, n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942, n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097, n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167, n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342, n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476, n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626, n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826, n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032, n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215, n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362, n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550, n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773, n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938, n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179, n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375, n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598, n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719, n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815, n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943, n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096, n27110, n27112, n27130, n27145, n27158, n27163, n27194);
input n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089, n27104, n27120, n27134, n27188;
output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298, n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548, n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819, n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984, n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196, n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518, n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703, n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891, n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105, n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374, n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555, n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703, n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929, n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125, n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332, n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555, n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755, n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932, n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103, n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173, n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340, n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552, n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770, n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952, n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120, n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325, n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564, n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742, n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911, n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084, n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271, n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407, n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558, n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655, n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802, n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983, n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236, n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349, n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558, n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643, n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834, n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031, n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149, n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339, n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519, n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744, n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911, n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129, n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308, n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451, n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633, n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767, n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919, n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101, n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295, n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387, n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525, n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653, n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851, n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078, n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138, n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326, n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398, n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515, n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710, n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843, n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157, n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304, n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397, n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540, n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665, n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783, n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904, n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043, n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168, n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407, n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501, n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754, n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059, n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190, n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342, n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475, n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763, n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944, n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052, n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180, n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353, n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470, n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573, n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793, n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889, n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062, n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215, n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350, n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433, n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527, n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656, n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841, n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075, n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202, n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344, n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450, n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592, n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855, n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976, n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152, n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310, n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414, n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515, n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679, n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830, n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919, n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141, n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233, n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385, n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523, n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749, n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923, n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086, n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330, n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441, n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602, n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691, n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761, n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936, n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154, n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238, n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404, n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665, n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874, n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076, n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157, n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484, n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714, n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903, n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014, n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289, n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433, n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619, n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719, n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942, n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097, n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167, n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342, n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476, n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626, n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826, n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032, n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215, n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362, n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550, n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773, n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938, n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179, n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375, n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598, n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719, n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815, n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943, n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096, n27110, n27112, n27130, n27145, n27158, n27163, n27194;
wire n0, n1, n2, n3, n4, n5, n6, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n19, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n236, n237, n238, n239, n240, n241, n244, n245, n246, n247, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n330, n331, n333, n334, n335, n336, n338, n339, n340, n341, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n423, n424, n425, n426, n427, n428, n429, n430, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n458, n459, n460, n461, n462, n464, n465, n466, n467, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n492, n493, n494, n495, n497, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n549, n550, n551, n552, n553, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n584, n585, n586, n587, n589, n590, n591, n592, n593, n594, n595, n596, n598, n599, n600, n601, n602, n603, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n638, n639, n640, n641, n642, n643, n644, n645, n648, n649, n650, n651, n652, n653, n654, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n810, n811, n812, n813, n814, n815, n816, n817, n818, n820, n821, n822, n823, n824, n825, n826, n827, n828, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n850, n851, n852, n853, n854, n855, n856, n857, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n874, n875, n876, n877, n878, n880, n881, n882, n883, n884, n885, n886, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n949, n950, n951, n952, n953, n954, n955, n956, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n981, n983, n985, n986, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1017, n1018, n1019, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1041, n1042, n1043, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1113, n1114, n1115, n1116, n1117, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1238, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1289, n1290, n1291, n1292, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1315, n1316, n1317, n1318, n1319, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1433, n1434, n1435, n1436, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1499, n1500, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1519, n1520, n1521, n1522, n1523, n1524, n1526, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1581, n1582, n1583, n1584, n1585, n1587, n1588, n1589, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1631, n1632, n1633, n1635, n1637, n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1663, n1664, n1665, n1666, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1683, n1685, n1686, n1687, n1688, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1702, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1739, n1740, n1741, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1943, n1944, n1945, n1946, n1947, n1948, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n2000, n2001, n2002, n2003, n2005, n2006, n2008, n2009, n2010, n2011, n2012, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2089, n2090, n2091, n2093, n2094, n2096, n2097, n2098, n2099, n2100, n2101, n2103, n2104, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2114, n2115, n2116, n2118, n2119, n2120, n2121, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2211, n2212, n2213, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2329, n2330, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2356, n2357, n2358, n2359, n2360, n2362, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2410, n2411, n2412, n2413, n2414, n2415, n2417, n2418, n2419, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2441, n2442, n2443, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2514, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2534, n2536, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2548, n2549, n2550, n2551, n2552, n2554, n2556, n2557, n2558, n2559, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2571, n2572, n2574, n2575, n2576, n2577, n2579, n2580, n2581, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2660, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2704, n2705, n2707, n2708, n2709, n2710, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2775, n2776, n2777, n2778, n2780, n2781, n2782, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2810, n2811, n2812, n2813, n2814, n2815, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2854, n2855, n2856, n2857, n2859, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2945, n2946, n2947, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2972, n2973, n2974, n2975, n2976, n2977, n2980, n2981, n2982, n2983, n2984, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3011, n3012, n3013, n3014, n3015, n3016, n3019, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3162, n3163, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3229, n3230, n3231, n3232, n3233, n3234, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3254, n3255, n3256, n3257, n3258, n3259, n3261, n3262, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3302, n3303, n3304, n3305, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3317, n3318, n3319, n3321, n3322, n3323, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3341, n3342, n3344, n3345, n3346, n3347, n3348, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3503, n3504, n3505, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3556, n3557, n3558, n3559, n3560, n3562, n3564, n3565, n3566, n3567, n3568, n3569, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3643, n3644, n3645, n3646, n3647, n3648, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3734, n3735, n3736, n3737, n3738, n3739, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3756, n3757, n3759, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3782, n3783, n3784, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3870, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3919, n3920, n3921, n3922, n3923, n3924, n3926, n3927, n3928, n3929, n3930, n3931, n3933, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3946, n3947, n3948, n3949, n3950, n3951, n3953, n3954, n3955, n3956, n3957, n3958, n3960, n3961, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4011, n4012, n4013, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4086, n4087, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4101, n4102, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4120, n4121, n4122, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4147, n4148, n4149, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4166, n4167, n4168, n4169, n4170, n4171, n4174, n4175, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4216, n4217, n4218, n4219, n4220, n4222, n4223, n4225, n4226, n4227, n4228, n4229, n4230, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4267, n4268, n4269, n4270, n4271, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4320, n4321, n4322, n4323, n4324, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4375, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4425, n4427, n4428, n4429, n4430, n4431, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4477, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4589, n4591, n4592, n4593, n4594, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4746, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4767, n4768, n4769, n4771, n4772, n4773, n4774, n4775, n4776, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4805, n4806, n4807, n4808, n4809, n4811, n4813, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4948, n4949, n4950, n4951, n4953, n4954, n4955, n4956, n4958, n4959, n4960, n4961, n4962, n4963, n4965, n4968, n4969, n4970, n4971, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5021, n5022, n5023, n5027, n5028, n5029, n5030, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5061, n5063, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5078, n5079, n5080, n5081, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5099, n5100, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5116, n5117, n5118, n5119, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5129, n5130, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5212, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5227, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5301, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5326, n5327, n5328, n5329, n5331, n5332, n5333, n5334, n5335, n5336, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5352, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5401, n5402, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5440, n5441, n5442, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5518, n5519, n5520, n5522, n5523, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5604, n5606, n5607, n5608, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5681, n5682, n5683, n5684, n5685, n5686, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5697, n5698, n5699, n5701, n5702, n5703, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5777, n5778, n5779, n5780, n5781, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5835, n5836, n5837, n5838, n5839, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5905, n5906, n5907, n5908, n5909, n5910, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5937, n5938, n5939, n5940, n5941, n5942, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6045, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6184, n6185, n6186, n6187, n6188, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6219, n6220, n6221, n6222, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6246, n6247, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6272, n6273, n6274, n6275, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6309, n6310, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6324, n6325, n6326, n6327, n6328, n6329, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6355, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6370, n6371, n6372, n6373, n6374, n6376, n6377, n6378, n6380, n6382, n6384, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6428, n6429, n6430, n6432, n6433, n6434, n6435, n6436, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6466, n6467, n6468, n6469, n6471, n6472, n6473, n6474, n6475, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6503, n6504, n6505, n6507, n6508, n6509, n6510, n6511, n6512, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6557, n6559, n6561, n6562, n6563, n6564, n6565, n6566, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6588, n6589, n6591, n6592, n6593, n6594, n6595, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6629, n6632, n6633, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6653, n6654, n6656, n6657, n6658, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6670, n6672, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6685, n6686, n6687, n6688, n6689, n6690, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6730, n6731, n6732, n6733, n6734, n6735, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6774, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6786, n6787, n6788, n6789, n6792, n6793, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6864, n6865, n6866, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6966, n6968, n6969, n6970, n6972, n6973, n6974, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6984, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7027, n7028, n7029, n7030, n7031, n7033, n7034, n7035, n7036, n7037, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7231, n7232, n7234, n7235, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7254, n7255, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7278, n7279, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7299, n7300, n7301, n7302, n7303, n7304, n7306, n7307, n7309, n7310, n7311, n7312, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7331, n7332, n7333, n7334, n7336, n7337, n7338, n7340, n7341, n7342, n7343, n7344, n7345, n7347, n7348, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7404, n7405, n7406, n7407, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7422, n7423, n7424, n7425, n7426, n7427, n7429, n7430, n7431, n7433, n7434, n7435, n7436, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7476, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7508, n7509, n7510, n7511, n7512, n7513, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7567, n7568, n7570, n7571, n7573, n7574, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7586, n7587, n7589, n7590, n7591, n7592, n7594, n7595, n7596, n7597, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7608, n7609, n7611, n7612, n7613, n7614, n7615, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7644, n7645, n7646, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7671, n7672, n7673, n7675, n7676, n7677, n7680, n7681, n7682, n7683, n7684, n7685, n7687, n7688, n7689, n7690, n7691, n7694, n7695, n7696, n7697, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7770, n7771, n7772, n7774, n7775, n7776, n7777, n7778, n7779, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7789, n7790, n7791, n7792, n7793, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7831, n7832, n7833, n7835, n7836, n7837, n7838, n7839, n7840, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7938, n7939, n7940, n7941, n7942, n7944, n7945, n7946, n7947, n7948, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7960, n7961, n7962, n7964, n7965, n7966, n7967, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7993, n7994, n7995, n7996, n7997, n7998, n8000, n8001, n8002, n8003, n8004, n8005, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8028, n8029, n8030, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8104, n8105, n8106, n8107, n8108, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8128, n8129, n8131, n8132, n8133, n8134, n8136, n8137, n8138, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8257, n8258, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8286, n8287, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8307, n8308, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8322, n8323, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8377, n8378, n8379, n8380, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8400, n8401, n8402, n8403, n8404, n8406, n8407, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8433, n8434, n8435, n8436, n8437, n8438, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8506, n8507, n8508, n8509, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8520, n8521, n8522, n8523, n8524, n8525, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8609, n8610, n8611, n8612, n8613, n8615, n8616, n8617, n8618, n8619, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8657, n8658, n8659, n8660, n8661, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8688, n8689, n8690, n8691, n8692, n8693, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8717, n8718, n8719, n8720, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8804, n8805, n8807, n8808, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8822, n8823, n8825, n8826, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8850, n8851, n8852, n8853, n8854, n8855, n8857, n8858, n8859, n8860, n8863, n8864, n8865, n8866, n8867, n8868, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8910, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8965, n8966, n8967, n8968, n8969, n8970, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9043, n9044, n9045, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9165, n9167, n9168, n9169, n9170, n9171, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9218, n9219, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9247, n9248, n9249, n9250, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9260, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9319, n9320, n9321, n9322, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9365, n9366, n9367, n9368, n9369, n9370, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9381, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9397, n9398, n9400, n9401, n9402, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9420, n9421, n9422, n9424, n9425, n9426, n9427, n9428, n9429, n9431, n9432, n9433, n9434, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9446, n9447, n9448, n9449, n9450, n9452, n9453, n9454, n9455, n9456, n9457, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9509, n9510, n9511, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9553, n9555, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9617, n9618, n9619, n9620, n9621, n9623, n9624, n9625, n9627, n9628, n9629, n9630, n9631, n9632, n9634, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9647, n9649, n9650, n9651, n9652, n9653, n9654, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9690, n9691, n9692, n9693, n9694, n9696, n9697, n9698, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9762, n9764, n9765, n9766, n9768, n9769, n9770, n9772, n9773, n9774, n9775, n9776, n9777, n9779, n9780, n9781, n9782, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9834, n9835, n9836, n9837, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9868, n9869, n9870, n9871, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9918, n9920, n9921, n9922, n9923, n9924, n9925, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9935, n9936, n9937, n9939, n9940, n9941, n9943, n9944, n9945, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10011, n10012, n10013, n10014, n10015, n10016, n10020, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10054, n10056, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10097, n10098, n10099, n10100, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10112, n10113, n10114, n10115, n10116, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10159, n10160, n10161, n10162, n10163, n10164, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10237, n10238, n10240, n10241, n10242, n10243, n10245, n10246, n10247, n10248, n10249, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10322, n10323, n10324, n10325, n10328, n10329, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10341, n10342, n10343, n10344, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10386, n10389, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10406, n10407, n10408, n10410, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10485, n10486, n10487, n10488, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10562, n10563, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10589, n10590, n10591, n10592, n10594, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10612, n10613, n10615, n10616, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10648, n10649, n10651, n10652, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10693, n10695, n10696, n10697, n10698, n10699, n10700, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10711, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10757, n10758, n10759, n10760, n10761, n10762, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10776, n10777, n10778, n10779, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11006, n11007, n11008, n11009, n11010, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11024, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11057, n11058, n11059, n11060, n11061, n11062, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11079, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11095, n11096, n11097, n11098, n11099, n11100, n11102, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11122, n11123, n11124, n11125, n11126, n11128, n11129, n11130, n11131, n11133, n11135, n11136, n11137, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11183, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11221, n11222, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11262, n11263, n11264, n11265, n11267, n11268, n11269, n11270, n11271, n11272, n11274, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11327, n11328, n11329, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11349, n11350, n11351, n11353, n11354, n11355, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11376, n11377, n11378, n11380, n11381, n11382, n11383, n11384, n11385, n11387, n11388, n11389, n11390, n11392, n11393, n11394, n11395, n11396, n11397, n11399, n11400, n11401, n11402, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11420, n11421, n11422, n11423, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11456, n11457, n11458, n11459, n11460, n11461, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11471, n11474, n11475, n11476, n11477, n11478, n11480, n11482, n11483, n11484, n11485, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11497, n11498, n11499, n11500, n11501, n11502, n11504, n11505, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11565, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11668, n11669, n11670, n11671, n11672, n11673, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11711, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11737, n11738, n11739, n11740, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11772, n11773, n11774, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11838, n11839, n11840, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11899, n11900, n11901, n11902, n11903, n11904, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12001, n12002, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12147, n12148, n12149, n12150, n12151, n12154, n12155, n12156, n12159, n12160, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12224, n12226, n12227, n12229, n12230, n12231, n12232, n12233, n12234, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12303, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12326, n12327, n12328, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12342, n12343, n12344, n12345, n12347, n12348, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12381, n12382, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12447, n12448, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12463, n12464, n12465, n12466, n12468, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12541, n12542, n12543, n12544, n12547, n12548, n12549, n12550, n12551, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12563, n12564, n12565, n12567, n12568, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12588, n12589, n12590, n12591, n12592, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12622, n12623, n12624, n12625, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12651, n12652, n12653, n12655, n12656, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12666, n12667, n12668, n12669, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12703, n12704, n12705, n12706, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12726, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12741, n12743, n12744, n12745, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12813, n12814, n12815, n12817, n12818, n12819, n12820, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12862, n12863, n12866, n12867, n12868, n12869, n12872, n12874, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12901, n12902, n12903, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12979, n12981, n12982, n12983, n12984, n12986, n12988, n12989, n12990, n12991, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13045, n13046, n13047, n13049, n13050, n13051, n13052, n13053, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13111, n13112, n13113, n13114, n13115, n13117, n13118, n13119, n13120, n13121, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13138, n13139, n13140, n13142, n13143, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13200, n13201, n13202, n13203, n13205, n13206, n13207, n13208, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13264, n13265, n13266, n13267, n13268, n13269, n13271, n13272, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13334, n13335, n13336, n13337, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13408, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13420, n13421, n13422, n13423, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13454, n13455, n13458, n13459, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13478, n13479, n13480, n13481, n13482, n13483, n13485, n13488, n13489, n13491, n13492, n13493, n13495, n13496, n13497, n13498, n13499, n13502, n13503, n13504, n13505, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13550, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13678, n13679, n13680, n13681, n13682, n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13709, n13711, n13712, n13713, n13715, n13716, n13717, n13718, n13720, n13721, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13776, n13777, n13778, n13779, n13780, n13782, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13913, n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14091, n14092, n14093, n14094, n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14122, n14123, n14124, n14125, n14127, n14128, n14129, n14131, n14132, n14133, n14134, n14135, n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14268, n14269, n14270, n14272, n14273, n14274, n14276, n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14324, n14325, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14343, n14344, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14413, n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14458, n14459, n14460, n14461, n14462, n14463, n14465, n14466, n14467, n14468, n14469, n14470, n14472, n14473, n14474, n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14542, n14543, n14544, n14545, n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14571, n14572, n14573, n14574, n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14634, n14635, n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14681, n14682, n14683, n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14703, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14820, n14821, n14822, n14823, n14824, n14825, n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15003, n15005, n15006, n15007, n15008, n15009, n15010, n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15032, n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15078, n15079, n15080, n15081, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15140, n15141, n15142, n15143, n15144, n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15166, n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15177, n15178, n15179, n15181, n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15256, n15257, n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15272, n15273, n15274, n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15301, n15302, n15303, n15304, n15305, n15306, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15328, n15329, n15330, n15331, n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15379, n15380, n15381, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15425, n15426, n15427, n15429, n15430, n15431, n15432, n15433, n15434, n15436, n15437, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15466, n15468, n15469, n15471, n15472, n15473, n15474, n15475, n15476, n15478, n15479, n15480, n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15491, n15492, n15493, n15494, n15495, n15497, n15498, n15499, n15500, n15502, n15503, n15504, n15505, n15507, n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15540, n15541, n15542, n15543, n15544, n15545, n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15556, n15557, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15571, n15572, n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15589, n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15599, n15600, n15601, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15744, n15745, n15746, n15747, n15748, n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15763, n15764, n15765, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15813, n15814, n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15886, n15887, n15888, n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15919, n15920, n15921, n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15957, n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15980, n15981, n15982, n15983, n15984, n15985, n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16061, n16063, n16064, n16065, n16066, n16067, n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16216, n16220, n16221, n16222, n16224, n16225, n16226, n16227, n16228, n16229, n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16244, n16245, n16246, n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16276, n16277, n16278, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16323, n16324, n16325, n16326, n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16377, n16378, n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16397, n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16420, n16421, n16422, n16423, n16425, n16426, n16427, n16429, n16430, n16431, n16432, n16434, n16435, n16436, n16437, n16438, n16441, n16442, n16443, n16444, n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16477, n16478, n16479, n16480, n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16503, n16504, n16505, n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16518, n16519, n16520, n16522, n16523, n16525, n16526, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16585, n16586, n16587, n16588, n16590, n16591, n16592, n16593, n16594, n16595, n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16683, n16685, n16686, n16687, n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16813, n16814, n16815, n16816, n16817, n16819, n16820, n16821, n16822, n16823, n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16835, n16836, n16838, n16839, n16840, n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16906, n16907, n16908, n16909, n16910, n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16952, n16953, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16969, n16970, n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16990, n16991, n16992, n16993, n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17036, n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17071, n17072, n17073, n17074, n17076, n17078, n17079, n17080, n17081, n17082, n17083, n17085, n17086, n17087, n17088, n17089, n17091, n17092, n17093, n17094, n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17105, n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17164, n17165, n17166, n17167, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17233, n17234, n17235, n17237, n17238, n17239, n17240, n17241, n17242, n17244, n17245, n17246, n17247, n17248, n17249, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17338, n17339, n17340, n17341, n17342, n17343, n17345, n17346, n17347, n17348, n17349, n17350, n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17388, n17389, n17390, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17433, n17434, n17435, n17437, n17438, n17439, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17459, n17460, n17462, n17463, n17464, n17465, n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17494, n17495, n17496, n17497, n17498, n17499, n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17525, n17526, n17527, n17528, n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17736, n17737, n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17747, n17748, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17928, n17929, n17930, n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17949, n17950, n17951, n17952, n17953, n17955, n17957, n17958, n17960, n17961, n17962, n17964, n17965, n17966, n17967, n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18044, n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18060, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18144, n18146, n18147, n18148, n18149, n18150, n18153, n18154, n18155, n18156, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18228, n18229, n18230, n18231, n18233, n18234, n18235, n18236, n18237, n18239, n18240, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18289, n18291, n18292, n18293, n18294, n18296, n18297, n18298, n18299, n18300, n18302, n18303, n18305, n18306, n18307, n18308, n18309, n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18344, n18346, n18347, n18348, n18349, n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18406, n18407, n18408, n18410, n18411, n18412, n18413, n18415, n18416, n18417, n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18438, n18440, n18441, n18442, n18443, n18446, n18447, n18448, n18449, n18450, n18451, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18510, n18511, n18512, n18514, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18573, n18575, n18577, n18579, n18580, n18581, n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18650, n18651, n18652, n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678, n18680, n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18691, n18692, n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18722, n18723, n18724, n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18746, n18747, n18748, n18749, n18750, n18752, n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18781, n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18832, n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18860, n18861, n18862, n18863, n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18881, n18882, n18883, n18884, n18885, n18888, n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18902, n18903, n18904, n18905, n18906, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18920, n18921, n18922, n18923, n18924, n18925, n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18941, n18942, n18943, n18944, n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18971, n18972, n18973, n18974, n18975, n18976, n18978, n18979, n18980, n18981, n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998, n19000, n19001, n19002, n19003, n19004, n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19043, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19142, n19143, n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19175, n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19197, n19198, n19199, n19200, n19201, n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19222, n19225, n19226, n19227, n19229, n19230, n19231, n19232, n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19324, n19325, n19326, n19328, n19329, n19330, n19331, n19332, n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19349, n19350, n19351, n19352, n19353, n19355, n19356, n19358, n19359, n19360, n19362, n19363, n19364, n19365, n19366, n19368, n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19386, n19387, n19388, n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19451, n19452, n19453, n19455, n19456, n19457, n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19468, n19469, n19470, n19471, n19473, n19474, n19475, n19476, n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19495, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19571, n19572, n19573, n19574, n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19603, n19604, n19605, n19606, n19607, n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19619, n19620, n19621, n19622, n19624, n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19642, n19643, n19644, n19645, n19646, n19647, n19649, n19650, n19651, n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19750, n19751, n19752, n19753, n19754, n19755, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766, n19768, n19769, n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19790, n19791, n19793, n19794, n19795, n19796, n19797, n19799, n19800, n19801, n19802, n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19906, n19907, n19908, n19910, n19912, n19913, n19914, n19915, n19917, n19918, n19919, n19920, n19921, n19924, n19925, n19926, n19927, n19928, n19929, n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20014, n20015, n20016, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20034, n20035, n20037, n20038, n20039, n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20097, n20098, n20099, n20100, n20101, n20102, n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20150, n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20331, n20332, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20350, n20351, n20352, n20353, n20354, n20356, n20357, n20358, n20360, n20361, n20362, n20363, n20364, n20365, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20386, n20387, n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20404, n20405, n20406, n20407, n20408, n20410, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, n20423, n20425, n20426, n20427, n20428, n20430, n20431, n20432, n20433, n20434, n20435, n20437, n20438, n20439, n20440, n20442, n20443, n20444, n20446, n20447, n20448, n20449, n20451, n20452, n20453, n20454, n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20491, n20492, n20493, n20494, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20603, n20605, n20606, n20607, n20608, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622, n20624, n20625, n20626, n20627, n20628, n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20659, n20660, n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20674, n20675, n20676, n20677, n20679, n20681, n20682, n20683, n20684, n20686, n20687, n20688, n20689, n20690, n20692, n20693, n20694, n20695, n20697, n20698, n20699, n20701, n20702, n20703, n20706, n20707, n20708, n20710, n20711, n20712, n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20789, n20790, n20791, n20792, n20793, n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20924, n20925, n20926, n20927, n20928, n20930, n20931, n20932, n20933, n20934, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21135, n21136, n21137, n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21155, n21156, n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21169, n21170, n21171, n21172, n21174, n21175, n21177, n21178, n21179, n21180, n21181, n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21223, n21224, n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21277, n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21299, n21300, n21301, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21366, n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395, n21397, n21400, n21401, n21402, n21403, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21616, n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21646, n21647, n21648, n21650, n21651, n21652, n21653, n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21675, n21676, n21677, n21678, n21679, n21681, n21682, n21683, n21684, n21686, n21688, n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21718, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21736, n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21751, n21752, n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21780, n21781, n21782, n21783, n21785, n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819, n21821, n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830, n21831, n21833, n21834, n21835, n21836, n21837, n21838, n21840, n21841, n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21899, n21900, n21901, n21902, n21903, n21904, n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21958, n21959, n21961, n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974, n21975, n21977, n21978, n21979, n21980, n21982, n21983, n21984, n21985, n21987, n21988, n21989, n21990, n21991, n21992, n21994, n21995, n21996, n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22044, n22045, n22046, n22047, n22048, n22049, n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062, n22064, n22065, n22066, n22067, n22069, n22070, n22071, n22073, n22074, n22075, n22077, n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22108, n22109, n22110, n22111, n22112, n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22125, n22127, n22128, n22129, n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142, n22143, n22145, n22146, n22147, n22148, n22149, n22151, n22152, n22153, n22154, n22155, n22156, n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22199, n22200, n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22271, n22272, n22273, n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22284, n22285, n22286, n22287, n22288, n22289, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22310, n22312, n22313, n22314, n22315, n22316, n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331, n22333, n22334, n22336, n22337, n22338, n22339, n22340, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22354, n22355, n22356, n22357, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22443, n22445, n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22468, n22469, n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22485, n22486, n22487, n22488, n22490, n22491, n22493, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583, n22585, n22586, n22587, n22590, n22592, n22593, n22594, n22595, n22596, n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22621, n22622, n22624, n22625, n22627, n22628, n22629, n22630, n22632, n22633, n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659, n22661, n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22762, n22763, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22788, n22789, n22790, n22791, n22792, n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22880, n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22892, n22893, n22894, n22895, n22896, n22898, n22899, n22900, n22901, n22902, n22904, n22905, n22906, n22908, n22909, n22911, n22912, n22913, n22915, n22916, n22917, n22919, n22920, n22921, n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23008, n23010, n23011, n23012, n23013, n23015, n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23036, n23037, n23038, n23040, n23041, n23042, n23043, n23044, n23045, n23046, n23048, n23049, n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23059, n23060, n23061, n23062, n23063, n23064, n23069, n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118, n23119, n23121, n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159, n23161, n23162, n23163, n23164, n23165, n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198, n23199, n23201, n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246, n23249, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23271, n23273, n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303, n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23370, n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23431, n23432, n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462, n23464, n23465, n23466, n23467, n23468, n23469, n23470, n23472, n23473, n23474, n23475, n23476, n23477, n23478, n23479, n23481, n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23542, n23543, n23544, n23545, n23547, n23548, n23549, n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23587, n23589, n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23620, n23621, n23622, n23623, n23625, n23626, n23627, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23658, n23659, n23660, n23661, n23662, n23664, n23665, n23666, n23667, n23668, n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683, n23685, n23686, n23687, n23688, n23689, n23691, n23692, n23693, n23694, n23695, n23696, n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23715, n23716, n23718, n23720, n23721, n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747, n23749, n23750, n23751, n23752, n23753, n23754, n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774, n23776, n23777, n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830, n23832, n23833, n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23843, n23844, n23845, n23846, n23847, n23848, n23850, n23851, n23852, n23853, n23854, n23855, n23857, n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23884, n23885, n23886, n23887, n23889, n23890, n23891, n23892, n23893, n23894, n23896, n23897, n23898, n23900, n23901, n23902, n23904, n23905, n23906, n23907, n23908, n23909, n23910, n23911, n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934, n23936, n23937, n23938, n23939, n23940, n23941, n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23955, n23956, n23957, n23959, n23960, n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973, n23975, n23976, n23977, n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24003, n24005, n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24033, n24034, n24035, n24036, n24037, n24038, n24040, n24041, n24042, n24043, n24044, n24045, n24046, n24047, n24049, n24050, n24051, n24053, n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24086, n24087, n24088, n24089, n24090, n24091, n24094, n24095, n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117, n24118, n24120, n24121, n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24130, n24131, n24132, n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24142, n24143, n24144, n24147, n24148, n24149, n24151, n24152, n24153, n24154, n24156, n24157, n24158, n24159, n24161, n24162, n24163, n24164, n24165, n24166, n24168, n24169, n24171, n24173, n24174, n24175, n24176, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195, n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227, n24229, n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24259, n24261, n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318, n24320, n24321, n24322, n24324, n24325, n24326, n24328, n24329, n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24343, n24344, n24346, n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24416, n24417, n24418, n24419, n24420, n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430, n24432, n24433, n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470, n24471, n24473, n24474, n24475, n24477, n24478, n24479, n24480, n24481, n24482, n24484, n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510, n24511, n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575, n24577, n24578, n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24603, n24605, n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24619, n24621, n24622, n24623, n24624, n24625, n24627, n24628, n24630, n24631, n24632, n24633, n24634, n24635, n24637, n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731, n24733, n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757, n24759, n24760, n24761, n24762, n24763, n24764, n24765, n24766, n24767, n24769, n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781, n24782, n24783, n24785, n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805, n24806, n24808, n24809, n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24854, n24855, n24856, n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877, n24878, n24880, n24881, n24882, n24883, n24884, n24885, n24886, n24888, n24889, n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933, n24935, n24936, n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997, n24999, n25000, n25001, n25002, n25003, n25004, n25005, n25007, n25008, n25009, n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021, n25022, n25024, n25025, n25026, n25027, n25028, n25029, n25030, n25031, n25033, n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061, n25063, n25064, n25065, n25066, n25067, n25069, n25070, n25071, n25072, n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093, n25095, n25096, n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25121, n25122, n25123, n25124, n25125, n25127, n25128, n25129, n25130, n25131, n25132, n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165, n25166, n25167, n25169, n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25210, n25211, n25212, n25213, n25214, n25216, n25217, n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237, n25238, n25239, n25241, n25242, n25243, n25245, n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25255, n25257, n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25294, n25295, n25297, n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25317, n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326, n25327, n25329, n25330, n25333, n25334, n25335, n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355, n25357, n25358, n25359, n25360, n25361, n25363, n25364, n25366, n25367, n25368, n25369, n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411, n25413, n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25461, n25462, n25463, n25465, n25466, n25467, n25469, n25470, n25472, n25473, n25474, n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493, n25495, n25496, n25497, n25498, n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25514, n25515, n25516, n25517, n25519, n25520, n25521, n25522, n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25533, n25534, n25535, n25536, n25537, n25538, n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25551, n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25612, n25613, n25615, n25616, n25617, n25618, n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25630, n25631, n25632, n25633, n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715, n25716, n25717, n25718, n25720, n25721, n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25750, n25752, n25753, n25754, n25755, n25757, n25759, n25760, n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781, n25782, n25783, n25785, n25786, n25787, n25788, n25789, n25790, n25791, n25793, n25794, n25795, n25796, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814, n25815, n25817, n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837, n25838, n25841, n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869, n25870, n25871, n25874, n25875, n25876, n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25924, n25925, n25927, n25928, n25929, n25930, n25931, n25932, n25933, n25935, n25936, n25937, n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971, n25973, n25975, n25976, n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035, n26037, n26038, n26039, n26040, n26041, n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051, n26052, n26055, n26056, n26057, n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083, n26085, n26086, n26087, n26088, n26089, n26090, n26091, n26092, n26093, n26094, n26095, n26097, n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26108, n26109, n26110, n26112, n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155, n26157, n26158, n26160, n26161, n26162, n26163, n26164, n26165, n26166, n26168, n26169, n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26181, n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219, n26221, n26222, n26223, n26225, n26226, n26227, n26228, n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262, n26263, n26265, n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285, n26286, n26288, n26289, n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26319, n26320, n26321, n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371, n26372, n26373, n26374, n26376, n26377, n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395, n26397, n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26430, n26432, n26433, n26434, n26435, n26436, n26437, n26438, n26440, n26441, n26442, n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26453, n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491, n26493, n26494, n26495, n26496, n26497, n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509, n26511, n26513, n26514, n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563, n26564, n26566, n26567, n26568, n26569, n26570, n26571, n26573, n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589, n26591, n26592, n26593, n26594, n26595, n26596, n26597, n26599, n26600, n26601, n26602, n26603, n26604, n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653, n26654, n26655, n26657, n26658, n26659, n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26676, n26677, n26678, n26679, n26680, n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26697, n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717, n26718, n26720, n26721, n26722, n26723, n26724, n26726, n26728, n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742, n26743, n26746, n26747, n26749, n26750, n26751, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771, n26772, n26773, n26774, n26776, n26777, n26778, n26779, n26781, n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26796, n26798, n26799, n26800, n26802, n26803, n26804, n26805, n26806, n26807, n26809, n26810, n26811, n26812, n26813, n26814, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843, n26844, n26845, n26846, n26848, n26849, n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899, n26901, n26903, n26904, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26922, n26924, n26925, n26926, n26927, n26928, n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940, n26941, n26942, n26944, n26945, n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26980, n26981, n26982, n26983, n26984, n26985, n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27005, n27006, n27007, n27008, n27009, n27010, n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27032, n27033, n27034, n27035, n27036, n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27073, n27074, n27075, n27076, n27077, n27078, n27080, n27081, n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27090, n27091, n27092, n27093, n27094, n27095, n27097, n27098, n27099, n27100, n27101, n27102, n27103, n27105, n27106, n27107, n27108, n27109, n27111, n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27121, n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27131, n27132, n27133, n27135, n27136, n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157, n27159, n27160, n27161, n27162, n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187, n27189, n27190, n27191, n27192, n27193, n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205, n27206;
assign n25456 = n12222 | n17800;
assign n4950 = ~n24186;
assign n12724 = n24693 & n14425;
assign n5884 = n17333 | n19247;
assign n13231 = ~n1735;
assign n363 = n15446 | n2417;
assign n12601 = n3124 | n3018;
assign n54 = ~n21300;
assign n21820 = ~(n20820 ^ n14706);
assign n22318 = ~n12713;
assign n21745 = ~n21544;
assign n15177 = ~n13572;
assign n26507 = n22220 | n14118;
assign n11793 = n1963 | n21122;
assign n17152 = ~(n3747 ^ n21909);
assign n7943 = ~(n20710 ^ n21590);
assign n6658 = n22626 | n8583;
assign n7064 = n17471 | n6429;
assign n27148 = n11024 & n25179;
assign n20223 = n23276 | n5847;
assign n21320 = n16928 | n25210;
assign n5572 = ~n14089;
assign n21011 = n14363 | n1476;
assign n8578 = ~(n10709 ^ n18924);
assign n8495 = ~n20410;
assign n18595 = ~n12969;
assign n17670 = ~n4879;
assign n14512 = n9502 | n15705;
assign n3873 = ~(n24313 | n26728);
assign n11734 = ~(n3824 ^ n7395);
assign n3299 = ~(n23618 ^ n8329);
assign n17003 = ~(n21347 ^ n15280);
assign n2679 = n24317 & n6516;
assign n13649 = ~n3590;
assign n8887 = ~(n623 | n11195);
assign n25052 = ~(n18717 | n15155);
assign n24531 = n10568 | n18558;
assign n15082 = ~(n26753 ^ n7886);
assign n20173 = n2268 & n22417;
assign n12897 = n22856 & n10163;
assign n11091 = ~(n11016 ^ n9883);
assign n14307 = n9910 | n23272;
assign n22644 = ~n5060;
assign n21615 = ~(n7998 ^ n12883);
assign n23233 = ~n25902;
assign n8928 = n20833 | n9536;
assign n865 = n20401 | n2489;
assign n23890 = ~(n5059 ^ n14583);
assign n25890 = ~n1314;
assign n13709 = n8186 & n20797;
assign n12843 = n10218 & n4788;
assign n23844 = n5290 & n11851;
assign n16048 = n21071 | n2110;
assign n14394 = ~(n27148 ^ n18538);
assign n12328 = ~(n9594 | n8285);
assign n26628 = n17013 | n10611;
assign n21340 = ~n10493;
assign n23817 = n8105 | n14522;
assign n17139 = n8123 & n10975;
assign n18341 = ~(n3637 ^ n2783);
assign n5543 = n1522 | n14138;
assign n14935 = n20837 | n13470;
assign n1565 = ~n10660;
assign n20724 = n655 | n26253;
assign n21434 = ~n5196;
assign n4768 = n17860 & n16055;
assign n7011 = n1959 | n14473;
assign n756 = n21327 | n22876;
assign n18475 = n12342 | n16519;
assign n14183 = n14331 | n23294;
assign n15724 = n4638 & n49;
assign n4632 = ~(n1509 ^ n16521);
assign n16576 = ~(n20830 ^ n18596);
assign n4854 = ~(n19259 ^ n5749);
assign n14775 = n1176 | n3480;
assign n23867 = ~(n22278 | n7465);
assign n8044 = ~n11095;
assign n10635 = n15870 & n5748;
assign n24477 = ~(n6232 | n13472);
assign n14912 = n4494 | n19986;
assign n14542 = ~(n16065 | n26413);
assign n515 = ~(n575 ^ n3570);
assign n25252 = n22235 & n18699;
assign n10089 = n18505 & n8369;
assign n25395 = n8678 & n16500;
assign n21195 = n1041 & n13744;
assign n22762 = ~(n27037 | n20099);
assign n7811 = ~(n17890 ^ n18231);
assign n1933 = n10763 & n18799;
assign n19474 = n14744 & n17936;
assign n7927 = n13762 & n10110;
assign n9079 = n15575 & n14072;
assign n20192 = ~(n1084 ^ n21832);
assign n5519 = n2331 | n12546;
assign n21186 = n9493 | n15507;
assign n3755 = ~(n15690 ^ n14252);
assign n20468 = n9401 & n25042;
assign n13095 = ~(n12232 ^ n8526);
assign n23133 = ~(n26211 | n15583);
assign n1372 = n8309 | n24203;
assign n2668 = ~(n13137 | n7674);
assign n24057 = n161 | n24154;
assign n3922 = n22265 | n18194;
assign n2669 = ~(n7437 | n13367);
assign n2703 = ~(n11983 ^ n18667);
assign n16256 = n6341 & n23512;
assign n10723 = ~(n14032 ^ n14651);
assign n17620 = ~n1386;
assign n7046 = n18274 | n24202;
assign n16829 = ~(n17629 ^ n8317);
assign n14470 = n20566 | n18211;
assign n11876 = n4957 | n5034;
assign n14443 = n2435 & n11984;
assign n2431 = ~(n7107 ^ n5183);
assign n15706 = n23316 | n9122;
assign n5705 = n10620 | n17142;
assign n19749 = ~(n93 ^ n12777);
assign n13300 = ~(n5611 ^ n20600);
assign n5374 = ~(n26758 ^ n13026);
assign n8315 = ~(n813 ^ n19294);
assign n18433 = ~(n21479 ^ n22435);
assign n25431 = ~n25353;
assign n11971 = ~(n25146 ^ n13444);
assign n24147 = ~(n20595 ^ n2322);
assign n3882 = ~n461;
assign n10007 = n3862 | n10392;
assign n19603 = ~n4660;
assign n25904 = n21860 | n1513;
assign n7266 = n6442 | n8959;
assign n2551 = ~(n763 ^ n5222);
assign n16817 = n14465 | n23230;
assign n8805 = ~(n106 ^ n22516);
assign n10240 = ~(n21451 ^ n4893);
assign n1193 = n6054 | n16114;
assign n12210 = ~(n10113 | n11006);
assign n11367 = n9964 & n4880;
assign n3148 = ~(n14733 ^ n13453);
assign n25666 = n1363 & n13692;
assign n25180 = ~(n3349 ^ n25464);
assign n13307 = n6734 | n3;
assign n14050 = ~(n7149 ^ n16971);
assign n17242 = ~(n5160 ^ n5652);
assign n25351 = n18115 | n10837;
assign n14322 = n10557 | n8070;
assign n6900 = ~n20039;
assign n7028 = n8500 & n23716;
assign n23229 = ~(n12869 ^ n17277);
assign n9097 = n27185 | n4660;
assign n7665 = n11446 & n8831;
assign n5432 = ~(n16573 | n788);
assign n19127 = ~n7180;
assign n16090 = n11041 & n7112;
assign n13296 = ~(n12880 ^ n24684);
assign n19164 = ~(n18845 ^ n6021);
assign n14832 = ~(n6554 ^ n26205);
assign n4327 = n13590 | n1765;
assign n10396 = n23973 | n6738;
assign n22728 = n26642 | n3569;
assign n25020 = n2497 & n25695;
assign n5953 = n4760 | n24711;
assign n20039 = ~(n14219 ^ n12529);
assign n6290 = ~(n15519 ^ n5924);
assign n3398 = n17098 | n11510;
assign n23613 = ~(n11056 ^ n20250);
assign n21191 = ~(n23474 | n12333);
assign n21760 = ~(n4490 ^ n13167);
assign n948 = ~(n9641 ^ n11267);
assign n20705 = ~(n18839 ^ n22632);
assign n11480 = n24539 & n11709;
assign n3527 = n18851 & n5606;
assign n22908 = ~(n22139 ^ n19472);
assign n5001 = n17173 & n1906;
assign n7592 = ~(n22190 ^ n9243);
assign n17403 = ~(n8309 | n13158);
assign n20445 = ~(n26203 ^ n24681);
assign n14640 = n6872 & n16559;
assign n7897 = n4098 | n13323;
assign n20679 = n4218 | n26981;
assign n9531 = ~n13034;
assign n16875 = n15258 | n4588;
assign n4886 = ~(n19298 ^ n6611);
assign n11517 = n19939 & n26624;
assign n12118 = n18677 | n19416;
assign n7712 = ~(n10882 | n10760);
assign n13130 = n1796 | n21748;
assign n4765 = ~(n24460 ^ n23261);
assign n19631 = ~(n24364 | n21280);
assign n26458 = ~(n25622 | n11945);
assign n19423 = n11452 & n14689;
assign n5155 = ~(n11161 | n8281);
assign n15747 = n23039 & n12734;
assign n21163 = ~n25168;
assign n5754 = n1402 | n24675;
assign n4667 = ~n16502;
assign n4472 = n13314 & n15099;
assign n20715 = n8773 & n10610;
assign n15624 = ~(n17077 ^ n2289);
assign n4851 = ~(n26702 ^ n1172);
assign n20595 = ~(n11345 ^ n7045);
assign n21081 = ~(n13233 ^ n8944);
assign n6340 = n7084 & n15381;
assign n1981 = ~(n2765 ^ n15981);
assign n18154 = ~(n16697 ^ n20293);
assign n18047 = ~n11185;
assign n7317 = ~n22014;
assign n18727 = n2659 | n16619;
assign n5368 = n3062 & n18047;
assign n4347 = ~(n25872 | n20196);
assign n21838 = ~n7329;
assign n7302 = n4078 & n25281;
assign n22353 = ~(n4751 ^ n15406);
assign n11827 = ~(n19157 | n22379);
assign n15264 = n24610 | n8900;
assign n19781 = n13780 & n21949;
assign n11533 = ~n24609;
assign n22679 = ~(n11841 ^ n2479);
assign n9670 = ~(n1777 | n26724);
assign n8390 = n5712 | n16701;
assign n4145 = n22764 | n14448;
assign n3747 = n6395 | n1335;
assign n17073 = n6739 & n25488;
assign n11535 = ~n61;
assign n17782 = ~(n2268 | n11503);
assign n14931 = ~(n8901 ^ n14919);
assign n10150 = ~(n16366 ^ n3018);
assign n26798 = n1750 & n21321;
assign n21172 = n14979 & n14317;
assign n8454 = ~n2481;
assign n19713 = n16773 & n4219;
assign n716 = n4892 | n21466;
assign n3084 = n22312 & n3762;
assign n8790 = n7861 | n16401;
assign n22973 = ~(n19789 ^ n15424);
assign n22573 = n15809 | n4721;
assign n10803 = n18813 & n7219;
assign n16509 = ~(n23408 | n25643);
assign n7407 = ~(n12653 ^ n18965);
assign n9060 = ~(n21114 | n17814);
assign n14476 = n14149 | n2397;
assign n6291 = n21905 & n24481;
assign n12475 = ~n12920;
assign n12105 = ~n9731;
assign n21131 = ~(n19529 ^ n4049);
assign n23383 = ~(n20487 ^ n2968);
assign n7606 = ~(n8155 | n10763);
assign n21938 = n22479 & n18618;
assign n20221 = ~(n20235 ^ n6502);
assign n57 = ~(n5231 | n14048);
assign n20143 = n11891 | n18985;
assign n15550 = n2156 | n18931;
assign n26248 = ~(n18985 ^ n26931);
assign n1587 = ~n3785;
assign n7948 = ~n22043;
assign n21208 = ~n10899;
assign n20919 = ~(n7437 ^ n17077);
assign n4126 = n20801 | n6363;
assign n14123 = n20898 | n5110;
assign n16494 = n20658 | n6307;
assign n527 = ~(n13828 ^ n19905);
assign n2706 = ~(n18949 ^ n15725);
assign n11654 = n23487 & n18542;
assign n7595 = n4845 | n24624;
assign n16415 = n15041 & n13224;
assign n16276 = ~(n19067 ^ n17643);
assign n26105 = ~n9043;
assign n21053 = n20583 | n3298;
assign n10499 = ~n13333;
assign n3022 = ~(n856 | n11365);
assign n14956 = n3293 | n25189;
assign n24457 = ~(n7057 | n14570);
assign n16788 = ~(n15282 ^ n9859);
assign n12294 = n13106 | n21028;
assign n25063 = ~(n25066 ^ n8827);
assign n5963 = ~n14580;
assign n13726 = n10120 | n22629;
assign n11858 = n13712 & n6945;
assign n15324 = n10885 | n19276;
assign n9816 = n5255 | n25289;
assign n15325 = ~(n2436 ^ n11714);
assign n24407 = n1867 & n14308;
assign n9499 = ~(n7099 ^ n6691);
assign n1328 = n11634 & n3437;
assign n13504 = ~(n3840 ^ n24908);
assign n26668 = ~(n17141 ^ n494);
assign n4863 = n7974 | n24618;
assign n9086 = ~(n12050 ^ n19982);
assign n22543 = n12589 & n22979;
assign n11487 = n26312 | n13873;
assign n1966 = n6406 | n12100;
assign n13157 = ~(n14440 ^ n14130);
assign n12779 = n25890 | n25494;
assign n13836 = ~(n10951 ^ n13895);
assign n11275 = ~(n24719 ^ n26343);
assign n10284 = ~(n18724 ^ n6891);
assign n13539 = ~n7416;
assign n25658 = ~(n13459 | n15167);
assign n20563 = n342 & n26789;
assign n22920 = n4687 | n19245;
assign n13898 = ~n9399;
assign n1271 = n22459 | n9662;
assign n20838 = ~(n12341 ^ n15053);
assign n17975 = ~(n7112 ^ n20919);
assign n6683 = ~(n26499 ^ n25604);
assign n7757 = ~(n6173 | n12917);
assign n19576 = ~(n9557 ^ n16158);
assign n6412 = ~(n4469 ^ n25071);
assign n8569 = ~(n16377 ^ n4269);
assign n25816 = ~(n16538 ^ n4506);
assign n7005 = ~n24557;
assign n1377 = n18980 & n22096;
assign n16007 = n2342 & n12984;
assign n10161 = n4419 & n8291;
assign n7063 = n13563 | n26889;
assign n4764 = ~(n18286 ^ n1884);
assign n12884 = n10995 ^ n6397;
assign n25784 = ~(n17067 ^ n2946);
assign n6744 = ~(n6698 | n20556);
assign n17836 = ~(n10169 | n7133);
assign n24561 = ~(n10188 ^ n25738);
assign n13660 = ~(n6794 ^ n14090);
assign n35 = n24337 & n11954;
assign n12736 = n3988 & n8686;
assign n25985 = ~(n2475 ^ n1419);
assign n6568 = ~n1710;
assign n17409 = ~n12137;
assign n13119 = ~(n5741 ^ n15081);
assign n3031 = n120 | n21687;
assign n22493 = ~(n6731 ^ n5066);
assign n18996 = n17826 | n23878;
assign n8137 = n13786 | n10242;
assign n14675 = ~(n14400 ^ n6857);
assign n972 = ~(n18178 ^ n18840);
assign n27090 = n7300 & n6793;
assign n24135 = ~(n27081 ^ n1622);
assign n6620 = ~(n7871 ^ n5696);
assign n9790 = n15944 | n2783;
assign n15845 = ~n6719;
assign n24339 = n15651 | n3613;
assign n25571 = ~(n1835 | n2645);
assign n83 = ~(n3009 | n1288);
assign n15405 = ~n2868;
assign n20630 = ~n11941;
assign n13085 = n8518 | n231;
assign n26538 = ~(n3658 ^ n23325);
assign n21224 = ~n21291;
assign n25867 = ~(n8609 ^ n9584);
assign n6067 = ~(n746 | n27078);
assign n11805 = n12446 & n966;
assign n24508 = ~(n23876 ^ n14477);
assign n24891 = n20667 | n14151;
assign n19204 = ~(n56 ^ n17590);
assign n3494 = n11989 | n2981;
assign n7513 = n5364 | n22653;
assign n20318 = n17110 | n17502;
assign n21806 = n1848 | n5421;
assign n5980 = ~(n21920 ^ n6210);
assign n15458 = ~(n9504 ^ n26524);
assign n6756 = ~(n20210 ^ n19144);
assign n1600 = n23793 | n12004;
assign n6946 = ~n25947;
assign n18713 = n24126 | n18359;
assign n17626 = ~n13621;
assign n10442 = ~(n12423 ^ n9259);
assign n18123 = ~(n3128 ^ n4566);
assign n14973 = ~(n19446 ^ n3931);
assign n15408 = ~(n5858 ^ n10127);
assign n12950 = ~(n2333 ^ n5161);
assign n7087 = n4920 | n26664;
assign n3768 = n3654 | n23601;
assign n15544 = n23267 & n25005;
assign n11914 = n13186 | n11611;
assign n12440 = ~(n9251 ^ n2387);
assign n17092 = ~(n17184 | n18587);
assign n7482 = n24304 | n7425;
assign n16546 = n11731 | n16991;
assign n16539 = n3395 & n11939;
assign n21077 = n12963 & n6797;
assign n12548 = n17409 ^ n26000;
assign n21540 = ~(n1256 ^ n11281);
assign n19621 = n5140 | n14158;
assign n4099 = n1432 & n2852;
assign n9518 = n23000 | n24908;
assign n838 = n21593 | n7787;
assign n6999 = ~(n17647 ^ n20146);
assign n14815 = n20922 & n17950;
assign n4354 = n26129 | n22292;
assign n11856 = ~(n21969 | n5949);
assign n27198 = n913 | n6390;
assign n16206 = ~(n13191 ^ n12913);
assign n21009 = n19272 | n25541;
assign n16517 = ~(n17914 ^ n4596);
assign n26581 = n397 & n5177;
assign n18861 = ~n22511;
assign n26762 = n6551 & n5527;
assign n24673 = n17812 | n4675;
assign n4421 = n5575 | n13019;
assign n16813 = n14440 & n7523;
assign n6439 = n21174 | n4065;
assign n16938 = ~(n6658 ^ n1980);
assign n15148 = n7953 | n6397;
assign n22181 = n23178 & n3418;
assign n25444 = ~(n5547 | n3241);
assign n20481 = n14963 | n12379;
assign n25873 = ~(n5008 ^ n24433);
assign n11434 = n1176 | n26913;
assign n16334 = n17645 & n10945;
assign n7564 = n3681 | n18510;
assign n4676 = ~(n19163 | n13945);
assign n13098 = ~(n4212 ^ n15679);
assign n10079 = n21314 & n23051;
assign n15029 = n15935 | n22738;
assign n3252 = ~(n16183 | n5283);
assign n20936 = ~(n15811 ^ n1943);
assign n11594 = n19386 | n6561;
assign n24130 = ~n10514;
assign n1871 = n22558 | n5733;
assign n24229 = ~(n16524 | n13668);
assign n21341 = ~(n24969 | n13124);
assign n4540 = ~(n23688 ^ n12697);
assign n15284 = ~(n1756 ^ n4464);
assign n13147 = n18239 & n11541;
assign n19595 = n16812 | n21688;
assign n6506 = ~(n7239 ^ n4064);
assign n25463 = ~(n21222 | n26752);
assign n10700 = ~(n9244 | n6303);
assign n3440 = ~(n8356 ^ n5853);
assign n18183 = ~(n15810 ^ n17306);
assign n5542 = n20186 & n15844;
assign n18569 = ~(n25484 ^ n22586);
assign n18445 = ~(n16306 ^ n1857);
assign n14962 = n2336 | n6842;
assign n1606 = n103 & n16388;
assign n3079 = n11152 | n22880;
assign n20542 = ~n10403;
assign n18161 = n20020 | n448;
assign n11587 = ~(n7494 ^ n19483);
assign n14780 = n17030 & n20547;
assign n16427 = ~(n3375 ^ n8033);
assign n15136 = ~(n3603 | n455);
assign n23400 = ~n5648;
assign n10970 = ~(n8043 ^ n26699);
assign n18213 = ~(n24506 ^ n1681);
assign n3880 = ~(n5767 ^ n22440);
assign n25111 = n1474 & n3032;
assign n17131 = ~(n19674 ^ n5131);
assign n16456 = ~(n22820 ^ n8244);
assign n24544 = n25564 | n25390;
assign n11338 = ~(n20826 | n835);
assign n8949 = ~(n2559 | n26255);
assign n10910 = ~(n7351 ^ n6464);
assign n25894 = n24680 | n4931;
assign n5395 = n7597 | n17156;
assign n19587 = n21035 | n9696;
assign n14169 = n9439 | n24624;
assign n22303 = n16708 & n10518;
assign n4928 = n774 & n25145;
assign n17305 = ~(n23966 ^ n18770);
assign n7191 = n23312 & n18920;
assign n23574 = n12522 | n12674;
assign n22163 = n6565 | n12310;
assign n23479 = ~(n24890 | n19150);
assign n20448 = n22675 | n15810;
assign n2168 = ~n6911;
assign n21360 = n3009 | n24031;
assign n17018 = n9988 & n21667;
assign n1740 = n18598 | n20946;
assign n10444 = n17230 & n26747;
assign n7118 = ~(n3556 ^ n21434);
assign n7148 = n26224 | n8672;
assign n3935 = ~(n11486 ^ n20138);
assign n1646 = ~n12380;
assign n20003 = n3458 | n2001;
assign n13362 = n13730 & n18019;
assign n2238 = ~(n2925 ^ n5810);
assign n16322 = n201 | n15877;
assign n9444 = n1269 | n18416;
assign n18774 = n17846 & n12488;
assign n1101 = n1979 | n16245;
assign n21509 = ~(n8942 ^ n15516);
assign n19038 = n10379 & n13772;
assign n17925 = n11228 | n10821;
assign n19464 = ~n12767;
assign n12403 = n1216 | n26887;
assign n25257 = n10092 & n11477;
assign n7747 = ~(n8285 | n20036);
assign n7325 = ~n477;
assign n18924 = ~(n22587 ^ n16681);
assign n1514 = n1151 | n16111;
assign n13156 = ~n17108;
assign n232 = n26859 & n8590;
assign n6936 = ~(n1252 | n6204);
assign n23454 = ~(n17552 ^ n7337);
assign n11500 = n26188 | n10652;
assign n20237 = n26508 | n20945;
assign n4896 = ~n22455;
assign n26846 = n19052 & n16826;
assign n3096 = ~(n19616 | n18558);
assign n12162 = ~(n747 | n20164);
assign n10363 = n24089 | n1233;
assign n9482 = n15408 | n19158;
assign n5859 = n20291 | n27027;
assign n3739 = ~(n7853 ^ n22407);
assign n14253 = n26778 | n22520;
assign n225 = ~(n15519 | n5924);
assign n4113 = n18975 & n8411;
assign n19800 = n13741 | n3841;
assign n21602 = ~(n23304 ^ n17069);
assign n25207 = n5557 | n23013;
assign n3850 = ~(n6410 ^ n17651);
assign n5464 = n13591 | n24156;
assign n26704 = ~(n21974 | n20437);
assign n15737 = ~(n11898 ^ n23166);
assign n25725 = n15338 | n20280;
assign n17119 = ~(n397 ^ n26076);
assign n6801 = n12055 | n25855;
assign n14122 = n19243 & n9776;
assign n26138 = n16582 & n8945;
assign n18262 = ~n13112;
assign n9274 = ~(n11202 ^ n15304);
assign n2785 = ~(n1831 ^ n10250);
assign n16188 = n2724 | n9399;
assign n11215 = ~n2898;
assign n2240 = ~(n2908 ^ n17771);
assign n7857 = ~(n9825 ^ n133);
assign n6799 = ~(n23254 ^ n6204);
assign n5666 = n19682 & n7041;
assign n15521 = ~(n532 ^ n18272);
assign n20666 = ~(n2980 | n4781);
assign n26807 = ~n8518;
assign n24657 = n14510 | n8994;
assign n22100 = n22554 | n1414;
assign n18392 = n1424 | n6810;
assign n18539 = ~n13133;
assign n3667 = n25013 & n25965;
assign n14085 = ~n13538;
assign n6110 = n17447 | n22380;
assign n21752 = n20520 & n2859;
assign n3034 = ~n1947;
assign n7382 = ~(n21235 | n19241);
assign n9956 = ~(n11393 | n19875);
assign n15913 = n7593 & n17415;
assign n8708 = n3206 | n21931;
assign n19240 = n20698 & n3157;
assign n20611 = ~(n11308 ^ n26205);
assign n14714 = ~(n22660 | n26823);
assign n16834 = ~(n3250 ^ n22831);
assign n5459 = n24942 | n8789;
assign n4030 = n18290 | n26888;
assign n25477 = n13381 | n10063;
assign n1603 = ~(n22322 ^ n468);
assign n6488 = n23974 & n26085;
assign n2806 = n14328 & n5720;
assign n24689 = n9091 | n1607;
assign n26833 = ~(n17250 | n10125);
assign n9203 = n5484 | n18484;
assign n26152 = n8273 & n3292;
assign n19650 = ~(n27074 | n19391);
assign n25800 = ~(n17660 | n1704);
assign n7691 = ~n2612;
assign n3688 = n19002 | n18340;
assign n9614 = n1319 | n3769;
assign n26039 = n11816 & n24954;
assign n17332 = n2449 & n19470;
assign n16274 = ~(n18426 ^ n25168);
assign n15806 = n15167 & n20948;
assign n22389 = ~(n4718 | n16715);
assign n8412 = n23076 | n18950;
assign n6997 = n11732 | n13219;
assign n26673 = ~n24278;
assign n26193 = ~(n10676 ^ n5556);
assign n2525 = ~n7426;
assign n17375 = n3975 | n22303;
assign n3657 = n14409 | n7806;
assign n21627 = ~(n4466 ^ n15346);
assign n18904 = n2576 & n1325;
assign n10510 = n14571 & n26818;
assign n5118 = n16623 | n26060;
assign n13581 = ~(n25043 ^ n25612);
assign n25828 = n3811 | n17139;
assign n6424 = n26036 | n1505;
assign n3129 = n22585 | n8680;
assign n4202 = ~(n1466 ^ n7996);
assign n14243 = ~(n23089 ^ n12877);
assign n10310 = n26506 | n26248;
assign n1476 = n13598 & n3467;
assign n19386 = ~(n11003 ^ n22721);
assign n25874 = n9158 & n10223;
assign n18258 = ~n462;
assign n11632 = ~(n23591 ^ n24690);
assign n6741 = ~(n21839 ^ n19282);
assign n14247 = n21761 & n26083;
assign n14099 = ~(n5145 | n25486);
assign n19841 = ~n1986;
assign n22877 = ~(n11321 | n8933);
assign n6243 = ~(n20937 | n13435);
assign n2746 = ~(n23529 | n20700);
assign n3199 = ~(n17090 ^ n6773);
assign n18446 = ~(n701 ^ n23960);
assign n24554 = ~(n1220 ^ n13573);
assign n1675 = ~n4768;
assign n12630 = ~(n15073 ^ n15827);
assign n20091 = n21846 | n22861;
assign n2293 = n13978 & n21332;
assign n14155 = ~n15490;
assign n5198 = n1811 | n13994;
assign n27035 = n921 | n10590;
assign n15481 = ~(n5116 ^ n15617);
assign n13127 = n21485 | n6445;
assign n16295 = ~(n19606 ^ n13735);
assign n18683 = ~(n17430 ^ n23852);
assign n560 = ~(n16502 ^ n21654);
assign n4027 = n14860 | n7030;
assign n2281 = ~n8084;
assign n17372 = ~(n8773 ^ n11476);
assign n12389 = n24990 | n22321;
assign n24155 = ~(n21220 ^ n11987);
assign n74 = n729 | n25813;
assign n3681 = ~n25738;
assign n20753 = n21828 | n7177;
assign n9175 = ~(n1405 ^ n9067);
assign n12556 = ~(n21915 ^ n7674);
assign n18625 = ~(n3485 | n24070);
assign n19205 = ~(n6369 | n3164);
assign n1668 = n5809 | n25176;
assign n15211 = n10944 | n720;
assign n4844 = ~n24618;
assign n20506 = ~n4375;
assign n27008 = n11070;
assign n9671 = ~n23586;
assign n23830 = ~(n1181 | n5708);
assign n16420 = ~n21693;
assign n16612 = ~(n3587 ^ n15766);
assign n7819 = n16745 & n12828;
assign n8268 = ~n9506;
assign n17673 = n3345 | n10375;
assign n8284 = n7057 | n16729;
assign n23763 = ~(n23531 ^ n8036);
assign n11661 = n24437 | n21738;
assign n13254 = n17542 | n6185;
assign n2349 = ~(n19911 ^ n24278);
assign n18489 = ~(n12513 ^ n14106);
assign n6465 = ~(n12803 ^ n807);
assign n20847 = n3079 & n20143;
assign n8097 = ~n14600;
assign n25682 = ~(n2899 | n24731);
assign n27040 = n5831 | n3181;
assign n572 = n11011 & n1019;
assign n8328 = ~n16993;
assign n12770 = ~n15808;
assign n25499 = ~(n24871 ^ n7867);
assign n22411 = ~(n8675 | n26541);
assign n21215 = n10535 & n10172;
assign n24633 = n23102 | n11677;
assign n17169 = n22926 | n23866;
assign n3826 = n10402 & n22570;
assign n851 = ~(n368 ^ n19925);
assign n24188 = ~(n3003 ^ n17172);
assign n13006 = n16168 | n11757;
assign n24391 = n15613 & n8157;
assign n9675 = n17091 & n9711;
assign n6800 = ~(n20667 | n19616);
assign n11660 = n487 | n1919;
assign n25203 = ~(n12871 ^ n20411);
assign n22044 = n8904 | n25978;
assign n20033 = ~(n21445 ^ n10829);
assign n14771 = n11679 | n24509;
assign n12986 = ~(n6595 | n23681);
assign n18502 = ~(n24897 ^ n24040);
assign n2037 = n13709 | n3302;
assign n17512 = n22370 | n22332;
assign n2671 = n24403 | n8850;
assign n9652 = n4722 | n6403;
assign n14873 = n22919 | n8794;
assign n11597 = ~n26528;
assign n13569 = ~(n13319 ^ n25435);
assign n22319 = ~(n19057 | n26292);
assign n1931 = n20081 & n20846;
assign n12989 = n328 | n22173;
assign n8563 = ~(n1494 ^ n13235);
assign n25160 = ~n3220;
assign n20284 = ~n6444;
assign n18303 = n16937 & n5488;
assign n22425 = ~n17954;
assign n3052 = ~(n25330 | n13518);
assign n6715 = n24992 | n22139;
assign n17391 = n3958 & n18354;
assign n23879 = ~(n6561 ^ n19386);
assign n7945 = n10459 | n13243;
assign n2952 = ~(n20138 ^ n9251);
assign n4916 = n4900 | n10215;
assign n19897 = n6435 | n9245;
assign n14671 = ~n1065;
assign n12643 = n1164 | n4388;
assign n20714 = ~(n17536 ^ n11201);
assign n18033 = n3096 | n17775;
assign n1187 = n6404 & n23349;
assign n6905 = n17580 & n11008;
assign n17140 = ~(n9770 ^ n25054);
assign n6033 = n8307 & n18616;
assign n19839 = n14341 & n10398;
assign n23555 = ~n25877;
assign n25044 = ~(n17077 ^ n4256);
assign n16179 = ~(n8013 | n27147);
assign n17862 = ~(n3338 ^ n20647);
assign n8641 = n7102 & n280;
assign n26770 = ~(n21687 | n6606);
assign n711 = n639 & n16132;
assign n8780 = n19527 | n7808;
assign n24124 = n23768 | n8353;
assign n17348 = n6104 & n19985;
assign n17126 = n16679 | n7341;
assign n9779 = ~n26224;
assign n15883 = ~(n8864 ^ n6334);
assign n25204 = ~(n25573 ^ n18592);
assign n25459 = n12002 | n11382;
assign n19740 = ~(n1562 ^ n2422);
assign n21622 = ~(n9611 ^ n24834);
assign n12967 = ~(n199 ^ n8587);
assign n21946 = n15030 & n17231;
assign n2195 = n570 | n19701;
assign n14984 = ~(n22469 ^ n12358);
assign n16123 = n11856 | n2070;
assign n458 = n26810 | n12797;
assign n16903 = ~n21378;
assign n12028 = n21063 | n7164;
assign n6727 = ~(n2165 ^ n664);
assign n5795 = ~(n1296 ^ n16758);
assign n3192 = n24974 | n7460;
assign n1478 = n20565 & n14644;
assign n18837 = ~(n18921 | n17926);
assign n23942 = ~(n16578 ^ n3897);
assign n15878 = n6916 | n7160;
assign n6019 = ~(n21793 ^ n3352);
assign n13638 = ~(n13443 | n6580);
assign n5246 = ~(n19446 ^ n11980);
assign n20976 = ~n14484;
assign n25899 = n5309 & n15523;
assign n11335 = ~(n4980 ^ n6436);
assign n17459 = n14528 | n3552;
assign n21110 = n5838 | n13399;
assign n9561 = ~n15242;
assign n24771 = n14728 | n8570;
assign n6995 = ~(n19711 | n11697);
assign n20195 = n24389 | n3650;
assign n18725 = ~(n20386 ^ n13001);
assign n1028 = ~(n14908 ^ n23405);
assign n12101 = n24149 & n9933;
assign n19846 = n2487 | n15834;
assign n21338 = n991 & n1659;
assign n5157 = ~(n11410 | n18706);
assign n1532 = ~n1484;
assign n6364 = ~(n6814 ^ n23463);
assign n5909 = n12988 | n24854;
assign n20026 = n796 | n24197;
assign n24134 = ~n15277;
assign n25706 = ~(n6415 ^ n23060);
assign n10334 = ~(n1467 | n18113);
assign n22540 = ~(n8964 | n18539);
assign n21086 = n2469 | n21946;
assign n12673 = ~n5768;
assign n24954 = n16561 & n23596;
assign n6509 = ~(n11901 | n27089);
assign n17480 = n2178 | n16329;
assign n899 = n2332 | n19532;
assign n14549 = n2516 & n25638;
assign n25989 = ~n11693;
assign n22225 = ~(n4534 ^ n13522);
assign n16312 = n7026 | n21165;
assign n24402 = ~n18326;
assign n19683 = ~(n10281 ^ n24638);
assign n27098 = ~(n11481 ^ n23493);
assign n16970 = n21512 | n23988;
assign n11016 = n4534 | n13522;
assign n1546 = n8709 | n17787;
assign n16406 = ~(n462 ^ n23495);
assign n2148 = ~(n1403 ^ n12898);
assign n13241 = n4683 | n23926;
assign n7038 = ~(n11925 ^ n25964);
assign n11995 = n18451 ^ n12278;
assign n18092 = ~(n20425 ^ n15170);
assign n22064 = ~(n21073 ^ n3472);
assign n7960 = n18869 | n22548;
assign n5683 = ~n24452;
assign n13990 = ~n10133;
assign n4656 = ~(n16722 ^ n8381);
assign n25225 = ~(n17360 ^ n19680);
assign n14051 = ~(n2146 | n19144);
assign n4331 = ~(n11533 ^ n11095);
assign n4084 = n2174 | n11455;
assign n9125 = ~n24121;
assign n23395 = n12220 & n14553;
assign n3854 = n6806 & n18722;
assign n19225 = ~(n24728 ^ n24161);
assign n19329 = n5437 | n3205;
assign n22725 = n12644 & n18314;
assign n17718 = ~n22480;
assign n7486 = ~(n1408 ^ n23643);
assign n9026 = ~n19378;
assign n3712 = n6936 | n19182;
assign n5636 = ~(n23923 ^ n16608);
assign n107 = ~(n11670 ^ n7281);
assign n25183 = n5185 | n18444;
assign n11100 = ~n9646;
assign n3180 = n4834 & n23823;
assign n23919 = n26687 & n25830;
assign n21035 = ~(n14680 | n20359);
assign n24981 = n11193 | n9135;
assign n8676 = n11270 & n11976;
assign n8645 = n20089 & n21216;
assign n23481 = ~(n8302 ^ n16840);
assign n21071 = ~n16582;
assign n4724 = n26257 & n9205;
assign n8069 = n10112 | n21849;
assign n13966 = n10138 | n10105;
assign n17553 = n8161 ^ n4232;
assign n12949 = n2685 & n26426;
assign n15662 = ~(n13609 ^ n5597);
assign n15601 = ~(n22101 | n17553);
assign n10094 = ~(n9770 ^ n24612);
assign n22156 = ~(n17982 ^ n8028);
assign n14922 = n3909 | n17045;
assign n15380 = ~n10642;
assign n4061 = ~n3018;
assign n12077 = n3664 | n21830;
assign n20749 = ~n12658;
assign n25670 = ~(n744 ^ n13714);
assign n15547 = ~(n15834 ^ n22433);
assign n11279 = n1151 | n20536;
assign n5273 = ~(n7789 ^ n8871);
assign n23159 = ~(n5440 | n11503);
assign n6671 = ~(n10724 ^ n24965);
assign n20862 = ~n17640;
assign n14949 = ~(n4652 ^ n1573);
assign n15699 = n14153 | n21894;
assign n16727 = ~n21850;
assign n22963 = n987 & n11871;
assign n12789 = ~n18690;
assign n13470 = n25295 & n25774;
assign n6114 = n4339 | n6286;
assign n8892 = n8917 & n24753;
assign n2702 = n4733 | n7497;
assign n26976 = n11877 | n21824;
assign n21903 = n15886 & n5459;
assign n16568 = n21822 & n2462;
assign n4942 = ~(n7134 | n9830);
assign n5995 = n8218 | n3854;
assign n20932 = ~(n14899 ^ n7026);
assign n4110 = n10659 | n23586;
assign n25869 = ~(n17028 ^ n18444);
assign n4647 = ~(n10760 ^ n801);
assign n17368 = ~n1279;
assign n22246 = n6282 & n15387;
assign n21033 = n7286 | n12030;
assign n4291 = n9294 | n4319;
assign n5390 = n4159 | n14776;
assign n10943 = ~(n17882 ^ n10456);
assign n12801 = ~(n24380 ^ n17476);
assign n26592 = ~(n23581 | n4572);
assign n9389 = n10768 | n17821;
assign n7010 = ~(n14911 ^ n20494);
assign n24522 = n15905 | n14996;
assign n5840 = ~(n1210 ^ n21579);
assign n17244 = ~(n19608 ^ n4426);
assign n17396 = n1845 | n7169;
assign n11334 = n15902 | n23605;
assign n20361 = ~(n6680 ^ n7667);
assign n6353 = n18141 & n8870;
assign n6210 = ~(n21740 ^ n12547);
assign n15607 = ~(n11533 ^ n4100);
assign n22919 = ~n1681;
assign n21030 = ~(n26414 ^ n3506);
assign n26758 = ~n13369;
assign n17833 = ~(n9125 ^ n22472);
assign n239 = n19829 & n18441;
assign n10035 = ~(n14040 ^ n8477);
assign n24734 = ~n5944;
assign n16181 = n14962 & n26308;
assign n9748 = ~(n4817 ^ n25605);
assign n21260 = ~n22472;
assign n21461 = n24299 | n630;
assign n19852 = ~n23657;
assign n14697 = n7522 & n18824;
assign n287 = n4460 & n25217;
assign n17377 = n3545 | n25889;
assign n15257 = ~n13318;
assign n10744 = n8455 & n24835;
assign n19964 = n2287 | n26176;
assign n22106 = ~(n25565 ^ n24374);
assign n13246 = n1463 & n17053;
assign n20023 = ~(n2539 ^ n1279);
assign n14535 = n7294 & n8171;
assign n15354 = n12996 | n19196;
assign n18462 = ~(n14440 ^ n17911);
assign n453 = n13653 | n25051;
assign n15017 = ~n20633;
assign n17310 = ~n281;
assign n3792 = ~(n7841 ^ n9445);
assign n9462 = ~n7473;
assign n17816 = ~n790;
assign n5083 = n6096 | n278;
assign n5113 = ~n3097;
assign n6454 = n10025 | n24456;
assign n22527 = ~n22173;
assign n24839 = ~n5178;
assign n23528 = ~n8721;
assign n20308 = ~(n11764 ^ n26946);
assign n8402 = n1583 ^ n1648;
assign n23624 = ~(n7016 ^ n7729);
assign n14872 = ~(n12052 ^ n19590);
assign n9454 = ~(n20138 ^ n19494);
assign n23362 = n12513 & n8395;
assign n2850 = ~(n27064 ^ n25850);
assign n8407 = n25108 & n7064;
assign n10933 = n13695 | n26056;
assign n22141 = n23004 | n14913;
assign n18068 = ~(n6377 ^ n987);
assign n20232 = n8071 | n26851;
assign n18159 = n136 & n15982;
assign n19535 = ~(n10167 | n24104);
assign n7329 = n9979 | n1227;
assign n18026 = n18705 | n8083;
assign n8589 = ~(n7375 ^ n5454);
assign n18472 = n12732 & n15250;
assign n11647 = ~(n22543 ^ n4540);
assign n20820 = n9289 & n17309;
assign n2565 = ~(n13930 ^ n6105);
assign n26661 = ~n24732;
assign n1736 = n13278 | n23372;
assign n12513 = n24249 & n3058;
assign n17078 = ~(n15490 ^ n7339);
assign n6332 = n26892 | n11623;
assign n25144 = ~(n3952 ^ n12315);
assign n14079 = n9964 | n5067;
assign n18849 = n25324 & n5951;
assign n12893 = ~(n10763 | n5696);
assign n17865 = ~(n6726 ^ n22934);
assign n19023 = n26661 | n19371;
assign n5825 = ~(n9180 | n8006);
assign n1242 = ~(n23692 | n15236);
assign n280 = ~(n2855 ^ n2002);
assign n10804 = ~n7284;
assign n17297 = n21641 & n7383;
assign n25389 = ~n12562;
assign n4638 = n17162 | n868;
assign n15485 = n5371 | n22539;
assign n5561 = ~(n13328 ^ n16439);
assign n8183 = n4210 | n17628;
assign n11379 = ~(n24584 ^ n6873);
assign n7347 = ~n8858;
assign n7508 = n2098 | n606;
assign n12682 = ~(n3540 | n10885);
assign n22781 = ~(n8520 | n18338);
assign n8606 = ~(n11201 | n14366);
assign n18726 = ~(n11575 ^ n16703);
assign n25901 = n25163 & n9354;
assign n12447 = ~(n18947 | n10331);
assign n4333 = ~(n21638 ^ n7567);
assign n24564 = n3827 | n5055;
assign n18228 = ~(n16261 | n24188);
assign n16043 = n2348 | n25064;
assign n18470 = n23527 | n18275;
assign n900 = n1866 | n17656;
assign n16654 = ~(n13441 ^ n13094);
assign n14251 = ~n2429;
assign n22366 = ~(n7319 | n17458);
assign n6400 = ~n21138;
assign n23251 = ~(n25119 ^ n21934);
assign n13185 = n13674 | n14316;
assign n16799 = n8146 & n5285;
assign n26495 = ~n2829;
assign n26027 = n12811 & n11822;
assign n4773 = n14831 & n21415;
assign n6802 = ~(n7140 ^ n26934);
assign n20243 = ~(n387 | n9300);
assign n6797 = n26607 | n13840;
assign n8401 = ~(n12436 ^ n24937);
assign n13225 = n18058 | n3828;
assign n2641 = n18527 | n1991;
assign n16331 = ~n1320;
assign n849 = ~(n2221 ^ n26917);
assign n19735 = n13430 & n1056;
assign n24534 = n8134 | n27005;
assign n22846 = n10195 & n14889;
assign n16591 = ~(n19474 | n151);
assign n1814 = n6686 | n2163;
assign n4051 = ~(n25068 ^ n6790);
assign n11288 = n4586 | n3381;
assign n18244 = n21841 | n14110;
assign n14357 = n20167 & n19826;
assign n15439 = ~(n19110 | n5467);
assign n26690 = n4398 | n12694;
assign n3652 = ~(n2424 | n84);
assign n17835 = ~n31;
assign n22466 = n20918 | n7874;
assign n6825 = n13731 | n6195;
assign n5078 = n2762 & n17868;
assign n5585 = ~n837;
assign n8835 = ~n1878;
assign n17519 = ~(n20671 ^ n26963);
assign n26401 = n19260 | n8830;
assign n777 = ~(n5498 | n12928);
assign n172 = ~n6988;
assign n20552 = ~n22918;
assign n22828 = ~(n23186 ^ n24047);
assign n20215 = ~(n6389 ^ n14350);
assign n15773 = ~n18569;
assign n2874 = n10710 | n26510;
assign n1707 = n23922 & n2843;
assign n13017 = ~(n19094 | n1197);
assign n12464 = ~n26823;
assign n1856 = n15329 | n7528;
assign n12888 = ~n25017;
assign n12590 = n19568 | n162;
assign n5048 = ~(n7383 ^ n19576);
assign n22566 = ~(n12573 | n19312);
assign n23534 = ~(n18035 ^ n3279);
assign n27142 = ~n6230;
assign n18230 = n3874 & n1485;
assign n20094 = ~n21567;
assign n18803 = n2812 | n18812;
assign n16128 = ~(n658 | n27120);
assign n25615 = ~(n6744 | n18568);
assign n14883 = ~(n16856 ^ n21081);
assign n26219 = ~(n22378 ^ n5026);
assign n17015 = ~n23765;
assign n24335 = ~(n24511 ^ n10096);
assign n19400 = n5303 & n7508;
assign n4935 = ~(n23832 ^ n3161);
assign n12312 = n11270 | n11976;
assign n4861 = ~(n1426 ^ n12419);
assign n166 = ~n19080;
assign n8196 = ~(n2979 | n9554);
assign n6044 = ~(n1564 ^ n2050);
assign n6550 = ~(n12422 ^ n1780);
assign n27097 = n3021 | n16308;
assign n26174 = ~(n24668 ^ n23671);
assign n1885 = ~(n15090 ^ n12209);
assign n4693 = ~(n4907 ^ n1012);
assign n6914 = ~(n10405 ^ n25370);
assign n6662 = ~(n22153 ^ n3984);
assign n19397 = n13058 | n7749;
assign n24492 = n7195 | n12861;
assign n7683 = ~(n9498 | n12494);
assign n10331 = ~n21444;
assign n4700 = n21730 & n18464;
assign n25181 = ~(n12450 ^ n5876);
assign n24334 = n24885 & n20381;
assign n8129 = n19444 | n20689;
assign n5923 = ~n10735;
assign n18929 = ~(n12475 | n18263);
assign n20959 = ~(n1365 ^ n10158);
assign n24064 = n23703 & n2344;
assign n11270 = n8436 & n4886;
assign n2711 = ~(n2375 ^ n6453);
assign n7856 = n14307 & n6629;
assign n23275 = n17486 & n25662;
assign n22030 = ~(n12112 | n20444);
assign n3168 = n5137 & n9762;
assign n798 = n25090 & n3182;
assign n7431 = n27006 & n7197;
assign n26938 = n14559 | n4290;
assign n9388 = ~(n18398 ^ n1605);
assign n10528 = n9857 | n27148;
assign n24436 = n21153 & n11907;
assign n17667 = ~(n13490 ^ n7751);
assign n598 = ~n25360;
assign n12449 = ~(n11969 ^ n25279);
assign n13750 = n7191 | n25697;
assign n1256 = n16049 | n18199;
assign n7615 = ~n20183;
assign n26856 = ~(n12861 ^ n1255);
assign n13661 = n25354 & n16936;
assign n15552 = n36 & n23127;
assign n15314 = ~(n14774 ^ n23200);
assign n6011 = ~n3274;
assign n15192 = ~(n8230 | n10454);
assign n17134 = n6880 & n775;
assign n15631 = n329 & n6541;
assign n13527 = n23852 & n17430;
assign n16442 = n3043 | n3861;
assign n3900 = n15734 & n18664;
assign n19762 = ~(n556 ^ n26348);
assign n6009 = n19804 | n14311;
assign n194 = n14775 & n14925;
assign n4301 = ~(n8739 | n23655);
assign n20300 = ~(n15942 | n17499);
assign n8406 = ~(n27128 ^ n12275);
assign n21963 = ~(n7330 ^ n2479);
assign n14340 = n25722 & n16004;
assign n11325 = ~(n8341 ^ n4443);
assign n2481 = ~(n5130 ^ n24419);
assign n13903 = ~(n23459 | n10603);
assign n11512 = ~(n26875 ^ n5530);
assign n17860 = n12143 | n20215;
assign n10907 = n5501 | n23824;
assign n9884 = n2453 | n26318;
assign n14188 = n22167 | n11373;
assign n25238 = ~n13774;
assign n26552 = ~(n16653 ^ n16558);
assign n8242 = ~(n7439 ^ n15182);
assign n9868 = n12822 | n10231;
assign n3073 = n12368 | n14670;
assign n62 = n14542 | n23147;
assign n16438 = n19097 | n5333;
assign n21210 = ~(n2085 ^ n21361);
assign n5082 = ~(n25807 ^ n9388);
assign n9335 = ~n19544;
assign n20684 = ~(n337 | n17902);
assign n12281 = ~(n25056 ^ n23192);
assign n11193 = ~n9940;
assign n993 = n16152 | n1377;
assign n1530 = n22072 & n7529;
assign n11727 = n18218 | n7430;
assign n26398 = n4119 | n24746;
assign n21668 = ~n9575;
assign n9310 = ~n1525;
assign n15985 = ~(n5124 ^ n14675);
assign n15384 = n752 | n4105;
assign n20144 = ~(n10191 ^ n23279);
assign n26242 = n1179 | n6579;
assign n13121 = n15347 & n1774;
assign n10892 = n22236 & n3399;
assign n22420 = ~(n494 | n17141);
assign n6001 = ~(n20777 ^ n13848);
assign n3155 = ~(n9586 | n24196);
assign n22757 = n1771 | n17033;
assign n2423 = ~n161;
assign n18835 = n5206 | n2937;
assign n12484 = ~(n16091 ^ n16602);
assign n22496 = ~(n17536 ^ n19060);
assign n26835 = ~(n24473 ^ n19472);
assign n426 = n4514 & n21162;
assign n10297 = n1870 | n18701;
assign n21497 = ~(n12379 ^ n1434);
assign n1323 = n2414 & n5754;
assign n10699 = ~(n4724 ^ n6418);
assign n20142 = ~(n18639 | n20771);
assign n2012 = n3018 | n16366;
assign n11310 = n786 | n24281;
assign n16026 = ~(n7619 ^ n16446);
assign n6575 = ~(n18754 ^ n5211);
assign n16333 = ~n1601;
assign n9160 = ~(n19507 ^ n17798);
assign n25760 = n3403 & n3271;
assign n26023 = ~n8164;
assign n7387 = ~(n14741 ^ n25454);
assign n6120 = ~(n1525 | n11018);
assign n10957 = n7523 | n8385;
assign n18205 = ~n10963;
assign n21864 = n5174 & n24336;
assign n10153 = n15290 & n25734;
assign n23945 = n23144 | n10306;
assign n8151 = n4939 & n120;
assign n26999 = ~n5206;
assign n12907 = ~(n24493 ^ n22198);
assign n686 = n9905 & n20174;
assign n8586 = n22964 | n19924;
assign n11672 = n12017 & n8169;
assign n16393 = ~(n10523 ^ n25203);
assign n7141 = ~(n1896 | n27104);
assign n2496 = n15911 | n26939;
assign n11593 = ~(n11840 ^ n15423);
assign n6075 = n26450 | n22958;
assign n5928 = n6268 | n1218;
assign n16702 = n7322 & n15689;
assign n16754 = n19432 | n11337;
assign n2865 = n13274 | n8524;
assign n18177 = ~(n2035 ^ n26054);
assign n16752 = ~(n26974 ^ n10305);
assign n19855 = n19018 | n20910;
assign n15263 = n20303 | n14598;
assign n24438 = n4539 | n368;
assign n23698 = ~(n4963 ^ n24796);
assign n19942 = n15989 | n7665;
assign n22881 = ~(n6122 ^ n678);
assign n1302 = ~(n10891 ^ n10367);
assign n22959 = ~(n16163 | n15932);
assign n25752 = ~(n24902 | n25572);
assign n17289 = n4164 & n9865;
assign n22852 = ~(n9615 ^ n21055);
assign n17210 = ~n563;
assign n19180 = n27088 & n10031;
assign n22965 = n23490 | n15048;
assign n10132 = n751 | n14788;
assign n21546 = n22534 | n12577;
assign n22893 = n3769 | n4485;
assign n5732 = ~(n8346 ^ n6344);
assign n6142 = ~(n24480 ^ n14634);
assign n20121 = n11246 & n14974;
assign n18391 = n13709 | n15696;
assign n26766 = ~(n1398 | n20548);
assign n10878 = ~(n8679 ^ n14516);
assign n3597 = n25470 | n3307;
assign n9632 = n3849 & n10750;
assign n10207 = ~n16197;
assign n20514 = n15326 | n21875;
assign n7462 = ~(n18537 | n4376);
assign n5506 = ~n5288;
assign n1798 = ~n23337;
assign n3648 = ~(n22795 | n2100);
assign n25633 = n25428 | n22412;
assign n19370 = n10290 & n3824;
assign n20511 = n14415 | n8032;
assign n10644 = ~(n3967 ^ n27054);
assign n8438 = n14764 & n13836;
assign n1608 = n4344 & n13849;
assign n18736 = ~(n14795 ^ n14189);
assign n24709 = ~(n19454 | n15042);
assign n26042 = ~(n1192 | n5743);
assign n22977 = ~n21;
assign n26784 = ~(n12944 ^ n6864);
assign n20269 = ~(n18444 ^ n13719);
assign n15738 = n26299 & n25208;
assign n9613 = n3648 | n5405;
assign n1285 = n667 & n15372;
assign n8821 = ~(n25583 ^ n15286);
assign n3979 = ~(n2783 ^ n1667);
assign n17156 = ~n24009;
assign n7476 = ~(n16330 ^ n14597);
assign n18286 = n27080 & n24515;
assign n1985 = n12024 | n18622;
assign n10082 = n23945 & n21411;
assign n22589 = ~(n14829 | n21889);
assign n22349 = ~n3143;
assign n9976 = n4733 & n7497;
assign n12165 = n16869 & n14908;
assign n1317 = n23873 | n21726;
assign n10395 = n25038 | n12639;
assign n14066 = n13795 & n17404;
assign n2566 = ~n24072;
assign n9836 = n15766 | n3587;
assign n22179 = ~(n21226 | n2906);
assign n25019 = n7166 & n9271;
assign n8383 = ~(n21134 ^ n11356);
assign n7638 = ~(n7170 ^ n24606);
assign n13160 = n22942 | n712;
assign n3492 = ~(n17369 ^ n26512);
assign n11905 = ~(n3913 ^ n8140);
assign n26732 = n23089 | n9830;
assign n24031 = ~n7674;
assign n22467 = ~(n3631 ^ n14493);
assign n14918 = n25434 | n22086;
assign n1446 = ~(n9542 ^ n12773);
assign n5217 = n15493 & n21345;
assign n4493 = n25923 & n24184;
assign n25326 = ~(n21134 | n11356);
assign n12344 = n14813 & n16863;
assign n13942 = n7012 | n24830;
assign n6747 = ~(n10486 ^ n19584);
assign n1554 = ~n23523;
assign n13387 = ~(n20957 ^ n21897);
assign n15219 = n12284 & n363;
assign n17084 = ~(n9304 ^ n6345);
assign n26662 = n5783 & n11432;
assign n14012 = n22743 | n2346;
assign n26022 = ~n14031;
assign n13934 = ~(n3770 ^ n24801);
assign n27176 = n26211 | n15333;
assign n19405 = n8285 | n14480;
assign n794 = ~(n11235 ^ n10352);
assign n25723 = n21805 & n13937;
assign n21402 = ~(n19005 ^ n19144);
assign n20918 = ~(n10629 | n6660);
assign n2206 = n1948 & n16250;
assign n24379 = ~n15141;
assign n26041 = n15625 | n2049;
assign n18431 = ~n17663;
assign n14336 = ~n22433;
assign n2515 = ~(n5027 ^ n21335);
assign n2782 = ~n4520;
assign n12260 = n24903 | n26466;
assign n19611 = ~(n19594 | n6235);
assign n11464 = n16784 | n15500;
assign n26894 = ~n20171;
assign n250 = n27062 | n12805;
assign n21465 = ~n18809;
assign n2003 = ~n13291;
assign n9468 = ~(n22875 ^ n5813);
assign n21180 = ~(n23264 ^ n27120);
assign n4500 = ~(n4031 | n24560);
assign n9599 = ~n22780;
assign n17062 = ~n25483;
assign n6436 = ~(n8241 ^ n11566);
assign n22136 = ~(n9748 ^ n6915);
assign n9874 = n11464 & n16425;
assign n24915 = n8999 | n1122;
assign n1859 = ~(n14112 ^ n22639);
assign n5772 = ~(n15294 | n15270);
assign n23654 = n6651 & n12037;
assign n4390 = n8186 | n3425;
assign n6567 = ~(n22551 ^ n6020);
assign n9305 = n22860 & n21494;
assign n19384 = n7237 & n2813;
assign n12948 = n26309 | n11726;
assign n3985 = ~n1610;
assign n17678 = ~(n14048 | n4467);
assign n23011 = n16302 | n2489;
assign n24151 = ~(n26249 ^ n4129);
assign n22633 = ~(n21849 ^ n5954);
assign n7307 = n6411 | n5649;
assign n75 = ~(n10702 ^ n12776);
assign n14211 = ~(n6188 ^ n17117);
assign n11048 = ~(n25560 ^ n13914);
assign n10467 = ~(n7673 ^ n3176);
assign n14196 = ~(n19797 ^ n4559);
assign n10670 = n1405 | n27181;
assign n1084 = n15426 & n22521;
assign n20607 = ~(n16874 ^ n530);
assign n11534 = n5025 & n12771;
assign n25795 = ~n11008;
assign n17257 = n26844 & n18964;
assign n1216 = n23150 & n2183;
assign n6640 = ~(n2809 ^ n15508);
assign n16204 = ~n12885;
assign n23201 = n17871 & n15067;
assign n20893 = n6750 | n13328;
assign n26967 = n26627 & n6577;
assign n2413 = n23901 & n16038;
assign n8075 = n14939 | n25449;
assign n7024 = n3192 & n15388;
assign n24723 = ~(n21553 ^ n7660);
assign n16982 = ~n6003;
assign n10291 = n24263 & n3608;
assign n15123 = n14198 | n12902;
assign n10195 = n10018 | n513;
assign n5693 = n4998 & n4888;
assign n26392 = n17540 & n14987;
assign n10657 = n25355 | n5110;
assign n25570 = ~(n9211 | n24394);
assign n25482 = n2227 & n24079;
assign n16031 = n21474 | n19865;
assign n219 = n1447 | n22482;
assign n2933 = n5696 | n23463;
assign n16551 = ~n7609;
assign n19807 = n13203 & n2430;
assign n5790 = ~n24609;
assign n16590 = ~n21509;
assign n21352 = ~(n12428 ^ n18215);
assign n3687 = ~n18674;
assign n22462 = ~(n1587 | n22977);
assign n4637 = n20467 | n13615;
assign n18314 = n11090 & n26267;
assign n24601 = ~n3829;
assign n12150 = n9906 | n22349;
assign n4781 = ~n26403;
assign n19600 = n19195 | n177;
assign n11177 = ~n1288;
assign n14062 = n25022 | n7441;
assign n23399 = ~(n25318 ^ n3955);
assign n6355 = ~(n19839 | n6518);
assign n3202 = ~(n2145 ^ n5521);
assign n20161 = ~(n6032 ^ n13623);
assign n20532 = ~(n149 ^ n15243);
assign n13624 = n9850 | n1162;
assign n1496 = n14523 | n19419;
assign n23571 = n23367 & n1856;
assign n19212 = n2084 | n17135;
assign n20564 = ~(n1801 ^ n18906);
assign n15615 = n22373 & n5009;
assign n15429 = n15894 | n10560;
assign n6560 = ~(n7385 ^ n11493);
assign n18979 = n6962 | n5119;
assign n10619 = ~(n15204 | n14122);
assign n6416 = ~(n2939 | n6366);
assign n23858 = n25888 | n19149;
assign n1077 = n22197 & n5927;
assign n21507 = n17173 | n21644;
assign n24719 = n8923 & n26175;
assign n8248 = n15454 | n2171;
assign n24625 = ~n252;
assign n18602 = n10763 | n18799;
assign n7065 = ~(n7099 | n6691);
assign n17999 = n218 | n25327;
assign n7985 = n5375 & n18267;
assign n4877 = ~(n11198 ^ n4391);
assign n8637 = ~(n3866 ^ n7491);
assign n13033 = ~n18901;
assign n16363 = n17676 | n25404;
assign n16811 = ~(n17846 ^ n12488);
assign n3439 = ~(n21380 | n11592);
assign n11028 = ~n17652;
assign n10261 = ~(n25145 ^ n14423);
assign n18594 = n23234 & n1688;
assign n26214 = n14920 | n8591;
assign n729 = ~n15339;
assign n14484 = ~(n23493 ^ n8405);
assign n7107 = ~n4448;
assign n26729 = ~(n9984 ^ n25526);
assign n19283 = ~(n2979 ^ n11898);
assign n24872 = ~(n23352 ^ n25659);
assign n15040 = n6702 | n14893;
assign n6056 = n6368 & n8879;
assign n6058 = n21438 & n2291;
assign n26550 = n20777 & n2461;
assign n23625 = n21828 & n7177;
assign n17971 = ~(n14411 ^ n16983);
assign n14160 = n5438 & n9964;
assign n825 = ~(n24908 ^ n23000);
assign n24106 = ~(n44 ^ n26290);
assign n26128 = ~(n3097 ^ n3764);
assign n17308 = n23804 | n21422;
assign n1553 = n24440;
assign n16269 = n5582 | n24842;
assign n20492 = n1372 & n16414;
assign n26961 = ~n5128;
assign n12615 = ~(n13367 ^ n13074);
assign n6198 = n6946 | n11136;
assign n16412 = n4802 & n25725;
assign n9591 = ~(n11603 ^ n16399);
assign n2025 = n19346 & n1985;
assign n26119 = ~(n15264 ^ n19720);
assign n24288 = n10700 | n23468;
assign n20875 = ~(n6704 | n21878);
assign n20290 = ~(n6832 ^ n11898);
assign n15972 = ~(n20627 ^ n12036);
assign n25883 = ~(n4858 ^ n26752);
assign n783 = ~(n12622 ^ n26289);
assign n21972 = ~n13783;
assign n11110 = ~n6224;
assign n1836 = n9712 | n9214;
assign n18515 = ~(n24507 ^ n12809);
assign n14659 = n27116 & n10170;
assign n18260 = ~(n8827 ^ n4306);
assign n3469 = n20472 | n2181;
assign n5 = ~n5625;
assign n12459 = ~(n10131 | n8507);
assign n24990 = ~(n14376 ^ n9608);
assign n15755 = ~n11823;
assign n12342 = ~(n23395 ^ n8950);
assign n8885 = n1403 | n16176;
assign n8310 = n20290 & n21577;
assign n15062 = ~(n9367 ^ n12353);
assign n11296 = ~(n456 ^ n24479);
assign n13097 = n7141 | n7654;
assign n24866 = ~(n11229 | n17195);
assign n17683 = n18604 & n4912;
assign n11771 = ~(n938 ^ n4524);
assign n18196 = ~n4068;
assign n889 = ~(n15217 | n14695);
assign n14884 = n26918 | n18827;
assign n27193 = ~(n19408 ^ n6879);
assign n22767 = ~(n27111 | n25265);
assign n1876 = ~n11482;
assign n4636 = n14053 & n12253;
assign n4203 = ~n5051;
assign n15987 = n13360 | n16392;
assign n5799 = n2903 | n4570;
assign n17300 = ~(n7731 | n13109);
assign n14481 = n15903 & n10802;
assign n21418 = n11334 & n8696;
assign n13161 = ~(n14695 ^ n15473);
assign n25510 = ~(n23234 | n20235);
assign n15172 = n19663 & n8025;
assign n26134 = ~n10932;
assign n9365 = ~n19234;
assign n24185 = n23555 | n26443;
assign n7855 = n10026 | n18432;
assign n5186 = ~(n15409 | n1145);
assign n19630 = n22729 & n18744;
assign n3906 = ~(n7826 ^ n26600);
assign n12234 = ~(n14723 ^ n24560);
assign n20120 = ~n10908;
assign n15902 = ~(n12025 ^ n21198);
assign n25011 = n19619 | n2625;
assign n1114 = ~(n15261 ^ n16902);
assign n9762 = n955 | n13509;
assign n4884 = n4143 | n19184;
assign n21456 = ~n11382;
assign n18668 = ~(n6283 ^ n19081);
assign n10098 = n14139 & n14838;
assign n18006 = ~(n5893 ^ n22488);
assign n18417 = n7618 & n22560;
assign n8340 = n17578 & n8653;
assign n12231 = ~(n21114 ^ n14477);
assign n19836 = ~(n3144 ^ n1683);
assign n6923 = ~(n5355 | n19094);
assign n26111 = ~(n7656 ^ n24176);
assign n7668 = n8468 & n24026;
assign n15694 = n17602 | n8644;
assign n19333 = ~(n18211 ^ n8674);
assign n3551 = ~(n2666 | n14739);
assign n99 = n12236 | n11589;
assign n5814 = n25036 | n18498;
assign n5981 = ~(n1267 ^ n12507);
assign n10728 = ~(n18650 ^ n17206);
assign n9453 = ~n25069;
assign n19080 = ~(n374 ^ n10483);
assign n9875 = ~(n23083 | n17858);
assign n15058 = ~(n7626 ^ n13691);
assign n7772 = n19790 & n19151;
assign n18507 = n3161 | n16888;
assign n26169 = ~(n6353 ^ n8434);
assign n822 = ~(n14743 ^ n2990);
assign n14850 = n15789 & n261;
assign n23261 = ~n25490;
assign n663 = ~n26102;
assign n4439 = n25759 | n25224;
assign n13655 = n14840 | n12489;
assign n18547 = ~n25594;
assign n4618 = ~(n10890 ^ n14157);
assign n17570 = n26644 | n15403;
assign n14972 = ~(n12335 ^ n11148);
assign n866 = n23912 | n25601;
assign n10844 = n24241 & n23713;
assign n3444 = n18268 | n15526;
assign n19524 = ~(n7397 ^ n14196);
assign n21786 = ~(n25291 ^ n7061);
assign n13060 = ~(n6164 ^ n22850);
assign n25256 = ~(n15247 ^ n19403);
assign n123 = ~(n12281 | n15007);
assign n26654 = ~n5682;
assign n26779 = n3120 | n14361;
assign n27091 = ~(n12291 | n25689);
assign n11946 = n16234 | n25069;
assign n6580 = ~n2210;
assign n19294 = ~(n2919 ^ n27037);
assign n4979 = n15895 | n16222;
assign n21424 = ~(n9589 ^ n18427);
assign n4633 = ~(n26472 | n7359);
assign n16357 = n4145 & n20725;
assign n1901 = n11052 | n21691;
assign n14432 = n21669 & n11836;
assign n17962 = n12444 | n25048;
assign n416 = n17212 | n16627;
assign n5489 = n17549 | n1657;
assign n17552 = n15344 & n4264;
assign n7859 = ~(n14899 ^ n18496);
assign n24466 = n16587 & n9501;
assign n21869 = n25877 & n6393;
assign n8816 = ~n11543;
assign n8525 = ~(n16576 | n10581);
assign n3538 = n12900 & n16547;
assign n9451 = ~(n22611 ^ n16979);
assign n11569 = ~(n20470 | n4590);
assign n23757 = ~(n5413 ^ n2185);
assign n227 = ~(n22964 ^ n19907);
assign n3242 = n3430 & n12994;
assign n26316 = ~n19765;
assign n13107 = n17981 | n7125;
assign n12437 = n16022 & n1519;
assign n7315 = n5432 | n12092;
assign n19371 = ~n26808;
assign n23861 = ~(n12734 ^ n23039);
assign n1060 = ~(n877 ^ n13202);
assign n26231 = ~(n21070 | n27078);
assign n23562 = n3198 & n18766;
assign n16225 = n21896 | n12494;
assign n20579 = ~(n15636 ^ n11615);
assign n21183 = n19242 & n3215;
assign n14632 = ~(n4181 | n2194);
assign n3413 = n14336 & n18149;
assign n14240 = n15819 & n3763;
assign n22423 = n9692 | n6761;
assign n11392 = ~(n3843 | n1336);
assign n12715 = n14818 & n26491;
assign n23557 = n3828 | n10392;
assign n6222 = ~n11273;
assign n11968 = ~(n23996 | n5685);
assign n12099 = ~(n19110 ^ n5467);
assign n24869 = n867 | n21430;
assign n4474 = n20180 & n26616;
assign n1382 = n25070 | n20637;
assign n7140 = n24223 & n14259;
assign n10825 = n23901 | n16038;
assign n6347 = n25846 | n5874;
assign n18030 = n2235 | n3556;
assign n25271 = ~n19357;
assign n27191 = ~(n8402 | n10987);
assign n14623 = n27131 | n473;
assign n9151 = ~(n20175 ^ n4514);
assign n2800 = n10530 & n21500;
assign n21818 = ~(n14016 ^ n22282);
assign n12240 = n20777 | n4712;
assign n16519 = ~(n18196 ^ n25380);
assign n2454 = ~(n12229 ^ n442);
assign n151 = ~n11971;
assign n15905 = ~n7678;
assign n15503 = ~(n3959 | n5855);
assign n17433 = ~n9997;
assign n10215 = n20097 & n11934;
assign n7153 = n20864 | n25262;
assign n1883 = ~(n21577 ^ n20290);
assign n13305 = ~n1160;
assign n9027 = ~(n2453 | n23095);
assign n5619 = ~(n24018 | n10499);
assign n5608 = ~(n9493 ^ n4426);
assign n16437 = n27061 & n8617;
assign n284 = n11590 & n21690;
assign n5690 = ~(n20259 | n22043);
assign n22001 = n24014 | n12728;
assign n19862 = ~n6385;
assign n10685 = ~(n13945 ^ n19163);
assign n11494 = ~(n25688 ^ n27104);
assign n154 = ~(n2982 ^ n21120);
assign n25544 = n987 | n11871;
assign n13192 = n20522 & n17007;
assign n22418 = ~(n24879 | n3687);
assign n20060 = ~(n17886 ^ n20219);
assign n10468 = ~(n20374 ^ n1266);
assign n14802 = n7119 | n25171;
assign n25035 = n15276 | n21659;
assign n26699 = ~(n10995 ^ n13894);
assign n2948 = ~(n19343 ^ n7958);
assign n7411 = n16417 | n2924;
assign n12571 = n13514 & n5492;
assign n19956 = ~n16833;
assign n22458 = ~(n20754 ^ n24786);
assign n23321 = ~n22909;
assign n3422 = ~(n20036 | n23537);
assign n16741 = n14909 | n2601;
assign n4708 = n18554 | n4497;
assign n14604 = n20489 | n26913;
assign n7733 = ~(n25015 | n1850);
assign n21709 = n3160 | n9414;
assign n12831 = ~(n446 | n12650);
assign n642 = ~n17780;
assign n21616 = n4584 & n11916;
assign n25102 = ~(n24561 ^ n8782);
assign n18277 = ~(n2601 ^ n10304);
assign n22523 = ~(n23114 | n3454);
assign n12331 = n15620 | n7977;
assign n21608 = ~n376;
assign n15004 = ~(n23201 ^ n23151);
assign n7903 = n10648 & n18392;
assign n8876 = n12169 | n6414;
assign n19543 = ~n9376;
assign n21279 = n15217 | n17542;
assign n16955 = n22424 & n25417;
assign n12524 = ~(n16543 | n22862);
assign n25022 = n23913 & n8144;
assign n26044 = ~(n6848 ^ n23920);
assign n14016 = ~n25436;
assign n2296 = ~(n16536 | n13492);
assign n23765 = n592 | n3347;
assign n15245 = n21138 & n23804;
assign n10738 = ~(n25021 | n21997);
assign n8965 = ~(n14635 ^ n15773);
assign n11984 = n27001 | n12263;
assign n5108 = ~n1658;
assign n19646 = ~(n13077 ^ n7702);
assign n25953 = ~n25490;
assign n23730 = n17240 & n4355;
assign n11887 = n6995 | n8452;
assign n5966 = n1819 | n19709;
assign n19458 = n7501 | n14717;
assign n668 = n19887 | n22246;
assign n15098 = n7382 | n20018;
assign n5686 = n26830 | n19707;
assign n16326 = ~(n18123 | n4569);
assign n21445 = n18185 & n19801;
assign n15348 = n22480 | n17703;
assign n17353 = ~(n26124 ^ n6379);
assign n3737 = ~(n4859 | n25972);
assign n25311 = n8735 | n2055;
assign n21019 = n11337 | n12430;
assign n24571 = ~(n27113 | n16704);
assign n5164 = n25249 ^ n25795;
assign n17952 = n9690 & n24036;
assign n21145 = n18382 | n24216;
assign n5017 = n18101 | n12550;
assign n13005 = ~(n2074 ^ n2390);
assign n26430 = n26266 | n22785;
assign n13063 = n9138 | n10896;
assign n173 = ~n24129;
assign n6384 = n20617 | n26977;
assign n3212 = n3142 | n12937;
assign n3561 = ~(n16776 | n25386);
assign n164 = n3473 | n20580;
assign n15953 = n26592 | n21932;
assign n9181 = n5295 | n9812;
assign n12693 = ~n14110;
assign n17602 = n26636 & n19661;
assign n24936 = ~n18833;
assign n5770 = ~(n17350 ^ n8784);
assign n2049 = ~n16896;
assign n20856 = n18916 | n1974;
assign n24181 = ~(n22191 | n265);
assign n364 = n1118 & n6477;
assign n25043 = ~(n8708 ^ n21047);
assign n450 = ~(n14337 ^ n7876);
assign n8504 = n6659 & n12991;
assign n20558 = ~n13743;
assign n14008 = ~(n928 ^ n21384);
assign n18669 = ~(n16029 | n19228);
assign n15622 = ~(n12405 | n19489);
assign n2795 = n2371 | n19255;
assign n8499 = n19867 | n27191;
assign n22205 = n15066 | n6970;
assign n16200 = ~n16312;
assign n981 = n7049 | n18877;
assign n21277 = n13944 | n23871;
assign n17428 = ~n18281;
assign n15942 = ~(n15167 | n23921);
assign n13552 = n18138 & n14743;
assign n22784 = n7129 & n8211;
assign n21044 = ~(n12658 ^ n26618);
assign n20762 = n24867 | n5310;
assign n10233 = ~(n26748 ^ n12161);
assign n1544 = n12866 & n24713;
assign n12976 = ~(n11669 | n11366);
assign n10683 = ~n3161;
assign n24629 = ~(n11240 ^ n24271);
assign n18918 = n16580 & n19587;
assign n21005 = ~(n13282 ^ n14685);
assign n24890 = ~n18558;
assign n3605 = n15167 | n25330;
assign n22220 = ~(n17979 | n11158);
assign n6959 = ~(n27100 | n25637);
assign n17794 = ~(n7817 | n23036);
assign n6129 = ~(n16474 ^ n15491);
assign n17054 = n20040 & n23983;
assign n2907 = n25409 | n23154;
assign n19844 = ~n4296;
assign n15220 = ~(n18049 ^ n2365);
assign n9236 = n26263 & n77;
assign n5534 = n14163 | n921;
assign n19914 = ~n4446;
assign n3452 = ~(n23168 | n13028);
assign n17075 = ~(n2687 ^ n6346);
assign n20486 = ~(n2141 | n23851);
assign n12776 = ~(n106 ^ n26882);
assign n26175 = n15665 | n1033;
assign n19827 = ~(n3124 | n5516);
assign n7894 = ~(n10303 ^ n1136);
assign n24700 = ~(n21415 ^ n924);
assign n12899 = n22918 | n20719;
assign n4504 = n13781 & n24358;
assign n13887 = ~(n10051 | n3526);
assign n19181 = ~n26936;
assign n5419 = ~(n10981 ^ n6517);
assign n8623 = ~n23181;
assign n3323 = n18442 & n12611;
assign n1804 = ~(n25021 | n19025);
assign n19339 = n11159 & n10186;
assign n20815 = n26779 & n5588;
assign n14219 = n1825 | n15095;
assign n26680 = ~n3846;
assign n13826 = ~(n18707 ^ n19618);
assign n21525 = ~(n25780 ^ n26969);
assign n7655 = n17300 | n12466;
assign n4813 = ~(n1398 ^ n1552);
assign n16112 = n18857 | n5242;
assign n4080 = n18080 & n24398;
assign n23907 = n13385 & n8618;
assign n20870 = n26571 | n21791;
assign n19088 = ~(n11425 | n12657);
assign n39 = n9193 & n12854;
assign n1151 = ~n6218;
assign n9463 = ~(n11062 ^ n21489);
assign n15186 = ~(n18814 | n8645);
assign n25075 = n8685 & n21283;
assign n16617 = ~(n18359 ^ n1052);
assign n16077 = ~(n5570 ^ n17667);
assign n13896 = n17523 & n5671;
assign n19559 = n5885 | n17686;
assign n8450 = n9011 | n19143;
assign n4424 = ~(n18706 ^ n11744);
assign n18884 = n9679 | n4319;
assign n19073 = n744 | n18630;
assign n23921 = ~n3786;
assign n14176 = ~(n16743 ^ n5882);
assign n25481 = n25291 | n13743;
assign n7179 = n22039 & n1520;
assign n23498 = ~(n5165 ^ n6834);
assign n14660 = n23990 | n14184;
assign n24249 = n8827 | n26142;
assign n26343 = ~(n11390 ^ n26705);
assign n26253 = n18145 | n12168;
assign n25105 = n20411 | n17212;
assign n20609 = ~(n378 ^ n23743);
assign n11490 = n5624 | n21632;
assign n14557 = ~n17152;
assign n6467 = ~(n26584 ^ n14830);
assign n9805 = ~(n12446 | n6553);
assign n6582 = n15070 & n25672;
assign n10885 = ~n24292;
assign n11539 = ~(n21121 ^ n22692);
assign n25287 = n27183 | n2150;
assign n8301 = n25218 & n5527;
assign n8350 = n5491 | n4664;
assign n17260 = n3791 | n24301;
assign n12444 = ~(n22425 | n4461);
assign n21736 = ~(n14758 ^ n25636);
assign n16068 = ~(n22648 ^ n8530);
assign n20358 = ~n23104;
assign n13742 = n24639 & n7663;
assign n13142 = ~(n2289 ^ n20946);
assign n5617 = ~(n9236 ^ n17157);
assign n20903 = n20532 | n7416;
assign n21650 = n24402 | n13123;
assign n25646 = n15882 & n25039;
assign n2723 = ~(n1846 ^ n22502);
assign n25237 = ~n5669;
assign n22528 = n16020 & n10907;
assign n5431 = n16476 & n19146;
assign n662 = n10721 | n7845;
assign n1748 = n22186 | n11657;
assign n23314 = ~(n23864 | n17994);
assign n3408 = ~(n1262 | n1777);
assign n3343 = ~(n18298 ^ n14952);
assign n334 = n6984 & n3954;
assign n6927 = n8244 & n22820;
assign n11084 = n19764 & n8114;
assign n20364 = ~(n4299 ^ n10843);
assign n25028 = n12217 | n5701;
assign n21120 = ~(n4870 ^ n2857);
assign n26073 = ~(n3783 ^ n11630);
assign n8851 = ~n20794;
assign n6407 = ~(n2554 ^ n14949);
assign n15695 = ~n22843;
assign n7143 = ~n400;
assign n3214 = n13859 & n26276;
assign n7660 = ~(n12217 ^ n23798);
assign n13877 = ~(n8107 ^ n18363);
assign n23279 = ~(n26983 ^ n24076);
assign n8735 = ~n23559;
assign n18184 = n9705 | n12448;
assign n6588 = n16464 | n16223;
assign n13172 = ~n8827;
assign n26287 = ~(n18757 ^ n5162);
assign n715 = n23494 & n14812;
assign n26993 = ~n18805;
assign n4837 = n6442 & n8959;
assign n9951 = n8101 | n3019;
assign n26684 = n12624 & n15735;
assign n7162 = ~(n14815 ^ n18958);
assign n17825 = n24264 | n7178;
assign n11835 = ~n10651;
assign n18292 = n18765 | n21975;
assign n8325 = n25502 | n1545;
assign n2756 = ~n20477;
assign n779 = n8345 | n24628;
assign n739 = ~n25814;
assign n11349 = n27183 & n2150;
assign n17435 = n25748 | n3751;
assign n7404 = n15676 | n21116;
assign n11939 = n1656 | n11397;
assign n22709 = n12709 | n8085;
assign n20147 = n4352 & n11683;
assign n23650 = ~(n20134 ^ n15237);
assign n5702 = n24229 | n5801;
assign n20598 = n7644 & n11235;
assign n18019 = n19848 | n6979;
assign n3644 = n14431 & n25739;
assign n25407 = ~(n3840 | n11254);
assign n18401 = n14655 | n9565;
assign n16330 = n15061 & n14892;
assign n8415 = ~n19707;
assign n24356 = n9417 & n11558;
assign n17364 = n2520 | n2267;
assign n6838 = ~(n22119 ^ n9252);
assign n3421 = ~(n1163 ^ n24620);
assign n23084 = ~n6246;
assign n5637 = ~(n19005 ^ n24618);
assign n6252 = n524 | n14736;
assign n10697 = n13590 | n22370;
assign n15224 = ~(n19616 | n26673);
assign n7291 = n5015 & n18246;
assign n23032 = ~(n19156 ^ n24706);
assign n7611 = n6111 | n16868;
assign n22904 = n11331 & n17988;
assign n3728 = ~(n19594 ^ n25627);
assign n13290 = ~(n10184 | n22470);
assign n10766 = ~(n20151 ^ n19042);
assign n15919 = ~(n8974 ^ n14289);
assign n18772 = n16819 | n5017;
assign n7699 = n9732 | n26441;
assign n5738 = n569 & n8110;
assign n1135 = n27068 | n10505;
assign n8215 = ~(n7220 ^ n17920);
assign n5212 = ~n12168;
assign n9487 = ~(n4602 ^ n12402);
assign n24103 = ~(n16544 | n2160);
assign n1239 = ~(n22397 ^ n12191);
assign n21027 = n18384 | n12952;
assign n13650 = ~(n1688 ^ n3544);
assign n23859 = n27125 & n26595;
assign n14941 = ~(n4973 ^ n17563);
assign n14300 = ~(n21140 ^ n24456);
assign n17812 = ~n12145;
assign n20808 = ~n22748;
assign n5341 = ~n14066;
assign n17813 = ~(n26724 ^ n1777);
assign n24977 = ~(n26875 ^ n6131);
assign n10196 = ~(n6442 ^ n6828);
assign n11738 = ~(n8828 ^ n6443);
assign n3832 = ~(n6797 ^ n22568);
assign n8762 = ~(n6895 ^ n4858);
assign n13126 = ~(n23317 | n38);
assign n20789 = ~(n26982 | n2679);
assign n12125 = ~(n5657 ^ n5704);
assign n12427 = ~(n5914 | n790);
assign n26357 = n26059 | n7672;
assign n2354 = n18274 & n24383;
assign n22 = ~(n3743 | n3038);
assign n4473 = ~(n19680 | n18341);
assign n10232 = n8064 & n449;
assign n13841 = ~(n8030 ^ n4050);
assign n18888 = ~(n22690 ^ n4736);
assign n19580 = n26547 & n15163;
assign n22968 = ~n17277;
assign n25548 = ~(n9069 | n22169);
assign n5024 = ~(n23764 ^ n21533);
assign n8029 = n122 | n15227;
assign n2616 = ~(n23146 | n21585);
assign n16370 = n14186 | n27170;
assign n24133 = ~(n12370 ^ n11613);
assign n10090 = ~(n25370 | n23819);
assign n13230 = ~(n4502 ^ n13760);
assign n401 = ~n19905;
assign n25647 = n11707 ^ n14829;
assign n17702 = n2735 & n5628;
assign n13553 = ~n18632;
assign n8469 = n9361 | n2947;
assign n2470 = ~(n21333 ^ n232);
assign n13982 = ~n13006;
assign n17233 = n9257 | n5798;
assign n17802 = n26797 & n14654;
assign n8142 = n27038 | n19374;
assign n9726 = ~(n10196 ^ n20741);
assign n14687 = ~(n1802 ^ n6038);
assign n116 = n20023 | n12734;
assign n1776 = n17954 | n23767;
assign n13233 = n21188 | n10011;
assign n14173 = n19277 | n6327;
assign n8349 = ~(n18664 ^ n9077);
assign n22155 = ~(n20966 | n17938);
assign n8357 = n8212 | n1782;
assign n24332 = n3594 | n1504;
assign n115 = ~(n16723 ^ n24618);
assign n4284 = ~(n1380 ^ n11220);
assign n2975 = ~(n2750 | n7543);
assign n15119 = n6348 & n6116;
assign n24813 = ~n11817;
assign n18787 = ~n7775;
assign n7406 = ~(n16821 ^ n21545);
assign n14996 = ~(n22956 ^ n11952);
assign n3632 = ~n26311;
assign n20768 = ~(n1690 | n1000);
assign n14485 = n12940 | n6157;
assign n10409 = ~(n11214 ^ n2078);
assign n8296 = ~(n22892 ^ n24298);
assign n1733 = ~(n24091 ^ n2272);
assign n9383 = n18151 & n6414;
assign n5327 = n10494 | n26304;
assign n11287 = ~(n14826 ^ n17458);
assign n23327 = n17780 | n12430;
assign n20202 = n22626 & n18765;
assign n18302 = ~(n8571 ^ n10872);
assign n20969 = n25680 | n14348;
assign n19378 = ~(n10837 ^ n1576);
assign n13062 = ~n23432;
assign n13537 = n20777 | n2461;
assign n14255 = ~n17064;
assign n9991 = ~(n19588 | n13329);
assign n10147 = ~(n4479 | n23724);
assign n14001 = n19361 & n15918;
assign n6930 = ~(n16932 | n6913);
assign n21947 = n17999 | n17982;
assign n25154 = n25506 | n14237;
assign n15190 = ~(n25880 ^ n18609);
assign n542 = n1144 & n9299;
assign n22876 = n15550 & n2347;
assign n185 = ~(n24862 ^ n3906);
assign n4352 = n4085 | n16547;
assign n15966 = n8845 | n22773;
assign n237 = n24004 | n12900;
assign n2386 = n160 & n25275;
assign n16759 = ~(n17881 ^ n25068);
assign n5761 = n2409 | n25057;
assign n11610 = n18737 | n2328;
assign n3944 = n12997 & n13532;
assign n1219 = n16319 | n19170;
assign n23527 = n94 & n9476;
assign n339 = ~n9926;
assign n26977 = n2527 & n23507;
assign n16746 = ~(n10650 ^ n22253);
assign n5900 = n9883 | n13885;
assign n3794 = ~(n18390 ^ n13587);
assign n3750 = ~(n16880 | n21734);
assign n6418 = ~(n12911 ^ n1222);
assign n8034 = n3466 & n19917;
assign n7052 = ~(n2085 ^ n5169);
assign n20089 = ~n12384;
assign n23815 = n10043 | n25252;
assign n5569 = ~n26216;
assign n12052 = n25445 | n244;
assign n26889 = n21588 & n15449;
assign n8722 = ~(n6931 ^ n17612);
assign n9290 = ~n9460;
assign n11341 = n12923 & n204;
assign n2695 = ~(n2155 ^ n16938);
assign n12577 = n689 & n19627;
assign n17610 = ~n26752;
assign n10690 = n25841 | n3053;
assign n8672 = ~(n26886 ^ n1099);
assign n19229 = ~n2146;
assign n19293 = n19797 | n3903;
assign n2071 = ~n14480;
assign n2182 = n10696 | n72;
assign n25162 = n11804 | n17755;
assign n14807 = n17248 | n21020;
assign n16319 = ~(n25030 ^ n1549);
assign n25534 = n26036 | n7832;
assign n10210 = ~(n2432 ^ n15017);
assign n23175 = ~n8850;
assign n24050 = ~(n22550 | n7465);
assign n4410 = ~(n25081 ^ n17560);
assign n18432 = n3493 & n24087;
assign n2603 = n10313 | n26932;
assign n17234 = ~(n3405 | n9665);
assign n3939 = ~n17204;
assign n14141 = n3915 | n17411;
assign n18369 = n1879 | n670;
assign n14700 = ~n6734;
assign n5197 = n5061 & n6016;
assign n23496 = n5567 | n19152;
assign n23754 = ~(n12310 ^ n6575);
assign n13882 = n6805 | n8679;
assign n8829 = n19890 | n12810;
assign n18970 = ~(n26663 ^ n20087);
assign n15 = ~n21143;
assign n20287 = ~(n11802 ^ n9112);
assign n23100 = ~(n9765 ^ n20213);
assign n21756 = ~(n6032 | n13623);
assign n11408 = ~(n27016 ^ n14947);
assign n11787 = ~(n8363 ^ n2816);
assign n22071 = ~n1752;
assign n4157 = n18207 | n25511;
assign n18573 = n15636 & n25139;
assign n9522 = n25628 | n27129;
assign n9348 = n2176 | n19561;
assign n8203 = ~(n25470 | n12898);
assign n21919 = ~(n19222 ^ n6691);
assign n9404 = ~n25441;
assign n20435 = n23011 & n23971;
assign n23145 = ~(n27109 ^ n3884);
assign n10397 = ~(n24247 | n558);
assign n19918 = n20497 | n16482;
assign n1091 = ~n14323;
assign n8104 = n18734 | n14870;
assign n6445 = ~(n15457 ^ n15997);
assign n21910 = ~n1278;
assign n19047 = ~n14648;
assign n11187 = ~(n20151 | n22428);
assign n26171 = n995 & n229;
assign n17081 = ~(n12950 ^ n8083);
assign n12841 = ~(n801 | n10760);
assign n12817 = n22725 | n11480;
assign n12336 = n13777 & n15370;
assign n26831 = n23430 | n20628;
assign n2546 = ~(n19702 ^ n19270);
assign n3960 = ~(n4236 ^ n22846);
assign n2791 = n5993 | n13104;
assign n13931 = n10209 | n19442;
assign n4805 = n20831 & n26690;
assign n26300 = ~n21210;
assign n2685 = n22820 | n19137;
assign n13515 = ~(n11302 | n20948);
assign n14000 = ~(n26255 | n27102);
assign n14843 = ~(n15603 ^ n15901);
assign n21372 = n26895 | n13543;
assign n2085 = ~n4759;
assign n12725 = ~(n3654 ^ n20996);
assign n23499 = n4390 & n2381;
assign n17360 = ~n23890;
assign n8963 = n5397 & n17825;
assign n14489 = n4144 | n25634;
assign n26377 = ~(n10903 | n24584);
assign n20766 = n3428 | n25216;
assign n1891 = ~(n19008 ^ n2524);
assign n3114 = ~(n12265 | n5728);
assign n6470 = ~(n13055 ^ n20172);
assign n21829 = ~(n5374 | n23002);
assign n14159 = n3736 | n4790;
assign n10797 = ~(n12717 ^ n25679);
assign n22355 = ~(n7628 ^ n23982);
assign n21746 = ~(n4749 ^ n12385);
assign n19642 = ~(n10590 ^ n3677);
assign n1812 = n12107 & n10853;
assign n5172 = ~n6379;
assign n3226 = n15861 & n4887;
assign n15406 = ~(n20937 ^ n21596);
assign n25418 = ~(n13748 ^ n24923);
assign n8517 = n9614 & n6890;
assign n24035 = ~(n26495 ^ n5789);
assign n26769 = ~n26935;
assign n4159 = ~(n2713 | n25271);
assign n18693 = ~(n2584 ^ n10698);
assign n20594 = ~(n10198 ^ n6119);
assign n18214 = n20112 | n26102;
assign n1785 = ~(n8196 | n3992);
assign n6772 = ~(n15389 ^ n23913);
assign n13902 = n8647 | n26226;
assign n23957 = ~(n14761 | n26460);
assign n3065 = n1556 & n13974;
assign n5062 = ~(n4934 ^ n18279);
assign n22935 = n19586 & n18147;
assign n6277 = n13666 & n1131;
assign n16155 = ~(n13668 | n835);
assign n7565 = n21979 | n23135;
assign n25909 = n24311 | n17430;
assign n17853 = ~(n22378 ^ n22619);
assign n138 = n26648 & n8817;
assign n3607 = n7066 & n9413;
assign n4699 = n3506 & n26414;
assign n14921 = n7396 | n27178;
assign n10209 = ~(n12650 | n11220);
assign n8660 = ~(n20638 ^ n10512);
assign n8320 = ~(n16100 ^ n23139);
assign n11313 = ~(n4663 ^ n8409);
assign n18063 = n8129 & n8972;
assign n25335 = n647 | n1773;
assign n18842 = n6209 | n2597;
assign n8227 = ~n2111;
assign n15509 = n15920 & n13545;
assign n19982 = ~(n19411 ^ n5978);
assign n15480 = n10319 | n23812;
assign n7086 = ~(n26008 ^ n17201);
assign n24205 = n2102 | n19560;
assign n5907 = ~(n19406 | n21905);
assign n20152 = n26870 & n7902;
assign n2586 = ~(n26011 ^ n4154);
assign n25106 = ~(n20999 ^ n3353);
assign n18221 = ~(n20137 | n17077);
assign n13991 = ~(n11525 | n11258);
assign n23485 = n17896 & n1475;
assign n18144 = n20375 & n16075;
assign n25104 = ~(n18047 ^ n22933);
assign n6479 = n16910 | n502;
assign n23906 = n10190 | n5478;
assign n23667 = ~(n7604 ^ n11580);
assign n23112 = n5406 | n11145;
assign n25852 = ~(n20011 ^ n17953);
assign n7271 = ~(n23352 ^ n22953);
assign n14249 = ~n10765;
assign n14426 = n2979 | n23258;
assign n3434 = n22867 | n12334;
assign n15369 = ~(n26654 | n3554);
assign n4451 = ~(n1675 ^ n20220);
assign n25881 = n1571 & n23833;
assign n3423 = ~(n19888 | n13308);
assign n13648 = ~(n10152 ^ n10581);
assign n21274 = n13173 & n10006;
assign n16749 = n11328 | n21255;
assign n24579 = ~(n19219 ^ n27197);
assign n9725 = ~(n7674 | n16468);
assign n26123 = ~(n2057 | n19603);
assign n10524 = n23021 & n4690;
assign n7953 = ~n13775;
assign n15897 = ~n3012;
assign n8487 = ~(n1542 ^ n12916);
assign n20281 = n13822 | n767;
assign n11466 = n23114 | n6362;
assign n5422 = n11188 | n21316;
assign n17541 = n6185 & n11646;
assign n20979 = n26284 & n12403;
assign n12040 = ~n2732;
assign n23614 = n4085 | n3211;
assign n12431 = n10274 | n17636;
assign n17978 = ~(n24717 ^ n2979);
assign n20884 = n26899 | n4743;
assign n11095 = ~(n24985 ^ n185);
assign n15103 = n3984 | n22153;
assign n18012 = ~(n2341 | n2967);
assign n22261 = ~n3306;
assign n3558 = n20224 | n23881;
assign n5523 = ~n24474;
assign n8492 = n15931;
assign n7779 = ~(n13745 ^ n26460);
assign n19363 = ~(n10710 ^ n23529);
assign n11626 = n25129 | n9446;
assign n4762 = ~(n14507 ^ n17488);
assign n4890 = ~(n10081 ^ n890);
assign n5178 = ~(n12633 ^ n9900);
assign n19499 = n1203 | n24556;
assign n22556 = n9045 & n4437;
assign n24721 = ~(n21644 ^ n18555);
assign n12074 = n12458 | n26373;
assign n547 = n9258 & n19250;
assign n1345 = n1615 & n20856;
assign n3663 = ~(n24291 ^ n17196);
assign n839 = ~n12342;
assign n15758 = ~(n10468 ^ n20770);
assign n27177 = ~(n12513 ^ n25568);
assign n19168 = ~(n23313 | n16345);
assign n1626 = ~n8391;
assign n23453 = ~(n7785 ^ n7817);
assign n6394 = ~(n24665 ^ n5704);
assign n20895 = n26258 & n10154;
assign n27055 = ~(n1365 ^ n23333);
assign n2435 = n8016 | n21911;
assign n5939 = ~(n14230 | n10185);
assign n22451 = n3599 | n5366;
assign n20212 = n25726 | n5200;
assign n5804 = ~(n23084 ^ n3253);
assign n13849 = n2970 | n3793;
assign n9653 = ~(n20295 ^ n23659);
assign n22294 = ~(n1686 ^ n1292);
assign n17755 = ~n3031;
assign n2763 = n21324 | n1446;
assign n14020 = n10794 | n10400;
assign n18855 = n1003 & n8931;
assign n14033 = ~n1414;
assign n20289 = ~n387;
assign n1955 = n17768 | n8517;
assign n16565 = n18749 & n4156;
assign n20090 = n5572 | n7684;
assign n18127 = n14560 | n4267;
assign n19355 = ~(n20828 ^ n6751);
assign n7684 = ~(n2398 ^ n107);
assign n22933 = ~(n8938 ^ n4255);
assign n11051 = n405 & n4561;
assign n16858 = ~(n23878 ^ n2035);
assign n9415 = ~(n19863 ^ n2210);
assign n16856 = ~n24488;
assign n21992 = n25914 | n20359;
assign n17902 = ~(n15957 ^ n23697);
assign n8543 = n821 | n17584;
assign n18582 = ~(n11215 ^ n19533);
assign n26085 = ~n23235;
assign n11983 = n21831 & n25448;
assign n23102 = n13480 & n22769;
assign n8719 = ~n8406;
assign n17735 = ~(n16132 ^ n22857);
assign n26792 = n3629 & n10474;
assign n18403 = n16903 | n17061;
assign n25159 = n5068 | n14715;
assign n15105 = ~(n2980 ^ n12514);
assign n26261 = n24321 & n18885;
assign n24501 = ~(n18229 ^ n25509);
assign n21532 = ~(n1437 ^ n17784);
assign n20764 = n6608 & n19654;
assign n23389 = n17603 & n22608;
assign n25195 = ~(n8713 ^ n24736);
assign n21715 = ~(n3937 | n21295);
assign n5769 = ~(n2355 ^ n16223);
assign n11381 = n10777;
assign n11686 = n24848 | n23972;
assign n11327 = n2562 & n5823;
assign n11870 = ~(n13136 | n26065);
assign n24701 = ~n1162;
assign n4653 = n17376 | n8842;
assign n15006 = ~(n7769 | n26625);
assign n11746 = ~(n15512 ^ n22607);
assign n7603 = n19068 | n9925;
assign n15174 = n18027 & n4866;
assign n19547 = n13982 & n15092;
assign n17023 = ~(n6381 ^ n13914);
assign n26721 = n22896 & n26345;
assign n12417 = ~(n22449 ^ n7157);
assign n17047 = ~n4537;
assign n20960 = n16919 & n7628;
assign n22541 = n19822 & n17760;
assign n10466 = ~(n10882 ^ n8406);
assign n21916 = n3366 | n15670;
assign n13120 = n9001 & n20995;
assign n3535 = n2315 & n17375;
assign n543 = ~(n7888 ^ n5500);
assign n18810 = ~(n13884 ^ n7917);
assign n20267 = ~(n20796 ^ n5140);
assign n22052 = n12811 | n11822;
assign n10067 = ~(n19106 | n2680);
assign n22635 = ~(n22093 ^ n26743);
assign n15796 = ~n13490;
assign n18554 = ~n14230;
assign n9750 = ~(n15241 ^ n15146);
assign n26502 = n7338 | n10899;
assign n23780 = n3797 & n2203;
assign n7922 = n26577 | n3052;
assign n1167 = n16743 | n16875;
assign n6137 = ~n3477;
assign n26648 = ~n12440;
assign n8049 = n20409 | n19117;
assign n21514 = n16743 & n24485;
assign n17382 = ~(n25089 ^ n10253);
assign n2624 = n13459 | n593;
assign n22724 = ~n21222;
assign n7078 = n8547 | n22045;
assign n6463 = ~(n16162 ^ n10251);
assign n23086 = ~(n18551 ^ n8632);
assign n20772 = ~(n20131 ^ n17418);
assign n12329 = ~(n13431 ^ n13943);
assign n4182 = ~(n26830 ^ n8415);
assign n19615 = ~n26803;
assign n4109 = ~n7706;
assign n741 = n18485 | n2731;
assign n8977 = n6204 | n5065;
assign n25373 = ~(n16482 ^ n13333);
assign n22082 = ~(n1271 ^ n26647);
assign n1103 = ~(n8847 | n3993);
assign n6003 = ~(n9212 ^ n3456);
assign n16618 = ~n24901;
assign n4443 = ~(n6259 ^ n24152);
assign n2594 = n20326 | n5694;
assign n22190 = n22882 | n21572;
assign n19195 = ~(n10557 | n12381);
assign n23864 = ~(n23501 ^ n10563);
assign n1257 = n1709 & n24961;
assign n4550 = n22031 & n20824;
assign n20574 = ~(n20542 ^ n9575);
assign n18002 = ~(n26277 ^ n23778);
assign n157 = n26510 & n11246;
assign n14593 = ~(n23017 ^ n23853);
assign n22761 = ~(n4244 ^ n7345);
assign n9711 = ~n1845;
assign n1329 = ~n5438;
assign n16516 = ~(n8838 ^ n4828);
assign n11125 = n21867 & n8557;
assign n38 = n13886 & n17242;
assign n9029 = n22250 | n1071;
assign n7640 = ~(n3885 ^ n19208);
assign n16854 = ~(n12398 | n23586);
assign n2091 = n12622 & n26289;
assign n13795 = n9053 | n22015;
assign n3879 = ~(n23895 | n13976);
assign n7950 = ~(n19528 ^ n24782);
assign n23884 = ~(n17004 | n24496);
assign n11316 = ~(n23099 | n17517);
assign n1964 = n6168 | n4537;
assign n23500 = ~(n22849 | n16824);
assign n19318 = n21528 & n7488;
assign n23196 = ~(n19905 ^ n3030);
assign n7910 = ~n24203;
assign n8684 = n20379 | n10677;
assign n6452 = n932 & n2666;
assign n21798 = n15103 & n25325;
assign n8592 = n13052 & n4635;
assign n14189 = ~(n5441 ^ n2426);
assign n2371 = ~(n19213 ^ n25730);
assign n13943 = ~(n25049 ^ n23451);
assign n23093 = n24582 | n14116;
assign n18599 = ~(n9272 ^ n16764);
assign n2227 = n8451 | n7555;
assign n8968 = n18514 | n15182;
assign n5629 = ~n8297;
assign n6258 = n26725 | n24292;
assign n10908 = ~(n26622 ^ n11471);
assign n24952 = n18014 | n20619;
assign n3702 = n23030 | n8381;
assign n8282 = ~(n4665 ^ n24278);
assign n6268 = ~(n25913 | n15568);
assign n16945 = n19339 | n21770;
assign n19456 = ~(n5739 ^ n4293);
assign n6359 = ~(n16313 ^ n25736);
assign n6071 = ~n20417;
assign n5861 = n787 | n9973;
assign n3916 = ~(n18145 ^ n19196);
assign n6027 = ~(n14153 | n16466);
assign n5936 = ~(n10914 ^ n11892);
assign n24993 = ~(n14765 ^ n12650);
assign n21428 = ~(n2651 | n4400);
assign n11826 = ~(n481 | n11220);
assign n12144 = ~(n1444 ^ n15239);
assign n11403 = ~(n6297 ^ n17016);
assign n17676 = ~(n17277 | n12869);
assign n3127 = ~(n9445 | n5812);
assign n13335 = n10277 | n1082;
assign n19053 = n16806 | n16005;
assign n19959 = n15244 | n23952;
assign n11405 = n17581 & n4330;
assign n22559 = n8101 & n9468;
assign n15137 = ~n3071;
assign n23332 = n19083 | n7450;
assign n8644 = ~(n20059 | n15603);
assign n708 = ~(n15580 | n4913);
assign n3211 = ~(n11549 ^ n14223);
assign n18501 = n9863 | n19480;
assign n17191 = n8069 & n4044;
assign n18064 = n9607 & n14935;
assign n20427 = ~(n1197 ^ n25061);
assign n5522 = ~(n9206 ^ n23792);
assign n5365 = ~(n13359 ^ n4665);
assign n2516 = n18814 | n802;
assign n22235 = n726 | n26849;
assign n24443 = n10382 & n24001;
assign n19556 = ~n26248;
assign n1770 = n23574 & n18923;
assign n24515 = n23182 | n5542;
assign n15646 = n11884 | n13313;
assign n14925 = n23687 | n12025;
assign n18786 = ~n2565;
assign n5934 = ~n2900;
assign n4368 = ~(n14549 ^ n25861);
assign n18581 = ~n11048;
assign n21721 = ~n22395;
assign n16264 = ~(n6792 ^ n410);
assign n1281 = ~(n7682 | n3952);
assign n26124 = ~n3040;
assign n11268 = ~n11383;
assign n9545 = n23937 | n282;
assign n12063 = ~(n2570 ^ n7569);
assign n17021 = n16594 | n23250;
assign n27000 = n19372 | n25902;
assign n985 = ~(n13574 ^ n9341);
assign n102 = ~(n14079 ^ n19670);
assign n15339 = ~(n23827 ^ n27070);
assign n2576 = ~n18157;
assign n1680 = ~(n4877 | n11135);
assign n4468 = ~n23974;
assign n23992 = n8066 | n23340;
assign n14393 = ~(n20110 ^ n1147);
assign n14391 = ~(n9188 ^ n10612);
assign n1591 = ~(n21740 | n12547);
assign n21932 = n3941 & n2701;
assign n27123 = n14882 | n21072;
assign n5450 = n23390 | n1411;
assign n6535 = ~n7073;
assign n14994 = n9698 & n1818;
assign n7256 = ~(n13706 ^ n2033);
assign n19092 = n19161 | n22405;
assign n5832 = ~(n13820 ^ n5541);
assign n1287 = n2458 & n1732;
assign n23373 = n11229 & n9741;
assign n22219 = ~n3721;
assign n3157 = n23920 | n25920;
assign n6784 = n7521 | n9871;
assign n17346 = n3349 | n10501;
assign n9960 = n5538 & n24111;
assign n19520 = ~n27170;
assign n19968 = ~(n16089 ^ n9316);
assign n22690 = n4839 & n17133;
assign n4131 = n14228 | n14770;
assign n6383 = ~(n22936 ^ n10596);
assign n22827 = n8010 | n19086;
assign n15969 = ~(n7307 ^ n9728);
assign n2609 = n24103 | n2025;
assign n3229 = ~(n2545 ^ n3740);
assign n17436 = ~(n872 ^ n10214);
assign n2967 = ~n23068;
assign n12388 = n25741 & n19942;
assign n2234 = ~(n10098 | n263);
assign n3798 = n3313 & n4367;
assign n24381 = n22290 & n13018;
assign n18385 = ~(n17351 | n21850);
assign n6584 = n24417 & n4719;
assign n13391 = ~n9850;
assign n5560 = n19618 & n18707;
assign n8560 = n18088 | n11173;
assign n1578 = n1802 & n7331;
assign n20129 = ~n25384;
assign n24075 = n8199 | n22638;
assign n21036 = ~(n18880 | n15456);
assign n11025 = ~(n5490 ^ n7599);
assign n8744 = ~(n4135 ^ n13610);
assign n17053 = n25187 | n23728;
assign n9093 = ~(n23368 ^ n19793);
assign n16023 = n19024 | n5893;
assign n4070 = ~(n25603 | n14389);
assign n2555 = ~(n17332 ^ n9759);
assign n16074 = ~(n24170 ^ n24085);
assign n26558 = n12196 | n18289;
assign n2024 = n11915 | n21864;
assign n4738 = ~(n7827 ^ n9505);
assign n4897 = ~(n19010 ^ n10212);
assign n11117 = n21171 & n10121;
assign n25218 = ~(n13505 ^ n10895);
assign n7163 = ~(n19608 ^ n15378);
assign n20602 = ~(n26351 ^ n26225);
assign n13938 = n8820 & n13197;
assign n12734 = ~(n14918 ^ n16694);
assign n14452 = n8266 | n7538;
assign n27042 = ~(n10852 ^ n9898);
assign n608 = ~(n20076 ^ n21082);
assign n8090 = ~(n20437 ^ n20151);
assign n18609 = ~(n21287 ^ n9967);
assign n17327 = n23069 | n18153;
assign n93 = n13006 & n20266;
assign n21601 = n11392 | n6654;
assign n4220 = n2576 | n13853;
assign n6242 = ~n17132;
assign n2309 = ~(n1895 | n20972);
assign n12928 = ~n18486;
assign n1027 = ~(n16972 ^ n2895);
assign n17800 = ~(n12655 | n11214);
assign n20578 = ~(n10522 ^ n23024);
assign n13757 = ~(n1333 | n19051);
assign n10769 = n5302 | n19116;
assign n24908 = ~(n6153 ^ n19775);
assign n21722 = n14011 & n17309;
assign n20828 = n10697 & n7075;
assign n6016 = n15302 | n12912;
assign n18718 = n18086 & n24777;
assign n16298 = n5134 & n2830;
assign n9640 = n10392 | n20897;
assign n24976 = n20894 | n18022;
assign n20295 = n1460 & n20783;
assign n23429 = ~(n23889 ^ n20616);
assign n17937 = n6750 & n19058;
assign n14514 = ~n16092;
assign n1636 = ~(n2820 ^ n13973);
assign n18981 = ~n26334;
assign n482 = n25976 & n4292;
assign n11251 = ~(n19033 ^ n17037);
assign n9035 = ~n20192;
assign n11558 = n4667 | n21654;
assign n26329 = n2279 & n21232;
assign n11891 = ~(n20604 | n23331);
assign n26144 = ~n1822;
assign n17607 = ~n22537;
assign n12936 = n8703 & n25290;
assign n2057 = ~n27185;
assign n17522 = n4858 | n6895;
assign n8899 = n9135 | n24194;
assign n12753 = n6572 & n20710;
assign n20617 = n10207 & n20084;
assign n7297 = ~n860;
assign n18964 = n10976 | n9757;
assign n476 = ~(n1689 ^ n20036);
assign n21894 = ~(n13512 ^ n10934);
assign n24526 = n2047 | n1048;
assign n11351 = ~(n27087 ^ n24274);
assign n1628 = n1750 | n21321;
assign n16458 = ~n15564;
assign n11248 = ~n12119;
assign n1976 = ~(n2242 ^ n6449);
assign n4856 = ~(n21843 ^ n14998);
assign n7808 = ~n16025;
assign n13683 = ~(n9115 ^ n18586);
assign n3980 = n11917 & n22193;
assign n13933 = ~(n11919 | n26510);
assign n10004 = n10992 | n25438;
assign n26706 = ~(n13688 ^ n25462);
assign n9136 = n2268 | n19153;
assign n7823 = ~n17180;
assign n13001 = ~(n22363 ^ n11848);
assign n21170 = n3278 & n12710;
assign n552 = ~n15090;
assign n13401 = ~n22771;
assign n2446 = n25620 | n17407;
assign n14257 = ~(n10567 ^ n14421);
assign n19908 = ~(n21774 ^ n20980);
assign n22807 = ~n15654;
assign n23507 = n25599 | n7232;
assign n11974 = ~(n3397 ^ n2889);
assign n24995 = n9945 | n22227;
assign n369 = ~(n8244 ^ n21226);
assign n26802 = n17296 | n21181;
assign n16283 = ~n21385;
assign n5373 = n18290 | n12875;
assign n16321 = ~(n16276 ^ n1348);
assign n16020 = n8079 | n21736;
assign n14948 = n19119 | n21833;
assign n6197 = n4703 | n10926;
assign n9278 = n18561 & n1488;
assign n18085 = n22688 & n3474;
assign n17996 = n26618 & n12658;
assign n11243 = ~n12379;
assign n25361 = n20780 | n7819;
assign n27160 = ~n4196;
assign n25927 = ~(n6724 ^ n22405);
assign n25948 = ~(n11429 ^ n12315);
assign n5912 = n26186 | n1028;
assign n22621 = n24057 & n2910;
assign n563 = ~(n15896 ^ n12295);
assign n9567 = ~(n13925 ^ n21538);
assign n21605 = ~n10614;
assign n25802 = ~(n16825 ^ n7020);
assign n12026 = n11777 & n16644;
assign n20396 = n26264 | n19454;
assign n20734 = ~n22414;
assign n10535 = n11455 | n14870;
assign n24781 = n8922 | n10553;
assign n8530 = ~(n8520 ^ n20506);
assign n11079 = ~n23303;
assign n15434 = n26273 | n7186;
assign n21697 = ~(n5318 | n7439);
assign n620 = n19897 & n26987;
assign n8163 = ~(n25992 ^ n17298);
assign n13665 = n4913 | n17525;
assign n21422 = ~n3246;
assign n14187 = ~(n26426 ^ n12205);
assign n15168 = ~(n19952 | n17444);
assign n8761 = ~(n12863 | n13046);
assign n8846 = ~(n24488 ^ n24996);
assign n11606 = n6758 & n24361;
assign n15478 = n17884 & n24010;
assign n14195 = ~(n1822 ^ n1813);
assign n21846 = ~n4426;
assign n2813 = ~(n20387 ^ n7077);
assign n20685 = n12327 | n14447;
assign n23694 = ~(n8389 ^ n17454);
assign n24159 = n7671 | n8354;
assign n25703 = n17737 | n7744;
assign n16588 = n4963 & n2818;
assign n9893 = ~(n23272 | n14826);
assign n12276 = n23250 & n11209;
assign n8023 = n11652 | n12639;
assign n2490 = ~n24884;
assign n2228 = ~(n5946 ^ n2445);
assign n26087 = n19652 & n22610;
assign n19933 = ~(n14195 ^ n13533);
assign n1940 = n21010 & n22678;
assign n20510 = n25775 | n1397;
assign n10349 = ~(n24450 ^ n14533);
assign n15787 = ~n8380;
assign n12245 = ~(n10964 | n3314);
assign n9406 = ~(n15268 ^ n18737);
assign n21564 = ~n4908;
assign n21250 = n1858 & n24921;
assign n7453 = ~(n2210 | n19863);
assign n24039 = ~(n1812 ^ n3233);
assign n8764 = n19682 | n7041;
assign n23852 = ~(n939 ^ n2283);
assign n27022 = ~(n17345 ^ n11935);
assign n6468 = ~n22772;
assign n15691 = ~(n2723 ^ n5806);
assign n2912 = n22007 | n67;
assign n4559 = ~n21497;
assign n21254 = ~(n9128 ^ n16816);
assign n3842 = ~(n13521 ^ n9420);
assign n9887 = ~(n17447 | n12968);
assign n25718 = n17977 | n11875;
assign n4873 = ~(n17986 ^ n3947);
assign n7185 = n328 | n15490;
assign n7298 = ~(n19326 ^ n4855);
assign n10217 = ~(n4125 ^ n19477);
assign n23000 = ~(n12489 ^ n15753);
assign n4567 = n8146 | n5285;
assign n25267 = ~(n663 ^ n24327);
assign n18146 = n416 & n10981;
assign n17773 = n16259 & n4394;
assign n7392 = ~(n17606 | n24936);
assign n17839 = n5948 | n15415;
assign n10997 = ~n17371;
assign n13967 = ~n23849;
assign n3514 = ~(n17120 | n26510);
assign n27028 = ~(n3161 ^ n11630);
assign n13212 = ~(n22637 | n12837);
assign n1251 = n19898 | n8319;
assign n7631 = n20342 | n4570;
assign n20832 = ~(n2415 ^ n19514);
assign n2762 = n13975 | n14163;
assign n8179 = ~(n22776 ^ n15305);
assign n19018 = ~(n11936 | n9531);
assign n6746 = ~(n9194 ^ n16913);
assign n8879 = n13814 | n5815;
assign n21534 = n17136 & n12662;
assign n1260 = n6551 | n5527;
assign n2653 = ~n4016;
assign n25590 = n11764 & n10349;
assign n22892 = ~(n22549 ^ n16722);
assign n21278 = n7961 & n20561;
assign n11745 = ~n5026;
assign n26793 = ~n9251;
assign n14011 = ~(n9964 ^ n5438);
assign n10664 = n22051 & n22649;
assign n10920 = ~n11592;
assign n9728 = ~(n3271 ^ n2757);
assign n13416 = n26019 | n21407;
assign n2839 = n19961 & n13077;
assign n590 = ~n7304;
assign n6607 = ~(n6243 | n4751);
assign n15216 = ~(n8614 ^ n23895);
assign n1188 = n14495 & n25251;
assign n19773 = n27026 & n351;
assign n20709 = ~(n4079 ^ n2758);
assign n2007 = ~(n3057 | n7054);
assign n1755 = n24513 & n845;
assign n24042 = ~(n12785 ^ n21762);
assign n18925 = ~n7725;
assign n9628 = ~(n23126 | n17369);
assign n20912 = n23454 | n8647;
assign n13530 = ~n14489;
assign n2217 = ~(n1739 ^ n4913);
assign n12351 = ~(n18621 ^ n4957);
assign n10407 = ~(n16362 ^ n6296);
assign n13646 = ~(n2314 | n5407);
assign n8653 = ~(n21143 ^ n1842);
assign n19966 = n16386 | n5739;
assign n2104 = ~(n9693 | n12457);
assign n16787 = ~(n23974 | n8309);
assign n14778 = ~(n17906 | n4372);
assign n4396 = ~(n12869 ^ n822);
assign n19338 = ~(n8952 ^ n25240);
assign n7029 = n26151 & n3221;
assign n312 = ~n16906;
assign n23851 = ~(n17744 ^ n19033);
assign n10995 = ~n18006;
assign n25067 = ~n22309;
assign n19471 = ~(n19618 | n18707);
assign n13602 = ~(n562 ^ n8219);
assign n14144 = n22040 | n24707;
assign n13759 = ~(n9108 ^ n8873);
assign n24742 = ~(n20102 ^ n23751);
assign n21299 = ~(n12733 ^ n25972);
assign n4146 = ~(n4046 ^ n20668);
assign n8976 = n21644 | n4426;
assign n18605 = n1273 | n1070;
assign n7150 = n24851 | n10711;
assign n25426 = ~(n13097 ^ n17225);
assign n24058 = ~n19981;
assign n17859 = ~(n3914 ^ n23962);
assign n8373 = n710 | n8398;
assign n21930 = ~n15240;
assign n14327 = ~n3920;
assign n19085 = ~n6712;
assign n20220 = ~(n20777 ^ n2461);
assign n13293 = ~(n26464 ^ n20057);
assign n24506 = ~(n24323 ^ n8581);
assign n13616 = n3439 | n1995;
assign n17658 = ~n11329;
assign n14446 = ~(n11989 ^ n3526);
assign n26533 = n21847 | n4980;
assign n6551 = ~(n19160 ^ n14835);
assign n2966 = ~(n13627 ^ n4847);
assign n10827 = n26404 | n9751;
assign n3601 = ~n16496;
assign n15313 = ~n14314;
assign n3575 = n8448 & n15892;
assign n26098 = ~(n2029 ^ n13776);
assign n11652 = ~n9934;
assign n5430 = ~(n13878 ^ n2942);
assign n20030 = ~n5340;
assign n2068 = n14953 | n1581;
assign n5007 = ~(n8232 | n20749);
assign n10273 = n24653 & n10746;
assign n24621 = n17959 | n25221;
assign n12550 = ~n20499;
assign n26173 = n15878 & n21011;
assign n7849 = ~(n1009 | n18145);
assign n20906 = ~(n7855 ^ n20161);
assign n17401 = n5796 & n25856;
assign n11034 = ~(n2994 ^ n25872);
assign n5533 = n2432 | n20633;
assign n1926 = n23916 & n6827;
assign n7781 = ~(n4887 ^ n6298);
assign n12869 = ~n17186;
assign n21298 = ~(n12934 ^ n6349);
assign n3025 = ~(n5624 | n13490);
assign n4268 = n18368 & n12428;
assign n23502 = ~(n11302 | n17213);
assign n25010 = n21527 | n20509;
assign n18767 = ~n2499;
assign n8040 = n20345 | n9320;
assign n25764 = ~n19741;
assign n14849 = ~(n632 ^ n23955);
assign n1641 = n14000 | n7816;
assign n16631 = n9365 | n13543;
assign n2545 = ~(n27041 ^ n3582);
assign n19634 = ~n4812;
assign n20476 = ~(n26876 | n3730);
assign n2322 = ~n10728;
assign n12720 = ~n24919;
assign n10893 = ~(n17995 | n4222);
assign n13554 = n294 | n23020;
assign n884 = n26510 | n11246;
assign n1902 = n24375 | n9942;
assign n22454 = ~n9372;
assign n23343 = n5790 & n14398;
assign n7189 = ~(n2151 | n26425);
assign n4433 = n574 & n24689;
assign n21333 = n2979 | n24764;
assign n11725 = ~(n3173 | n25393);
assign n18633 = n4625 & n9523;
assign n1962 = n27012 | n1737;
assign n19619 = ~(n839 | n15709);
assign n3404 = n13292 | n21911;
assign n26855 = n19076 | n3903;
assign n21758 = n4351 & n25153;
assign n23037 = n23227 & n16315;
assign n18077 = ~(n11314 | n7689);
assign n19503 = n9157 | n23931;
assign n10979 = ~(n6353 ^ n12391);
assign n25396 = n26628 & n26960;
assign n5080 = n23658 | n17121;
assign n12405 = ~n2841;
assign n2074 = n23416 | n18597;
assign n14725 = ~n2394;
assign n11146 = ~n26713;
assign n23516 = n14066 | n23432;
assign n20088 = ~(n9490 | n23693);
assign n26935 = ~(n26837 ^ n13251);
assign n1994 = ~n7652;
assign n16030 = ~(n5960 | n13490);
assign n5209 = n17965 & n1744;
assign n2257 = ~(n6841 | n8439);
assign n25981 = n21606 & n26422;
assign n13690 = n23573 | n6637;
assign n246 = ~n626;
assign n27092 = ~(n9940 | n8013);
assign n11438 = ~(n15432 | n18883);
assign n6391 = n15905 & n27118;
assign n9384 = ~(n9497 | n23751);
assign n16942 = ~n23220;
assign n14302 = ~(n12042 | n11308);
assign n13389 = ~n7692;
assign n21576 = n11460 & n27056;
assign n10246 = ~(n655 ^ n6397);
assign n6626 = ~(n22198 ^ n5337);
assign n6876 = ~(n3373 ^ n2892);
assign n13839 = n24355 & n21935;
assign n15435 = ~(n9058 ^ n20286);
assign n7055 = ~(n15220 | n3846);
assign n302 = ~n23277;
assign n6874 = n3170 & n23699;
assign n2070 = n18658 & n15035;
assign n19561 = n17861 & n24190;
assign n26082 = n25855 & n26461;
assign n26949 = n13783 & n13590;
assign n20392 = n2621 & n2364;
assign n14353 = ~(n25020 ^ n14607);
assign n21048 = n1815 | n26735;
assign n26460 = n5703;
assign n11501 = ~n18229;
assign n3182 = n2384 | n18873;
assign n13776 = ~(n18765 ^ n21975);
assign n9589 = n24462 | n6748;
assign n7932 = n1497 & n4184;
assign n20216 = ~n8540;
assign n20793 = n19531 | n26872;
assign n25728 = n10761 | n3985;
assign n22228 = n12955 | n5220;
assign n25339 = n7923 | n5998;
assign n23299 = ~(n16687 ^ n6449);
assign n3787 = n18192 | n9473;
assign n12462 = n6650 | n11260;
assign n6195 = ~n18630;
assign n3683 = n26738 | n6666;
assign n470 = ~(n11136 ^ n6435);
assign n16086 = n7092 & n24486;
assign n8852 = n11425 | n9967;
assign n809 = ~(n23077 ^ n12266);
assign n6979 = n8275 & n7220;
assign n7114 = n21450 | n24821;
assign n11874 = n682 | n14811;
assign n11645 = n3853 | n23372;
assign n242 = ~(n5477 ^ n6433);
assign n19493 = ~n16261;
assign n4140 = n26564 & n7471;
assign n12916 = ~(n20065 ^ n2184);
assign n22557 = ~(n9354 ^ n3722);
assign n4449 = ~(n21537 ^ n18274);
assign n15063 = n22261 | n10117;
assign n14524 = n19494 | n2387;
assign n4703 = ~(n26536 | n19607);
assign n19651 = n4887 | n5045;
assign n25887 = ~(n6122 ^ n23200);
assign n21083 = ~n8399;
assign n13035 = ~n17982;
assign n18994 = ~n5582;
assign n23735 = ~(n2320 ^ n26053);
assign n4771 = ~(n3472 | n15790);
assign n9870 = n11542 | n7057;
assign n2462 = ~n25617;
assign n22941 = n11171 | n26026;
assign n10540 = ~(n4430 ^ n3218);
assign n3630 = ~(n25074 ^ n12956);
assign n18399 = ~(n10666 ^ n19856);
assign n25552 = n16105 & n6118;
assign n11789 = n8094 & n11051;
assign n1394 = ~(n10611 ^ n24879);
assign n20010 = n18203 | n15910;
assign n12937 = n6110 & n16990;
assign n26221 = n1783 | n2587;
assign n12733 = ~(n3028 ^ n13965);
assign n5811 = n8614 & n21162;
assign n18522 = ~(n22554 ^ n25381);
assign n21610 = n2743 & n1584;
assign n1386 = n13032 ^ n12188;
assign n7027 = ~(n1777 | n4812);
assign n19014 = n4039 | n8742;
assign n1470 = ~(n15041 ^ n26553);
assign n11825 = n21936 | n46;
assign n17698 = n10191 | n26463;
assign n8478 = n13370 | n25644;
assign n3012 = ~(n3071 ^ n1305);
assign n805 = n23090 & n3353;
assign n2848 = n13909 | n520;
assign n15863 = n23441 | n9926;
assign n4775 = ~(n25187 ^ n11619);
assign n17149 = ~(n15073 ^ n19814);
assign n16593 = ~(n14114 | n14111);
assign n4880 = n16033 & n7121;
assign n3341 = n1969 & n20729;
assign n2730 = n1689 | n9450;
assign n27049 = ~(n20077 ^ n19494);
assign n2401 = ~(n4706 ^ n905);
assign n12394 = n24461 | n26095;
assign n10308 = n6845 & n4211;
assign n16650 = n1138 | n17000;
assign n9690 = n9110 | n25442;
assign n26500 = n18521 | n3802;
assign n12807 = n11445 & n25587;
assign n24946 = n3013 | n19436;
assign n4958 = ~(n2718 ^ n9291);
assign n1645 = n19675 & n24173;
assign n66 = n6677 | n25026;
assign n25722 = n24650 | n13033;
assign n3362 = n25524 | n16234;
assign n2268 = ~n12593;
assign n16157 = n15827 | n15073;
assign n9824 = ~(n15251 | n4422);
assign n9921 = n19321 | n19737;
assign n803 = ~(n19311 ^ n992);
assign n6492 = ~(n24789 ^ n19252);
assign n20456 = n18155 & n16027;
assign n9827 = ~(n8142 ^ n22835);
assign n8330 = ~(n6631 ^ n7339);
assign n16534 = ~(n13577 | n12341);
assign n18965 = ~(n19905 ^ n2547);
assign n22507 = ~n19425;
assign n8077 = ~n9240;
assign n5674 = ~(n6041 ^ n14550);
assign n11235 = ~(n3401 ^ n1249);
assign n7485 = n16635 | n24450;
assign n22790 = n25916 | n18570;
assign n4789 = n5029 & n23263;
assign n9190 = ~(n13912 ^ n11980);
assign n18106 = n8 | n19678;
assign n16839 = ~(n21713 ^ n26835);
assign n13803 = ~n8479;
assign n13727 = ~(n9974 ^ n24138);
assign n16054 = ~(n5542 ^ n22372);
assign n4148 = ~(n23039 ^ n4590);
assign n2253 = ~(n21508 ^ n10183);
assign n17527 = n17018 | n26968;
assign n25559 = n8678 | n3882;
assign n14757 = ~n22864;
assign n4482 = ~(n8456 ^ n5605);
assign n14383 = ~(n22247 | n21126);
assign n1350 = ~(n16970 ^ n11287);
assign n27024 = n9729 & n4985;
assign n20755 = ~(n1149 ^ n8349);
assign n22522 = n25119 | n3719;
assign n9773 = n20245 | n8006;
assign n753 = n20479 | n9222;
assign n2911 = ~n19285;
assign n22307 = n22565 & n5656;
assign n23316 = n20040 & n16555;
assign n26519 = n5400 & n9512;
assign n7378 = ~(n2659 | n1941);
assign n12326 = n725 | n24804;
assign n24921 = n4279 | n13566;
assign n14461 = n1515 & n19207;
assign n9081 = ~(n1689 | n17095);
assign n20234 = n5075 | n25768;
assign n18028 = ~(n23359 | n15454);
assign n6699 = n26998 & n3592;
assign n17072 = n2104 | n10609;
assign n14767 = ~(n18015 ^ n3027);
assign n10280 = ~(n23996 ^ n5685);
assign n733 = ~n5704;
assign n17071 = ~(n19048 ^ n25007);
assign n26421 = ~n2383;
assign n21263 = n12211;
assign n7789 = n9583 | n15566;
assign n13837 = ~(n22342 ^ n16993);
assign n1879 = n23304 & n1465;
assign n9167 = n21481 | n14867;
assign n4209 = n5230 | n9682;
assign n21831 = n9924 | n26216;
assign n586 = ~n3614;
assign n15609 = n12636 | n4633;
assign n991 = n778 | n23769;
assign n5515 = n19630 | n3361;
assign n14710 = ~n22764;
assign n1119 = ~(n18605 ^ n24144);
assign n10194 = n11100 & n22513;
assign n6650 = ~(n25781 | n2155);
assign n15894 = ~(n12019 ^ n17585);
assign n6764 = ~n15780;
assign n18173 = ~n6659;
assign n18056 = n17160 & n5927;
assign n3196 = n13882 & n8058;
assign n4930 = ~(n11309 ^ n26452);
assign n1907 = ~(n13951 ^ n12507);
assign n26567 = n13497 | n22631;
assign n21253 = ~(n17124 ^ n15979);
assign n15305 = n27 | n25973;
assign n9864 = ~(n4256 ^ n20946);
assign n9667 = n4383 | n3808;
assign n26330 = ~(n21544 ^ n18924);
assign n4269 = ~(n23819 ^ n25370);
assign n27036 = ~(n5156 ^ n13460);
assign n797 = n1103 | n18389;
assign n18524 = n19105 & n9010;
assign n333 = ~n2568;
assign n7495 = n4893 | n21451;
assign n14088 = n405 | n13842;
assign n25885 = n23327 & n25945;
assign n12206 = n1680 | n479;
assign n14167 = n11536 & n8684;
assign n23380 = n21599 & n26324;
assign n3116 = ~n8638;
assign n16751 = ~n16426;
assign n21064 = n600 & n12497;
assign n14490 = n19551 | n2705;
assign n9686 = ~(n23580 ^ n26350);
assign n18879 = n7338 | n22355;
assign n21518 = n24649 | n14719;
assign n6960 = n13061 | n23552;
assign n14041 = n17394 & n9727;
assign n16531 = ~n4514;
assign n20100 = ~n8687;
assign n5196 = n16485 & n14745;
assign n14553 = n3139 | n23037;
assign n18109 = n18775 | n20825;
assign n13447 = ~(n20950 ^ n15376);
assign n4985 = n57 | n7539;
assign n14479 = ~(n5521 | n1803);
assign n15027 = n15602 | n3690;
assign n24388 = n23832 & n19238;
assign n4185 = ~n23939;
assign n1373 = ~(n27175 | n5474);
assign n12062 = n19006 | n22180;
assign n23223 = n12612 | n14048;
assign n2647 = n22148 & n10566;
assign n9276 = n11368 & n8939;
assign n24167 = ~(n24817 ^ n8896);
assign n15526 = n12114 & n25796;
assign n9232 = n23895 | n8491;
assign n25078 = n17558 | n26403;
assign n14930 = n16654 & n7824;
assign n12610 = ~(n15023 ^ n13113);
assign n11868 = n1373 | n1080;
assign n23488 = ~(n21817 ^ n9057);
assign n15282 = ~(n3798 ^ n23140);
assign n26907 = ~(n18079 | n21460);
assign n2225 = n6499 | n5002;
assign n10078 = ~(n18792 | n15417);
assign n25672 = n24310 | n16116;
assign n12376 = n19899 | n18608;
assign n15496 = ~(n26737 ^ n12975);
assign n15249 = ~(n7457 | n32);
assign n12761 = ~(n1685 ^ n3785);
assign n21229 = ~(n9888 | n3827);
assign n18896 = n18274 & n24202;
assign n6325 = n10422 & n19383;
assign n15507 = ~n12236;
assign n16092 = ~(n14197 ^ n12808);
assign n4666 = n5612 | n3144;
assign n3132 = ~(n2941 ^ n655);
assign n12769 = ~n19219;
assign n6199 = ~n16423;
assign n5665 = n19992 & n3427;
assign n4447 = n19640 | n13916;
assign n7790 = n17234 | n7993;
assign n51 = n25943 & n12118;
assign n7283 = n19616 | n13359;
assign n23628 = ~(n24357 ^ n16346);
assign n19498 = n15348 & n9722;
assign n6974 = ~(n4753 ^ n3366);
assign n19376 = ~(n23061 ^ n7305);
assign n19693 = n3685 | n19821;
assign n16662 = ~(n7019 ^ n10665);
assign n17064 = ~(n20987 ^ n7635);
assign n21772 = ~n8763;
assign n25449 = ~(n8230 ^ n21024);
assign n13737 = ~n23170;
assign n13303 = ~(n17374 ^ n9006);
assign n6487 = n24168 | n1617;
assign n20275 = ~n16832;
assign n4600 = n8384 & n11067;
assign n18894 = ~(n16830 | n20032);
assign n4296 = n13402 & n20322;
assign n5054 = ~(n23290 | n20185);
assign n21859 = ~(n20575 ^ n23725);
assign n22184 = n8098 | n22344;
assign n13874 = ~(n22183 | n25595);
assign n9442 = ~(n8952 ^ n7841);
assign n1230 = ~n13123;
assign n24947 = ~n3909;
assign n11116 = ~(n7304 ^ n10095);
assign n17429 = n27052 | n4944;
assign n23655 = ~(n16831 ^ n10582);
assign n885 = ~(n7593 ^ n5101);
assign n3973 = ~(n12592 ^ n10267);
assign n5701 = ~(n16150 ^ n14010);
assign n16073 = ~(n22012 ^ n8688);
assign n11694 = ~n7008;
assign n15047 = n18613 | n5526;
assign n26317 = ~(n24858 ^ n18763);
assign n27139 = ~(n18795 ^ n18854);
assign n17559 = ~n26098;
assign n22153 = ~(n21836 ^ n18020);
assign n21464 = n12132 | n239;
assign n18816 = n21895 & n4303;
assign n15112 = n14995 | n11430;
assign n7720 = n6601 | n3600;
assign n5957 = n24136 & n18806;
assign n10111 = ~(n10566 ^ n16108);
assign n25958 = ~(n16609 ^ n7949);
assign n13422 = ~n25586;
assign n7627 = ~n15975;
assign n13357 = ~n5386;
assign n16176 = ~(n130 ^ n5247);
assign n16069 = n25037 | n9183;
assign n20471 = ~(n2145 | n5521);
assign n9909 = ~n20361;
assign n957 = ~(n7957 ^ n12412);
assign n12335 = n26158 & n8262;
assign n282 = n1235 & n23700;
assign n7582 = n709 & n3337;
assign n7098 = n3522 & n25338;
assign n26944 = n7434 & n23025;
assign n18587 = ~n13885;
assign n19039 = ~(n16094 ^ n26660);
assign n26247 = n21777 & n4685;
assign n3384 = n2420 & n23807;
assign n13197 = ~(n1606 ^ n13607);
assign n8544 = n17252 | n22338;
assign n14681 = n1283 & n2427;
assign n14929 = n8180 | n5734;
assign n4670 = ~(n21285 ^ n12907);
assign n6017 = n15361 | n3044;
assign n2532 = ~(n5244 ^ n255);
assign n516 = n10796 & n15653;
assign n6955 = n17617 | n16426;
assign n8797 = n16427 & n17888;
assign n14544 = ~(n10664 ^ n14606);
assign n7334 = n8835 | n19544;
assign n6854 = n26892 | n17200;
assign n1178 = ~(n7072 | n9851);
assign n11710 = ~(n6322 ^ n16422);
assign n25133 = ~(n4637 ^ n17074);
assign n14209 = n8459 & n404;
assign n24819 = ~(n21469 | n16017);
assign n20813 = n9716 | n1495;
assign n22693 = n21373 | n13182;
assign n10222 = ~(n148 ^ n2113);
assign n20050 = n13256 & n25780;
assign n18148 = ~(n15091 ^ n26693);
assign n728 = ~n21155;
assign n11104 = ~(n12470 ^ n11455);
assign n6520 = n24377 & n20514;
assign n9759 = ~(n23835 ^ n2950);
assign n15291 = ~(n11609 ^ n26386);
assign n1289 = ~(n10357 | n20284);
assign n19738 = ~n10228;
assign n14029 = n24490 & n3930;
assign n9227 = ~n21723;
assign n13272 = n23156 | n26813;
assign n4503 = ~(n23290 | n15742);
assign n8739 = ~n23755;
assign n6847 = ~(n18824 ^ n2596);
assign n19206 = n1958 | n1187;
assign n11144 = ~n18105;
assign n396 = ~n9396;
assign n7577 = n6659 | n20384;
assign n18872 = n21984 & n6255;
assign n11765 = ~(n21850 ^ n17351);
assign n9183 = n9573 & n17480;
assign n1956 = ~n337;
assign n25006 = ~(n26148 ^ n26323);
assign n19780 = ~(n7165 ^ n16099);
assign n9807 = ~(n6925 ^ n10505);
assign n12644 = ~n18672;
assign n7923 = ~n9380;
assign n9465 = n7237 & n15087;
assign n26256 = n25333 & n3847;
assign n22606 = ~(n7566 | n586);
assign n29 = ~(n16738 | n12860);
assign n12847 = n3460 & n11452;
assign n21165 = n13719 | n6710;
assign n20366 = ~(n23381 ^ n21417);
assign n10069 = n9697 & n19251;
assign n14339 = ~(n14710 | n2416);
assign n22374 = n709 | n3337;
assign n13096 = ~(n9334 ^ n13045);
assign n16750 = ~n20072;
assign n14198 = ~(n4080 ^ n16394);
assign n11602 = n3977 | n4136;
assign n14036 = ~(n15526 ^ n4382);
assign n15126 = ~(n20254 ^ n14687);
assign n16051 = ~(n23837 ^ n22092);
assign n4469 = n19838 | n11083;
assign n14113 = ~(n14923 | n12050);
assign n20775 = ~(n5976 | n2694);
assign n13295 = n206 & n13020;
assign n18312 = ~(n18068 ^ n20826);
assign n14968 = ~(n18496 ^ n25331);
assign n637 = ~(n11108 ^ n18988);
assign n21969 = n12417;
assign n1031 = n1186 | n12317;
assign n6619 = n31 | n16065;
assign n5716 = ~n20958;
assign n3039 = n22179 | n1944;
assign n4862 = ~n20336;
assign n22109 = n8984 & n62;
assign n26814 = ~(n7974 | n8399);
assign n15994 = n12925 & n8919;
assign n25341 = n26580 | n5428;
assign n24636 = ~(n12796 ^ n21809);
assign n257 = n1270 & n4428;
assign n4486 = ~(n19277 | n23430);
assign n7612 = n16495 & n12401;
assign n14165 = n8433 & n2292;
assign n25928 = ~(n22215 | n26350);
assign n13519 = n16709 | n22771;
assign n27152 = n3155 | n14697;
assign n25621 = ~(n16910 | n15975);
assign n10381 = ~(n27199 | n4003);
assign n16379 = ~(n8460 ^ n10064);
assign n22555 = n23298 | n19131;
assign n9209 = n12341 | n5727;
assign n19613 = ~(n187 | n10549);
assign n4121 = ~(n14680 ^ n20359);
assign n24961 = ~(n7480 ^ n13347);
assign n19813 = ~(n21876 | n18121);
assign n11751 = ~(n19049 ^ n14097);
assign n20199 = ~(n8052 ^ n24618);
assign n8429 = n10499 | n2248;
assign n2842 = ~n6678;
assign n14723 = ~(n6954 ^ n17730);
assign n20076 = ~(n16891 ^ n21602);
assign n11699 = n20334 | n13493;
assign n7498 = n8213 & n26657;
assign n10733 = ~(n2291 ^ n25629);
assign n27079 = ~(n9153 ^ n11053);
assign n7451 = n18516 | n26714;
assign n6281 = ~(n26691 ^ n7563);
assign n4943 = ~(n11088 ^ n22843);
assign n13498 = ~n14299;
assign n11336 = ~(n14346 ^ n26797);
assign n26442 = ~(n21929 | n9575);
assign n2041 = ~(n648 ^ n7271);
assign n13511 = n8163 ^ n13752;
assign n3397 = ~n1455;
assign n22077 = ~n15894;
assign n23720 = ~n822;
assign n3612 = n20009 & n23980;
assign n999 = n4602 | n8250;
assign n25508 = n24949 | n789;
assign n18190 = ~(n6372 | n11784);
assign n273 = ~(n12652 ^ n21309);
assign n3217 = n6993 | n15706;
assign n25233 = n21350 | n18049;
assign n13594 = n5934 & n25517;
assign n1728 = ~n21956;
assign n21727 = n4502 | n16618;
assign n13758 = n16678 | n25384;
assign n14455 = ~n13521;
assign n25190 = ~(n18585 | n12993);
assign n7744 = n24505 & n12460;
assign n5829 = n16609 & n22666;
assign n11134 = ~(n13147 ^ n12730);
assign n10633 = ~(n3562 ^ n19694);
assign n23284 = ~(n3846 ^ n15220);
assign n9770 = ~n9222;
assign n20399 = ~(n25846 | n4800);
assign n2337 = n6557 & n17673;
assign n10469 = ~n4245;
assign n18570 = ~(n22378 ^ n24630);
assign n11337 = ~n11070;
assign n3898 = n18476 & n27042;
assign n12216 = ~(n23083 ^ n8724);
assign n21513 = ~(n25036 ^ n9983);
assign n16234 = ~n3959;
assign n25461 = ~n2191;
assign n12838 = ~(n17333 ^ n19247);
assign n1341 = n21674 | n5090;
assign n8435 = n13459 | n17183;
assign n10770 = ~(n14408 | n3486);
assign n9235 = n21538 | n11335;
assign n6315 = n11378 ^ n3515;
assign n20069 = ~(n8124 ^ n24100);
assign n12738 = n329 | n21735;
assign n21379 = n25854 | n9379;
assign n8228 = ~(n13490 | n7751);
assign n21761 = n4752 | n7674;
assign n20156 = n6273 | n21206;
assign n6101 = n10687 | n5910;
assign n21055 = ~n13031;
assign n4385 = n8928 & n9231;
assign n3365 = ~n17003;
assign n14789 = n658 & n25339;
assign n18952 = ~(n20205 | n2218);
assign n19925 = ~(n8774 ^ n22198);
assign n16491 = n6537 & n21311;
assign n20928 = n7770 & n13413;
assign n4888 = n13681 | n17307;
assign n24514 = ~(n15127 ^ n3846);
assign n19892 = n976 | n17050;
assign n17752 = n25299 & n17907;
assign n8111 = ~(n2858 ^ n5521);
assign n9774 = n15939 | n18927;
assign n24459 = n3275 | n2800;
assign n17004 = n11113 & n5917;
assign n3176 = ~(n16291 ^ n13044);
assign n6032 = n12035 & n2609;
assign n11147 = ~(n17826 | n10554);
assign n421 = ~(n4469 | n5987);
assign n16638 = ~(n9912 ^ n7547);
assign n20008 = ~(n11615 ^ n8052);
assign n23645 = ~n7460;
assign n3119 = n891 & n17364;
assign n11583 = ~n20151;
assign n17444 = ~n9219;
assign n22686 = n18625 | n17249;
assign n12142 = n6100 & n19965;
assign n17247 = n19743 & n2683;
assign n6124 = ~(n3577 | n25171);
assign n12438 = ~(n851 ^ n5255);
assign n11075 = ~(n21749 | n26744);
assign n23008 = ~n20296;
assign n1406 = ~n20235;
assign n12540 = ~(n10726 ^ n23481);
assign n10172 = n9424 | n15413;
assign n21112 = n19144 | n9170;
assign n7553 = n26722 & n15074;
assign n20194 = n2792 | n21113;
assign n26534 = n20134 | n9192;
assign n16060 = ~(n25219 ^ n21425);
assign n19627 = ~(n7184 ^ n23107);
assign n18203 = ~n19245;
assign n16533 = n8231 & n13565;
assign n22766 = ~n8774;
assign n7408 = ~(n7029 ^ n18372);
assign n4527 = n10837 | n23890;
assign n24712 = ~(n26235 ^ n22439);
assign n21419 = n8334 | n19946;
assign n1527 = ~(n20683 ^ n17882);
assign n10454 = ~(n23590 ^ n510);
assign n20134 = ~n5337;
assign n20285 = ~(n4626 ^ n604);
assign n6836 = n17256 | n14693;
assign n13496 = n7586 | n2467;
assign n16602 = ~n6422;
assign n18728 = ~(n17052 | n439);
assign n12298 = n22309 & n10711;
assign n6157 = n24060 & n11345;
assign n1008 = ~(n9468 ^ n15241);
assign n1149 = n20865 | n517;
assign n14798 = n22987 | n13357;
assign n8849 = ~(n26468 ^ n12838);
assign n3435 = n26825 & n1271;
assign n26975 = n6023 | n20649;
assign n149 = n19462 | n8131;
assign n7260 = ~(n25367 ^ n20163);
assign n19149 = ~n3366;
assign n11863 = n3268 & n14062;
assign n8240 = ~(n1720 ^ n6543);
assign n6062 = ~(n8827 ^ n1881);
assign n27033 = ~(n4199 | n11118);
assign n8210 = ~n619;
assign n22120 = n15891 ^ n9493;
assign n7223 = ~n20291;
assign n20683 = n24174 & n22145;
assign n17621 = n22094 & n21920;
assign n15625 = ~(n6222 ^ n9744);
assign n15423 = ~n5416;
assign n8751 = ~(n10228 ^ n11473);
assign n13193 = n25151 & n214;
assign n24645 = ~n4834;
assign n10565 = ~(n19975 ^ n3121);
assign n25033 = ~(n13360 ^ n13124);
assign n4842 = n15604 | n18001;
assign n16423 = ~(n20499 ^ n18689);
assign n19492 = n10894 | n11484;
assign n16365 = n878 & n2123;
assign n1850 = ~n10970;
assign n4635 = n18789 | n1535;
assign n4225 = ~(n14974 ^ n11246);
assign n11511 = n975 | n25618;
assign n776 = ~n18880;
assign n13467 = n26493 & n4842;
assign n7802 = ~(n20544 ^ n12071);
assign n24315 = ~(n17760 ^ n25373);
assign n23445 = n21232 & n7471;
assign n7883 = n13286 | n26080;
assign n16255 = n19449 & n22757;
assign n15839 = ~(n26399 ^ n3710);
assign n11136 = ~(n9545 ^ n2232);
assign n3729 = n2644 & n289;
assign n3734 = n1278 & n22695;
assign n11202 = n15293 | n24644;
assign n22413 = ~(n12646 ^ n19725);
assign n26402 = n13734 & n6019;
assign n3375 = n18013 | n12926;
assign n11762 = n4227 | n11050;
assign n10807 = ~n3827;
assign n19510 = n5822 | n7963;
assign n11842 = ~(n16857 ^ n26131);
assign n25216 = n19506 & n1897;
assign n6750 = ~n16439;
assign n6890 = n2380 | n25253;
assign n15674 = n23406 | n20962;
assign n23559 = ~(n19601 ^ n10800);
assign n7967 = ~(n8526 | n12232);
assign n6121 = ~(n17183 ^ n20036);
assign n12338 = n12085 & n9277;
assign n9661 = ~(n11924 | n10986);
assign n13705 = n24769 & n25401;
assign n25388 = n24008 | n5;
assign n331 = ~(n1045 ^ n1603);
assign n26678 = ~(n658 | n21095);
assign n4587 = n22631 | n1167;
assign n18706 = n3567 & n8137;
assign n3464 = n5355 & n5000;
assign n15571 = n5140 | n20796;
assign n26934 = ~(n7102 ^ n12249);
assign n20866 = n18485 | n19228;
assign n565 = ~(n22379 ^ n767);
assign n2488 = ~(n19989 ^ n18639);
assign n5481 = n18808 & n1874;
assign n19120 = ~(n15696 ^ n23545);
assign n17710 = ~(n21539 | n6200);
assign n9895 = n13855 | n1246;
assign n15554 = n25041 | n16205;
assign n5188 = n18573 | n15830;
assign n18368 = n21386 | n21287;
assign n3227 = n9039 | n12286;
assign n3092 = ~(n17940 | n111);
assign n14190 = ~(n9224 ^ n21449);
assign n1629 = ~(n7413 ^ n15285);
assign n1456 = n11302 | n19876;
assign n11862 = n23709 & n14268;
assign n3442 = n11370 | n3837;
assign n6906 = n13584 | n1830;
assign n3588 = ~(n15892 ^ n3739);
assign n20549 = n27086 & n5504;
assign n17526 = ~(n4435 ^ n8533);
assign n16236 = ~(n19540 | n25637);
assign n4613 = ~(n13214 ^ n19144);
assign n16017 = ~(n9713 | n1471);
assign n398 = ~(n10117 ^ n23250);
assign n16410 = n4884 & n8091;
assign n3603 = ~(n12061 ^ n1887);
assign n7618 = n14293 | n20409;
assign n18936 = n15294 & n15270;
assign n12786 = n25527 | n16171;
assign n23137 = n14569 | n20658;
assign n23634 = ~n25504;
assign n18531 = ~(n2409 ^ n14071);
assign n16006 = n5965 & n9200;
assign n472 = ~n4858;
assign n22675 = ~(n9655 | n20946);
assign n16717 = ~(n24048 | n19683);
assign n19569 = ~(n1199 ^ n11698);
assign n9818 = ~(n20359 | n23704);
assign n1584 = ~n10949;
assign n367 = n25914 & n198;
assign n11261 = ~(n18796 ^ n2667);
assign n7343 = ~n16794;
assign n24274 = ~(n18880 ^ n2978);
assign n3355 = ~(n22247 ^ n21126);
assign n21091 = n2252 | n22020;
assign n14690 = n6218 | n7669;
assign n1678 = n24367 | n15991;
assign n3493 = n16267 | n4299;
assign n12363 = ~(n3967 | n8338);
assign n24131 = ~n21848;
assign n18868 = n5672 & n21086;
assign n5587 = ~(n17587 ^ n25958);
assign n25535 = n12272 | n16709;
assign n14856 = ~n22274;
assign n7703 = ~(n6727 ^ n5182);
assign n14094 = ~n25781;
assign n18583 = ~(n6409 ^ n4477);
assign n25352 = n19634 & n27184;
assign n26482 = n13944 & n23871;
assign n6724 = ~n19161;
assign n11065 = n13689 | n19004;
assign n16117 = ~(n2089 ^ n25094);
assign n21914 = n13976 ^ n10250;
assign n19157 = ~n15077;
assign n26948 = n25269 | n23641;
assign n22659 = ~n13150;
assign n9615 = ~n25924;
assign n18008 = ~n26167;
assign n26334 = ~(n9061 ^ n314);
assign n8611 = n7893 | n19701;
assign n15862 = n21023 & n19537;
assign n8808 = n6347 & n10589;
assign n754 = n13662 & n7589;
assign n10119 = ~(n12673 | n25220);
assign n21535 = n15411 | n1079;
assign n9472 = n6912 | n18488;
assign n20635 = n19662 | n5930;
assign n5409 = ~(n5329 ^ n1);
assign n13816 = n22631 | n21078;
assign n23113 = n4137 & n7789;
assign n9593 = ~(n726 ^ n25749);
assign n1108 = ~(n3770 | n24801);
assign n19372 = ~(n12289 ^ n12892);
assign n22569 = ~(n25228 ^ n5337);
assign n19029 = n27043 | n27170;
assign n18121 = ~(n6919 | n1755);
assign n15782 = n22290 | n12878;
assign n9122 = n8698 & n22788;
assign n8510 = ~(n12190 ^ n21368);
assign n21679 = ~(n2191 ^ n26053);
assign n22096 = n25707 | n10510;
assign n15739 = ~(n24495 ^ n22764);
assign n5243 = ~(n6399 ^ n14738);
assign n23814 = ~n22625;
assign n16545 = n6313 | n25529;
assign n11285 = ~(n4512 ^ n24201);
assign n10785 = ~(n11729 ^ n10718);
assign n11936 = ~(n9250 ^ n885);
assign n1993 = ~(n5213 ^ n4812);
assign n8235 = ~(n9627 | n8712);
assign n14995 = ~(n25021 | n11841);
assign n12461 = ~(n14820 ^ n6257);
assign n17719 = n19511 | n8857;
assign n25991 = n8316 & n18284;
assign n16939 = n7640 & n3509;
assign n5989 = ~(n2565 | n25490);
assign n10471 = n2226 & n17146;
assign n23691 = ~(n8661 ^ n24786);
assign n7134 = ~(n22296 ^ n4936);
assign n13573 = ~(n10017 ^ n20349);
assign n25253 = n5534 & n19693;
assign n2619 = ~(n10149 ^ n12047);
assign n122 = ~(n8964 | n11764);
assign n3572 = n4565 & n2600;
assign n21858 = ~(n14808 ^ n25358);
assign n5586 = n710 & n8398;
assign n17141 = ~n9440;
assign n4826 = ~(n25475 ^ n23697);
assign n7254 = ~n5752;
assign n20939 = ~n18358;
assign n20189 = n5302 | n19484;
assign n20370 = n4957 | n22688;
assign n12024 = ~(n6814 | n10763);
assign n10293 = n24572 | n95;
assign n19415 = n15916 & n392;
assign n11990 = n15466 & n3969;
assign n15187 = n24134 | n8164;
assign n21586 = ~(n12018 ^ n19453);
assign n10435 = n8513 & n10709;
assign n21442 = ~n21458;
assign n21808 = n13924 | n22449;
assign n7241 = n11100 | n22513;
assign n2558 = n7208 | n23968;
assign n26768 = ~n13667;
assign n16594 = ~n16507;
assign n25593 = n3251 & n3530;
assign n3764 = ~n4294;
assign n19275 = n1075 | n137;
assign n11207 = ~(n7657 ^ n25926);
assign n1633 = n11855 | n25366;
assign n22596 = ~(n4562 ^ n3136);
assign n12487 = ~(n8451 ^ n4537);
assign n2400 = n2722 | n9390;
assign n18280 = n20056 & n17692;
assign n6714 = ~(n18319 ^ n6267);
assign n14221 = n15553 | n16883;
assign n11492 = n11177 | n13137;
assign n11722 = n9386 & n17691;
assign n1165 = n7082 | n23466;
assign n4003 = ~n25221;
assign n17338 = ~(n20862 ^ n6876);
assign n23714 = ~(n20900 ^ n9350);
assign n10600 = n11081 | n12023;
assign n20380 = n12387 | n6057;
assign n11912 = n19584 | n6279;
assign n7970 = ~n26705;
assign n12466 = n11530 & n11545;
assign n10149 = n21635 | n13295;
assign n17864 = ~n3187;
assign n6505 = n11780 & n12254;
assign n26104 = ~(n23907 ^ n25731);
assign n17473 = n18814 | n9037;
assign n5240 = ~n19665;
assign n8987 = ~(n21984 | n4440);
assign n12005 = n6426 | n2362;
assign n1295 = n26543 | n26244;
assign n3354 = ~n21175;
assign n5836 = ~(n21066 | n23789);
assign n22958 = ~n26797;
assign n23626 = n18096 & n14377;
assign n9651 = n18855 & n20925;
assign n6564 = ~(n4338 | n24430);
assign n6827 = n437 | n26945;
assign n7571 = ~(n6038 | n12171);
assign n16292 = n18952 | n16966;
assign n11004 = n604 & n4626;
assign n26810 = ~(n2503 ^ n20929);
assign n2214 = ~(n16076 ^ n13660);
assign n3033 = ~(n5260 | n16130);
assign n19379 = ~(n16274 ^ n23849);
assign n19254 = ~n485;
assign n8791 = n2955 & n6191;
assign n23889 = n7842 | n23989;
assign n8500 = n22442 | n3131;
assign n25745 = n14695 | n847;
assign n12096 = ~(n1497 | n4184);
assign n1420 = ~(n7143 ^ n3625);
assign n10460 = n24248 & n10640;
assign n3731 = ~(n27068 | n8508);
assign n18493 = n26564 | n7471;
assign n518 = n6860 & n10539;
assign n18001 = n2011 & n18845;
assign n26170 = ~n5750;
assign n27096 = ~(n17309 ^ n1909);
assign n20561 = n3831 | n21366;
assign n4751 = n19999 & n26561;
assign n11753 = ~(n2815 | n10455);
assign n3309 = n401 | n17410;
assign n13762 = n6039 | n9394;
assign n6944 = ~(n8876 ^ n4975);
assign n4033 = ~n19108;
assign n21681 = n12947 & n24449;
assign n22884 = ~(n4775 ^ n20235);
assign n24083 = ~(n13357 | n506);
assign n22579 = n9600 | n19701;
assign n15044 = n20555 & n17246;
assign n5085 = ~(n5696 ^ n23463);
assign n12365 = n24486 | n7092;
assign n21542 = n4169 & n25300;
assign n16887 = ~(n22862 ^ n16543);
assign n22417 = n13731 | n21038;
assign n3853 = ~n12265;
assign n9630 = n18018 | n1337;
assign n11649 = ~n26726;
assign n84 = n22486 & n14266;
assign n17148 = n17951 | n14084;
assign n19671 = n5779 | n2103;
assign n23337 = ~(n19610 ^ n9159);
assign n24440 = n10066 | n18565;
assign n4285 = ~(n25797 | n10611);
assign n18650 = n6092 | n26261;
assign n10824 = n6247 | n11867;
assign n12867 = n11826 | n7205;
assign n6722 = n16389 | n13700;
assign n6178 = ~(n2430 ^ n16550);
assign n17619 = n21486 | n12338;
assign n4981 = n18637 & n9916;
assign n7413 = n4728 | n969;
assign n11592 = ~(n10806 ^ n21160);
assign n16501 = n17904 & n683;
assign n14293 = ~n1099;
assign n4934 = ~(n7876 ^ n25435);
assign n26505 = ~n3700;
assign n8775 = ~(n9469 | n3237);
assign n2066 = n24850 & n22706;
assign n17985 = n3626 & n21099;
assign n23330 = ~(n11121 | n19494);
assign n19586 = n21867 | n19155;
assign n4135 = n3948 | n4551;
assign n22428 = ~n18416;
assign n21708 = ~(n21556 | n23068);
assign n25108 = n12576 | n17287;
assign n24385 = n1522 & n14138;
assign n7736 = n25778 | n7223;
assign n3024 = n16654 | n7824;
assign n19856 = ~n6458;
assign n970 = ~(n3069 | n18485);
assign n15489 = ~(n578 ^ n24622);
assign n12795 = ~(n24327 | n25967);
assign n14727 = n24362 & n10007;
assign n23620 = ~n26853;
assign n4382 = ~(n5360 ^ n10493);
assign n21733 = ~(n24763 ^ n18089);
assign n3467 = n27182 | n9033;
assign n100 = n9107 & n18008;
assign n3295 = n6488 | n10521;
assign n22818 = ~(n18318 ^ n3946);
assign n9409 = ~(n19368 ^ n24828);
assign n7067 = n24432 | n14327;
assign n5785 = n6299 & n7096;
assign n15487 = ~n11036;
assign n25871 = ~(n13839 ^ n2575);
assign n22947 = n24614 | n5830;
assign n15682 = ~(n5580 | n3359);
assign n18761 = ~(n24990 | n19502);
assign n2818 = ~n24796;
assign n7351 = ~(n26865 ^ n15839);
assign n474 = n7000 | n19535;
assign n21872 = n14496 | n14552;
assign n6366 = ~n14184;
assign n25307 = n17641 & n8336;
assign n22260 = ~n5387;
assign n7696 = n24062 | n4911;
assign n26955 = n6231 & n13107;
assign n311 = ~n13465;
assign n3281 = ~(n5743 ^ n17967);
assign n1096 = ~(n9873 | n20558);
assign n674 = ~(n6698 ^ n21295);
assign n3706 = n7974 & n2759;
assign n20627 = n14483 & n18747;
assign n14683 = ~(n19460 | n12586);
assign n21141 = ~(n8322 | n3468);
assign n13150 = n26744 | n16240;
assign n22123 = ~n18578;
assign n16486 = ~n26619;
assign n19259 = n13701 & n14270;
assign n8022 = ~(n11657 ^ n12426);
assign n7126 = n21016 | n19254;
assign n22550 = ~n11605;
assign n14742 = n8396 | n12539;
assign n73 = ~(n18451 | n27034);
assign n25420 = n22261 | n20094;
assign n24224 = n22418 | n23443;
assign n87 = n4757 & n3598;
assign n3188 = n9701 | n6076;
assign n22087 = n26093 & n10529;
assign n13842 = ~n23775;
assign n18806 = ~(n8197 ^ n1927);
assign n17307 = n12899 & n3534;
assign n19753 = n3620 | n14753;
assign n24788 = ~(n19942 ^ n11387);
assign n23597 = ~(n654 ^ n13932);
assign n23599 = n13180 & n10103;
assign n4338 = ~n20980;
assign n12722 = n21066 | n11497;
assign n6956 = ~(n6899 ^ n1883);
assign n17605 = ~n25355;
assign n4809 = n874 | n9043;
assign n20822 = ~(n25110 ^ n2570);
assign n13545 = n1559 | n4348;
assign n10112 = ~n5954;
assign n933 = ~(n17943 ^ n4306);
assign n5228 = ~(n9312 ^ n3336);
assign n8218 = ~(n26344 | n1433);
assign n1672 = ~n5206;
assign n10393 = n6221 | n14287;
assign n8618 = n5223 | n23136;
assign n12353 = ~(n15146 ^ n10125);
assign n13540 = ~(n3256 | n16300);
assign n21631 = ~(n23591 | n24690);
assign n24690 = ~n20624;
assign n13336 = ~(n1143 ^ n12817);
assign n15908 = ~(n18452 ^ n6397);
assign n26630 = ~(n24202 ^ n9595);
assign n7326 = ~n22355;
assign n9039 = ~(n3319 | n10255);
assign n582 = n15865 | n3415;
assign n23165 = ~(n14391 ^ n6293);
assign n3445 = ~(n6077 ^ n24767);
assign n5597 = ~(n5722 ^ n402);
assign n3724 = ~n12319;
assign n18070 = ~n8302;
assign n21744 = n1654 & n24245;
assign n24265 = ~(n12208 ^ n12522);
assign n22727 = ~(n3680 ^ n2697);
assign n871 = n24116 | n19797;
assign n8211 = n24545 | n26364;
assign n4875 = n649 | n16374;
assign n3955 = ~(n14349 ^ n19142);
assign n5173 = n10307 | n23633;
assign n12474 = ~n3984;
assign n8788 = n23444 & n15561;
assign n25759 = ~(n21634 | n7930);
assign n25178 = ~(n3031 ^ n8017);
assign n678 = ~n25413;
assign n9752 = ~(n22043 ^ n12121);
assign n20892 = n24471 | n5209;
assign n21765 = ~(n5937 ^ n18719);
assign n9804 = n12714 | n18584;
assign n3871 = ~(n6040 ^ n26280);
assign n16231 = n14569 | n26661;
assign n20164 = n8829 & n4452;
assign n26131 = ~(n5974 ^ n19313);
assign n20778 = n25314 | n19335;
assign n18142 = ~(n7083 ^ n18037);
assign n15860 = ~n10351;
assign n6367 = ~(n4288 ^ n24646);
assign n1601 = n4759 & n4818;
assign n18240 = ~(n3311 | n1139);
assign n7269 = n20134 & n15237;
assign n10572 = n21826 | n17670;
assign n12820 = n20383 | n3341;
assign n4672 = n12312 & n16107;
assign n6117 = ~(n1956 | n16594);
assign n12034 = ~(n16672 ^ n2252);
assign n15542 = n5767 & n23435;
assign n21984 = ~n16906;
assign n7644 = ~n10352;
assign n9525 = ~n4639;
assign n18710 = ~n26007;
assign n11321 = n19499;
assign n12255 = n12069 & n16115;
assign n23941 = n3273 & n20414;
assign n26209 = n4371 & n11849;
assign n6313 = n24072 & n14312;
assign n13872 = n13081 & n18451;
assign n22840 = n5326 & n15669;
assign n6855 = ~(n8851 | n9944);
assign n2249 = ~(n22693 ^ n19722);
assign n24692 = n21933 & n668;
assign n16560 = ~n10377;
assign n6493 = n4807 | n5059;
assign n4630 = n12650 | n18486;
assign n26019 = ~(n23589 | n12891);
assign n20975 = ~(n21613 | n6242);
assign n13469 = ~(n45 | n15657);
assign n11002 = ~(n42 ^ n5348);
assign n4494 = n21242 & n6167;
assign n11297 = ~(n23161 ^ n3383);
assign n6961 = ~(n16158 ^ n24085);
assign n4963 = ~(n24293 ^ n12765);
assign n18201 = ~(n5571 ^ n9672);
assign n4544 = ~(n20213 | n9765);
assign n5692 = n22281 & n8537;
assign n19837 = n22420 | n15862;
assign n22021 = ~n18812;
assign n12653 = n27039 | n18656;
assign n23303 = ~(n22176 ^ n12384);
assign n197 = ~(n24635 ^ n11800);
assign n3364 = n23895 | n4446;
assign n21420 = ~n18934;
assign n15586 = ~(n12828 ^ n3602);
assign n7432 = ~(n18984 ^ n5856);
assign n10204 = ~(n19113 ^ n2731);
assign n21365 = ~(n16005 ^ n17081);
assign n3654 = n3255 & n18169;
assign n23506 = ~n4978;
assign n13312 = n4868 | n10993;
assign n19138 = n22924 | n15745;
assign n3441 = n11652 & n5047;
assign n9860 = ~(n22049 ^ n24196);
assign n19938 = ~(n14932 ^ n17623);
assign n12302 = ~(n18670 ^ n135);
assign n25581 = n2906 & n14187;
assign n26573 = ~(n7128 ^ n24030);
assign n25172 = ~(n25007 | n24286);
assign n377 = ~(n11172 | n7325);
assign n10497 = n10650 | n17978;
assign n9681 = ~(n8186 | n20040);
assign n16756 = n13637 | n2622;
assign n20957 = n4155 & n13031;
assign n21552 = n21621 | n813;
assign n27170 = ~(n15084 ^ n16615);
assign n18521 = ~(n17641 | n12198);
assign n23595 = n7306 | n8374;
assign n8213 = n11583 | n20544;
assign n20748 = ~(n4950 ^ n97);
assign n2121 = ~n19454;
assign n22348 = n21599 | n26324;
assign n22833 = n10886 & n9542;
assign n8298 = n6857 & n14400;
assign n12783 = ~(n2911 ^ n9072);
assign n14975 = ~(n25120 ^ n3582);
assign n4233 = n7224 | n26663;
assign n19920 = ~(n20455 ^ n3828);
assign n5578 = ~(n1558 | n3918);
assign n25079 = ~(n6218 ^ n25464);
assign n27060 = ~(n866 ^ n17155);
assign n22080 = ~(n3839 ^ n21774);
assign n26088 = ~(n17381 | n13649);
assign n10266 = ~n14524;
assign n2294 = n3290 | n5873;
assign n14261 = n8543 & n12028;
assign n6234 = n10761 & n3985;
assign n15392 = n8147 & n9650;
assign n3761 = n11141 & n9189;
assign n21494 = n22760 | n7576;
assign n23673 = ~(n10767 ^ n15062);
assign n2236 = ~(n13443 | n23923);
assign n15804 = n6136 | n10708;
assign n11409 = ~n15670;
assign n8889 = ~(n13468 ^ n3705);
assign n8731 = ~(n15693 ^ n3391);
assign n3358 = n18029 & n16779;
assign n26674 = ~(n26038 ^ n5522);
assign n24294 = n8284 & n25361;
assign n24687 = n4295 | n11151;
assign n20585 = n153 | n26301;
assign n6538 = n21592 & n14709;
assign n16290 = ~(n18885 ^ n2116);
assign n7737 = n21578 & n1295;
assign n7208 = n16722 & n21101;
assign n25755 = n15117 & n13716;
assign n10880 = n11402 | n7854;
assign n27045 = n10443 | n25537;
assign n21032 = ~(n13098 ^ n3056);
assign n6215 = ~(n16449 | n4185);
assign n6753 = ~n18290;
assign n15642 = ~(n21508 ^ n19393);
assign n15928 = ~(n11938 | n25126);
assign n16101 = ~(n6138 | n3317);
assign n5358 = n11046 & n18890;
assign n12533 = n19234 & n1365;
assign n16251 = ~(n2044 ^ n7130);
assign n25210 = ~(n22913 ^ n441);
assign n22128 = n13731 | n8920;
assign n1147 = ~(n10405 ^ n7731);
assign n19114 = ~(n23862 ^ n14538);
assign n8423 = ~(n20075 | n18158);
assign n11882 = ~(n2979 ^ n9554);
assign n17080 = n10740 | n17564;
assign n25822 = n12576 | n25475;
assign n1580 = ~(n5294 ^ n17279);
assign n16390 = n5808 & n7696;
assign n17875 = n25101 | n15174;
assign n18153 = n15673 & n21003;
assign n9503 = ~(n643 ^ n17804);
assign n20162 = ~(n24705 ^ n26444);
assign n19961 = n932 | n10739;
assign n6545 = n23092 & n22228;
assign n19337 = ~(n7925 ^ n15926);
assign n8178 = ~(n26495 ^ n19701);
assign n20858 = n23957 | n3825;
assign n7687 = n21921 & n14214;
assign n21308 = ~(n12351 ^ n6503);
assign n16794 = ~(n21662 ^ n6773);
assign n8634 = n18333 | n12509;
assign n26584 = ~(n4377 ^ n18961);
assign n4010 = ~(n19755 ^ n6367);
assign n26092 = n16524 & n17539;
assign n3017 = ~(n4600 ^ n9981);
assign n21824 = ~(n17127 ^ n17731);
assign n12288 = ~(n5951 ^ n17383);
assign n21620 = ~(n24448 ^ n9534);
assign n23932 = ~n8656;
assign n1130 = n23296 | n5413;
assign n25851 = n13358 & n25453;
assign n27052 = ~(n4692 | n21469);
assign n4273 = ~(n14620 ^ n17077);
assign n20085 = n12821 | n6596;
assign n24970 = ~n6699;
assign n23663 = ~(n1033 ^ n8619);
assign n22983 = ~(n21138 | n3187);
assign n10581 = ~n1700;
assign n17111 = n20165 | n5721;
assign n20829 = ~n1738;
assign n4954 = ~(n26553 ^ n23775);
assign n6377 = n10181 & n2066;
assign n12906 = ~n4108;
assign n7935 = ~(n1874 ^ n1313);
assign n14564 = ~n21492;
assign n22831 = ~(n5354 ^ n14972);
assign n19408 = n7564 & n10952;
assign n6417 = n23063 | n15265;
assign n16197 = n1816 | n19013;
assign n9917 = ~(n1758 ^ n10878);
assign n3579 = n14002 | n16396;
assign n26486 = ~n12531;
assign n17460 = n18663 & n11820;
assign n10022 = ~(n19729 ^ n10745);
assign n16640 = ~(n6955 ^ n22457);
assign n10772 = ~(n15086 ^ n17971);
assign n8362 = ~(n23884 | n17289);
assign n5499 = n22727 & n17411;
assign n774 = n16582 | n17808;
assign n16335 = n16983 | n14411;
assign n21545 = ~(n18203 ^ n16366);
assign n7878 = n2916 | n24559;
assign n17824 = n808 & n12102;
assign n23291 = n22231 & n24640;
assign n23344 = n13502 | n11224;
assign n8462 = ~n26763;
assign n25406 = ~(n20478 ^ n1204);
assign n6700 = ~(n17640 ^ n13217);
assign n11098 = ~n9653;
assign n6730 = n11405 | n18305;
assign n1739 = ~n17525;
assign n7135 = n24836 | n10329;
assign n6005 = n23278 & n7493;
assign n21247 = n5178;
assign n23259 = ~(n2421 ^ n5337);
assign n7576 = n2138 & n5035;
assign n25999 = ~(n15229 ^ n8050);
assign n16385 = n19701 | n13074;
assign n9049 = ~(n21608 | n7721);
assign n13744 = n13102 | n14199;
assign n27027 = ~n16285;
assign n14830 = ~(n10688 ^ n1169);
assign n8480 = ~(n4684 ^ n2471);
assign n27119 = n22585 | n23226;
assign n26879 = n19911 | n10472;
assign n24373 = ~(n26357 ^ n7976);
assign n25911 = n10102 | n12661;
assign n21677 = n11166 | n5358;
assign n7616 = ~(n1508 ^ n13928);
assign n10949 = ~(n18220 ^ n20634);
assign n15355 = ~(n16260 ^ n26804);
assign n7380 = n19371 | n15960;
assign n13215 = ~(n13953 ^ n18950);
assign n19590 = ~(n16477 ^ n11697);
assign n23524 = n9836 & n16676;
assign n9588 = n20489 & n26913;
assign n19594 = ~n8422;
assign n24212 = ~n21112;
assign n6401 = ~n18703;
assign n27015 = ~(n8141 ^ n18094);
assign n17076 = n14246 & n13272;
assign n8119 = ~(n22560 ^ n23575);
assign n27102 = ~(n3182 ^ n21854);
assign n27053 = n24358 | n24665;
assign n20055 = n11651 & n12906;
assign n17509 = n7330 | n2479;
assign n6086 = ~(n88 | n14453);
assign n18086 = n17479 | n12821;
assign n22925 = ~(n15189 | n1364);
assign n1217 = n2350 | n19487;
assign n9718 = n2915 & n10224;
assign n22634 = ~(n6045 ^ n16690);
assign n2905 = n24478 | n1623;
assign n14601 = ~(n17664 | n5115);
assign n12813 = ~(n22332 ^ n21934);
assign n24795 = ~(n15258 ^ n11775);
assign n4219 = n6932 | n5973;
assign n8027 = ~(n16000 ^ n16692);
assign n7874 = n3105 & n27097;
assign n24676 = n27046 | n14282;
assign n11212 = n7935 | n18608;
assign n9565 = ~n13258;
assign n21187 = n9380 & n24686;
assign n4478 = ~(n3462 ^ n7703);
assign n7395 = ~(n7466 ^ n21721);
assign n18980 = n8672 | n5296;
assign n11852 = n26654 | n9538;
assign n16586 = ~n9250;
assign n18982 = ~(n1094 ^ n10644);
assign n15580 = ~n17251;
assign n12410 = ~(n8721 | n1040);
assign n17226 = ~(n15910 | n8609);
assign n13916 = n10544 & n6163;
assign n14104 = ~(n1163 | n18901);
assign n2123 = n8208 | n18718;
assign n13341 = n14798 & n10162;
assign n10398 = ~n23212;
assign n4054 = n23514 | n15132;
assign n21673 = ~(n12734 ^ n20023);
assign n13512 = n14284 | n4276;
assign n10809 = n8542 | n7029;
assign n8991 = ~n10633;
assign n5475 = ~n22404;
assign n1258 = n2688 & n8163;
assign n16997 = n10416 | n5107;
assign n6898 = ~(n18472 | n20745);
assign n25765 = ~(n21606 ^ n26786);
assign n231 = n10083 & n7762;
assign n10041 = ~(n14513 ^ n12063);
assign n18281 = n24978 | n17278;
assign n21933 = n2903 | n25120;
assign n18833 = n26310 & n14799;
assign n26490 = n26470 | n21654;
assign n7714 = ~(n17101 | n552);
assign n25298 = ~(n24074 | n23464);
assign n17692 = ~(n12017 ^ n8169);
assign n578 = n19405 & n15115;
assign n10306 = ~(n9028 ^ n25240);
assign n5265 = ~(n4034 ^ n3291);
assign n8302 = ~(n24831 ^ n4349);
assign n20948 = ~n3786;
assign n24372 = ~(n17408 ^ n20235);
assign n9927 = n14692 | n9387;
assign n23886 = n15992 & n6093;
assign n7457 = ~(n19207 ^ n12424);
assign n18111 = n16633 & n9923;
assign n5662 = n4778 & n1787;
assign n16855 = n3449 & n22195;
assign n9358 = ~(n21692 ^ n24812);
assign n25750 = n7712 | n13972;
assign n10427 = ~(n13976 ^ n16903);
assign n4134 = ~(n9116 ^ n10466);
assign n8811 = n22244 | n12834;
assign n14149 = ~(n8001 | n20516);
assign n22292 = n2835 & n26262;
assign n10447 = ~(n3280 ^ n8117);
assign n16222 = ~(n19816 | n9421);
assign n13359 = n17180;
assign n23569 = n15513 | n6690;
assign n6696 = n24718 | n22677;
assign n25978 = n26198 & n2982;
assign n20924 = ~(n18496 | n25331);
assign n1315 = n759 | n22848;
assign n1870 = ~(n11363 | n6590);
assign n20246 = n17305 | n7817;
assign n3070 = n22814 | n26355;
assign n1161 = ~(n3837 | n12184);
assign n2633 = ~n23432;
assign n1519 = ~(n19235 ^ n6799);
assign n16408 = n20581 | n24109;
assign n2583 = ~(n12946 ^ n21067);
assign n1735 = ~(n20507 ^ n25086);
assign n22376 = ~(n644 ^ n12868);
assign n25866 = n20921 & n25106;
assign n20991 = ~(n14539 | n12878);
assign n22976 = n4555 | n11736;
assign n16991 = n18856 & n7413;
assign n17343 = ~(n22021 ^ n1441);
assign n23495 = ~(n22655 ^ n13189);
assign n11350 = ~n19863;
assign n18966 = ~(n302 | n16672);
assign n10102 = ~(n23170 | n20655);
assign n3926 = n21414 & n24577;
assign n19757 = ~n25977;
assign n20229 = ~(n15688 | n26912);
assign n19436 = n12519 & n21571;
assign n18733 = n7106 | n12750;
assign n25980 = n21937 & n17431;
assign n20140 = ~(n12098 | n21522);
assign n18500 = ~(n13724 ^ n17398);
assign n9918 = n2281 | n17343;
assign n5410 = ~n26189;
assign n16976 = n26319 | n9610;
assign n8274 = ~(n18947 ^ n10331);
assign n1272 = ~(n24031 | n19033);
assign n27064 = n17341 & n2672;
assign n23149 = n5019 | n25851;
assign n17764 = n13118 & n4694;
assign n13439 = ~(n21066 ^ n12509);
assign n3526 = ~n2981;
assign n26965 = ~(n23089 ^ n9830);
assign n26407 = ~(n20011 | n5697);
assign n14178 = n780 & n15811;
assign n705 = n11455 | n9940;
assign n24530 = ~(n19509 | n4924);
assign n16819 = n11378 | n9754;
assign n21950 = n18684 & n3688;
assign n19218 = ~n15764;
assign n24578 = ~(n4251 ^ n23361);
assign n6693 = ~n19647;
assign n6483 = ~(n5983 ^ n2265);
assign n9685 = ~(n18371 ^ n7933);
assign n5176 = ~(n16638 ^ n12380);
assign n19057 = ~n8629;
assign n9476 = ~(n9319 ^ n1810);
assign n12251 = ~n24137;
assign n7167 = ~n25430;
assign n5116 = n25010 & n7087;
assign n10430 = ~(n12338 ^ n26856);
assign n11695 = ~n13479;
assign n12334 = n9209 & n25992;
assign n12527 = n6609 & n21220;
assign n8474 = n18593 | n1544;
assign n19950 = ~(n7818 | n7320);
assign n23740 = ~n18727;
assign n23589 = ~n23203;
assign n8902 = n23795 & n22883;
assign n15900 = n25043 & n17901;
assign n17543 = ~(n24417 | n15271);
assign n22703 = ~(n26999 | n3990);
assign n5599 = n7074 ^ n3559;
assign n8714 = ~n10797;
assign n20997 = ~(n644 ^ n154);
assign n3035 = n20700 | n26240;
assign n15386 = n5368 | n3360;
assign n4183 = n23845 | n20548;
assign n10337 = n20613 & n14138;
assign n10850 = n561 | n16278;
assign n2752 = n19673 | n22743;
assign n12748 = n4365 | n16303;
assign n3908 = ~(n25164 | n10689);
assign n6499 = ~(n11893 | n11337);
assign n2456 = ~(n14251 ^ n1742);
assign n10787 = n3959 | n11810;
assign n1267 = ~(n17265 ^ n17458);
assign n26289 = ~n15883;
assign n15061 = n19163 | n10513;
assign n15444 = n7237 | n16351;
assign n23773 = n22447 | n7047;
assign n13824 = n18410 & n11762;
assign n8068 = ~n21095;
assign n3863 = n9752 | n4467;
assign n816 = ~n5794;
assign n20132 = ~(n26529 | n3939);
assign n8059 = n2121 & n4213;
assign n14245 = n24866 | n3826;
assign n19011 = n10346 | n2163;
assign n17099 = ~(n16022 | n18575);
assign n10183 = ~(n9207 ^ n19577);
assign n20812 = n4483 & n3566;
assign n23209 = ~n3769;
assign n965 = n8144 | n17792;
assign n2878 = ~(n5996 ^ n2528);
assign n18618 = n3666 | n3926;
assign n26933 = n20924 | n7869;
assign n25038 = ~n3324;
assign n22625 = ~(n7609 ^ n21496);
assign n4727 = n18814 & n9037;
assign n11635 = n21867 | n22248;
assign n11152 = ~n20604;
assign n13988 = ~(n6566 ^ n9509);
assign n17883 = ~n197;
assign n5548 = ~(n6025 ^ n13941);
assign n11330 = ~(n6771 ^ n5074);
assign n9250 = n6117 | n25901;
assign n17421 = ~(n2364 ^ n803);
assign n21329 = n6742 & n7510;
assign n10952 = n13268 | n11729;
assign n5269 = n192 & n12706;
assign n2712 = n20575 | n11933;
assign n15005 = n19973 | n14794;
assign n17223 = n2566 & n4894;
assign n24884 = n11763 & n2888;
assign n10894 = ~(n14016 | n22282);
assign n24475 = ~(n13289 ^ n14927);
assign n19659 = n15826 | n20438;
assign n11123 = n4589 & n6370;
assign n24098 = ~n10117;
assign n210 = n22708 & n3757;
assign n7908 = n7537 | n21724;
assign n5367 = ~(n2878 ^ n13775);
assign n25402 = n15447 & n24951;
assign n5224 = ~(n8745 ^ n26913);
assign n6462 = ~(n22219 ^ n12514);
assign n14947 = ~(n16396 ^ n18295);
assign n16474 = ~n11926;
assign n18561 = n8101 | n9468;
assign n2859 = n16568 | n183;
assign n2864 = ~n12679;
assign n937 = n10554 | n330;
assign n7846 = n1355 & n20363;
assign n325 = ~(n23235 ^ n8253);
assign n7499 = n2006 & n22453;
assign n22101 = n13569 & n7374;
assign n20693 = ~(n8695 ^ n19932);
assign n17616 = ~n81;
assign n19873 = ~(n14611 ^ n742);
assign n15477 = ~(n20561 ^ n3735);
assign n23043 = ~(n11615 | n23018);
assign n262 = n15717 | n15611;
assign n23676 = n19 | n24875;
assign n12393 = n2309 | n15845;
assign n4558 = ~n25656;
assign n1572 = ~(n24481 ^ n21905);
assign n7775 = ~(n13068 ^ n826);
assign n1206 = n16761 & n19169;
assign n14937 = ~n23475;
assign n16367 = n8513 | n415;
assign n20971 = n19430 & n20337;
assign n9775 = ~(n2071 ^ n8285);
assign n21433 = ~n26185;
assign n16080 = ~(n171 ^ n10260);
assign n15643 = ~(n13363 ^ n2828);
assign n19063 = ~(n1631 ^ n21247);
assign n16958 = n7088 | n20393;
assign n23970 = ~n20564;
assign n20938 = n11692 & n16710;
assign n6666 = n1871 & n18083;
assign n20345 = ~(n13967 | n9655);
assign n15945 = n13309 | n24278;
assign n13244 = ~(n10441 | n6727);
assign n10450 = n6275 | n2075;
assign n4526 = n140 & n22354;
assign n1238 = ~(n1145 ^ n11794);
assign n1292 = ~(n14761 ^ n26460);
assign n3841 = n16387 & n507;
assign n3457 = n643 | n17804;
assign n3866 = n19398 | n20050;
assign n12857 = ~(n17458 | n23064);
assign n14059 = ~(n2714 ^ n24837);
assign n8000 = ~n17999;
assign n351 = n269 | n24719;
assign n8496 = ~n6281;
assign n2801 = ~n650;
assign n25545 = n7292 | n546;
assign n12422 = ~n14444;
assign n8924 = n10863 | n16581;
assign n25410 = n9661 | n14850;
assign n11777 = n4045 | n23688;
assign n12211 = ~(n27083 ^ n3508);
assign n26461 = ~(n21681 ^ n256);
assign n8041 = ~(n23626 ^ n16149);
assign n18707 = ~(n1343 ^ n26748);
assign n8713 = ~n26583;
assign n23244 = ~n1639;
assign n18694 = ~(n16427 ^ n17888);
assign n4031 = ~n14723;
assign n4430 = n25136 & n15005;
assign n18565 = n8953 & n6594;
assign n5600 = n1294 & n1585;
assign n795 = n2483 | n6079;
assign n11726 = n1064 & n11436;
assign n17611 = n12682 | n817;
assign n18082 = n10655 | n18064;
assign n16684 = ~(n22967 ^ n24542);
assign n23103 = ~(n13197 ^ n17674);
assign n4286 = ~(n18514 | n11597);
assign n14643 = ~n19158;
assign n23378 = n19830 | n21457;
assign n5076 = n21764 | n16026;
assign n14227 = n12920 | n18557;
assign n10829 = ~(n12744 ^ n816);
assign n15226 = ~(n26215 ^ n22083);
assign n10029 = ~(n10918 | n5633);
assign n766 = n25168 | n17094;
assign n11218 = n1327 | n13201;
assign n9428 = n11554 | n2964;
assign n25090 = n17013 | n23974;
assign n20420 = n22841 | n9935;
assign n24730 = n22963 | n7110;
assign n17879 = n23084 | n3870;
assign n8425 = ~(n25074 | n10053);
assign n17142 = ~(n17483 ^ n24573);
assign n7845 = n24906 & n8397;
assign n13855 = n8100 & n2481;
assign n15395 = ~(n23359 | n19444);
assign n14465 = ~n12956;
assign n8459 = n11186 | n26054;
assign n3937 = n571 | n23499;
assign n26297 = n19282 | n23709;
assign n11142 = n22462 | n10994;
assign n4154 = ~(n7149 ^ n22871);
assign n16567 = ~(n14230 | n19922);
assign n23824 = n13871 & n20746;
assign n17725 = ~n11751;
assign n19814 = ~n11539;
assign n4965 = n15055 | n5270;
assign n2556 = ~(n9247 | n18715);
assign n8140 = ~(n8569 ^ n13119);
assign n3827 = ~(n24777 ^ n5940);
assign n16782 = n13346 & n15592;
assign n2018 = n5775 & n15934;
assign n14959 = n18069 & n1130;
assign n12133 = n25661 & n25182;
assign n7605 = ~n6175;
assign n22182 = ~n25251;
assign n24785 = ~(n26209 | n10462);
assign n8262 = n5204 | n1761;
assign n3948 = n17333 & n14783;
assign n15577 = ~(n23095 | n22332);
assign n10184 = ~n11736;
assign n22651 = ~n16722;
assign n17687 = ~(n764 ^ n8798);
assign n22121 = ~(n16119 ^ n4739);
assign n26457 = n21691 | n16158;
assign n26284 = n3968 | n6070;
assign n14267 = ~(n22109 ^ n18168);
assign n15529 = ~(n12446 | n1112);
assign n19010 = n5761 & n7955;
assign n9880 = ~n18151;
assign n4232 = ~(n15743 ^ n2809);
assign n7186 = n4414 & n17019;
assign n13378 = ~n8285;
assign n3158 = ~(n20250 ^ n1682);
assign n12322 = ~(n16412 ^ n25214);
assign n10256 = n25259 | n14757;
assign n2902 = n2155 & n7097;
assign n13584 = n12126 & n7023;
assign n427 = ~n14424;
assign n9207 = n22931 & n3701;
assign n19686 = ~(n24802 ^ n9359);
assign n4569 = ~n3247;
assign n7364 = ~n19560;
assign n19924 = ~(n4866 ^ n1809);
assign n14128 = n10146 | n21753;
assign n22407 = ~(n24202 ^ n18274);
assign n25340 = n12197 & n10068;
assign n20961 = n16783 | n21891;
assign n930 = ~(n22527 | n19820);
assign n18511 = ~(n24066 ^ n12555);
assign n23719 = ~(n23547 | n25569);
assign n21426 = ~(n2360 ^ n22764);
assign n22094 = n8261 | n18905;
assign n21066 = ~n18333;
assign n8937 = ~n5696;
assign n11813 = n12918 | n1758;
assign n5828 = n15684 | n1852;
assign n14578 = ~(n115 | n22859);
assign n25013 = n18485 | n12811;
assign n20011 = ~n7825;
assign n17589 = ~(n2093 ^ n18520);
assign n14800 = ~(n5714 | n1222);
assign n2484 = n3537 & n7542;
assign n21209 = ~n2953;
assign n48 = ~(n17034 ^ n23951);
assign n25031 = n7929 & n24581;
assign n18007 = n4707 & n19622;
assign n10725 = ~(n25120 ^ n23272);
assign n20836 = ~(n25514 | n13696);
assign n16582 = ~(n14489 ^ n18317);
assign n13219 = n3259 & n21720;
assign n24994 = n9466 | n21798;
assign n17729 = ~(n4542 ^ n18295);
assign n16261 = ~(n1990 ^ n14548);
assign n8696 = n29 | n14372;
assign n10264 = n18746 | n26452;
assign n15043 = n10061 | n5027;
assign n6768 = ~(n21333 | n20098);
assign n517 = n18564 & n9562;
assign n20390 = n9755 | n18048;
assign n24733 = n16839 & n19030;
assign n20075 = ~n24051;
assign n1228 = n7768 | n1345;
assign n14364 = ~(n3839 ^ n10363);
assign n4869 = ~(n12298 ^ n22400);
assign n817 = n6258 & n18801;
assign n12974 = n9310 | n24115;
assign n3059 = n10622 | n501;
assign n14217 = ~(n11662 ^ n11775);
assign n2167 = n20991 | n20699;
assign n11254 = ~(n1241 ^ n11803);
assign n4937 = ~(n8656 ^ n9380);
assign n17848 = ~(n6051 | n15053);
assign n134 = n16393 & n16627;
assign n709 = ~(n14959 ^ n3183);
assign n10083 = n26901 | n22807;
assign n1900 = n7812 & n495;
assign n6344 = ~(n12673 ^ n25220);
assign n16431 = n11513 | n4111;
assign n14866 = ~(n22173 | n12593);
assign n7480 = n25143 & n25988;
assign n1471 = n2079 | n12095;
assign n14048 = ~(n22128 ^ n3151);
assign n8867 = n25628 | n23432;
assign n16816 = ~(n3608 ^ n24263);
assign n9699 = ~(n26440 ^ n7990);
assign n18915 = n23081 & n6205;
assign n14497 = n16680 | n15692;
assign n1875 = n26071 & n1425;
assign n15337 = ~n10915;
assign n8424 = n15217 | n15241;
assign n23090 = n2080 | n1319;
assign n18351 = n8910 | n19321;
assign n11866 = ~(n6127 ^ n4642);
assign n18130 = ~n18479;
assign n14042 = ~n22031;
assign n21754 = n1390 & n7495;
assign n16863 = n1161 | n377;
assign n18715 = ~n3663;
assign n5797 = n6788 | n18590;
assign n19323 = ~(n16603 ^ n11300);
assign n13267 = n26777 | n17;
assign n18418 = ~(n1390 ^ n10240);
assign n12386 = ~(n5823 ^ n6513);
assign n15382 = ~(n3820 ^ n3684);
assign n18957 = n22017 | n22671;
assign n19416 = n26916 & n24288;
assign n11135 = ~n13356;
assign n23504 = n5740 & n14653;
assign n16867 = n6872 | n16559;
assign n27082 = n12418 & n21959;
assign n16205 = ~n18907;
assign n9088 = ~(n8614 ^ n25972);
assign n18188 = n11099 & n26751;
assign n4056 = ~(n11457 | n15636);
assign n25451 = ~n9889;
assign n6574 = ~(n11938 | n19472);
assign n23702 = n21915 | n2509;
assign n3334 = ~(n17125 | n10532);
assign n24861 = ~(n4957 ^ n7421);
assign n25182 = n3408 | n2484;
assign n9933 = n6039 | n10199;
assign n10936 = n17732 & n20823;
assign n829 = ~(n13063 ^ n6278);
assign n27013 = n11750 | n9270;
assign n16596 = ~(n26293 ^ n26128);
assign n18335 = ~n7773;
assign n19596 = ~(n4230 | n8378);
assign n1719 = ~n3705;
assign n9707 = ~(n20169 ^ n1949);
assign n16947 = ~(n23487 | n6556);
assign n9263 = n21124 & n3295;
assign n18488 = ~(n16204 ^ n26117);
assign n19702 = ~n18972;
assign n4053 = n22743 & n2346;
assign n23619 = ~(n9785 ^ n16199);
assign n6547 = ~(n10602 | n21721);
assign n22812 = ~n4491;
assign n11357 = n16211 | n4256;
assign n16664 = n21937 | n14007;
assign n18396 = n8903 & n3950;
assign n20188 = n862 | n20386;
assign n10121 = n25161 | n8287;
assign n18116 = ~(n12446 ^ n1112);
assign n8206 = ~(n16478 ^ n3461);
assign n15788 = n15148 & n452;
assign n7299 = n18499 | n19009;
assign n23695 = ~(n21276 | n23061);
assign n24221 = ~n5718;
assign n3197 = ~(n3908 | n16490);
assign n3517 = n3016 | n7827;
assign n7700 = n26495 | n5789;
assign n5199 = n22060 & n594;
assign n6667 = n2708 & n12528;
assign n25269 = n6781 & n25477;
assign n14069 = n5373 & n14558;
assign n19118 = ~(n19245 ^ n9584);
assign n12441 = ~n21184;
assign n5014 = n21649 | n20192;
assign n5427 = ~(n6180 ^ n25487);
assign n1309 = ~(n23583 ^ n22531);
assign n11970 = ~(n22938 ^ n13732);
assign n10168 = n8910 | n19201;
assign n17235 = ~(n16042 ^ n11955);
assign n9833 = ~(n25350 ^ n3889);
assign n2229 = ~(n10372 ^ n12152);
assign n13547 = ~(n13569 | n7374);
assign n19486 = ~(n25804 ^ n13350);
assign n23091 = ~n14393;
assign n1299 = ~(n7566 | n22640);
assign n3359 = ~n1528;
assign n14388 = n21610 | n6151;
assign n4226 = n14884 & n18533;
assign n19271 = ~(n4495 ^ n15666);
assign n5195 = ~(n2152 ^ n25156);
assign n17452 = ~(n7913 ^ n23541);
assign n20695 = ~(n8411 | n945);
assign n5460 = n16034 & n10451;
assign n2264 = ~(n23864 | n12693);
assign n17523 = n12474 | n23109;
assign n24909 = n20416 | n12563;
assign n8636 = ~(n3515 | n93);
assign n22650 = n6264 | n3804;
assign n17680 = n22672 & n16404;
assign n3417 = n6981 & n11825;
assign n15463 = ~(n23529 | n9124);
assign n2692 = ~(n24615 | n1742);
assign n8017 = ~(n6729 ^ n10792);
assign n1724 = ~(n18715 ^ n6178);
assign n3508 = ~(n1019 ^ n11011);
assign n20613 = ~(n13019 ^ n10108);
assign n9426 = ~(n19312 ^ n17928);
assign n13032 = n24674 & n19846;
assign n6 = n24004 & n12900;
assign n8045 = n18220 | n8420;
assign n20584 = n8372 | n20378;
assign n1864 = ~n19515;
assign n14080 = n7704 & n21318;
assign n3974 = n771 | n23383;
assign n2513 = n15110 & n19292;
assign n18654 = n26926 & n22245;
assign n25274 = n18473 | n4812;
assign n4395 = ~n18895;
assign n26926 = n25250 | n18793;
assign n7608 = ~(n22895 ^ n27200);
assign n14413 = n19359 | n9781;
assign n3063 = ~(n23559 ^ n11481);
assign n27162 = n1030 | n19240;
assign n21431 = n19770 & n12022;
assign n13203 = n16205 | n26823;
assign n19056 = n2915 | n10224;
assign n18908 = ~(n11792 | n22571);
assign n26395 = n2986 | n25422;
assign n3189 = ~(n3568 ^ n22934);
assign n925 = ~(n16064 ^ n19460);
assign n5124 = n14436 & n8992;
assign n22587 = n22919 | n24506;
assign n18639 = n3223;
assign n12866 = n25208 | n26299;
assign n26303 = ~(n24037 ^ n13812);
assign n17661 = n7043 | n10616;
assign n25371 = n23555 | n18269;
assign n16572 = ~n16302;
assign n3133 = ~n2408;
assign n22548 = ~(n7972 ^ n12659);
assign n17217 = ~(n12019 | n2512);
assign n6717 = n17160 | n5927;
assign n2987 = n8023 & n19447;
assign n19756 = ~(n17594 ^ n4738);
assign n16221 = ~(n23012 ^ n1851);
assign n17159 = ~(n6226 ^ n4564);
assign n11869 = n21807 & n1417;
assign n15543 = n5145 | n9886;
assign n2213 = n10570 & n13374;
assign n12658 = ~(n4981 ^ n15152);
assign n21393 = n13781 & n26793;
assign n8605 = ~(n13480 | n16544);
assign n15237 = n246 & n17401;
assign n23828 = n13503 | n25575;
assign n13259 = n15107 & n15954;
assign n8629 = ~(n17645 ^ n10945);
assign n14342 = ~(n26679 ^ n26419);
assign n13092 = ~(n25514 | n4361);
assign n24382 = n6834 & n5165;
assign n20233 = ~(n19127 ^ n21727);
assign n6263 = ~(n27183 ^ n4185);
assign n12691 = n22149 | n23134;
assign n16975 = ~n22686;
assign n2000 = ~n13158;
assign n14162 = ~(n14907 | n25238);
assign n18533 = n2446 | n15969;
assign n26244 = n18702 & n22668;
assign n3743 = ~(n10918 ^ n9731);
assign n4835 = ~(n20489 ^ n26913);
assign n11562 = n25054 | n10138;
assign n6938 = n4722 & n6403;
assign n24458 = ~(n7903 ^ n6450);
assign n4918 = n7335 & n11578;
assign n24056 = ~(n19444 ^ n2979);
assign n2480 = ~(n24924 | n20876);
assign n26026 = n2153 & n5018;
assign n4274 = n6492 | n17718;
assign n26689 = ~(n25431 ^ n16824);
assign n7875 = n12619 & n20115;
assign n6668 = n18320 & n12653;
assign n7308 = ~(n20130 ^ n10599);
assign n24235 = n20481 & n2620;
assign n17671 = ~(n6295 ^ n9709);
assign n669 = n13647 & n18109;
assign n19248 = ~(n15739 ^ n12507);
assign n17472 = ~(n5685 ^ n189);
assign n6767 = n4604 & n8116;
assign n649 = ~(n13645 ^ n12001);
assign n4753 = ~(n22066 ^ n25130);
assign n7165 = n25391 & n19855;
assign n22373 = n2821 | n13594;
assign n20882 = n14910 | n21250;
assign n19331 = ~(n3920 ^ n1993);
assign n23875 = ~(n13360 ^ n26544);
assign n18178 = n4309 | n14727;
assign n20247 = ~(n26186 ^ n19556);
assign n505 = ~n3037;
assign n1622 = ~(n26180 ^ n10650);
assign n16737 = n7662 | n16616;
assign n25949 = ~(n15064 ^ n12861);
assign n25517 = n14564 | n9809;
assign n218 = ~n12125;
assign n4717 = ~(n22724 | n19614);
assign n7219 = n1257 | n1369;
assign n1828 = n7584 | n13221;
assign n23480 = ~(n10600 ^ n18683);
assign n8127 = n23347 | n23452;
assign n19061 = ~n25693;
assign n16244 = n15972;
assign n18771 = ~(n13018 ^ n22290);
assign n12963 = n22631 | n8819;
assign n72 = n25301 & n26679;
assign n9133 = ~(n23948 ^ n3193);
assign n14788 = n17284 & n7896;
assign n24955 = ~(n24600 ^ n3641);
assign n26125 = n26722 | n15074;
assign n13380 = n7948 | n1583;
assign n18844 = n2077 | n11749;
assign n5649 = n23038 & n23286;
assign n3200 = n4190 & n10328;
assign n23588 = ~(n15674 ^ n25503);
assign n12136 = ~(n3276 | n268);
assign n17271 = n25436 | n8162;
assign n12616 = ~(n20934 ^ n2306);
assign n14782 = ~(n8369 ^ n15120);
assign n12572 = ~(n17900 | n16459);
assign n17397 = ~n18139;
assign n4716 = n10381 | n1772;
assign n5820 = n25650 | n7177;
assign n15705 = ~(n14165 ^ n17729);
assign n2125 = ~n2886;
assign n7187 = ~(n15309 | n3846);
assign n17174 = n24752 | n4082;
assign n4887 = ~(n5698 ^ n27173);
assign n21161 = ~(n22433 | n10158);
assign n25862 = n3571 & n4607;
assign n23806 = ~n8317;
assign n10990 = ~(n10201 | n11336);
assign n19879 = n12240 & n14833;
assign n15372 = n22485 | n1100;
assign n9881 = ~(n17545 ^ n8750);
assign n11435 = n12533 | n7942;
assign n4023 = n1298 | n8203;
assign n13576 = ~(n14251 | n26946);
assign n23760 = ~n3552;
assign n8220 = ~n12094;
assign n21510 = n24131 & n25260;
assign n24691 = ~(n26417 | n6789);
assign n18397 = n24031 | n17993;
assign n13715 = ~n2987;
assign n1651 = n94 | n9476;
assign n24175 = n8747 & n3212;
assign n16555 = ~(n11341 ^ n25365);
assign n9558 = ~(n6743 ^ n23152);
assign n10401 = n15125 & n11929;
assign n10718 = ~(n11314 ^ n25738);
assign n23553 = n24018 | n1654;
assign n25786 = ~(n23497 ^ n21004);
assign n13117 = ~n17606;
assign n1033 = n19612 & n24459;
assign n4277 = ~(n22292 ^ n14589);
assign n21413 = n9618 & n14629;
assign n13987 = ~(n9151 ^ n7569);
assign n21347 = n20128 | n7862;
assign n24451 = ~(n21973 ^ n24916);
assign n585 = ~(n12702 ^ n12507);
assign n1683 = ~(n24638 ^ n442);
assign n9307 = n5908 | n792;
assign n4779 = n7431 | n26178;
assign n3801 = ~(n14528 | n16019);
assign n16151 = n15622 | n633;
assign n18513 = ~(n4864 ^ n13266);
assign n9489 = n5760 & n13954;
assign n19599 = n12554 | n21083;
assign n12768 = ~(n8773 | n10610);
assign n24321 = n7892 | n15734;
assign n27109 = n23868 | n2154;
assign n26246 = n18220 | n21577;
assign n23104 = n21812 & n14568;
assign n12845 = ~n14996;
assign n7471 = ~n22744;
assign n8080 = n7551 | n20535;
assign n13535 = ~n22824;
assign n16536 = ~(n25824 ^ n2349);
assign n5411 = ~(n25313 ^ n24859);
assign n12666 = ~(n24788 | n6025);
assign n4883 = ~n9431;
assign n59 = n19395 & n5497;
assign n21702 = ~(n10514 | n6105);
assign n11230 = n21775 & n2793;
assign n2698 = ~(n20738 ^ n3158);
assign n13287 = n27120 & n25504;
assign n23789 = ~(n6594 ^ n6559);
assign n13805 = n7453 | n20847;
assign n17028 = ~(n125 ^ n2659);
assign n16670 = ~(n26629 | n19904);
assign n13892 = n24947 | n19277;
assign n25520 = ~(n3258 ^ n12108);
assign n6426 = n12513 & n25568;
assign n1311 = n20053 | n6887;
assign n16936 = n24193 | n10977;
assign n16548 = ~n11336;
assign n4052 = n20028 & n18087;
assign n3144 = n3372 & n2451;
assign n2092 = ~(n5973 ^ n26838);
assign n3251 = n4858 | n602;
assign n17361 = n24181 | n21938;
assign n9469 = n3051;
assign n20980 = n12831 | n8554;
assign n5516 = ~n16158;
assign n10428 = n18297 | n22378;
assign n24216 = ~(n23791 | n7083);
assign n25550 = ~(n7076 ^ n14005);
assign n24565 = ~(n13839 | n14218);
assign n13751 = ~(n15761 | n12445);
assign n813 = n25492 & n8029;
assign n15330 = n12768 | n18508;
assign n11397 = n26434 & n18543;
assign n5735 = n3945 | n21998;
assign n21751 = ~(n17499 ^ n11474);
assign n24230 = ~(n24164 | n23475);
assign n20556 = ~n21295;
assign n10425 = ~n5706;
assign n14466 = ~(n26362 ^ n17827);
assign n6718 = ~(n6112 ^ n16797);
assign n13492 = ~n20005;
assign n12808 = ~(n4409 ^ n10125);
assign n9198 = ~(n20045 | n14510);
assign n16542 = n22662 & n16762;
assign n20469 = n13816 & n14997;
assign n20981 = ~(n19404 | n14700);
assign n628 = n13641 | n16000;
assign n14527 = ~(n6446 ^ n20060);
assign n4255 = ~(n3136 ^ n2409);
assign n12612 = ~n20959;
assign n24358 = ~n12495;
assign n24227 = n27104 & n13317;
assign n25805 = ~(n25297 ^ n23857);
assign n15078 = n11498 | n6316;
assign n1014 = n23112 & n2;
assign n12269 = ~(n13990 | n3744);
assign n6429 = n1098 & n20448;
assign n7888 = n26548 | n14658;
assign n23230 = ~n1118;
assign n6916 = ~n14902;
assign n8138 = ~(n12341 | n13945);
assign n16377 = n460 & n26666;
assign n77 = n15292 | n15752;
assign n12068 = ~n6912;
assign n12488 = ~(n114 ^ n16093);
assign n4270 = ~(n25021 | n10593);
assign n27062 = ~(n16705 | n14244);
assign n4710 = ~(n14963 | n11579);
assign n26819 = ~n8772;
assign n21193 = ~(n20542 ^ n13697);
assign n5575 = n21749 & n2298;
assign n26959 = n8782 | n18643;
assign n10532 = n15402 & n7309;
assign n7738 = n3818 & n9795;
assign n26540 = n6521 | n6659;
assign n5610 = n23402 & n9283;
assign n5903 = ~(n17849 ^ n22136);
assign n1794 = ~n23779;
assign n13207 = n9301 & n7718;
assign n9163 = n11385 & n5422;
assign n43 = n2592 & n20882;
assign n3172 = n12454 | n11481;
assign n25474 = ~(n6369 ^ n3164);
assign n4797 = ~(n13319 | n15490);
assign n25993 = n21388 & n1228;
assign n24330 = ~(n26233 ^ n21561);
assign n21698 = ~n513;
assign n26492 = ~(n14495 ^ n4271);
assign n2402 = ~(n15405 ^ n3940);
assign n11703 = n15564 & n11499;
assign n23117 = n24673 & n20451;
assign n12840 = n3150 | n25439;
assign n16905 = ~(n479 ^ n8701);
assign n7804 = n23200 | n16077;
assign n1358 = n2113 & n148;
assign n15365 = ~(n287 ^ n26160);
assign n414 = ~(n11220 ^ n12507);
assign n16345 = ~n8805;
assign n255 = ~n16373;
assign n9268 = ~(n24237 ^ n19592);
assign n9637 = ~(n63 | n13671);
assign n12408 = ~(n12429 ^ n23424);
assign n14770 = n1135 & n11839;
assign n14194 = ~(n6232 ^ n13472);
assign n11271 = ~(n4626 ^ n21509);
assign n7376 = ~(n26101 ^ n14046);
assign n22970 = n21436 | n22983;
assign n3966 = n23776 | n7417;
assign n23353 = ~n348;
assign n26873 = n621 | n18688;
assign n22658 = ~(n20011 | n17953);
assign n6601 = n24031 & n17993;
assign n5308 = n18837 | n1321;
assign n16941 = n20022 | n15141;
assign n13008 = ~(n23160 ^ n7678);
assign n11668 = ~(n23209 | n11755);
assign n6309 = ~n2324;
assign n22118 = n13766 | n6297;
assign n3430 = n12657 | n10092;
assign n9185 = n3480 | n7850;
assign n20752 = n18218 & n7430;
assign n17594 = n1479 | n16032;
assign n26274 = ~(n14175 ^ n13658);
assign n22210 = n2424 & n84;
assign n13884 = ~(n6737 ^ n17544);
assign n441 = ~(n22662 ^ n5048);
assign n16652 = n11226 | n15893;
assign n5889 = n6687 & n9837;
assign n18562 = ~(n23141 | n2035);
assign n21788 = ~(n16197 ^ n24936);
assign n18791 = ~(n3138 ^ n24245);
assign n24575 = ~n11099;
assign n17951 = ~(n24868 | n23268);
assign n21524 = n15628 | n21722;
assign n22200 = ~n11289;
assign n3620 = ~(n9671 | n4858);
assign n23411 = ~(n7350 ^ n1480);
assign n13084 = n7237 | n4873;
assign n23075 = n5159 & n11377;
assign n5363 = ~(n13953 | n17323);
assign n5323 = n24949 | n16423;
assign n10141 = ~(n8557 ^ n24739);
assign n8015 = ~(n18598 | n17077);
assign n7786 = n8885 & n4023;
assign n22006 = ~(n848 ^ n7864);
assign n5601 = ~n5713;
assign n7422 = ~n16413;
assign n11234 = ~(n22874 ^ n25765);
assign n21373 = ~(n19258 | n10919);
assign n4830 = n26798 | n6951;
assign n23122 = n13591 & n22114;
assign n21728 = ~(n4570 ^ n17591);
assign n25794 = n6169 & n26302;
assign n1046 = ~n3804;
assign n10013 = n14125;
assign n26260 = n10951 & n13372;
assign n2849 = ~(n3530 ^ n15857);
assign n22737 = n11922 & n13639;
assign n7229 = ~(n19622 ^ n19322);
assign n25977 = n13707 & n14854;
assign n14916 = n21429 & n9083;
assign n5850 = ~(n15732 ^ n9075);
assign n12930 = n23261 & n24460;
assign n10341 = n18880 & n26594;
assign n11024 = n6393 | n7948;
assign n4831 = n14556 & n1442;
assign n7899 = n24537 & n11210;
assign n19169 = n22733 | n16403;
assign n14786 = ~(n23709 ^ n14268);
assign n7669 = ~(n6749 ^ n1589);
assign n15707 = ~(n8386 | n3217);
assign n2138 = n2409 | n14071;
assign n15566 = n16805 & n6906;
assign n24910 = ~(n17485 ^ n17555);
assign n15057 = ~(n11210 ^ n24537);
assign n11708 = ~(n726 ^ n26849);
assign n24833 = n12594 & n21452;
assign n1137 = n24116 | n21556;
assign n8794 = ~n13372;
assign n18069 = n9671 | n5205;
assign n15067 = ~(n8436 ^ n14677);
assign n21045 = ~(n20896 ^ n6435);
assign n24199 = n8979 | n9856;
assign n11012 = n14708 | n19257;
assign n18814 = ~n20986;
assign n14869 = n21127 | n4588;
assign n12964 = ~(n14142 ^ n10766);
assign n18380 = n7342 | n5372;
assign n22208 = ~(n13775 | n11830);
assign n26652 = n13427 & n16646;
assign n9840 = n23218 & n22266;
assign n23816 = ~(n647 ^ n26408);
assign n293 = n22732 | n3887;
assign n17398 = ~(n1685 ^ n15633);
assign n15620 = ~(n2432 | n11137);
assign n12319 = ~(n3119 ^ n7534);
assign n916 = n2217 | n15038;
assign n5591 = ~(n7689 ^ n11314);
assign n24711 = ~(n2847 ^ n16);
assign n4688 = ~(n9485 ^ n16839);
assign n17682 = n14736 | n15274;
assign n17856 = ~(n21457 ^ n20790);
assign n6594 = n23425 | n12560;
assign n11373 = n19306 & n14235;
assign n16278 = ~(n23157 ^ n1863);
assign n21158 = ~(n25929 ^ n10013);
assign n13413 = n26172 | n8938;
assign n17977 = ~(n22651 | n24552);
assign n23370 = n5297 | n6697;
assign n13146 = n5131 & n19674;
assign n9629 = n20405 | n23113;
assign n5753 = n22197 | n5927;
assign n17146 = ~(n2894 ^ n82);
assign n22308 = n22442 & n22253;
assign n5987 = ~n960;
assign n15812 = ~(n8342 ^ n10906);
assign n7249 = n20596 | n8771;
assign n15024 = n14076 & n8901;
assign n25796 = n16193 | n16001;
assign n3995 = n17664 & n5115;
assign n13978 = n26717 | n20020;
assign n2344 = n5079 | n5008;
assign n19046 = n4490 & n13167;
assign n6055 = ~(n20597 ^ n21623);
assign n26269 = ~(n2312 ^ n25891);
assign n15469 = ~(n11089 ^ n4955);
assign n3793 = n15013 & n17961;
assign n11133 = ~(n23161 | n22237);
assign n22816 = n6750 | n19058;
assign n2873 = n23676 & n5287;
assign n3418 = n5688 | n6680;
assign n1473 = n21674 | n22597;
assign n24349 = n1841 | n25127;
assign n18332 = ~(n25496 ^ n26566);
assign n1938 = n22743 & n4708;
assign n8217 = ~(n11028 ^ n7817);
assign n7680 = ~n12766;
assign n14412 = ~(n25497 ^ n470);
assign n13738 = n11927 & n14876;
assign n17639 = ~(n20052 ^ n4182);
assign n21118 = ~n22879;
assign n16892 = n840 | n24620;
assign n12719 = n24375 | n25119;
assign n5008 = n2936 & n20430;
assign n14472 = ~(n20053 | n18395);
assign n854 = n9082 & n24346;
assign n24245 = ~(n18461 ^ n11841);
assign n20977 = n25142 | n3828;
assign n269 = n11390 & n7970;
assign n14213 = n21133 | n25387;
assign n27195 = ~(n9509 ^ n9554);
assign n25506 = ~(n4901 | n20051);
assign n24 = n24143 & n12420;
assign n23186 = n445 & n10142;
assign n4230 = ~n3878;
assign n12219 = ~(n14684 ^ n1667);
assign n16626 = ~(n26936 ^ n20718);
assign n857 = ~(n21081 ^ n24004);
assign n8836 = ~(n6658 | n20141);
assign n21325 = ~n4937;
assign n10790 = ~(n12751 ^ n20982);
assign n19385 = ~(n6994 ^ n19542);
assign n6709 = n8958 & n21014;
assign n5291 = n19516 | n16412;
assign n13667 = ~(n17259 ^ n7211);
assign n10580 = n14336 | n7952;
assign n2067 = n11656 | n1970;
assign n7093 = n25024 | n25681;
assign n13041 = n26756 & n26862;
assign n3389 = n5379 & n3703;
assign n432 = n14747 | n21445;
assign n16693 = ~n23509;
assign n8326 = n19446 | n3931;
assign n8803 = ~(n8995 ^ n25925);
assign n6269 = n17378 | n16603;
assign n8270 = ~(n9180 | n15884);
assign n9484 = n7130 | n12851;
assign n6935 = ~n20413;
assign n15672 = ~(n24821 ^ n5706);
assign n26474 = n14936 | n20423;
assign n24148 = ~(n2482 ^ n26149);
assign n3102 = n11912 & n11421;
assign n3540 = ~n26725;
assign n24703 = n20173 | n7829;
assign n16700 = n18922 & n4455;
assign n26325 = ~(n14140 | n20822);
assign n16691 = n4657 | n26617;
assign n19433 = ~n19388;
assign n673 = n11126 & n23906;
assign n21301 = n12342 | n4811;
assign n12390 = ~(n16521 ^ n7139);
assign n14329 = n1406 | n6502;
assign n9208 = ~(n19058 ^ n16439);
assign n9835 = ~(n4434 ^ n13453);
assign n6984 = n2790 | n5517;
assign n901 = n3490 | n666;
assign n25152 = n13253 & n22276;
assign n20557 = ~(n16018 ^ n1435);
assign n16796 = n5036 | n23882;
assign n23289 = ~(n21461 ^ n26169);
assign n10854 = ~(n22436 ^ n100);
assign n25277 = ~(n14719 ^ n24215);
assign n3711 = ~(n12626 ^ n4272);
assign n1189 = n16712 | n17664;
assign n4595 = ~(n9338 ^ n4585);
assign n24084 = n11312 | n2568;
assign n25524 = ~n9832;
assign n15433 = ~n17664;
assign n23742 = n18710 | n15355;
assign n23818 = ~(n8266 | n13495);
assign n12179 = ~(n10892 ^ n721);
assign n22774 = ~n21763;
assign n1620 = ~(n22640 ^ n2013);
assign n10784 = n12354 | n22392;
assign n15852 = ~(n4964 | n8259);
assign n12084 = n15084 | n21161;
assign n3013 = ~(n26805 | n18404);
assign n17357 = n10131 | n3690;
assign n17299 = ~(n3500 ^ n12905);
assign n16063 = n20471 | n15308;
assign n19422 = ~(n9605 | n11806);
assign n24844 = ~(n15901 | n10220);
assign n3553 = n21580 & n16229;
assign n6630 = ~(n16990 ^ n20480);
assign n882 = n25094 | n3049;
assign n5279 = ~(n15153 ^ n9340);
assign n18504 = ~(n918 ^ n11356);
assign n9492 = ~(n21606 | n26422);
assign n16960 = ~n2316;
assign n13577 = ~n11302;
assign n19232 = n16101 | n8034;
assign n13346 = n13561 | n12593;
assign n22609 = ~n25196;
assign n18653 = ~(n16021 ^ n6550);
assign n2112 = ~(n3606 ^ n24643);
assign n10536 = n12576 | n18563;
assign n22498 = ~(n26050 ^ n10372);
assign n8906 = ~(n23470 ^ n2021);
assign n2500 = ~(n20923 | n11871);
assign n1589 = ~(n655 ^ n5386);
assign n9990 = ~(n23427 ^ n3795);
assign n8599 = n535 & n2705;
assign n11967 = ~(n20972 ^ n1895);
assign n24183 = ~n27100;
assign n7079 = ~(n24209 ^ n18339);
assign n22443 = ~(n27099 | n24367);
assign n24519 = ~n24886;
assign n8978 = n4479 | n11986;
assign n14691 = ~(n7373 ^ n3480);
assign n19208 = ~(n7693 ^ n7566);
assign n23376 = n15209 | n5952;
assign n14328 = n8569 | n10791;
assign n9114 = ~n26741;
assign n25659 = ~(n26446 ^ n12433);
assign n1296 = n12238 | n11518;
assign n26918 = ~(n12944 | n6864);
assign n4129 = ~(n1654 ^ n4256);
assign n9467 = ~(n1532 ^ n15058);
assign n11267 = ~(n9494 ^ n9227);
assign n7514 = ~(n13526 ^ n17713);
assign n13152 = ~n3828;
assign n1779 = ~n9151;
assign n17474 = n11098 & n15175;
assign n7120 = n26344 | n27146;
assign n18484 = n3863 & n21204;
assign n7965 = n10028 | n20682;
assign n8711 = ~(n15114 | n25389);
assign n25249 = ~(n12241 ^ n3986);
assign n25364 = n13127 & n1828;
assign n18954 = ~(n23200 | n6122);
assign n23802 = n4212 & n549;
assign n22329 = n24638 & n12057;
assign n12603 = ~(n3037 | n14385);
assign n23426 = n3097 & n3764;
assign n10231 = n14248 & n24108;
assign n23724 = ~n1991;
assign n12778 = n2914 & n13449;
assign n17700 = ~(n2894 ^ n12675);
assign n23432 = n18028 | n1785;
assign n7971 = n8099 | n17426;
assign n16110 = ~(n16363 ^ n19396);
assign n21924 = ~(n3102 ^ n16574);
assign n4607 = n14369 | n4549;
assign n13129 = ~n15142;
assign n24992 = ~(n14736 ^ n3529);
assign n8501 = ~(n4715 | n16507);
assign n15202 = ~n15979;
assign n18193 = ~(n19764 ^ n722);
assign n24671 = ~n14637;
assign n2959 = n22105 | n23277;
assign n14362 = ~(n24351 | n12113);
assign n7085 = n11413 | n15509;
assign n24720 = n16881 | n4167;
assign n17983 = n8948 | n14680;
assign n23583 = ~n25609;
assign n18732 = n12093 | n3535;
assign n9850 = n11112 | n26817;
assign n344 = n19754 | n11308;
assign n9226 = ~n3623;
assign n15558 = ~(n9265 ^ n14355);
assign n22839 = n10659 | n23126;
assign n18946 = n19161 | n19254;
assign n17689 = ~(n14148 ^ n11503);
assign n23868 = n17605 & n4263;
assign n9292 = n23720 | n17186;
assign n3901 = ~(n25533 ^ n23854);
assign n12479 = ~(n18290 ^ n12875);
assign n14268 = ~n10843;
assign n23953 = ~(n19330 | n19703);
assign n22519 = n16465 & n5449;
assign n15973 = n23339 & n16950;
assign n20084 = ~(n22747 ^ n26438);
assign n22229 = n11690 | n1914;
assign n3872 = ~(n23512 ^ n6341);
assign n21647 = ~(n11441 | n7688);
assign n21802 = n24791 | n2291;
assign n294 = ~(n26334 | n8792);
assign n16995 = ~(n6218 | n25464);
assign n22909 = ~(n24104 ^ n3344);
assign n5607 = ~(n4609 ^ n170);
assign n22435 = ~(n13471 ^ n15879);
assign n23701 = n7259 & n2019;
assign n3642 = ~(n10396 ^ n7526);
assign n193 = ~(n10274 | n8052);
assign n22795 = ~(n24663 ^ n26224);
assign n15729 = n8713 | n54;
assign n16282 = n13083 & n4131;
assign n9301 = n12002 | n27102;
assign n10185 = n15977 | n5638;
assign n10695 = n8621 & n7760;
assign n11345 = n16030 | n14916;
assign n8065 = ~(n5728 ^ n12265);
assign n24713 = n15738 | n17490;
assign n19842 = ~(n11427 ^ n17972);
assign n19358 = ~(n15813 ^ n15671);
assign n22110 = ~n800;
assign n400 = ~(n23701 ^ n23100);
assign n7671 = ~(n24163 ^ n7138);
assign n320 = ~(n16937 | n16971);
assign n1003 = ~n19372;
assign n25838 = ~n8643;
assign n7358 = ~(n4436 ^ n13297);
assign n14205 = n8367 | n5203;
assign n2784 = ~(n17301 ^ n27132);
assign n17333 = ~(n313 ^ n11463);
assign n13804 = n446 | n21839;
assign n3665 = ~(n2634 ^ n4163);
assign n15879 = ~(n1662 ^ n20946);
assign n24000 = n11455 & n14870;
assign n16462 = n8568 & n1600;
assign n16503 = ~(n19646 ^ n19770);
assign n1243 = ~(n11119 ^ n26863);
assign n2862 = ~n2355;
assign n56 = ~n6478;
assign n3138 = ~n5789;
assign n2708 = n22724 | n24939;
assign n5163 = ~n3445;
assign n15635 = ~(n17982 ^ n20986);
assign n14703 = n21 & n23513;
assign n6787 = ~(n11006 ^ n23457);
assign n24302 = ~n8371;
assign n5712 = n25144 & n5972;
assign n15657 = n1769 & n11076;
assign n2173 = ~(n18440 ^ n21914);
assign n20761 = ~(n22257 ^ n17859);
assign n21013 = ~(n7341 ^ n11254);
assign n19831 = n9294 | n11351;
assign n24922 = n26452 | n21025;
assign n5493 = ~(n16642 ^ n19630);
assign n8886 = ~(n17854 | n23724);
assign n5318 = ~n2184;
assign n15740 = ~(n987 | n626);
assign n2863 = n21021 | n18355;
assign n1354 = ~(n11121 ^ n19494);
assign n7095 = n644 & n12868;
assign n13435 = ~n21596;
assign n6145 = ~(n16476 ^ n15539);
assign n26050 = ~(n864 ^ n17684);
assign n24547 = n20112 | n847;
assign n23140 = ~(n18341 ^ n19680);
assign n6816 = n16784 & n15500;
assign n21020 = n8872 & n17443;
assign n15501 = ~(n4636 ^ n6263);
assign n10129 = ~(n26946 ^ n978);
assign n21177 = n8244 & n8431;
assign n17688 = ~(n17536 | n19060);
assign n24336 = n17949 | n22033;
assign n14358 = n3836 | n4459;
assign n12623 = ~(n20429 ^ n12587);
assign n6448 = ~(n17088 | n5241);
assign n584 = n221 & n10523;
assign n7281 = ~n690;
assign n10203 = n24222 & n15091;
assign n1745 = n4230 | n16290;
assign n12203 = ~(n1243 ^ n6698);
assign n3721 = n13804 & n26759;
assign n17691 = n16241 | n3885;
assign n12579 = ~(n16924 | n8624);
assign n1388 = n21351 & n20587;
assign n7918 = ~(n19392 ^ n18901);
assign n25243 = ~(n23286 ^ n13004);
assign n17479 = ~n5579;
assign n10575 = n13967 | n9788;
assign n19447 = n20518 | n10922;
assign n2487 = n14336 & n9349;
assign n16445 = ~(n21601 ^ n26776);
assign n25563 = n4066 & n23439;
assign n16564 = n1037 | n233;
assign n8281 = n3734 & n14257;
assign n15619 = n1508 | n23314;
assign n19729 = n6075 & n23733;
assign n11681 = n13016 | n13226;
assign n22730 = ~(n19862 | n10155);
assign n20824 = ~(n12286 ^ n6525);
assign n3403 = ~n2757;
assign n23579 = n26904 | n10250;
assign n15555 = ~(n27030 ^ n15057);
assign n12395 = ~(n7098 ^ n7820);
assign n23002 = n11416;
assign n9368 = n1278 & n19956;
assign n23570 = n14816 | n12744;
assign n15222 = n11454 | n19364;
assign n22304 = ~(n4108 ^ n18148);
assign n24639 = n1181 | n14458;
assign n1743 = n5165 | n12889;
assign n170 = ~(n23529 ^ n20700);
assign n9013 = n20201 | n20231;
assign n12763 = ~n23683;
assign n12296 = ~n15047;
assign n14552 = n12703 & n5959;
assign n14545 = ~n5549;
assign n13373 = ~(n13853 ^ n18157);
assign n6941 = n738 & n1920;
assign n7983 = ~n18904;
assign n14265 = ~(n13977 ^ n20148);
assign n4772 = n25886 | n2862;
assign n19380 = n2038 | n2574;
assign n9830 = ~n25918;
assign n24287 = n15248 | n1014;
assign n18550 = n18946 & n6322;
assign n9679 = ~n8856;
assign n19325 = n8269 & n21757;
assign n14040 = ~(n21872 ^ n3041);
assign n25604 = ~n15867;
assign n17746 = ~(n1046 ^ n9213);
assign n16249 = ~(n25860 ^ n4961);
assign n14086 = ~(n22247 | n19502);
assign n5102 = n17226 | n2984;
assign n11783 = n27159 & n19929;
assign n9170 = n12593 | n13714;
assign n24978 = n5025 & n23162;
assign n8668 = ~n2664;
assign n9517 = n13474 | n20462;
assign n360 = ~n1842;
assign n22199 = n12443 | n10664;
assign n8773 = ~(n8304 ^ n18771);
assign n2822 = n18891 | n16364;
assign n24780 = n2597 | n10682;
assign n12708 = ~(n16092 | n2279);
assign n8511 = ~(n6570 ^ n25684);
assign n7531 = n8311 & n8062;
assign n7444 = n17598 & n17926;
assign n15594 = ~(n10092 ^ n12657);
assign n15895 = ~(n15826 | n21585);
assign n4987 = n8916 & n25473;
assign n26020 = n17118 | n23730;
assign n1121 = ~(n17311 ^ n14172);
assign n19087 = ~(n25378 ^ n26630);
assign n16360 = ~(n26091 ^ n12667);
assign n18337 = ~(n4246 ^ n14511);
assign n24254 = n4889 & n8263;
assign n2645 = ~n21728;
assign n13755 = ~(n7587 ^ n18745);
assign n13051 = n14915 & n22997;
assign n23712 = n2549 & n3998;
assign n8409 = ~(n9200 ^ n2540);
assign n26459 = n7146 & n3549;
assign n26551 = ~(n4715 | n10117);
assign n15176 = ~(n18205 ^ n80);
assign n15907 = n7742 | n11853;
assign n2315 = n13858 | n5445;
assign n17373 = ~(n19350 | n24331);
assign n8336 = n537 & n21221;
assign n10008 = ~n22335;
assign n12436 = ~(n23699 ^ n11844);
assign n9131 = n12351 | n6503;
assign n6613 = n14627 | n21259;
assign n9095 = ~n23541;
assign n7689 = ~n9888;
assign n24572 = n15905 & n2510;
assign n26277 = n19351 | n11863;
assign n13071 = ~n2109;
assign n6763 = n2500 | n11718;
assign n7681 = ~(n13027 | n24929);
assign n6440 = n23739 & n24498;
assign n22783 = ~n82;
assign n1113 = ~(n26914 ^ n14620);
assign n18152 = ~(n7315 ^ n12705);
assign n528 = ~n23842;
assign n11467 = ~(n10823 ^ n11194);
assign n9683 = ~n10919;
assign n12202 = n19361 & n20060;
assign n15183 = n8525 | n4754;
assign n21797 = ~(n14365 ^ n25516);
assign n20996 = ~(n27200 ^ n2583);
assign n1959 = ~(n10500 | n12493);
assign n295 = ~n25252;
assign n1824 = n5757 & n20818;
assign n3520 = n6204 | n23254;
assign n17867 = ~n5779;
assign n2563 = ~(n2242 | n12810);
assign n11658 = ~(n23936 ^ n17620);
assign n7231 = ~(n2418 ^ n6303);
assign n10362 = ~(n21929 ^ n9575);
assign n21460 = ~n21736;
assign n12003 = ~(n3427 ^ n24793);
assign n4624 = ~(n22245 ^ n9268);
assign n6872 = ~(n17604 ^ n25102);
assign n10140 = n2272 | n26927;
assign n21825 = ~(n18978 ^ n25576);
assign n2899 = ~(n372 ^ n5085);
assign n13176 = ~(n18113 ^ n10557);
assign n23449 = n12845 | n3623;
assign n8463 = n2421 | n11243;
assign n2464 = n26130 | n3661;
assign n10704 = ~(n21693 | n15875);
assign n18372 = ~(n8455 ^ n13727);
assign n9130 = ~n16240;
assign n16675 = ~(n7731 ^ n2328);
assign n26773 = n12480 | n7318;
assign n13199 = ~(n18536 ^ n8577);
assign n17290 = n21764 | n23900;
assign n2812 = ~n2145;
assign n9534 = ~n7340;
assign n23807 = ~n8906;
assign n3461 = ~(n16547 ^ n19872);
assign n7477 = ~(n24137 ^ n18943);
assign n1570 = ~(n9246 ^ n7139);
assign n19235 = n4545 | n1297;
assign n10989 = ~n34;
assign n22642 = ~n20374;
assign n22065 = n21336 & n5536;
assign n5117 = ~(n24318 ^ n2013);
assign n16002 = ~n6104;
assign n20710 = n10971 | n17241;
assign n3670 = n24245 & n3138;
assign n2438 = ~(n17035 ^ n2680);
assign n19910 = n1565 | n1893;
assign n4359 = ~(n22634 | n26942);
assign n5281 = n17507 | n6277;
assign n8834 = ~(n16707 ^ n21749);
assign n19932 = ~(n10168 ^ n7267);
assign n11531 = n11404 | n12804;
assign n17061 = ~n14584;
assign n26608 = ~(n5538 ^ n20234);
assign n2544 = n13618 | n2213;
assign n2745 = n13734 | n6019;
assign n1018 = n12301 & n26467;
assign n22738 = ~(n8499 ^ n17314);
assign n11977 = n23133 | n23252;
assign n5968 = ~(n22210 | n24496);
assign n23616 = ~n25059;
assign n5553 = ~(n14163 | n15512);
assign n12378 = n10181 | n11056;
assign n19159 = ~n12912;
assign n8297 = ~(n6538 ^ n9847);
assign n7295 = ~(n6079 ^ n26168);
assign n6873 = ~(n10903 ^ n4767);
assign n3865 = ~(n12631 | n2867);
assign n5322 = n7642 | n25907;
assign n3420 = n14612 & n1400;
assign n22917 = ~(n23187 | n20031);
assign n12407 = ~(n6955 | n19390);
assign n13876 = n25271 | n21649;
assign n19438 = n23974 & n17013;
assign n23547 = n4505 | n24757;
assign n17147 = ~(n4775 ^ n49);
assign n3813 = ~(n12639 | n24091);
assign n6473 = n892 & n10888;
assign n4867 = ~(n8446 ^ n21940);
assign n1503 = ~(n25063 ^ n11898);
assign n15468 = n6146 & n4456;
assign n8663 = n2640 | n3476;
assign n20989 = n15891 & n9319;
assign n21135 = n23896 | n11595;
assign n17347 = n10117 & n19825;
assign n24755 = ~(n12797 | n22327);
assign n25686 = n951 | n7498;
assign n7794 = ~(n18436 ^ n13759);
assign n461 = ~(n14425 ^ n10638);
assign n8988 = ~(n11371 ^ n3370);
assign n16218 = ~(n16636 ^ n1114);
assign n501 = ~(n23482 ^ n3616);
assign n19239 = ~n12281;
assign n21974 = ~n1269;
assign n4852 = ~(n2856 | n15798);
assign n15752 = n6821 & n17527;
assign n13141 = ~(n14447 ^ n1604);
assign n5446 = ~(n7837 | n1973);
assign n5824 = n14853 & n5423;
assign n1160 = n22937 & n1676;
assign n343 = ~(n21747 | n26422);
assign n209 = ~n10254;
assign n3578 = n3936 | n16328;
assign n26695 = ~n14684;
assign n13501 = ~(n23518 ^ n6902);
assign n13149 = n26341 | n11204;
assign n23565 = ~(n6935 ^ n25194);
assign n1837 = ~(n5149 ^ n26024);
assign n2016 = n356 | n1606;
assign n2290 = ~(n14680 ^ n5031);
assign n26072 = ~(n17379 ^ n12421);
assign n10632 = n23160 & n13863;
assign n18316 = n12880 | n16229;
assign n24748 = n11011 | n10217;
assign n4870 = ~(n18948 ^ n5096);
assign n25792 = ~(n10879 ^ n12413);
assign n1659 = n15748 | n21882;
assign n21596 = n18893 | n2913;
assign n23633 = n15069 & n20157;
assign n17739 = ~(n5565 ^ n20500);
assign n9325 = n13263 & n22596;
assign n6695 = n24590 | n20835;
assign n23787 = ~(n6711 ^ n2117);
assign n5638 = ~(n25926 | n9646);
assign n7522 = n14654 | n10577;
assign n872 = n25088 | n5837;
assign n15617 = ~(n21580 ^ n18446);
assign n22102 = n11733 | n14215;
assign n3357 = n6416 | n9229;
assign n19851 = ~(n23076 ^ n17511);
assign n25485 = ~n25547;
assign n2118 = n21083 | n25974;
assign n6819 = ~(n12807 ^ n12966);
assign n23841 = n16848 | n11356;
assign n16820 = ~(n5905 | n8167);
assign n16805 = n12553 | n14872;
assign n15114 = ~n22290;
assign n24745 = ~(n24800 ^ n22463);
assign n7183 = ~n2471;
assign n26535 = n24583 & n9063;
assign n3106 = n10526 & n14512;
assign n14834 = n20836 | n13961;
assign n23484 = n5400 & n3149;
assign n9721 = n23237 | n9551;
assign n14405 = ~n22885;
assign n4924 = n16865 & n8470;
assign n15838 = n26433 | n690;
assign n3613 = n25286 & n9769;
assign n12521 = n16573 | n1714;
assign n16413 = n24006 & n25363;
assign n3003 = n322 & n23934;
assign n4681 = n17584 | n3425;
assign n18024 = ~(n18184 ^ n19572);
assign n18770 = ~n6725;
assign n11880 = ~(n12161 | n3072);
assign n12212 = ~n8645;
assign n11172 = n3837 & n12184;
assign n26549 = n2170 & n9811;
assign n4997 = n15577 | n13552;
assign n12307 = ~(n12363 | n18468);
assign n4404 = ~(n7821 ^ n25128);
assign n567 = ~(n10016 ^ n2401);
assign n5216 = n20371 | n8445;
assign n2140 = ~(n20937 ^ n424);
assign n11106 = n25523 | n25455;
assign n14338 = n619 | n14880;
assign n13879 = n8867 & n18411;
assign n15262 = n12961 | n2551;
assign n7142 = n24311 & n17430;
assign n15645 = ~(n10710 ^ n9372);
assign n5236 = ~(n5438 ^ n13714);
assign n2549 = n4941 | n9749;
assign n3791 = ~n1662;
assign n14819 = ~(n9543 ^ n6480);
assign n1927 = ~(n8431 ^ n21547);
assign n12453 = ~n7030;
assign n14049 = n23489 | n20134;
assign n24350 = n11523 | n6380;
assign n9382 = n12565 & n9280;
assign n16171 = n6978 & n6740;
assign n24166 = ~(n10320 ^ n3924);
assign n3207 = ~(n18797 ^ n24280);
assign n1069 = ~(n17821 ^ n2295);
assign n2408 = n15331 & n18638;
assign n19985 = ~(n818 ^ n9942);
assign n21891 = ~n4981;
assign n24375 = ~n23923;
assign n21144 = ~(n20060 ^ n19361);
assign n25411 = n15146 | n5532;
assign n7172 = ~(n5598 ^ n19728);
assign n6569 = ~(n5266 | n3724);
assign n2277 = n2056 | n14615;
assign n26206 = ~(n1803 ^ n5521);
assign n20163 = ~(n25972 ^ n10250);
assign n12443 = ~(n10125 | n18326);
assign n26723 = n12090 & n8487;
assign n12304 = ~(n21938 ^ n8072);
assign n13996 = n25669 | n1453;
assign n19847 = n16547 & n15;
assign n6266 = n21994 | n20465;
assign n16050 = n26230 | n19101;
assign n1166 = n11246 | n14974;
assign n21836 = n26034 & n13726;
assign n25998 = ~n21522;
assign n16354 = ~(n6204 ^ n7674);
assign n16899 = n895 & n5565;
assign n14655 = n6743 ^ n20385;
assign n5999 = n26064 & n10930;
assign n16327 = ~(n26033 ^ n5126);
assign n6098 = ~(n12673 ^ n2300);
assign n4437 = n3085 | n24747;
assign n5757 = n17539 | n16524;
assign n6952 = n12525 | n20928;
assign n22672 = n1099 | n3379;
assign n17371 = ~(n7913 ^ n14090);
assign n8455 = ~(n7875 ^ n3063);
assign n6267 = ~n12964;
assign n18556 = n6206 | n9708;
assign n20439 = n10438 | n23947;
assign n12721 = ~(n9615 ^ n19737);
assign n18194 = n16754 & n9374;
assign n23325 = ~(n19218 ^ n14957);
assign n13712 = n19588 | n19549;
assign n13676 = n8743 | n11468;
assign n18160 = n26891 | n8613;
assign n13375 = ~(n20271 ^ n10229);
assign n27169 = n18992 | n7454;
assign n4420 = n11938 | n3614;
assign n6253 = n19429 & n14610;
assign n5976 = ~(n26218 ^ n3480);
assign n25380 = ~(n16117 ^ n8891);
assign n20330 = n13918 & n20810;
assign n10046 = n7631 & n2673;
assign n5421 = n1713 & n14445;
assign n25912 = n3601 | n22456;
assign n18172 = n20700 & n26240;
assign n7430 = ~(n8211 ^ n16811);
assign n1951 = ~n11893;
assign n7443 = n26649 | n3980;
assign n12183 = n14580 & n14195;
assign n14045 = ~(n15106 ^ n10508);
assign n8786 = n22365 & n23122;
assign n22837 = n2342 | n5213;
assign n5223 = ~(n11736 | n10995);
assign n13739 = ~n10875;
assign n14447 = n21334 & n18399;
assign n9391 = ~(n24074 ^ n21969);
assign n23195 = n18632 | n2608;
assign n23779 = ~(n2530 ^ n26572);
assign n15522 = n16856 & n21081;
assign n14673 = n14703 | n9221;
assign n10621 = n9014 | n16208;
assign n15834 = ~(n11667 ^ n21398);
assign n21574 = n8466 | n10082;
assign n9815 = n11074 & n21872;
assign n7996 = ~(n8153 ^ n19355);
assign n16848 = ~n2999;
assign n13283 = ~(n12811 | n3260);
assign n7534 = ~(n1799 ^ n11580);
assign n4372 = n5043 & n24726;
assign n26257 = n25914 | n4941;
assign n7233 = ~(n26049 ^ n15642);
assign n4780 = ~n11775;
assign n22782 = ~(n9037 ^ n23188);
assign n15223 = ~(n12278 | n73);
assign n549 = n7524 | n10314;
assign n3641 = ~(n10410 ^ n5493);
assign n17205 = ~(n5006 | n9372);
assign n3231 = ~(n20595 | n2322);
assign n21655 = n23979 | n2690;
assign n7690 = n6923 | n21647;
assign n16831 = n21902 & n7154;
assign n71 = ~(n14486 ^ n16744);
assign n1701 = ~(n4805 ^ n25416);
assign n23965 = ~(n24617 ^ n6988);
assign n24818 = ~n20092;
assign n14292 = n14958 & n23822;
assign n24875 = ~(n13829 ^ n6145);
assign n428 = ~n22122;
assign n3247 = ~(n22520 ^ n6974);
assign n520 = n4678 & n17377;
assign n21354 = n17728 ^ n23586;
assign n22936 = n8628 & n1035;
assign n12076 = ~n19768;
assign n19778 = n10839 | n22293;
assign n24411 = n11745 | n6825;
assign n2537 = ~(n11620 ^ n17796);
assign n3953 = n13389 | n20536;
assign n3550 = n2247 & n19715;
assign n12751 = ~(n23376 ^ n19882);
assign n17106 = ~(n16300 ^ n5392);
assign n10137 = n22743 | n4708;
assign n24708 = ~(n7693 ^ n19472);
assign n25158 = n13417 | n23026;
assign n10312 = ~n9314;
assign n26143 = n2871 & n18376;
assign n3669 = ~(n25629 ^ n3795);
assign n22081 = n23650 | n25115;
assign n17181 = n14683 | n26010;
assign n14024 = n23065 & n27055;
assign n15867 = ~(n16570 ^ n8214);
assign n24053 = n19941 | n9345;
assign n19574 = n24638 | n12057;
assign n6126 = ~n17426;
assign n20937 = ~n25772;
assign n19516 = ~(n4409 | n25967);
assign n5768 = ~(n14116 ^ n12012);
assign n2254 = n26452 | n2999;
assign n21126 = ~n14782;
assign n648 = n26063 & n14115;
assign n26621 = n1293 | n15921;
assign n11522 = n26725 & n17212;
assign n11416 = ~(n3093 ^ n25264);
assign n4808 = n714 & n25357;
assign n15783 = ~(n24929 ^ n13027);
assign n480 = n12979 & n986;
assign n20807 = n5650 | n16360;
assign n19771 = n15850 | n22206;
assign n22975 = n11600 & n16843;
assign n26000 = n2743 | n16312;
assign n20278 = ~(n2659 ^ n11926);
assign n4604 = n13671 | n10275;
assign n27136 = ~(n11152 | n21735);
assign n15921 = ~n27193;
assign n6331 = n22475 | n22794;
assign n2739 = n8450 & n23042;
assign n23153 = ~(n9096 | n25937);
assign n7068 = n3878 | n20755;
assign n23892 = ~(n10153 ^ n15737);
assign n9296 = ~n14761;
assign n1227 = ~(n5208 ^ n2387);
assign n22988 = ~(n25581 | n1210);
assign n26583 = ~(n12669 ^ n10233);
assign n15345 = ~(n17668 ^ n6392);
assign n20720 = ~(n19061 ^ n9935);
assign n26411 = ~(n19393 | n21508);
assign n20408 = n11519 & n2681;
assign n439 = n23621 & n23260;
assign n13603 = n9136 & n7136;
assign n15688 = n834 | n4106;
assign n2681 = n27106 | n8264;
assign n9768 = n7353 & n3830;
assign n11756 = ~n12078;
assign n26636 = n14495 | n25251;
assign n4118 = n18681 & n12135;
assign n23464 = ~n12417;
assign n22436 = ~n17095;
assign n14056 = n10522 & n19110;
assign n7169 = ~n10980;
assign n25804 = n19847 | n11878;
assign n22016 = ~(n5301 ^ n23319);
assign n4663 = n16426 & n16774;
assign n23286 = n13938 | n17489;
assign n4552 = ~(n19600 ^ n14278);
assign n13009 = n1793 | n10702;
assign n4898 = ~(n27143 ^ n4371);
assign n20044 = ~(n8715 ^ n10611);
assign n9424 = n3945 & n3393;
assign n11186 = ~n2035;
assign n11404 = n20323 & n11118;
assign n8766 = n20425 | n12332;
assign n17383 = ~(n17408 ^ n4326);
assign n21584 = ~(n17397 ^ n5077);
assign n26901 = ~(n9251 ^ n22309);
assign n20336 = ~(n20244 ^ n27134);
assign n6921 = ~(n18451 ^ n13081);
assign n7559 = n11725 | n14075;
assign n7117 = ~(n11597 ^ n17351);
assign n14496 = n13453 & n4434;
assign n13976 = ~n14584;
assign n11197 = ~(n26363 ^ n1553);
assign n9851 = ~(n10742 ^ n25245);
assign n25739 = ~(n1566 ^ n18711);
assign n13113 = ~(n10383 ^ n2690);
assign n21284 = n13765 | n11540;
assign n19955 = ~(n24730 ^ n16277);
assign n4543 = ~(n7817 | n11028);
assign n13953 = ~n23076;
assign n10485 = ~n2043;
assign n24744 = ~(n18651 ^ n25307);
assign n24263 = ~(n17567 ^ n18628);
assign n23981 = n10117 & n22261;
assign n24957 = n26164 & n24770;
assign n23687 = ~(n13280 | n3136);
assign n21056 = n318 & n23770;
assign n12973 = ~(n24759 ^ n17930);
assign n10445 = n24185 & n12499;
assign n27032 = ~(n19446 ^ n17069);
assign n1460 = n10683 | n10109;
assign n15885 = ~(n4680 ^ n7478);
assign n16844 = ~(n7071 ^ n428);
assign n25695 = n18401 | n8289;
assign n22590 = n12950 | n19210;
assign n22934 = ~(n22001 ^ n4519);
assign n26199 = n21458 | n8891;
assign n10290 = n22395 | n12991;
assign n5414 = ~(n26947 ^ n5231);
assign n4060 = ~(n26706 ^ n21143);
assign n5471 = ~(n26256 ^ n3261);
assign n9129 = ~(n15253 ^ n9984);
assign n15687 = n21964 | n15961;
assign n1104 = ~(n26295 ^ n16896);
assign n22317 = ~(n13498 ^ n23240);
assign n18877 = ~(n18159 ^ n14716);
assign n22771 = ~(n20882 ^ n23685);
assign n5780 = ~(n10451 ^ n16034);
assign n6165 = n9615 & n12774;
assign n23791 = ~n18037;
assign n10223 = n19371 | n18;
assign n5461 = n7226 & n23727;
assign n26910 = n20775 | n20808;
assign n69 = n11133 | n430;
assign n2370 = ~(n14345 ^ n25381);
assign n7549 = n8521 | n4652;
assign n9498 = ~(n23446 ^ n2623);
assign n23517 = ~(n23226 ^ n26150);
assign n26985 = n15296 & n9478;
assign n6057 = n16987 & n11807;
assign n11776 = n17975 & n4202;
assign n22132 = n6814 | n23463;
assign n5713 = n22332 | n4104;
assign n22092 = n8464 & n5248;
assign n26413 = ~n7554;
assign n4786 = n19844 & n12299;
assign n1754 = ~(n13846 ^ n15652);
assign n13514 = n1997 | n11981;
assign n16350 = ~(n18082 ^ n23915);
assign n3259 = n13237 | n14394;
assign n22989 = n26074 & n19753;
assign n929 = n2485 | n1625;
assign n12470 = ~(n634 ^ n4334);
assign n12374 = n1077 | n18731;
assign n19412 = n9907 & n18243;
assign n419 = ~(n22557 | n1952);
assign n10376 = n4368 | n17660;
assign n7929 = n19258 | n9683;
assign n5333 = ~(n4108 ^ n11013);
assign n25455 = n5579 | n26831;
assign n1389 = n8358 & n24344;
assign n2663 = n16261 & n23013;
assign n4675 = ~(n11320 ^ n11252);
assign n11006 = n8442 & n249;
assign n21628 = ~(n12832 ^ n8238);
assign n10464 = ~n2072;
assign n14175 = n6382 | n25577;
assign n15142 = ~(n23961 ^ n7310);
assign n10227 = ~(n25931 | n13053);
assign n8230 = ~n3180;
assign n13606 = n531 | n18769;
assign n7316 = ~n23535;
assign n18871 = n10452 | n25558;
assign n17967 = ~n13518;
assign n18951 = n2731 | n26879;
assign n22789 = ~(n11477 ^ n13915);
assign n5630 = n18334 | n4433;
assign n6472 = n13454 | n20789;
assign n6045 = n17328 | n6947;
assign n12705 = ~(n10509 ^ n26417);
assign n4195 = ~n4499;
assign n15949 = n6474 & n16750;
assign n20383 = ~(n2035 | n2675);
assign n2602 = ~(n22901 ^ n861);
assign n12157 = ~(n20063 ^ n15036);
assign n17930 = ~(n14733 ^ n19905);
assign n23107 = ~(n20127 ^ n23970);
assign n16587 = n22943 | n24380;
assign n19335 = n4496 & n5369;
assign n17311 = ~(n18249 ^ n26219);
assign n9696 = ~n814;
assign n21192 = n23940 | n18541;
assign n26197 = ~n3228;
assign n17960 = ~n9768;
assign n16465 = ~(n4578 ^ n10411);
assign n21294 = ~(n5105 ^ n14790);
assign n23927 = ~n17914;
assign n27202 = n20072 & n3639;
assign n8466 = ~(n15077 | n6486);
assign n8323 = ~(n5596 | n2340);
assign n11328 = ~(n9244 | n10509);
assign n14408 = n4469 & n23545;
assign n14649 = ~(n6057 ^ n10679);
assign n4654 = ~(n14155 | n7339);
assign n9846 = n14574 & n9092;
assign n4978 = ~(n6520 ^ n6837);
assign n9018 = ~n22933;
assign n13848 = ~n4712;
assign n15713 = ~n18251;
assign n12178 = ~(n5337 | n25228);
assign n3000 = n2355 & n16223;
assign n11097 = n24388 | n23927;
assign n214 = n11191 | n4261;
assign n941 = ~(n11578 ^ n2261);
assign n8012 = n4940 | n18409;
assign n15111 = ~(n20084 ^ n13117);
assign n7568 = ~(n5998 ^ n16078);
assign n9509 = ~(n8278 ^ n23166);
assign n17501 = n20470 & n18634;
assign n19529 = ~n3147;
assign n20859 = ~(n16458 ^ n8685);
assign n723 = ~(n19666 ^ n6148);
assign n9789 = ~n21050;
assign n8986 = ~(n20358 ^ n3960);
assign n7785 = ~n17305;
assign n26633 = n16750 | n19828;
assign n23659 = ~(n25749 ^ n7377);
assign n13463 = ~(n4744 ^ n1999);
assign n4416 = n15863 & n5239;
assign n4303 = n743 | n20861;
assign n11339 = ~(n690 | n25700);
assign n4563 = n11294 | n24732;
assign n10127 = ~(n21749 ^ n26744);
assign n8498 = ~(n22083 | n26499);
assign n4695 = ~(n5167 ^ n6773);
assign n18857 = ~(n15767 | n19658);
assign n13857 = ~(n14148 | n14275);
assign n11143 = ~n632;
assign n25101 = ~n16239;
assign n14404 = ~(n5669 | n21575);
assign n20041 = n14631 | n19769;
assign n15793 = ~(n13836 ^ n15065);
assign n10622 = ~n22191;
assign n7209 = ~(n22197 ^ n16459);
assign n23352 = ~n12445;
assign n11931 = n9023 | n12307;
assign n18938 = n25068 | n8324;
assign n8522 = ~n19840;
assign n16849 = ~(n9789 ^ n19762);
assign n1316 = ~(n20151 ^ n17959);
assign n3232 = n3018 | n9185;
assign n19466 = n11694 & n18040;
assign n11941 = n22776 | n18767;
assign n371 = ~(n11736 | n2320);
assign n10944 = ~(n7060 | n13821);
assign n10887 = n12376 & n22967;
assign n10181 = ~n20478;
assign n8540 = ~(n3881 ^ n3964);
assign n189 = ~n24654;
assign n18492 = n25169 & n15078;
assign n4715 = ~n23250;
assign n26447 = ~n25249;
assign n25338 = n22745 | n10198;
assign n21216 = ~(n26895 ^ n12315);
assign n1791 = ~(n17793 ^ n24881);
assign n12314 = ~(n23913 ^ n16376);
assign n5387 = ~(n950 ^ n22789);
assign n9314 = ~(n473 ^ n6430);
assign n4187 = n3542 | n2014;
assign n23637 = ~(n4668 ^ n18373);
assign n5424 = ~(n18739 ^ n3911);
assign n20441 = ~(n2953 ^ n10996);
assign n4289 = n3294 & n14177;
assign n10446 = ~n10383;
assign n26232 = ~(n4719 ^ n23582);
assign n4754 = n14034 & n24546;
assign n10192 = ~(n401 | n3030);
assign n5250 = n9352 & n6269;
assign n2241 = n8851 | n15212;
assign n15473 = n22254 & n22699;
assign n10508 = ~(n14130 ^ n12861);
assign n23505 = ~(n16738 ^ n12860);
assign n6557 = n16351 | n2721;
assign n136 = n3199 | n3373;
assign n18664 = ~(n13185 ^ n1450);
assign n25876 = ~(n13154 | n15891);
assign n27145 = ~(n6197 ^ n2149);
assign n13961 = n17890 & n6009;
assign n20650 = n26417 | n11482;
assign n9223 = n19161 & n22405;
assign n3542 = n13171 & n13633;
assign n11940 = n15021 & n11663;
assign n2495 = ~(n16443 | n13166);
assign n3752 = ~n12274;
assign n23418 = n20367 & n13630;
assign n8652 = n20878 & n13024;
assign n7242 = ~n21860;
assign n1412 = n9854 | n14955;
assign n732 = ~(n15534 ^ n25572);
assign n10190 = ~(n14750 | n12470);
assign n12174 = n15416 & n13554;
assign n16598 = n13353 | n12317;
assign n10224 = ~(n13811 ^ n18454);
assign n1586 = ~(n12456 ^ n5404);
assign n1169 = ~(n15546 ^ n24937);
assign n26731 = n4119 & n9310;
assign n5093 = ~(n13303 ^ n12546);
assign n25842 = n21711 & n9630;
assign n24395 = n11111 | n286;
assign n8884 = ~(n23112 ^ n20443);
assign n26201 = ~n12502;
assign n26641 = ~(n19415 ^ n15874);
assign n14242 = n21649 | n17846;
assign n20581 = ~(n2481 | n23201);
assign n18199 = n23376 & n26108;
assign n8935 = ~n18002;
assign n14125 = ~(n3501 ^ n6152);
assign n21389 = n5329 | n2694;
assign n20268 = ~(n19911 ^ n14570);
assign n5849 = ~(n15182 | n21915);
assign n1333 = n10997 | n16486;
assign n8035 = n9517 & n18015;
assign n15353 = ~(n6598 ^ n14063);
assign n23319 = ~(n5238 ^ n9456);
assign n9929 = n8852 & n7888;
assign n27130 = ~(n8478 ^ n7905);
assign n24282 = ~(n8292 | n5916);
assign n17414 = ~n13089;
assign n13692 = n3423 | n21065;
assign n10719 = ~(n25505 | n23843);
assign n19058 = ~(n26182 ^ n12314);
assign n3459 = ~(n20769 ^ n4756);
assign n16888 = n9003 | n11876;
assign n19819 = n22141 & n6886;
assign n22614 = ~n2958;
assign n25574 = ~(n14557 ^ n16249);
assign n9063 = n23848 | n26792;
assign n24750 = ~n7186;
assign n26702 = n12572 | n8063;
assign n11206 = ~(n9096 ^ n6127);
assign n14744 = n940 | n25787;
assign n744 = ~n4588;
assign n14540 = n21937 | n7953;
assign n8384 = n15894 | n7329;
assign n23271 = ~n2111;
assign n20305 = n8680 | n11192;
assign n16908 = n4287 & n1670;
assign n8086 = n16896 | n781;
assign n898 = ~(n8875 | n18655);
assign n13693 = ~n16886;
assign n7709 = ~n25808;
assign n12110 = ~n26135;
assign n18158 = ~n15996;
assign n6008 = n4676 | n8980;
assign n2137 = n11455 & n9940;
assign n22777 = n6843 | n14871;
assign n23018 = ~n16696;
assign n18423 = n14818 | n16631;
assign n18404 = ~n21948;
assign n19654 = n3807 | n12536;
assign n15280 = ~(n5196 ^ n1878);
assign n6766 = n21557 & n14485;
assign n12913 = ~(n19170 ^ n3608);
assign n10679 = ~(n9142 ^ n26565);
assign n14774 = ~n16077;
assign n5141 = n13590 | n13783;
assign n11440 = n2377 & n12246;
assign n23247 = ~(n1538 ^ n8523);
assign n6527 = ~(n20151 ^ n20429);
assign n5244 = ~n20415;
assign n2705 = ~(n841 ^ n13718);
assign n2335 = n13330 & n7182;
assign n2267 = n4568 & n14023;
assign n8430 = ~n25043;
assign n26920 = n8569 & n10791;
assign n10958 = ~(n14718 | n468);
assign n16010 = n24684 | n12880;
assign n3205 = n21507 & n14037;
assign n26108 = n5330 | n1386;
assign n19719 = ~n19230;
assign n4698 = n1009 | n152;
assign n16778 = ~n8374;
assign n5709 = ~n13069;
assign n14030 = n4081 | n21810;
assign n26782 = ~n25926;
assign n447 = ~(n14033 ^ n22797);
assign n13637 = ~(n5211 | n12811);
assign n12602 = n15796 | n23095;
assign n23024 = n23837 & n7137;
assign n22289 = ~n7716;
assign n6349 = ~(n6043 ^ n4764);
assign n12760 = ~(n25749 | n7377);
assign n7510 = n21942 | n16908;
assign n4760 = ~(n25993 ^ n3421);
assign n12532 = n13382 & n13068;
assign n16209 = ~(n25038 | n23745);
assign n8334 = ~(n10712 | n26512);
assign n2738 = ~n12029;
assign n10325 = n3190 | n23141;
assign n16416 = n13753 | n16792;
assign n20894 = ~(n10650 | n22253);
assign n11890 = n1360 | n24257;
assign n4945 = n24000 | n21215;
assign n16513 = ~n23661;
assign n9145 = ~(n25917 ^ n3959);
assign n7826 = n21744 | n1900;
assign n18059 = ~(n25579 ^ n21032);
assign n15853 = n15629 | n18614;
assign n17055 = ~(n24358 | n20951);
assign n18963 = n16494 & n5486;
assign n6382 = n23486 & n11734;
assign n27046 = ~(n26575 ^ n11284);
assign n5567 = n528 & n13627;
assign n8153 = ~n24151;
assign n2399 = ~n3524;
assign n8600 = ~(n10562 ^ n4632);
assign n18876 = ~(n12968 ^ n16244);
assign n19667 = ~n12626;
assign n10553 = n444 & n8142;
assign n24423 = n8007 & n4244;
assign n16793 = ~(n12441 ^ n19379);
assign n10955 = n21375 | n16109;
assign n7708 = ~(n7011 ^ n11395);
assign n4847 = ~(n19152 ^ n23842);
assign n9101 = n9260 | n10093;
assign n14813 = n16609 | n22666;
assign n7221 = ~(n11406 ^ n15929);
assign n23665 = n20206 | n6105;
assign n3427 = n4073 | n17566;
assign n22951 = n12862 & n14503;
assign n6141 = ~(n7446 ^ n9691);
assign n21125 = ~(n11114 ^ n14345);
assign n7853 = n22323 | n24405;
assign n4614 = ~(n9167 ^ n14656);
assign n7273 = n26112 & n19207;
assign n22617 = n19200 | n26803;
assign n20873 = n16179 | n11164;
assign n19674 = ~(n5010 ^ n22481);
assign n4167 = n2441 & n806;
assign n10840 = ~(n20754 | n593);
assign n13626 = ~(n14834 ^ n24265);
assign n17599 = ~n21206;
assign n10043 = n18742 & n14319;
assign n5485 = ~(n4433 ^ n22508);
assign n1944 = n21217 & n697;
assign n10747 = n13166 | n22340;
assign n13632 = n10900 & n10087;
assign n10342 = ~(n23582 ^ n16738);
assign n1773 = ~(n19812 ^ n23652);
assign n4603 = ~n22476;
assign n22995 = n7266 & n17533;
assign n25500 = n14654 & n12664;
assign n4626 = ~(n25699 ^ n22290);
assign n15320 = n2022 | n1903;
assign n24285 = ~(n13405 | n22253);
assign n18704 = ~(n9741 | n11229);
assign n20338 = ~n11936;
assign n14288 = ~n8694;
assign n18416 = ~(n5525 ^ n25694);
assign n26070 = n20321 | n3861;
assign n11295 = ~(n26368 ^ n19118);
assign n4342 = ~n4957;
assign n1049 = ~(n12967 ^ n5028);
assign n7882 = ~n13685;
assign n1505 = ~(n16845 ^ n3228);
assign n9277 = n706 | n7771;
assign n11460 = n5611 | n25694;
assign n15413 = n23598 & n23604;
assign n886 = n21526 & n18732;
assign n2688 = ~(n14524 ^ n16223);
assign n24863 = n12004 & n12289;
assign n9244 = ~n2418;
assign n1462 = n6356 | n4665;
assign n18890 = n7606 | n25092;
assign n23641 = ~(n2049 | n9303);
assign n5453 = ~(n7788 ^ n20013);
assign n7613 = n13773 & n10778;
assign n10330 = ~(n20195 ^ n15336);
assign n12198 = ~n13578;
assign n13223 = ~(n4714 | n5030);
assign n2815 = ~n11416;
assign n8720 = ~n1592;
assign n23232 = ~(n15842 ^ n9665);
assign n21713 = n4620 & n26591;
assign n3124 = ~n9557;
assign n15746 = ~(n4792 ^ n10593);
assign n14720 = ~(n19086 ^ n18307);
assign n18665 = ~n3488;
assign n8880 = n14654 | n26797;
assign n18873 = n26612 & n21139;
assign n15519 = ~n5832;
assign n1286 = n9800 | n8905;
assign n12325 = ~(n24970 ^ n24913);
assign n785 = n10100 | n22898;
assign n25929 = ~n13695;
assign n3717 = n4520 | n10699;
assign n21350 = ~(n13459 | n24786);
assign n18917 = n1619 | n11684;
assign n18471 = ~(n1204 | n25701);
assign n17359 = ~(n3417 ^ n8934);
assign n22471 = ~(n11302 ^ n24786);
assign n24490 = n1458 | n1642;
assign n2632 = n12929 | n10691;
assign n21495 = n19282 & n23709;
assign n19476 = ~(n12507 | n15739);
assign n5355 = ~n25565;
assign n5204 = ~(n2453 | n20700);
assign n3283 = n20213 | n26725;
assign n23070 = n17416 & n1529;
assign n15156 = n24355 | n13951;
assign n15231 = n14759 & n24668;
assign n6148 = ~(n10527 ^ n3314);
assign n23116 = n12945 | n19160;
assign n11393 = ~n7057;
assign n17876 = n11147 | n12981;
assign n22242 = n10123 | n15557;
assign n12001 = ~(n3186 ^ n5834);
assign n21935 = ~n10107;
assign n3216 = ~(n8186 | n19282);
assign n14658 = n24071 & n22900;
assign n24410 = n4780 & n21922;
assign n25888 = ~n20470;
assign n1278 = ~(n8596 ^ n24732);
assign n16857 = n24691 | n10336;
assign n20001 = n23403 & n13880;
assign n13585 = n22694 & n15183;
assign n17810 = ~(n7072 ^ n6857);
assign n7111 = ~n24937;
assign n11157 = n6259 | n24152;
assign n3635 = ~n643;
assign n7532 = ~n24875;
assign n11448 = n9066 & n22894;
assign n14343 = n9953 & n4946;
assign n10625 = ~(n5975 ^ n21675);
assign n2363 = ~(n12016 ^ n11162);
assign n9564 = ~n11974;
assign n15251 = ~(n9259 | n12423);
assign n5988 = n20599 & n16450;
assign n6792 = n19593 | n7227;
assign n17408 = n9014 ^ n11567;
assign n4823 = n15284 | n26819;
assign n775 = n3022 | n7188;
assign n4025 = n4054 & n14820;
assign n11877 = ~(n26881 ^ n26651);
assign n5049 = ~(n18477 ^ n10629);
assign n17240 = n8315 | n26460;
assign n26298 = ~(n234 ^ n2755);
assign n2306 = ~(n2331 ^ n12546);
assign n15765 = ~(n3480 ^ n7057);
assign n1513 = ~(n758 ^ n14731);
assign n12607 = ~(n7772 ^ n2827);
assign n5389 = n6485 & n26265;
assign n25613 = n12989 & n23470;
assign n7084 = n15884 | n26001;
assign n18953 = ~(n18622 ^ n25893);
assign n26425 = ~(n1184 ^ n16657);
assign n13619 = n5796 | n1869;
assign n20444 = ~n22225;
assign n5538 = n2633 | n14058;
assign n22299 = n23769 | n13747;
assign n5654 = n14415 | n5822;
assign n3342 = n18550 | n22259;
assign n11886 = n18471 | n17706;
assign n16286 = ~(n24948 | n11322);
assign n23157 = n18078 | n10711;
assign n19904 = ~(n12200 ^ n13215);
assign n570 = ~n11841;
assign n5902 = ~(n17536 ^ n23799);
assign n12009 = n1314 & n20967;
assign n256 = ~(n20020 ^ n20145);
assign n19958 = n1988 & n2687;
assign n27138 = n9715 & n24527;
assign n16815 = n22515 | n10467;
assign n11808 = ~(n5620 | n23814);
assign n11611 = ~(n17161 ^ n8282);
assign n13369 = n2175 | n15384;
assign n9802 = ~n20349;
assign n1352 = ~(n20169 | n4426);
assign n1838 = ~n8732;
assign n13187 = n1348 | n9784;
assign n7247 = n13156 | n21321;
assign n22979 = n6569 | n6989;
assign n25430 = ~(n10275 ^ n22359);
assign n222 = n22 | n9674;
assign n1715 = ~n7339;
assign n25715 = ~n10650;
assign n22601 = ~(n11056 | n21276);
assign n19071 = ~(n26629 ^ n19904);
assign n4231 = ~(n5658 ^ n21682);
assign n13170 = ~(n19271 ^ n14045);
assign n7885 = ~(n8964 ^ n22554);
assign n17686 = n25997 & n24349;
assign n2655 = n4291 & n10823;
assign n13589 = n26199 & n14594;
assign n19305 = n17759 & n16391;
assign n27080 = n21317 | n8251;
assign n17892 = n19962 | n1570;
assign n18637 = n18786 | n25953;
assign n12088 = ~(n8683 ^ n15379);
assign n23013 = ~n15158;
assign n13045 = ~(n15482 ^ n5123);
assign n19461 = ~(n12535 | n15167);
assign n9496 = ~n20754;
assign n16422 = ~(n485 ^ n4642);
assign n5458 = n11727 & n25292;
assign n15744 = n25258 & n6838;
assign n6255 = ~n13623;
assign n25350 = n15116 | n15821;
assign n24876 = ~(n3740 | n12232);
assign n12585 = ~(n1558 ^ n3918);
assign n22637 = ~(n11976 | n11437);
assign n10151 = ~n1895;
assign n25099 = ~n5376;
assign n10843 = ~(n20368 ^ n6741);
assign n6947 = n7782 & n10688;
assign n3224 = n5531 | n22952;
assign n7770 = n11542 | n3136;
assign n6025 = ~n16752;
assign n23627 = n23068 & n13171;
assign n1712 = ~(n2633 ^ n5341);
assign n1688 = n7311 | n5657;
assign n2382 = ~(n15227 ^ n2794);
assign n19334 = ~(n9399 ^ n6502);
assign n21658 = ~(n23097 ^ n6082);
assign n15728 = ~(n16387 ^ n3673);
assign n22841 = ~(n7771 ^ n6885);
assign n21645 = ~(n6976 ^ n10035);
assign n13049 = ~(n23631 | n3365);
assign n17002 = ~n2328;
assign n6482 = n14979 | n19106;
assign n25321 = ~(n8819 ^ n16961);
assign n16013 = ~(n10569 ^ n5275);
assign n10086 = ~n13518;
assign n9362 = n10933 & n326;
assign n4536 = n10205 | n2538;
assign n4304 = n10285 & n471;
assign n19316 = n21042 & n13512;
assign n17910 = n6051 | n11302;
assign n23253 = ~(n4705 ^ n919);
assign n7958 = ~(n19377 ^ n23784);
assign n1184 = n5945 & n7067;
assign n8172 = n16238 & n22334;
assign n2232 = ~(n7092 ^ n20213);
assign n184 = n25055 & n4079;
assign n2472 = ~(n17035 ^ n19515);
assign n1122 = n21310 & n18620;
assign n3780 = ~n7636;
assign n25376 = ~n18452;
assign n24169 = n26388 & n702;
assign n22549 = ~n16165;
assign n9788 = ~n16274;
assign n9242 = ~n4259;
assign n1486 = n14711 & n20204;
assign n1564 = n4932 & n19969;
assign n11757 = n26540 & n8102;
assign n13177 = n19106 & n8715;
assign n19284 = ~(n20885 ^ n10537);
assign n17832 = ~n3671;
assign n24806 = ~n24948;
assign n6091 = n8679 | n8379;
assign n14369 = ~(n7670 | n10485);
assign n3581 = ~(n13981 ^ n6611);
assign n23497 = n21813 & n10133;
assign n25123 = n2415 | n172;
assign n1650 = n11014 | n23900;
assign n22195 = n23380 | n17008;
assign n7132 = ~(n7059 ^ n6202);
assign n15085 = ~n23636;
assign n4684 = ~(n9993 ^ n22201);
assign n17218 = ~(n15773 ^ n21997);
assign n23328 = ~(n16376 | n17467);
assign n2792 = ~(n21381 ^ n11507);
assign n4855 = ~(n7640 ^ n17511);
assign n9243 = ~(n21822 ^ n25617);
assign n3169 = n7982 & n8907;
assign n5620 = n6297 | n21587;
assign n433 = ~(n6200 ^ n12288);
assign n3308 = n18601 & n19874;
assign n12544 = ~(n20235 | n8259);
assign n10678 = n25444 | n6461;
assign n18824 = n12130 | n14894;
assign n7083 = ~(n21922 ^ n14217);
assign n20356 = ~(n14754 ^ n17366);
assign n4910 = n9821 | n11838;
assign n21106 = n15492 | n14478;
assign n19467 = ~(n16967 ^ n3080);
assign n5839 = n19901 & n8486;
assign n14719 = ~n15378;
assign n25635 = ~(n12650 ^ n16544);
assign n1453 = n23682 & n8404;
assign n781 = ~(n4763 ^ n22304);
assign n2004 = ~(n12549 ^ n23790);
assign n11969 = ~(n16642 ^ n964);
assign n8018 = n15905 & n14996;
assign n12542 = n10463 | n2647;
assign n24409 = n21819 & n26737;
assign n26177 = ~(n12662 ^ n11720);
assign n13680 = n16436 & n25849;
assign n24449 = n26231 | n11174;
assign n21127 = ~n27134;
assign n6716 = ~(n22613 ^ n18157);
assign n22966 = n10036 | n14360;
assign n23388 = ~(n27193 ^ n1293);
assign n1367 = n19299 & n4779;
assign n1782 = n15123 & n23017;
assign n2350 = n5462 ^ n14679;
assign n16758 = ~(n14923 ^ n7238);
assign n1613 = n23486 | n11734;
assign n3714 = ~n12567;
assign n13828 = ~n21501;
assign n14566 = ~n5451;
assign n20692 = n20425 ^ n3053;
assign n19262 = n20259 | n3925;
assign n25334 = ~(n12789 | n23180);
assign n5336 = ~(n5905 ^ n8167);
assign n404 = n18562 | n18195;
assign n16708 = n24744 | n14557;
assign n834 = ~n4943;
assign n466 = ~(n15062 ^ n12457);
assign n14462 = n3446 & n3267;
assign n16837 = ~(n20779 ^ n24910);
assign n5611 = ~n12398;
assign n8818 = ~n24312;
assign n7435 = ~(n22181 ^ n4284);
assign n613 = ~(n13152 | n167);
assign n8093 = n16286 | n13041;
assign n1236 = ~n25296;
assign n17544 = ~(n16731 ^ n26191);
assign n16550 = ~(n18907 ^ n26823);
assign n9269 = ~(n4979 ^ n9702);
assign n21881 = n10030 & n4557;
assign n17045 = n23974 | n281;
assign n1246 = ~(n9920 | n13650);
assign n13415 = n18394 | n26453;
assign n9205 = n7666 | n4914;
assign n14966 = ~(n21721 | n7466);
assign n12538 = ~(n11924 ^ n10986);
assign n21592 = n6904 | n26241;
assign n112 = ~n21905;
assign n19035 = n25674 | n19634;
assign n8799 = n15743 | n20658;
assign n5609 = ~(n2772 ^ n21131);
assign n13635 = ~(n9700 | n15482);
assign n19979 = n9961 ^ n8589;
assign n14077 = n13461 | n5746;
assign n6612 = ~(n23468 ^ n7231);
assign n3371 = n1509 & n16913;
assign n879 = ~(n25343 ^ n19261);
assign n5961 = ~(n22031 ^ n4923);
assign n14 = ~(n12522 | n12208);
assign n13278 = ~n24704;
assign n21196 = n5895 | n21817;
assign n8232 = ~n3179;
assign n17809 = n5014 & n18579;
assign n24783 = n21857 & n10861;
assign n1199 = ~n10231;
assign n1647 = n6478 | n4375;
assign n18271 = ~(n1186 ^ n26408);
assign n11318 = n9535 & n11846;
assign n12215 = n11184 | n6842;
assign n8026 = n25617 | n13448;
assign n8169 = n20502 | n19977;
assign n22171 = n4542 | n8805;
assign n10478 = ~(n5213 ^ n3468);
assign n21285 = n27186 | n15194;
assign n25337 = ~(n5774 ^ n5040);
assign n18851 = n25370 | n11603;
assign n6143 = ~n9450;
assign n9007 = ~(n2420 | n23807);
assign n18794 = ~(n18021 ^ n9486);
assign n5854 = n23250 | n11209;
assign n15157 = n13677 | n10451;
assign n629 = ~(n24727 ^ n7882);
assign n20053 = ~n19138;
assign n1567 = n26305 & n3657;
assign n18382 = n4862 & n25902;
assign n13627 = n8344 | n21804;
assign n3591 = ~n1773;
assign n3123 = n18602 & n20992;
assign n14375 = ~(n14188 ^ n4331);
assign n14406 = ~(n26797 | n15077);
assign n23324 = n26088 | n939;
assign n14672 = n23234 | n1688;
assign n25281 = n18321 | n20238;
assign n6586 = ~(n5862 ^ n18841);
assign n22445 = n22332 & n22370;
assign n5623 = n800 | n25547;
assign n1521 = ~(n1672 ^ n14244);
assign n24223 = n264 | n20344;
assign n23593 = ~(n4665 ^ n18558);
assign n15614 = ~(n19870 ^ n6495);
assign n7607 = ~(n7513 ^ n20431);
assign n15215 = n9520 & n26376;
assign n20377 = ~(n8227 ^ n11947);
assign n3113 = ~(n8161 | n6870);
assign n693 = ~(n23569 ^ n13139);
assign n18321 = ~(n16642 | n704);
assign n19523 = ~(n21103 ^ n629);
assign n15892 = ~(n22553 ^ n7891);
assign n14517 = n932 & n10739;
assign n16733 = ~(n1298 ^ n2148);
assign n4513 = ~(n26005 ^ n2742);
assign n9635 = ~(n11866 ^ n21356);
assign n16162 = ~(n7934 ^ n5608);
assign n14403 = n8340 | n4580;
assign n16739 = n411 & n22650;
assign n9071 = n6782 | n10498;
assign n8959 = n1268 & n23953;
assign n21849 = ~(n25159 ^ n24056);
assign n24553 = n19171 | n24293;
assign n545 = n3349 & n2919;
assign n17276 = ~n14811;
assign n21261 = ~n15135;
assign n13087 = n11685 | n21226;
assign n21927 = ~(n7115 ^ n3987);
assign n9224 = n12500 | n20930;
assign n15854 = n26660 & n26810;
assign n13974 = n19543 | n4618;
assign n9119 = ~(n17287 | n23697);
assign n11017 = ~(n7023 ^ n5942);
assign n9135 = ~(n18766 ^ n12186);
assign n13080 = ~(n26516 | n16052);
assign n10698 = ~(n12017 ^ n15807);
assign n12762 = ~n25355;
assign n8458 = n15395 | n15203;
assign n1058 = ~(n24301 | n4256);
assign n19732 = ~(n27175 | n7056);
assign n25299 = n23436 | n3276;
assign n6330 = ~(n6768 | n20412);
assign n17392 = ~(n1732 ^ n16887);
assign n2375 = n9329 & n11528;
assign n11361 = n2629 | n25124;
assign n16046 = ~(n25838 | n26935);
assign n23896 = n9393 & n24233;
assign n23270 = ~(n2397 ^ n4554);
assign n24474 = n27196 & n10393;
assign n11548 = ~(n17191 ^ n16104);
assign n818 = ~n13946;
assign n26838 = ~(n6154 ^ n23829);
assign n15613 = n2557 | n8441;
assign n23611 = n12493 | n16520;
assign n7258 = ~n1351;
assign n26309 = ~(n24937 | n12436);
assign n25579 = n660 & n22368;
assign n6791 = ~(n10457 ^ n11746);
assign n11470 = ~(n9189 ^ n14857);
assign n14321 = n19124 & n26381;
assign n13065 = n4579 | n511;
assign n23812 = n20640 & n13149;
assign n5947 = ~n3504;
assign n8378 = ~n20755;
assign n12589 = n12319 | n24745;
assign n10243 = ~(n20770 | n10468);
assign n9901 = ~(n11583 ^ n13538);
assign n7928 = ~(n2246 ^ n3668);
assign n23413 = ~(n14957 | n19218);
assign n15065 = ~n27117;
assign n8037 = ~n27202;
assign n7695 = ~(n26892 ^ n11623);
assign n2941 = ~n26253;
assign n5264 = ~n12142;
assign n5821 = n18221 | n16090;
assign n19553 = n17026 | n3078;
assign n20767 = ~(n93 ^ n3515);
assign n15749 = ~(n10434 ^ n3728);
assign n18029 = n14576 | n25069;
assign n13718 = ~(n4322 ^ n16029);
assign n22641 = n18758 | n12407;
assign n7968 = ~(n9299 ^ n17518);
assign n2870 = n10533 | n24117;
assign n15821 = n24549 | n26477;
assign n26122 = ~n9215;
assign n3600 = n13815 & n7449;
assign n27048 = ~(n25277 | n21860);
assign n11529 = n11175 & n18968;
assign n12560 = n11093 & n26400;
assign n9665 = ~n12606;
assign n2564 = n6104 & n2056;
assign n16049 = ~(n420 | n7365);
assign n11964 = n6206 & n17409;
assign n22472 = ~(n26843 ^ n18935);
assign n11433 = ~(n16524 ^ n3785);
assign n6231 = n16111 | n9219;
assign n3027 = ~(n5445 ^ n21759);
assign n21795 = ~n21599;
assign n15611 = n8014 & n26446;
assign n1810 = ~(n20075 ^ n15891);
assign n10507 = n6554 | n25060;
assign n14938 = n8370 | n6909;
assign n18674 = ~(n25035 ^ n16317);
assign n18009 = n16922 | n1486;
assign n23323 = ~(n9768 ^ n16321);
assign n17604 = n25395 | n17648;
assign n10038 = ~(n7621 | n2510);
assign n2634 = n17079 & n16556;
assign n22282 = ~(n90 ^ n22044);
assign n743 = n13190 & n15769;
assign n2162 = ~(n4469 ^ n23545);
assign n26822 = ~(n20825 ^ n17842);
assign n19635 = n26325 | n8892;
assign n6737 = n22446 & n24467;
assign n140 = n23168 | n8067;
assign n11907 = n23638 | n16271;
assign n12874 = ~(n24774 ^ n22660);
assign n9650 = ~(n18331 | n1415);
assign n2587 = n15549 & n22813;
assign n211 = n2682 & n5577;
assign n479 = n22168 & n5334;
assign n15331 = ~(n5640 | n3674);
assign n10345 = ~(n319 ^ n8226);
assign n8749 = ~(n17911 | n22207);
assign n12559 = n22029 | n10173;
assign n22714 = ~(n16245 ^ n21275);
assign n15630 = ~(n20883 ^ n5859);
assign n13299 = n17491 & n11977;
assign n16569 = n17423 | n14584;
assign n10703 = n22791 | n27064;
assign n9958 = ~(n15767 | n18973);
assign n23028 = n23555 | n11745;
assign n9456 = ~n26193;
assign n26839 = n12788 | n15808;
assign n25556 = ~(n12354 ^ n24323);
assign n16320 = ~(n10312 | n10013);
assign n15735 = n5849 | n2956;
assign n9304 = n12348 | n22603;
assign n5983 = n9475 & n22827;
assign n1892 = n12702 | n348;
assign n4657 = ~(n658 | n22274);
assign n5284 = ~n3307;
assign n10406 = ~n8881;
assign n2527 = n10207 | n20084;
assign n5484 = ~(n1844 | n54);
assign n6341 = ~(n7156 ^ n10710);
assign n20047 = n8658 | n6158;
assign n3050 = ~n23207;
assign n17109 = n20844 & n9059;
assign n3147 = ~(n1614 ^ n2771);
assign n10164 = n22176 | n7676;
assign n10431 = ~n11210;
assign n17705 = ~(n9083 ^ n21132);
assign n20659 = ~(n16994 | n4964);
assign n13945 = ~n26585;
assign n21793 = n5686 & n11773;
assign n23243 = n4453 & n12542;
assign n17981 = ~(n19652 | n17444);
assign n20763 = n16610 & n4793;
assign n2560 = ~(n27000 ^ n7181);
assign n9982 = n15984 | n26521;
assign n20071 = ~(n302 | n11975);
assign n4253 = ~(n11056 ^ n21276);
assign n14730 = ~n20153;
assign n12503 = n14965 & n25465;
assign n3210 = n2087 | n17986;
assign n23949 = n15760 | n23285;
assign n6037 = ~(n1886 ^ n10096);
assign n135 = ~(n4400 ^ n2651);
assign n577 = ~(n2509 ^ n22289);
assign n16878 = ~n9632;
assign n20754 = ~(n16691 ^ n476);
assign n19442 = ~n19745;
assign n2687 = n10816 | n23130;
assign n21607 = ~(n15389 | n24468);
assign n6510 = n4259;
assign n20073 = ~(n19215 ^ n395);
assign n7676 = ~n23065;
assign n11693 = n17677 & n17242;
assign n9450 = n22274 | n24129;
assign n2949 = n6122 & n1894;
assign n15829 = n11273 | n7949;
assign n20835 = ~(n14221 ^ n345);
assign n17905 = n13386 | n22305;
assign n13561 = ~n11503;
assign n1886 = n15427 & n19201;
assign n13740 = ~(n12837 ^ n6068);
assign n14663 = n11189 | n25666;
assign n19997 = n7889 & n17941;
assign n24273 = ~n7270;
assign n2579 = ~n23430;
assign n9438 = ~(n1834 | n3354);
assign n13186 = ~(n23241 ^ n24563);
assign n19109 = n23030 & n4333;
assign n368 = n21863 & n756;
assign n20931 = n10452 | n3785;
assign n16346 = ~(n9854 ^ n3056);
assign n11532 = n17957 | n30;
assign n3919 = n11747 | n5648;
assign n9673 = n4338 & n25106;
assign n24752 = ~(n12014 | n7215);
assign n5917 = ~n8160;
assign n12100 = n17399 & n16124;
assign n26155 = ~(n9254 | n25657);
assign n156 = n14452 & n21490;
assign n12729 = n24810 | n15898;
assign n13700 = n1788 & n16112;
assign n19532 = n14837 & n18093;
assign n17256 = ~(n17230 ^ n21687);
assign n14902 = ~(n6163 ^ n17829);
assign n17595 = n25004 | n18409;
assign n11040 = ~(n13569 ^ n4964);
assign n15101 = ~n6178;
assign n1371 = ~(n2844 ^ n20073);
assign n7881 = ~(n18869 ^ n13073);
assign n23181 = ~(n993 ^ n26479);
assign n11807 = n16634 | n12308;
assign n20970 = ~(n9669 ^ n20946);
assign n9698 = n19709 | n9806;
assign n15970 = ~(n25026 ^ n8669);
assign n11930 = n26559 & n24354;
assign n10422 = ~(n219 ^ n13450);
assign n10663 = n1678 & n6409;
assign n11222 = n20123 & n5909;
assign n13061 = n3480 & n7373;
assign n5650 = ~(n4869 | n15024);
assign n9474 = ~(n839 ^ n15709);
assign n8715 = n9570 & n3637;
assign n18174 = ~n19595;
assign n18795 = n6238 | n14664;
assign n1957 = ~(n11118 | n15442);
assign n20454 = ~(n14056 | n8915);
assign n17895 = n5304 | n15437;
assign n1140 = ~(n16336 | n16306);
assign n418 = n16924 | n22395;
assign n3162 = ~(n10758 | n14845);
assign n11624 = ~(n7284 | n7750);
assign n23038 = n23745 | n23053;
assign n2970 = ~(n8497 | n26914);
assign n23926 = n20010 & n26368;
assign n26091 = n26807 & n17677;
assign n15051 = ~(n19556 ^ n3483);
assign n18829 = n1757 & n11970;
assign n260 = ~n17345;
assign n7798 = ~n24847;
assign n12114 = n12967 | n11030;
assign n21477 = ~(n10053 ^ n19911);
assign n7596 = ~(n3468 ^ n23430);
assign n3429 = ~(n5442 ^ n19752);
assign n26953 = ~(n16396 ^ n22871);
assign n13664 = n26095 | n12939;
assign n23241 = n4772 & n25833;
assign n4217 = ~n17553;
assign n9044 = ~(n4917 | n23905);
assign n17987 = ~n14788;
assign n10104 = n15795 | n18606;
assign n20264 = ~(n5999 | n17762);
assign n3503 = ~(n7254 | n14071);
assign n21351 = n10096 | n26553;
assign n8934 = ~(n24949 ^ n23681);
assign n14877 = n4776 | n17420;
assign n9393 = n3958 | n10746;
assign n5682 = ~(n10445 ^ n1253);
assign n2904 = ~(n3570 ^ n8067);
assign n15832 = ~(n822 | n12869);
assign n5477 = n15855 & n11511;
assign n21990 = n12189 | n542;
assign n23307 = ~(n21147 ^ n25869);
assign n15374 = n11857 & n149;
assign n15441 = n2236 | n754;
assign n23144 = ~n3710;
assign n1961 = ~(n22274 ^ n11192);
assign n13184 = ~(n20314 | n10253);
assign n26974 = ~n23985;
assign n20335 = n11561 & n3732;
assign n6824 = n15454 & n26039;
assign n15194 = n1134 & n3876;
assign n6052 = n3479 | n11937;
assign n17863 = n16468 ^ n7674;
assign n25265 = n21495 | n23255;
assign n21642 = ~(n2782 ^ n5793);
assign n25720 = n5602 | n19179;
assign n14359 = n2108 & n1641;
assign n6704 = ~(n2355 | n115);
assign n22244 = ~(n14387 | n15007);
assign n8332 = ~(n3351 | n9842);
assign n25421 = n15041 | n13224;
assign n23320 = ~(n13033 | n19392);
assign n10379 = n21636 | n22154;
assign n12784 = n17250 & n26997;
assign n2920 = ~(n19368 ^ n5802);
assign n8861 = ~(n3852 ^ n2431);
assign n18723 = n19428 & n21553;
assign n9831 = n25516 & n16242;
assign n14515 = ~(n15693 | n24701);
assign n26892 = ~n15801;
assign n10131 = ~n15602;
assign n16723 = n1642 & n5512;
assign n4832 = n5957 | n19997;
assign n8807 = ~(n12143 ^ n20215);
assign n18779 = n1864 | n11835;
assign n4593 = n18444 | n26224;
assign n16922 = ~(n20641 | n3443);
assign n11281 = ~(n1533 ^ n5451);
assign n23751 = ~n2352;
assign n14456 = ~(n16213 ^ n14878);
assign n20416 = ~(n146 | n2979);
assign n20357 = n19949 | n16474;
assign n22584 = ~(n19034 ^ n26282);
assign n17695 = n6833 & n2040;
assign n3829 = ~(n5628 ^ n2054);
assign n8208 = ~(n21634 | n5579);
assign n3942 = n12002 & n11382;
assign n13745 = ~n8315;
assign n27159 = n2117 | n6711;
assign n13297 = ~(n16409 ^ n23861);
assign n26035 = ~(n27089 ^ n6814);
assign n17907 = n19205 | n11068;
assign n16706 = n17763 | n12908;
assign n12094 = ~(n17266 ^ n25239);
assign n26183 = n14193 | n16172;
assign n9354 = n10982 | n21560;
assign n18081 = n24107 & n14291;
assign n5091 = ~(n22426 ^ n20658);
assign n25046 = n11283 | n23128;
assign n22165 = n13770 | n12491;
assign n11917 = n2514 | n5213;
assign n13919 = ~n21047;
assign n9423 = ~(n22046 ^ n24268);
assign n18688 = n15990 & n2977;
assign n25799 = ~n11489;
assign n7865 = n9947 & n22726;
assign n20863 = n23838 & n24204;
assign n24072 = n20314 & n147;
assign n6765 = n3931 & n11596;
assign n127 = n10413 | n21881;
assign n1939 = ~(n19473 ^ n24372);
assign n3516 = ~(n12010 ^ n10624);
assign n24445 = n12478 | n3917;
assign n14610 = n11022 ^ n6890;
assign n9649 = n8983 & n21737;
assign n14444 = ~(n9965 ^ n26665);
assign n1753 = ~n21911;
assign n1783 = ~(n12 | n23725);
assign n19417 = n5932 & n5359;
assign n10732 = ~(n16107 ^ n6068);
assign n9479 = ~n2743;
assign n20034 = n25313 | n1212;
assign n15452 = ~(n17302 | n13784);
assign n1197 = n22426 | n20620;
assign n3156 = n26925 | n10199;
assign n20139 = ~n10072;
assign n12983 = ~(n17090 ^ n27120);
assign n24023 = n9472 & n7611;
assign n11272 = n20113 | n23930;
assign n17443 = n12651 | n24779;
assign n2302 = n26706 & n19872;
assign n18660 = n6604 & n24871;
assign n22954 = ~(n14507 | n18058);
assign n23009 = ~(n19713 ^ n10820);
assign n11151 = ~n20231;
assign n15104 = n17711 & n8398;
assign n11982 = n17879 & n15771;
assign n25743 = n6561 & n19386;
assign n15926 = ~(n8358 ^ n26189);
assign n21662 = ~(n25926 ^ n12384);
assign n408 = n7797 | n8925;
assign n14226 = ~n12861;
assign n26113 = ~(n9786 ^ n22217);
assign n19665 = n10436 | n16148;
assign n3382 = n3216 | n20591;
assign n20112 = ~n24327;
assign n10214 = ~(n3337 ^ n26552);
assign n26283 = n8424 & n26432;
assign n17341 = n14566 | n20378;
assign n14449 = n1494 & n7120;
assign n18348 = n19563 | n15045;
assign n16459 = ~n21164;
assign n9624 = n20152 | n13192;
assign n2142 = ~(n25156 | n2152);
assign n24982 = n19676 & n8812;
assign n500 = ~(n5675 ^ n1876);
assign n5915 = n13205 & n120;
assign n20258 = n19094 | n19156;
assign n22193 = n15527 | n3894;
assign n19921 = n19938 & n11623;
assign n9853 = ~(n5436 | n9972);
assign n3852 = n15540 & n23031;
assign n13797 = n13280 | n13309;
assign n21059 = n14040 | n24711;
assign n1979 = ~(n21622 | n15158);
assign n10429 = n4338 | n25106;
assign n19238 = ~(n15166 ^ n20377);
assign n4932 = n18797 | n11489;
assign n20225 = n4994 & n6447;
assign n3947 = ~(n25120 ^ n17458);
assign n14488 = ~(n21064 ^ n16397);
assign n13516 = n26997 | n17250;
assign n21900 = ~(n5889 ^ n6914);
assign n23049 = n19469 | n6209;
assign n16119 = n16649 & n6493;
assign n12159 = n15454 | n23892;
assign n11255 = n1814 & n5080;
assign n24705 = ~n8079;
assign n19935 = ~(n25048 ^ n22815);
assign n7716 = ~(n13088 ^ n18987);
assign n8011 = n7042 & n14159;
assign n16451 = ~(n19297 ^ n21248);
assign n13787 = n26093 | n20235;
assign n8844 = n20138 | n9251;
assign n833 = ~(n16911 ^ n7773);
assign n2601 = n23756 & n23194;
assign n10120 = ~(n26053 | n2320);
assign n13350 = ~(n17978 ^ n3134);
assign n1658 = ~(n24567 ^ n4366);
assign n3293 = ~(n4194 | n14643);
assign n3499 = ~(n10155 | n1738);
assign n24898 = ~(n6176 ^ n20849);
assign n22671 = ~n4202;
assign n23392 = n13343 ^ n1159;
assign n2501 = n1747 & n1078;
assign n5092 = n20100 & n17634;
assign n17562 = ~(n10333 | n9717);
assign n20797 = n11425 & n15957;
assign n13935 = ~n2479;
assign n10717 = n2833 | n7098;
assign n21371 = n25751 | n23190;
assign n6945 = n22024 | n23977;
assign n15464 = ~(n14845 ^ n23572);
assign n14038 = ~n16970;
assign n12741 = ~n17872;
assign n22533 = ~(n21003 ^ n16182);
assign n19150 = ~n6556;
assign n13403 = ~(n8600 ^ n19627);
assign n24852 = n9700 | n9969;
assign n10491 = n25974 | n6963;
assign n5237 = n21556 | n2035;
assign n22955 = n10206 & n22938;
assign n11713 = ~(n10191 ^ n20006);
assign n7659 = n24366 | n5438;
assign n13770 = ~(n23592 | n468);
assign n16266 = n26827 & n21303;
assign n10404 = ~(n17700 ^ n19089);
assign n24965 = ~(n24367 ^ n27099);
assign n19317 = ~(n7226 ^ n20693);
assign n1484 = ~(n3070 ^ n13568);
assign n7761 = ~n25555;
assign n10332 = n21697 | n1542;
assign n4669 = n8732 | n4651;
assign n27157 = n11694 | n14521;
assign n20422 = ~(n3791 | n7437);
assign n3297 = ~(n24590 | n22480);
assign n22412 = ~(n7049 | n21219);
assign n5234 = ~n13672;
assign n5044 = ~(n17415 | n16822);
assign n12047 = ~(n101 ^ n21643);
assign n26120 = ~(n3550 | n5171);
assign n23848 = ~(n5077 | n17397);
assign n25916 = ~(n4245 | n5599);
assign n5310 = n21178 & n8357;
assign n9216 = ~(n14536 | n1320);
assign n25250 = ~(n24235 ^ n2345);
assign n300 = ~n18068;
assign n20814 = ~(n26557 | n10048);
assign n26503 = n3721 | n1855;
assign n19975 = n22052 & n19231;
assign n26129 = ~(n8827 | n8176);
assign n8550 = ~(n6552 ^ n21045);
assign n5000 = n19962 | n19527;
assign n25886 = ~n25974;
assign n22763 = ~(n3710 | n26399);
assign n8118 = ~(n18300 | n13303);
assign n11014 = ~n26046;
assign n3482 = n21117 | n20700;
assign n15228 = n23483 & n26938;
assign n9794 = n16210 | n2731;
assign n10021 = ~(n24502 ^ n13617);
assign n13388 = n18926 & n2705;
assign n21307 = ~(n20271 | n11693);
assign n1485 = n19818 | n12388;
assign n23669 = ~(n23607 ^ n11812);
assign n12404 = n6255 | n8704;
assign n17644 = n8792 | n3764;
assign n16387 = ~(n10300 ^ n24829);
assign n12478 = ~(n13851 | n7010);
assign n18346 = ~(n2718 ^ n14981);
assign n23542 = n3892 & n6942;
assign n12625 = n24153 & n1445;
assign n8253 = ~n1245;
assign n20784 = n19340 | n7241;
assign n24573 = n23098 & n20550;
assign n25970 = n6571 | n12549;
assign n17647 = ~n23894;
assign n4444 = n10227 | n3102;
assign n20592 = ~(n26556 ^ n5438);
assign n22990 = n752 & n11504;
assign n10897 = ~(n24379 ^ n18810);
assign n14939 = ~(n11383 | n23558);
assign n4619 = n4436 | n21406;
assign n16088 = n8977 & n18821;
assign n20266 = ~n6933;
assign n19607 = ~n3751;
assign n18805 = n15182 | n2996;
assign n13411 = ~(n481 | n13951);
assign n9845 = ~(n14106 ^ n16880);
assign n10249 = ~n10454;
assign n21150 = n24804 & n17015;
assign n9587 = n18345 & n22700;
assign n11576 = ~(n15440 ^ n3147);
assign n15275 = ~(n15412 ^ n10731);
assign n6678 = ~(n21848 ^ n11230);
assign n24538 = ~(n21693 ^ n15875);
assign n12921 = ~n19618;
assign n11344 = ~(n25622 ^ n19186);
assign n20727 = ~(n25360 ^ n2102);
assign n3415 = ~n22782;
assign n13483 = ~(n5538 | n5772);
assign n17649 = ~(n22274 | n22591);
assign n15499 = ~(n14870 ^ n8888);
assign n25783 = ~(n18351 | n5690);
assign n6951 = n1628 & n24971;
assign n6392 = ~(n2168 ^ n9502);
assign n24914 = n22805 & n10297;
assign n22322 = ~(n21020 ^ n13703);
assign n18234 = n23913 | n7274;
assign n25060 = n8738 & n17700;
assign n2475 = n2130 | n16921;
assign n9654 = n15323 & n25177;
assign n8532 = ~(n20638 | n3540);
assign n17769 = n5321 | n22628;
assign n18695 = n23744 | n5380;
assign n531 = n1742 & n1798;
assign n22341 = ~(n8894 ^ n24441);
assign n23213 = ~(n5783 ^ n11432);
assign n23726 = n5440 | n4326;
assign n17352 = n1573 & n4652;
assign n24204 = n23228 | n10460;
assign n10302 = n4963 | n2818;
assign n5055 = ~(n23801 ^ n16646);
assign n15306 = n20860 & n15020;
assign n4036 = n4149 & n24799;
assign n11743 = ~(n22636 ^ n16971);
assign n5509 = n7334 & n5925;
assign n16351 = ~n14826;
assign n6375 = ~(n1171 ^ n5456);
assign n2622 = n16817 & n24401;
assign n20079 = ~(n20478 | n26030);
assign n25039 = n19422 | n14082;
assign n15701 = ~(n23272 ^ n14826);
assign n26642 = n23580 & n8925;
assign n3783 = ~n4007;
assign n5878 = n6261 | n292;
assign n23811 = n4530 | n14165;
assign n2981 = ~(n1244 ^ n11779);
assign n17083 = ~(n16483 | n18846);
assign n23439 = n12503 | n13362;
assign n15677 = n7247 & n6002;
assign n7124 = n9187 & n4870;
assign n24593 = ~n21894;
assign n6992 = n6847 | n2051;
assign n897 = ~(n7162 ^ n21226);
assign n17672 = n5933 | n625;
assign n14416 = n19481 & n12052;
assign n24823 = ~n15332;
assign n6832 = n25663 & n16721;
assign n27029 = n1702 & n2733;
assign n4297 = n4859 | n14584;
assign n12457 = ~n15985;
assign n2539 = n7621 & n7217;
assign n1327 = n20138 & n26093;
assign n15410 = n1340 | n16561;
assign n18796 = n18937 & n11942;
assign n16268 = n1472 | n14057;
assign n14751 = n6039 & n9394;
assign n19424 = ~(n5944 ^ n21231);
assign n7106 = ~(n3791 | n7330);
assign n2246 = ~n10114;
assign n16881 = ~(n10049 | n6790);
assign n1344 = ~(n18956 ^ n10427);
assign n1670 = n22053 | n1388;
assign n4907 = n26204 | n24360;
assign n8434 = ~n23630;
assign n21090 = n19493 | n25521;
assign n15610 = ~(n18203 ^ n18909);
assign n3236 = ~n7406;
assign n16729 = ~(n17468 ^ n20021);
assign n11305 = n23027 & n9734;
assign n205 = n21340 | n24266;
assign n21023 = n21306 | n9440;
assign n20149 = ~(n6419 ^ n20607);
assign n21965 = ~n27081;
assign n11759 = n19898 | n12531;
assign n26840 = n7148 & n23;
assign n13972 = n2763 & n15330;
assign n27201 = n13823 & n14166;
assign n26084 = n26603 | n6280;
assign n26911 = n10184 | n27037;
assign n3139 = ~(n1558 | n11566);
assign n21988 = ~n7486;
assign n10426 = n8006 | n19514;
assign n24807 = ~(n26516 ^ n10278);
assign n165 = n20750 | n24843;
assign n17554 = n12720 | n19192;
assign n21113 = ~n12367;
assign n4160 = ~(n18195 ^ n18177);
assign n8269 = n16712 | n24278;
assign n23853 = ~(n12902 ^ n14198);
assign n23345 = n19082 | n19321;
assign n17384 = n22631 & n22613;
assign n22315 = ~n9990;
assign n20567 = n23250 & n16856;
assign n26110 = n21304 | n15468;
assign n23161 = ~n16232;
assign n8945 = ~(n12466 ^ n5022);
assign n23405 = ~(n13171 ^ n23068);
assign n19875 = ~n16729;
assign n14998 = ~(n16994 ^ n4964);
assign n4487 = ~(n22021 ^ n2145);
assign n61 = ~(n5212 ^ n18145);
assign n12095 = n25205 & n6839;
assign n2868 = ~(n6667 ^ n22509);
assign n18999 = ~(n6370 ^ n13070);
assign n16809 = ~(n24711 ^ n4760);
assign n11920 = ~(n12660 ^ n27188);
assign n25114 = ~n8527;
assign n860 = ~(n3403 ^ n4193);
assign n22646 = ~(n15992 ^ n6093);
assign n16203 = ~n8280;
assign n26406 = ~(n24961 ^ n1709);
assign n18206 = n20674 | n5010;
assign n1935 = ~(n17959 | n17728);
assign n4905 = ~(n25318 ^ n16544);
assign n5680 = ~(n23904 ^ n9521);
assign n10504 = ~(n15628 ^ n18532);
assign n22536 = n20365 & n14127;
assign n2776 = ~n15902;
assign n6092 = ~(n9291 | n9077);
assign n17787 = n18182 & n9336;
assign n10054 = n18884 & n3224;
assign n6015 = n5003 & n22941;
assign n15774 = n26542 & n21403;
assign n25630 = ~(n11849 ^ n7191);
assign n22328 = n26864 | n18796;
assign n23477 = ~n14090;
assign n5892 = n9443 & n20188;
assign n477 = ~(n11441 ^ n22106);
assign n24460 = ~(n2325 ^ n19248);
assign n18330 = n6496 & n7307;
assign n7383 = n11899 | n27201;
assign n19578 = ~(n12022 ^ n8277);
assign n3142 = ~(n16244 | n18759);
assign n1378 = ~(n7871 ^ n8261);
assign n4517 = n24797 & n13063;
assign n10480 = n24135 & n3134;
assign n3149 = ~(n24779 ^ n21344);
assign n23074 = n23750 | n22254;
assign n24897 = ~(n2460 ^ n8439);
assign n25618 = n18449 & n12588;
assign n9279 = n11728 | n12641;
assign n23511 = n4701 & n25675;
assign n1717 = ~(n17751 ^ n23879);
assign n4696 = n4555 | n11455;
assign n5445 = ~n7387;
assign n17546 = n15059 | n13207;
assign n13981 = ~(n583 ^ n13714);
assign n1818 = n26407 | n3532;
assign n18421 = ~(n6358 ^ n8962);
assign n14513 = n9281 & n15621;
assign n6035 = n7018 | n6737;
assign n23490 = n7026 & n17835;
assign n11985 = n16141 & n7533;
assign n19864 = n11303 | n13133;
assign n20371 = ~(n21113 | n23760);
assign n11715 = n17192 | n26944;
assign n7066 = ~(n17611 ^ n2030);
assign n11650 = ~(n2188 ^ n2802);
assign n8304 = n25968 & n18242;
assign n1079 = ~n17555;
assign n18304 = ~(n295 ^ n27135);
assign n15129 = ~(n21912 | n9291);
assign n15868 = ~n19305;
assign n20228 = n914 & n139;
assign n24715 = ~(n6722 ^ n925);
assign n581 = ~(n22596 ^ n13263);
assign n16105 = n1672 | n14244;
assign n15018 = n17645 | n26405;
assign n9285 = ~n4651;
assign n5259 = ~(n20613 ^ n1599);
assign n6793 = n22269 | n20217;
assign n18378 = ~(n10152 | n7981);
assign n17656 = n12755 & n24438;
assign n16430 = ~(n7291 ^ n11128);
assign n17757 = ~(n22219 | n4781);
assign n10839 = n18737 & n2328;
assign n2247 = n17918 & n24669;
assign n10810 = n726 & n26849;
assign n2341 = ~n20929;
assign n21678 = ~(n26031 ^ n17154);
assign n20204 = n5514 | n24175;
assign n16027 = n13327 | n21401;
assign n22678 = n20776 | n18660;
assign n15133 = ~(n19701 | n2829);
assign n18652 = n26252 & n16765;
assign n14134 = n19944 | n5704;
assign n21001 = ~(n22338 ^ n1992);
assign n25964 = ~(n17388 ^ n13293);
assign n1097 = n16482 | n11293;
assign n7830 = ~(n16777 ^ n16788);
assign n18200 = ~(n6524 ^ n16851);
assign n26065 = ~n15534;
assign n434 = ~(n24630 ^ n8581);
assign n4735 = n22634 | n17816;
assign n20367 = n6262 | n8165;
assign n2910 = n9849 | n17039;
assign n17102 = ~(n10651 ^ n19515);
assign n24699 = n4147 | n20862;
assign n4566 = ~(n23352 ^ n15761);
assign n1906 = ~n1456;
assign n9179 = n25982 & n18262;
assign n8100 = n17871 & n6894;
assign n20304 = n8163 & n7173;
assign n17929 = ~(n19005 | n24618);
assign n12400 = n25905 & n17146;
assign n19550 = ~(n20721 | n2615);
assign n2890 = n25411 & n6977;
assign n12486 = n17474 | n16553;
assign n4461 = ~n23767;
assign n13224 = ~n23086;
assign n14398 = ~(n2834 ^ n8545);
assign n22013 = n15130 & n25567;
assign n16383 = ~(n2568 | n22091);
assign n18389 = n8586 & n23577;
assign n6402 = ~(n7837 ^ n26545);
assign n23293 = ~(n19127 ^ n18200);
assign n22439 = ~(n754 ^ n10547);
assign n4838 = n1068 | n22594;
assign n6852 = ~(n12291 ^ n24933);
assign n19843 = ~n13784;
assign n3126 = ~(n22570 ^ n22249);
assign n25986 = n4550 | n14379;
assign n11598 = n18341 | n18262;
assign n6880 = n6129 | n14749;
assign n8677 = ~n5532;
assign n20315 = n4040 & n16009;
assign n16573 = n3471;
assign n26364 = n5021 & n22553;
assign n6583 = ~(n15182 ^ n26797);
assign n10996 = ~(n5779 ^ n25001);
assign n10980 = n5160 & n8901;
assign n24456 = ~(n24855 ^ n21328);
assign n9983 = n5523 & n2653;
assign n16871 = ~(n20084 ^ n10207);
assign n1873 = n2576 | n8819;
assign n22119 = n5647 & n20320;
assign n5751 = ~(n8929 ^ n10012);
assign n4787 = n23477 | n6794;
assign n6862 = ~(n12372 ^ n15881);
assign n2082 = n19579 | n19729;
assign n12148 = ~(n17143 ^ n7566);
assign n19871 = n11904 & n11422;
assign n7740 = ~n14922;
assign n924 = ~(n10713 ^ n25494);
assign n254 = n24428 | n12450;
assign n4868 = ~n25475;
assign n25707 = n25624 & n9653;
assign n24822 = n4049 | n19529;
assign n10545 = n9264 | n19990;
assign n13371 = ~n13183;
assign n19406 = ~n26264;
assign n5801 = n16530 & n16735;
assign n1986 = n24566 & n17477;
assign n11514 = ~(n11308 ^ n3697);
assign n17751 = n24894 & n25433;
assign n21690 = n13527 | n16118;
assign n13271 = ~(n24624 ^ n13565);
assign n20182 = ~(n10481 ^ n3407);
assign n11659 = ~(n21071 | n7906);
assign n21633 = ~n1852;
assign n664 = ~(n23993 ^ n5640);
assign n17374 = n19438 | n798;
assign n2095 = ~(n12015 ^ n7840);
assign n23750 = ~n23160;
assign n16666 = ~(n16430 | n10915);
assign n4562 = ~n4423;
assign n3204 = ~n4272;
assign n16766 = n18676 | n6135;
assign n5941 = n15142 | n20120;
assign n19604 = ~(n20049 | n13806);
assign n3751 = ~(n11547 ^ n3713);
assign n7591 = n1054 | n6941;
assign n9052 = n6504 | n3618;
assign n1634 = ~(n25005 ^ n5195);
assign n12091 = ~(n7924 | n11333);
assign n1375 = n15430 | n25226;
assign n5740 = ~n8890;
assign n9058 = ~n4235;
assign n5535 = n18100 | n15743;
assign n13579 = n3822 & n26357;
assign n1549 = ~(n13460 ^ n22335);
assign n13370 = n22375 & n5722;
assign n24432 = ~(n5213 | n4812);
assign n10315 = ~(n12422 ^ n5616);
assign n1844 = ~(n17197 ^ n19618);
assign n13433 = n4254 | n21413;
assign n10108 = ~(n2298 ^ n21749);
assign n24013 = n12769 | n25405;
assign n10490 = n13104 & n5993;
assign n11952 = ~(n20929 ^ n6596);
assign n16118 = n4337 & n10600;
assign n2982 = n23491 | n14659;
assign n13031 = ~(n24366 ^ n18151);
assign n6209 = ~n1630;
assign n25147 = ~(n24496 ^ n22210);
assign n2319 = ~(n16938 | n8775);
assign n14411 = ~n26703;
assign n9764 = ~(n18173 | n25494);
assign n14746 = ~(n22864 ^ n23165);
assign n26924 = n25351 & n1331;
assign n17000 = ~(n547 ^ n8090);
assign n21313 = ~(n21222 | n26565);
assign n21156 = n7305 | n1204;
assign n7199 = n14137 & n4726;
assign n3195 = n20524 & n9571;
assign n18430 = ~(n10183 | n24824);
assign n23901 = ~(n6331 ^ n15822);
assign n8732 = ~(n14639 ^ n15663);
assign n23715 = ~(n17840 ^ n8834);
assign n12640 = ~n13263;
assign n10544 = n6904 | n3161;
assign n25234 = n4859 | n9793;
assign n20950 = n18530 | n12526;
assign n9808 = ~(n12811 ^ n19514);
assign n21536 = n19886 & n2391;
assign n3500 = n24547 & n15151;
assign n14278 = ~(n18655 ^ n8875);
assign n9486 = ~(n21693 ^ n20489);
assign n14608 = n7987 | n10911;
assign n9756 = ~(n20964 | n17077);
assign n26258 = n26717 | n16083;
assign n25504 = n14024 | n23568;
assign n17577 = n13760 | n8682;
assign n10967 = ~(n8815 ^ n946);
assign n22028 = n9117 & n20943;
assign n4606 = ~n24573;
assign n2 = n5243 | n24961;
assign n25810 = ~n14521;
assign n10239 = ~(n11568 ^ n13194);
assign n10371 = n6618 & n25911;
assign n7706 = n1692 & n13791;
assign n26118 = ~(n10138 ^ n12419);
assign n7667 = ~(n20920 ^ n22379);
assign n5012 = ~n4085;
assign n15003 = n22225 | n2842;
assign n23600 = n18900 & n23839;
assign n18616 = n24899 | n10160;
assign n23448 = n12390 & n9747;
assign n22819 = ~(n20451 ^ n19435);
assign n19718 = ~(n10964 | n22260);
assign n21609 = n2163 & n10346;
assign n9511 = n9079 | n26042;
assign n7418 = ~n16276;
assign n14445 = n22000 | n11572;
assign n11631 = n8819 | n10869;
assign n26179 = ~(n7863 ^ n25606);
assign n5103 = ~n15705;
assign n1011 = ~(n10357 ^ n6444);
assign n17542 = ~n10125;
assign n4227 = ~(n8571 | n25240);
assign n23536 = ~n23308;
assign n8231 = n24118 | n2525;
assign n13294 = n22642 | n17515;
assign n17213 = ~n23587;
assign n11728 = ~(n2597 | n13989);
assign n23462 = n8463 & n24730;
assign n1181 = n15339;
assign n16779 = n20222 | n4096;
assign n13731 = ~n8581;
assign n12122 = n26036 & n7832;
assign n10731 = ~(n18925 ^ n25150);
assign n3036 = n20981 | n20646;
assign n2582 = ~(n22064 ^ n21491);
assign n25001 = ~(n21880 ^ n11420);
assign n7502 = ~(n20249 ^ n21352);
assign n9200 = ~n26546;
assign n858 = ~(n138 ^ n10284);
assign n25987 = ~n11824;
assign n2887 = ~(n11319 ^ n13793);
assign n3515 = ~n9754;
assign n9316 = n15525 & n8145;
assign n22800 = n11268 | n13831;
assign n2893 = n26597 | n16296;
assign n12494 = ~n26942;
assign n22345 = ~n1886;
assign n18517 = ~(n15426 | n8745);
assign n20434 = n15858 | n14474;
assign n20706 = ~(n18846 ^ n16483);
assign n6147 = ~(n16470 ^ n755);
assign n18808 = n18227 | n21828;
assign n14989 = ~(n10058 ^ n10645);
assign n9647 = n25987 & n14122;
assign n15932 = ~n16541;
assign n22243 = n17978 & n7223;
assign n21511 = ~(n19218 ^ n985);
assign n4594 = ~(n19453 | n12018);
assign n26849 = ~(n16553 ^ n17112);
assign n143 = n15271 & n24850;
assign n15023 = n4878 & n12102;
assign n2364 = n14430 | n10887;
assign n17587 = n20258 & n3442;
assign n19266 = ~(n19742 ^ n19868);
assign n11428 = ~n18714;
assign n24886 = n5026 | n8581;
assign n4362 = ~(n808 ^ n23333);
assign n19597 = n19443 & n22799;
assign n101 = ~(n17480 ^ n22691);
assign n4445 = ~(n13152 | n20455);
assign n13410 = n2857 & n24821;
assign n835 = ~n7006;
assign n9796 = ~(n15113 ^ n24080);
assign n24017 = n26671 & n7790;
assign n17593 = ~(n1319 | n6864);
assign n17104 = ~(n15024 ^ n25631);
assign n19062 = ~(n4625 | n9523);
assign n11306 = n17128 & n26912;
assign n15527 = ~(n8322 | n12811);
assign n8922 = n26264 & n20326;
assign n20869 = ~(n25717 ^ n18700);
assign n20890 = n18726 | n11910;
assign n5474 = ~n20594;
assign n4012 = ~(n3878 | n22421);
assign n10451 = ~(n16170 ^ n6149);
assign n9551 = n4110 & n17283;
assign n24068 = n23484 | n19286;
assign n5348 = ~(n19816 ^ n7709);
assign n9763 = ~(n15953 ^ n3800);
assign n1234 = ~(n3776 | n12709);
assign n8106 = ~(n14494 ^ n13837);
assign n19362 = n10873 | n4572;
assign n23556 = n570 & n18461;
assign n22167 = ~(n15113 | n24080);
assign n17634 = n17286 & n20968;
assign n3392 = n14131 | n26680;
assign n24609 = ~(n22137 ^ n7887);
assign n6846 = n8516 & n7565;
assign n6094 = ~(n25092 ^ n10263);
assign n23147 = n23040 & n25782;
assign n18254 = ~(n17941 ^ n3082);
assign n18589 = ~(n17657 ^ n20546);
assign n848 = n15494 & n20046;
assign n12064 = ~n24166;
assign n14229 = ~(n24554 ^ n24032);
assign n3285 = n1406 | n11486;
assign n5006 = ~n10710;
assign n13932 = ~(n7832 ^ n7697);
assign n7981 = ~n10437;
assign n11639 = ~(n8338 ^ n15521);
assign n6184 = ~(n2052 ^ n13631);
assign n9539 = ~(n12802 | n3707);
assign n11772 = ~(n23710 ^ n5793);
assign n27084 = n10951 & n1577;
assign n10823 = n20759 | n6766;
assign n8888 = ~(n24110 ^ n27036);
assign n5810 = ~(n4801 ^ n20557);
assign n23300 = ~(n26170 ^ n23664);
assign n17128 = n21967 | n4106;
assign n24392 = ~(n9202 ^ n14790);
assign n6084 = ~(n19629 ^ n10520);
assign n9727 = n15585 | n13505;
assign n23198 = n14440 & n14718;
assign n4622 = ~n8806;
assign n20687 = ~(n10004 ^ n15701);
assign n1138 = ~(n26143 ^ n7388);
assign n22748 = n13921 | n16877;
assign n9166 = ~(n5620 ^ n1640);
assign n5084 = n8784 & n17350;
assign n14639 = n2115 | n4357;
assign n18898 = ~(n24217 ^ n15897);
assign n10317 = n3635 & n22635;
assign n6571 = ~(n9187 | n13368);
assign n15725 = ~(n21469 ^ n4692);
assign n14733 = ~n17410;
assign n19287 = n14633 | n20897;
assign n5863 = n13007 & n26401;
assign n4572 = ~n21502;
assign n21861 = ~(n21374 | n10891);
assign n11664 = ~(n21774 | n6564);
assign n9010 = n3326 | n334;
assign n21516 = n6841 | n1662;
assign n23924 = ~(n165 ^ n26874);
assign n18450 = ~n6015;
assign n14400 = ~(n3381 ^ n4816);
assign n4725 = ~(n10565 ^ n8317);
assign n12054 = ~(n14781 | n15703);
assign n7384 = n1558 & n5050;
assign n23258 = ~(n23520 ^ n21355);
assign n8705 = n10890 | n17510;
assign n17498 = n11359 & n26114;
assign n16623 = n23757 & n8195;
assign n5967 = n17255 | n24213;
assign n8734 = ~(n11302 ^ n12341);
assign n26356 = n6251 | n18972;
assign n24563 = ~(n1118 ^ n20489);
assign n7454 = n22132 & n1306;
assign n11816 = ~n26408;
assign n2385 = ~n12851;
assign n6034 = ~n18277;
assign n16810 = n7427 & n24113;
assign n3546 = n16015 | n21713;
assign n21206 = ~(n14590 ^ n12890);
assign n8036 = ~(n13263 ^ n18274);
assign n5166 = n7683 | n15774;
assign n15678 = ~(n14080 ^ n19319);
assign n19566 = n22442 & n3131;
assign n14297 = n2923 | n757;
assign n2626 = n21386 | n10763;
assign n7433 = n869 | n7601;
assign n15564 = n2263 ^ n2507;
assign n17934 = n143 | n8616;
assign n13028 = ~n3962;
assign n23515 = n9178 & n11549;
assign n1374 = n7341 | n8925;
assign n22048 = n6982 | n87;
assign n26271 = n14620 & n26914;
assign n3190 = ~n20429;
assign n24299 = n20973 & n13539;
assign n26038 = n22776 | n10353;
assign n15681 = ~(n5601 ^ n4256);
assign n5865 = ~(n12113 ^ n12917);
assign n20325 = n5140 & n14158;
assign n14696 = n8822 & n6459;
assign n20126 = ~(n5232 ^ n10289);
assign n3964 = ~(n5496 ^ n19144);
assign n13630 = n13991 | n5138;
assign n1942 = ~(n5289 ^ n26826);
assign n6390 = n2452 & n11007;
assign n19507 = n19347 | n13228;
assign n13818 = n23459 & n10603;
assign n18331 = n10918 & n5633;
assign n16959 = ~(n8358 ^ n24344);
assign n14017 = ~(n10369 | n599);
assign n27173 = ~(n15490 ^ n24032);
assign n3174 = ~(n10633 | n8378);
assign n11704 = n15623 | n13904;
assign n10364 = n3127 | n6060;
assign n3911 = ~(n25778 ^ n7223);
assign n13406 = ~(n12929 | n19005);
assign n15184 = n3253 | n6246;
assign n20048 = ~(n5934 ^ n12908);
assign n3057 = n9843 | n2024;
assign n4418 = ~(n15426 | n3136);
assign n356 = ~(n22558 | n17803);
assign n2779 = ~(n5588 ^ n9620);
assign n21989 = ~(n21021 ^ n15918);
assign n26263 = n21795 | n4762;
assign n14993 = ~(n12811 ^ n5213);
assign n17091 = n19459 & n5160;
assign n5905 = ~(n6363 ^ n16469);
assign n14163 = ~(n22246 ^ n14975);
assign n23046 = n22316 & n931;
assign n21259 = ~(n4577 | n9799);
assign n26448 = n7670 & n8227;
assign n10627 = n6691 | n21753;
assign n3694 = ~(n19423 ^ n1112);
assign n21666 = n14233 & n24082;
assign n14089 = ~(n1920 ^ n17023);
assign n24153 = n8827 | n4306;
assign n6410 = n10398 & n12629;
assign n8857 = n17046 & n18226;
assign n24503 = ~n14885;
assign n10077 = ~(n14351 ^ n18644);
assign n27144 = ~n14437;
assign n16332 = n8780 & n17622;
assign n52 = n20455 & n2884;
assign n23076 = ~(n5150 ^ n11433);
assign n8680 = ~n27120;
assign n3676 = n18125 | n10970;
assign n22093 = ~n21470;
assign n7934 = n25658 | n7379;
assign n24528 = n8777 | n10122;
assign n26683 = n11559 | n10405;
assign n6972 = ~n16888;
assign n20597 = ~n592;
assign n20110 = n17910 & n5546;
assign n8149 = ~(n12257 ^ n26718);
assign n3621 = n18797 | n11221;
assign n1716 = ~(n7099 ^ n2035);
assign n19644 = n26999 & n14244;
assign n65 = n8521 & n4652;
assign n19893 = n1677 | n20264;
assign n14486 = ~n20517;
assign n4240 = ~n21111;
assign n2087 = ~(n25120 | n17458);
assign n20632 = n2564 | n10695;
assign n10188 = ~n11265;
assign n1245 = ~(n10412 ^ n2992);
assign n15401 = ~(n2187 ^ n9572);
assign n26720 = n15436 & n7485;
assign n13281 = n22118 & n7058;
assign n5448 = n208 & n2496;
assign n26339 = n9999 & n9629;
assign n18815 = n15538 & n7971;
assign n15512 = ~n25243;
assign n14860 = ~n4719;
assign n6748 = n3933 & n21079;
assign n22999 = ~(n24245 ^ n1654);
assign n21696 = ~n3643;
assign n3066 = n21002 & n21906;
assign n21853 = ~n13453;
assign n15150 = ~(n24536 ^ n20150);
assign n10244 = ~(n20461 ^ n25952);
assign n22217 = ~(n7172 ^ n11738);
assign n10385 = ~(n26873 ^ n10680);
assign n10762 = n26093 | n10529;
assign n9662 = n26686 & n5571;
assign n23601 = ~(n2583 | n17845);
assign n17265 = n1222 | n15818;
assign n5324 = ~(n15215 ^ n10910);
assign n25756 = ~(n14742 ^ n13222);
assign n3699 = n9854 & n14955;
assign n22926 = ~n864;
assign n12758 = n3670 | n17199;
assign n8776 = ~(n19869 ^ n23805);
assign n10918 = ~n13580;
assign n5777 = n25096 | n6420;
assign n22502 = ~(n21095 ^ n25316);
assign n15708 = n7733 | n16549;
assign n6647 = n4713 & n14067;
assign n12671 = ~(n11211 | n3547);
assign n658 = ~n11192;
assign n21047 = n10339 & n3505;
assign n11131 = ~(n27143 | n15572);
assign n14701 = ~(n3168 ^ n3484);
assign n22856 = n18438 | n12081;
assign n11210 = ~(n3469 ^ n10354);
assign n5937 = n16926 & n18942;
assign n913 = ~(n15282 | n23268);
assign n11233 = n16890 | n18157;
assign n15628 = ~(n14160 ^ n17170);
assign n11599 = n20598 | n1491;
assign n5495 = ~n10534;
assign n9523 = ~n20835;
assign n8577 = ~(n25049 ^ n2872);
assign n4718 = ~(n26483 | n12088);
assign n8465 = n25421 & n6570;
assign n13526 = n5726 & n22578;
assign n435 = ~(n22342 | n16993);
assign n25511 = n26959 & n19687;
assign n5817 = ~(n4132 ^ n4282);
assign n16885 = ~(n3958 ^ n11002);
assign n20952 = ~(n19469 | n9399);
assign n11655 = ~(n2518 | n8272);
assign n10285 = n8343 | n8305;
assign n24589 = n730 | n7352;
assign n12528 = n21313 | n20230;
assign n19626 = n26516 & n16052;
assign n940 = n17211 ^ n4939;
assign n16022 = ~n5263;
assign n7439 = ~n23109;
assign n24546 = n9777 | n8502;
assign n2152 = ~n16808;
assign n18226 = n17944 | n24291;
assign n12829 = ~(n15998 ^ n12386);
assign n6280 = n5814 & n51;
assign n26161 = ~n15698;
assign n17287 = ~n9967;
assign n8509 = ~n5302;
assign n19354 = ~(n11793 ^ n9317);
assign n20049 = ~(n13169 ^ n17696);
assign n13058 = ~(n14680 | n25240);
assign n17851 = n20429 & n22365;
assign n21902 = n17095 | n26713;
assign n23331 = ~(n26488 ^ n18907);
assign n13174 = n19229 | n12929;
assign n26898 = n15734 | n18664;
assign n963 = n22015 & n16334;
assign n26829 = ~(n468 ^ n17911);
assign n704 = ~n3746;
assign n4290 = n22147 & n25720;
assign n1937 = ~(n11186 | n12464);
assign n1215 = ~n19584;
assign n2677 = n14537 & n25986;
assign n26568 = ~(n5752 | n22780);
assign n26638 = n3512 & n25970;
assign n24394 = n10140 & n26525;
assign n997 = ~(n9600 | n17613);
assign n10618 = ~(n16793 ^ n7089);
assign n5734 = n19808 & n562;
assign n26730 = n4434 | n23098;
assign n26383 = n12793 & n16352;
assign n26635 = n12495 & n24851;
assign n1190 = ~n14024;
assign n21979 = ~(n20907 | n18107);
assign n24164 = ~n13419;
assign n4156 = ~(n21082 ^ n8026);
assign n26902 = ~(n8221 ^ n3880);
assign n63 = ~n10275;
assign n4094 = ~(n4895 | n8393);
assign n19624 = ~n17069;
assign n15934 = n9852 | n10368;
assign n19888 = ~n8626;
assign n4178 = n12111 & n11217;
assign n23872 = ~(n12151 ^ n7496);
assign n5469 = ~(n2768 ^ n24327);
assign n23582 = ~n7030;
assign n8571 = ~n20359;
assign n19622 = n20695 | n5592;
assign n21096 = n180 | n6442;
assign n27023 = n16254 | n22988;
assign n15954 = n5007 | n22233;
assign n16603 = n2639 & n8257;
assign n11509 = ~(n11764 ^ n10349);
assign n27010 = ~(n10505 ^ n12153);
assign n26958 = ~(n2633 ^ n4181);
assign n10423 = ~(n14388 ^ n21575);
assign n10886 = n7285 | n14600;
assign n11605 = ~(n2219 ^ n8059);
assign n5646 = n9174 & n23991;
assign n25957 = ~(n24619 ^ n19115);
assign n14301 = ~n2715;
assign n12911 = ~n8292;
assign n12870 = ~(n1131 ^ n13412);
assign n24985 = n3410 | n388;
assign n14942 = ~(n9827 | n24280);
assign n22809 = n12871 & n20411;
assign n1300 = ~(n5012 | n17578);
assign n4037 = ~(n25126 ^ n19575);
assign n16448 = ~(n12509 ^ n7761);
assign n25452 = ~(n4343 ^ n14976);
assign n8048 = n2113 | n148;
assign n4238 = n19903 | n2020;
assign n22674 = n3356 | n26860;
assign n23749 = ~(n19444 ^ n20689);
assign n24257 = n6546 & n6694;
assign n26631 = n16155 | n5442;
assign n13366 = ~(n2540 | n24688);
assign n14315 = n3475 & n22949;
assign n22049 = ~n18519;
assign n654 = n6573 & n17719;
assign n14078 = n23094 & n18897;
assign n7688 = ~(n25565 | n24374);
assign n17841 = n24839 | n10219;
assign n12710 = n14645 | n14429;
assign n20562 = ~n23819;
assign n1685 = ~(n26163 ^ n6850);
assign n14521 = ~(n10635 ^ n6250);
assign n12785 = n1679 | n21913;
assign n15277 = ~(n854 ^ n15206);
assign n22664 = ~(n2926 | n17010);
assign n21519 = n19663 | n8025;
assign n14360 = n5717 & n4046;
assign n3931 = ~n21082;
assign n11180 = n19888 | n22414;
assign n26382 = n16044 | n10772;
assign n12321 = n20181 | n18037;
assign n17009 = n2142 | n15544;
assign n7062 = n2944 | n22270;
assign n26517 = n22817 | n22066;
assign n19440 = n11089 | n4955;
assign n2943 = ~(n5990 ^ n7326);
assign n7416 = ~(n9871 ^ n8240);
assign n27041 = n2812 & n5736;
assign n525 = n19271 & n22232;
assign n19948 = ~(n18883 ^ n21095);
assign n22410 = ~n26944;
assign n11730 = ~(n3882 ^ n22387);
assign n23917 = ~(n6946 ^ n20124);
assign n24622 = ~(n5261 ^ n20169);
assign n6111 = ~(n11840 | n15423);
assign n26834 = ~n7373;
assign n8883 = n26870 | n7902;
assign n6085 = ~n20635;
assign n11801 = ~(n2750 ^ n7543);
assign n10985 = ~(n682 | n3632);
assign n12922 = n26377 | n25076;
assign n10182 = n24523 | n22296;
assign n19245 = ~(n10778 ^ n22574);
assign n24001 = n21297 | n25993;
assign n3894 = n18364 & n13655;
assign n120 = ~n19922;
assign n13285 = ~(n46 ^ n26055);
assign n616 = ~(n2482 | n7448);
assign n23308 = n18444 | n25059;
assign n12858 = n17539 | n246;
assign n5442 = n21939 & n20298;
assign n13608 = n553 | n27200;
assign n3061 = ~(n15332 | n14792);
assign n23607 = n1412 & n9848;
assign n271 = ~(n11173 ^ n12874);
assign n2524 = ~(n12143 ^ n7258);
assign n22298 = ~(n5821 ^ n19698);
assign n15092 = n24230 | n7900;
assign n18882 = ~n22442;
assign n10661 = ~(n10527 | n4307);
assign n20353 = ~(n23568 ^ n1660);
assign n13081 = n19048 | n16955;
assign n10014 = n514 & n105;
assign n11176 = ~(n4076 | n13541);
assign n19681 = ~(n2423 ^ n24208);
assign n8820 = ~(n1306 ^ n6364);
assign n25744 = ~(n17959 | n13784);
assign n4580 = n15324 & n4795;
assign n9760 = ~(n25795 ^ n11587);
assign n3160 = ~(n24928 | n24510);
assign n26865 = n4463 & n11288;
assign n19148 = ~(n24972 ^ n5429);
assign n11008 = ~(n9921 ^ n9293);
assign n11991 = n17463 | n11115;
assign n6119 = ~(n20192 ^ n12481);
assign n1415 = ~(n10029 | n26004);
assign n16795 = ~(n4086 | n17858);
assign n8030 = n13888 | n19316;
assign n22878 = n23144 & n24371;
assign n10586 = n4469 & n5987;
assign n15785 = n22724 | n17610;
assign n18113 = ~n7119;
assign n25889 = n4427 & n4161;
assign n21015 = ~n11011;
assign n24338 = ~(n17173 | n7731);
assign n13090 = n168 & n20940;
assign n26399 = ~(n18174 ^ n7841);
assign n20662 = n24118 & n2525;
assign n13642 = ~(n354 ^ n19858);
assign n24642 = n15887 | n10153;
assign n7047 = n16467 | n26061;
assign n19593 = n1215 & n23715;
assign n4191 = ~n16638;
assign n6322 = n17355 | n19036;
assign n8942 = n16272 & n17024;
assign n18822 = n2486 | n20015;
assign n283 = n4243 | n15306;
assign n7393 = ~n1999;
assign n22475 = n7949 & n16609;
assign n2285 = ~(n7457 ^ n2615);
assign n18287 = ~(n2886 | n16609);
assign n16836 = n1904 | n26667;
assign n24820 = n13790 & n20679;
assign n10841 = n26408 & n1186;
assign n15996 = ~(n10126 ^ n11888);
assign n13079 = ~n19730;
assign n3078 = ~(n4716 ^ n15314);
assign n4853 = ~n23605;
assign n914 = ~(n13543 ^ n19234);
assign n9638 = n13190 & n23999;
assign n24718 = n4434 & n23098;
assign n801 = ~(n7542 ^ n2478);
assign n1381 = n25590 | n20800;
assign n1656 = ~(n17911 | n25331);
assign n1168 = ~(n22906 ^ n23369);
assign n18278 = n7226 | n23727;
assign n13878 = n20553 | n3165;
assign n2517 = ~(n20902 ^ n5991);
assign n13979 = ~n8844;
assign n26806 = n18327 | n24694;
assign n21232 = ~(n7505 ^ n25473);
assign n6206 = ~n21333;
assign n8804 = n18189 | n16590;
assign n23472 = n20470 | n18634;
assign n3617 = ~(n21539 ^ n13050);
assign n16949 = n20358 & n16560;
assign n5071 = ~(n9888 | n25115);
assign n1988 = n905 | n7435;
assign n26372 = n17302 | n18054;
assign n12498 = n26442 | n11524;
assign n26391 = ~(n9124 | n5483);
assign n2716 = n896 | n22915;
assign n6528 = n9509 & n6566;
assign n22259 = ~(n6724 | n485);
assign n24426 = n22987 | n6397;
assign n11284 = ~(n3783 ^ n26452);
assign n304 = ~n14330;
assign n12535 = ~n919;
assign n12891 = n19263;
assign n23514 = ~(n20047 ^ n9002);
assign n4387 = ~(n22700 ^ n18345);
assign n8443 = n23625 | n14101;
assign n864 = n19201 | n27189;
assign n15391 = n23913 | n8144;
assign n9657 = n7168 | n6068;
assign n8646 = ~(n12271 | n16233);
assign n23248 = ~(n20435 ^ n3281);
assign n25656 = ~(n27150 ^ n253);
assign n21691 = ~n24085;
assign n1192 = ~n8331;
assign n19267 = ~n16233;
assign n11096 = ~n11510;
assign n7626 = n10928 | n1616;
assign n19817 = ~(n24319 ^ n6971);
assign n3637 = n14155 & n12004;
assign n26669 = n21925 & n24763;
assign n11423 = n4837 | n22995;
assign n23834 = ~(n2100 ^ n22795);
assign n12237 = n9003 & n1735;
assign n7456 = n9097 & n16344;
assign n3956 = ~(n11745 | n10017);
assign n4414 = n14543 | n6988;
assign n18760 = ~(n24312 ^ n10847);
assign n10574 = ~(n24786 | n20754);
assign n12362 = ~(n19626 | n151);
assign n15809 = ~n15766;
assign n14543 = ~n17679;
assign n15517 = n26186 & n1028;
assign n17339 = ~n5599;
assign n21863 = n15560 | n300;
assign n4000 = ~(n26677 ^ n26330);
assign n22866 = n5394 | n19739;
assign n21335 = ~(n12902 ^ n26634);
assign n15340 = n18705 & n8083;
assign n24722 = ~(n3354 ^ n1834);
assign n14224 = n23832 | n19238;
assign n20274 = ~n14941;
assign n11394 = ~n19162;
assign n8408 = ~(n4786 | n4608);
assign n23741 = n25221 | n19425;
assign n22170 = ~n26452;
assign n7672 = n12958 & n14413;
assign n25303 = ~(n25877 ^ n5026);
assign n24340 = ~(n3295 ^ n12463);
assign n2833 = ~(n25289 | n4195);
assign n4124 = ~(n25877 ^ n10057);
assign n24759 = n24022 & n1043;
assign n5253 = ~(n21576 ^ n21559);
assign n7127 = n9469 | n14094;
assign n23881 = n8294 & n10476;
assign n3830 = ~(n12543 ^ n9090);
assign n4893 = ~(n5699 ^ n20025);
assign n25845 = n26871 | n15791;
assign n666 = n2855 & n19287;
assign n7101 = n10885 & n19276;
assign n2207 = ~(n26224 | n18483);
assign n12349 = ~(n27180 ^ n21511);
assign n19093 = n16718 | n22218;
assign n4065 = n5272 & n22526;
assign n9182 = ~(n6324 ^ n14531);
assign n21874 = ~(n7696 ^ n11017);
assign n1089 = ~(n26318 | n11248);
assign n8452 = n10310 & n14093;
assign n3658 = n10071 | n6490;
assign n8290 = n6508 | n13336;
assign n4756 = ~(n15437 ^ n8001);
assign n16694 = ~(n6553 ^ n12446);
assign n12882 = n18745 | n5510;
assign n17453 = ~n25972;
assign n4605 = ~n7828;
assign n3874 = n20733 | n3710;
assign n12065 = n6165 & n23183;
assign n1671 = ~(n3919 ^ n26105);
assign n2437 = n10418 | n19211;
assign n384 = ~(n23921 | n130);
assign n15775 = ~(n1122 ^ n5365);
assign n764 = n3243 | n17073;
assign n17170 = ~(n1630 ^ n4326);
assign n4742 = n16511 | n25825;
assign n1224 = ~(n5604 | n7026);
assign n19359 = ~(n20131 | n17418);
assign n25815 = ~(n1753 ^ n19457);
assign n14286 = n1359 | n7252;
assign n9458 = ~(n18910 ^ n4168);
assign n7992 = ~(n18401 ^ n12772);
assign n26820 = n958 | n9658;
assign n20059 = ~n5956;
assign n4919 = n12562 | n23978;
assign n20740 = ~(n15295 | n3195);
assign n7450 = n18475 & n15197;
assign n11617 = ~(n15743 ^ n13319);
assign n14919 = ~(n2646 ^ n22072);
assign n19734 = ~(n19806 ^ n24024);
assign n19160 = n20576 & n15349;
assign n26569 = n20137 | n17601;
assign n15686 = ~n10069;
assign n26659 = n21556 | n21207;
assign n24672 = n11816 | n8649;
assign n25649 = ~(n342 | n14570);
assign n8940 = n1379 & n9105;
assign n4197 = n20491 | n20769;
assign n21288 = ~n24440;
assign n19236 = ~(n11117 ^ n21980);
assign n3094 = ~n26053;
assign n18580 = ~(n24306 | n9116);
assign n1155 = ~n20966;
assign n16193 = n12967 & n11030;
assign n23839 = n1935 | n17552;
assign n3584 = ~(n16184 ^ n13247);
assign n10705 = ~(n25036 ^ n11016);
assign n2360 = ~n20687;
assign n24247 = n27111 & n3391;
assign n16692 = ~(n18861 ^ n10251);
assign n4057 = n26503 & n25702;
assign n25906 = n17770 & n12629;
assign n5959 = n1107 | n17257;
assign n5110 = ~(n24846 ^ n16714);
assign n9716 = n6508 & n21710;
assign n9957 = ~n11136;
assign n5602 = ~(n21502 | n4017);
assign n5056 = n823 | n19010;
assign n382 = ~(n2764 | n9789);
assign n16689 = ~(n19228 ^ n4812);
assign n7112 = n13933 | n24275;
assign n9549 = ~(n20117 | n9460);
assign n23236 = n3110 & n9902;
assign n3615 = n20688 | n3424;
assign n671 = ~(n21253 ^ n17664);
assign n25441 = ~(n4016 ^ n24474);
assign n16076 = ~(n17871 ^ n12675);
assign n16526 = n10870 & n8187;
assign n17724 = n205 & n22842;
assign n10751 = ~(n26410 ^ n23918);
assign n4971 = n9076 | n3727;
assign n18574 = ~(n7334 ^ n6728);
assign n8740 = n3827 & n5055;
assign n3054 = ~(n25120 ^ n8526);
assign n13261 = ~(n26625 ^ n14230);
assign n16338 = n5729 | n10308;
assign n3704 = n20874 | n13819;
assign n24539 = n21672 | n18314;
assign n4243 = ~(n5768 | n2300);
assign n18107 = n7311 & n20273;
assign n10855 = n12431 & n22189;
assign n5794 = ~(n7499 ^ n1223);
assign n10189 = n11544 | n2978;
assign n21942 = ~(n16349 | n8094);
assign n9102 = n16468 & n15511;
assign n24628 = n5043 & n18133;
assign n7893 = ~n21997;
assign n1596 = n1777 | n837;
assign n22392 = ~(n6775 ^ n12121);
assign n3969 = n19631 | n14449;
assign n25222 = ~(n6169 ^ n6944);
assign n24157 = ~(n3582 | n23064);
assign n17713 = ~(n18798 ^ n25486);
assign n5174 = n20358 | n3960;
assign n15012 = n20040 & n8186;
assign n16577 = n15262 & n15310;
assign n13505 = n22816 & n23576;
assign n8198 = ~(n22651 | n6385);
assign n11355 = n5774 & n960;
assign n1304 = ~(n7717 ^ n26313);
assign n3560 = n6776 | n17917;
assign n22005 = n4048 & n14433;
assign n26988 = ~(n7871 | n8261);
assign n20381 = n6592 | n19349;
assign n12377 = ~n6730;
assign n7370 = n16854 | n26143;
assign n11391 = ~(n2679 ^ n25592);
assign n19455 = ~(n6381 ^ n16376);
assign n8368 = n25622 & n11945;
assign n25476 = ~(n16948 ^ n6379);
assign n8950 = ~(n9832 ^ n3959);
assign n17410 = ~(n11068 ^ n25474);
assign n7146 = ~(n10107 ^ n12507);
assign n26869 = n12451 | n26880;
assign n6475 = n20409 | n429;
assign n9739 = n18032 | n9440;
assign n5767 = ~(n25965 ^ n9808);
assign n17846 = ~n5555;
assign n22067 = n5618 & n12786;
assign n21184 = n9844 & n16579;
assign n24640 = n13515 | n23961;
assign n7817 = n21858;
assign n3241 = ~n7759;
assign n24520 = n2717 | n10337;
assign n8053 = ~(n9412 | n17567);
assign n17150 = n328 & n15695;
assign n26513 = ~(n15427 | n16521);
assign n17931 = ~(n15754 ^ n3810);
assign n14546 = n8908 | n10047;
assign n20116 = ~(n21596 ^ n6352);
assign n23177 = n7870 | n24759;
assign n18458 = n24290 | n6526;
assign n2303 = ~(n9476 ^ n94);
assign n12271 = ~(n8910 ^ n22392);
assign n12089 = n3801 | n20440;
assign n19483 = n22349 ^ n15743;
assign n18661 = ~(n3659 ^ n17635);
assign n2079 = ~(n17366 | n14754);
assign n11089 = ~(n18964 ^ n20397);
assign n25302 = ~(n4644 ^ n4933);
assign n21332 = n11880 | n24218;
assign n26187 = ~n24536;
assign n19112 = ~n12501;
assign n25512 = ~(n56 | n4095);
assign n22214 = n11827 | n16471;
assign n22277 = n8156 | n24178;
assign n26304 = n10461 & n10132;
assign n25543 = n12181 & n14676;
assign n23381 = ~(n4878 ^ n12692);
assign n16382 = ~(n3823 ^ n21599);
assign n14007 = ~n23913;
assign n14035 = n11707 | n20926;
assign n2235 = ~n5196;
assign n22477 = ~n9806;
assign n6909 = n9660 & n10515;
assign n22872 = ~(n5582 ^ n9717);
assign n13418 = n4960 & n11427;
assign n15762 = ~(n17574 ^ n8335);
assign n26939 = ~(n23345 ^ n5381);
assign n13429 = ~n23731;
assign n4729 = ~n16824;
assign n20124 = ~n9245;
assign n206 = n14538 | n23862;
assign n1947 = n7034 & n20573;
assign n6745 = ~(n21014 ^ n9004);
assign n15498 = ~n15170;
assign n3924 = ~(n3019 ^ n1279);
assign n9427 = ~(n26443 ^ n10017);
assign n18349 = n19575 | n16126;
assign n26470 = ~n16968;
assign n17355 = ~(n27144 | n6774);
assign n20 = ~n19951;
assign n23420 = ~(n15167 ^ n919);
assign n12463 = ~(n20811 ^ n3909);
assign n15297 = ~(n16609 ^ n2886);
assign n5870 = n10237 & n23846;
assign n10011 = n16643 & n24110;
assign n17101 = n10135 & n24863;
assign n25492 = n11303 | n2429;
assign n24295 = n26138 | n17340;
assign n20572 = ~(n22977 | n23513);
assign n18497 = ~(n3346 ^ n19311);
assign n22394 = ~(n23353 ^ n14881);
assign n4701 = n26658 | n19911;
assign n20081 = n16755 | n18812;
assign n11818 = ~(n18248 ^ n16844);
assign n11299 = ~(n9990 ^ n18097);
assign n22662 = ~(n21494 ^ n16074);
assign n12594 = n18838 | n1484;
assign n12476 = ~(n20954 ^ n21263);
assign n5029 = n25258 | n6838;
assign n22131 = ~(n22191 | n12064);
assign n2894 = ~n22272;
assign n16712 = ~n15539;
assign n11648 = ~(n7924 ^ n4767);
assign n1987 = ~n14257;
assign n17578 = ~n3211;
assign n1703 = ~(n25618 ^ n16829);
assign n23670 = ~n4601;
assign n3989 = n12603 | n11983;
assign n26378 = n4843 & n872;
assign n7998 = n21108 | n8073;
assign n14075 = n11263 & n1538;
assign n2689 = ~(n26180 | n10650);
assign n22835 = ~(n12911 ^ n26264);
assign n16889 = ~n23166;
assign n22956 = n6421 | n23674;
assign n25387 = ~(n13244 | n3462);
assign n2404 = ~(n20053 | n23876);
assign n11061 = n559 & n11705;
assign n24478 = ~(n15291 | n13401);
assign n4411 = n17542 | n4409;
assign n6409 = n24469 | n9447;
assign n13093 = ~(n27005 ^ n27188);
assign n18538 = ~(n26882 ^ n19618);
assign n22829 = ~(n2320 ^ n11736);
assign n12093 = ~(n1798 | n8930);
assign n8167 = ~n14488;
assign n22154 = ~(n22932 ^ n10316);
assign n7986 = n22238 | n9036;
assign n14139 = ~n23773;
assign n13414 = n26691 | n20036;
assign n13949 = ~(n16994 ^ n9246);
assign n1612 = n6337 & n3686;
assign n11786 = n10207 | n18833;
assign n3264 = ~(n1662 ^ n7330);
assign n26778 = n3366 & n4753;
assign n23899 = ~(n14296 ^ n23374);
assign n11219 = n18257 | n23098;
assign n6530 = n20407 | n25093;
assign n4049 = ~(n10822 ^ n18462);
assign n16198 = n12414 | n16390;
assign n484 = n25548 | n3323;
assign n14676 = n8757 | n25383;
assign n18730 = n11786 & n6384;
assign n4996 = ~(n5960 | n9942);
assign n24569 = ~(n8491 ^ n23895);
assign n10434 = n11466 & n2393;
assign n23235 = ~(n16414 ^ n3902);
assign n5679 = n26106 & n23324;
assign n6042 = ~(n3740 | n3498);
assign n20332 = n16743 | n24485;
assign n24634 = ~(n1594 ^ n16602);
assign n3111 = n2953 | n10681;
assign n16951 = ~(n20164 ^ n23299);
assign n1369 = n8755 & n22923;
assign n17220 = ~(n7081 ^ n17597);
assign n20871 = n26529 & n3939;
assign n11103 = ~(n12400 ^ n14534);
assign n3310 = n16162 | n693;
assign n10356 = n18936 | n13483;
assign n12057 = ~(n4995 ^ n24327);
assign n18233 = n5913 & n4737;
assign n7999 = ~(n14877 ^ n26359);
assign n21664 = ~(n4397 | n26178);
assign n9410 = n21177 | n21534;
assign n25093 = n4192 & n15619;
assign n6713 = ~n21945;
assign n7554 = ~(n8171 ^ n4060);
assign n24428 = ~(n2036 | n8434);
assign n27110 = ~(n21546 ^ n17922);
assign n18122 = n17339 | n15564;
assign n1467 = ~n14544;
assign n1429 = ~(n22495 ^ n3789);
assign n1319 = n24692;
assign n15567 = n15631 | n4;
assign n1807 = ~(n14990 ^ n18526);
assign n2678 = ~(n9040 ^ n7769);
assign n5763 = ~(n16889 | n4306);
assign n2461 = ~(n810 ^ n23694);
assign n21272 = n1674;
assign n21880 = n9363 | n23044;
assign n21117 = ~n26510;
assign n4058 = n18100 & n16231;
assign n3834 = ~(n26152 ^ n21262);
assign n16436 = n10275 | n22359;
assign n9916 = n5989 | n15471;
assign n21179 = n19140 & n17148;
assign n15042 = ~n10625;
assign n7528 = ~(n7270 | n16902);
assign n599 = ~n14693;
assign n13780 = n12445 | n19255;
assign n24261 = ~(n11246 ^ n26510);
assign n1053 = ~(n15998 ^ n9723);
assign n13016 = ~(n5750 | n19884);
assign n8756 = ~(n20011 ^ n5697);
assign n15570 = ~(n12944 ^ n12614);
assign n21068 = n13529 | n14720;
assign n16242 = n22158 | n8717;
assign n2814 = n13263 | n22596;
assign n4147 = n11108 | n7327;
assign n26148 = n23398 & n8183;
assign n16711 = ~n22660;
assign n11965 = ~(n26238 ^ n24259);
assign n11463 = ~(n10485 ^ n7670);
assign n22124 = ~(n11211 ^ n17627);
assign n18485 = ~n19514;
assign n26414 = ~(n12763 ^ n3740);
assign n5699 = n7251 & n26057;
assign n23646 = n9290 | n196;
assign n22499 = n5465 | n11537;
assign n16764 = ~(n16637 ^ n2776);
assign n1602 = ~(n24527 ^ n12226);
assign n19172 = ~(n26689 | n22666);
assign n4568 = n20667 | n21927;
assign n9171 = n3402 | n18440;
assign n25627 = ~n12749;
assign n17888 = ~n5800;
assign n8913 = ~(n6218 ^ n19652);
assign n19645 = n18453 | n21657;
assign n22998 = ~(n11864 ^ n10279);
assign n25027 = n14822 & n2074;
assign n7427 = n3363 | n18506;
assign n7957 = ~n18941;
assign n21904 = n8344 | n6794;
assign n12932 = ~n19327;
assign n11938 = ~n21226;
assign n4538 = n22696 & n18167;
assign n6503 = ~n592;
assign n19119 = ~n18792;
assign n20696 = ~(n26496 ^ n1621);
assign n19504 = n22133 | n14598;
assign n22450 = ~(n7249 ^ n5182);
assign n8089 = ~(n26584 ^ n12204);
assign n16252 = ~n4306;
assign n19822 = n16482 | n13333;
assign n5440 = ~n14148;
assign n22194 = ~n3945;
assign n16554 = n7151 | n21427;
assign n14500 = ~n18827;
assign n13997 = n25425 & n20368;
assign n3910 = n21995 | n25789;
assign n18627 = n2259 | n10991;
assign n15283 = n19095 | n4783;
assign n11687 = n6394 | n9273;
assign n18959 = ~(n11056 ^ n18157);
assign n7797 = ~(n14732 ^ n10965);
assign n2972 = n104 | n20927;
assign n21588 = n15079 | n5752;
assign n18296 = ~(n24704 | n5728);
assign n23914 = n25972 & n3707;
assign n14252 = ~(n21502 ^ n4017);
assign n19808 = n6523 | n14298;
assign n2667 = ~(n25515 ^ n27066);
assign n13332 = ~(n26565 | n20437);
assign n23963 = n4658 | n11442;
assign n19288 = n3349 | n12762;
assign n9862 = n22059 | n25723;
assign n18381 = ~(n13231 | n27115);
assign n8529 = ~n15264;
assign n14911 = n22291 | n6874;
assign n22024 = ~(n15884 | n25602);
assign n938 = n9688 & n22466;
assign n20849 = ~(n8508 ^ n12153);
assign n9408 = n22523 | n24698;
assign n3650 = n89 & n10396;
assign n24207 = n4084 & n26051;
assign n7800 = n13657 | n15941;
assign n15734 = ~n9077;
assign n25855 = ~(n1032 ^ n19877);
assign n27113 = n24355 & n1267;
assign n8763 = ~(n22723 ^ n5692);
assign n4152 = ~(n10857 ^ n8133);
assign n6078 = ~(n329 ^ n21735);
assign n14368 = n382 | n10812;
assign n19755 = ~n1853;
assign n11450 = n12040 | n21459;
assign n17956 = ~(n9579 ^ n956);
assign n4549 = ~n313;
assign n10869 = ~(n11835 ^ n9179);
assign n17750 = n1537 | n13246;
assign n7017 = ~(n26046 | n23512);
assign n22252 = ~(n9631 | n18300);
assign n200 = n2422 & n1562;
assign n4248 = ~(n22346 | n23033);
assign n9156 = n6050 & n14898;
assign n16145 = n23752 | n26078;
assign n19030 = ~n9485;
assign n1941 = ~n15210;
assign n22231 = n13577 | n11944;
assign n24236 = n2915 | n23559;
assign n13038 = ~(n7380 ^ n24191);
assign n9375 = ~(n13359 ^ n7057);
assign n429 = n25749 | n18507;
assign n5576 = n23489 | n6733;
assign n23629 = ~(n17423 | n19914);
assign n18192 = ~(n17505 | n5465);
assign n19478 = ~(n23052 ^ n17038);
assign n9275 = n10008 | n13460;
assign n25209 = ~(n3237 ^ n2695);
assign n25967 = ~n847;
assign n5428 = ~(n2490 ^ n20447);
assign n22537 = ~(n18044 ^ n5383);
assign n21159 = ~(n19702 ^ n23849);
assign n21358 = ~(n10204 ^ n16158);
assign n24386 = n1382 & n4252;
assign n22640 = ~(n16450 ^ n18926);
assign n15170 = ~(n9008 ^ n23505);
assign n14372 = n9008 & n16145;
assign n23410 = ~(n4333 ^ n8869);
assign n4972 = ~(n26938 ^ n732);
assign n3965 = n17915 & n26049;
assign n1047 = ~(n7493 ^ n11860);
assign n15032 = n24250 & n22263;
assign n4194 = ~n15408;
assign n16827 = n524 | n24947;
assign n7942 = ~(n1365 | n19234);
assign n7920 = n9637 | n13680;
assign n12109 = ~(n18003 | n26013);
assign n16747 = ~(n13459 | n1689);
assign n1916 = ~n10344;
assign n9045 = n21957 | n14410;
assign n21318 = n4833 | n24221;
assign n26451 = ~(n9883 | n11016);
assign n13245 = ~n5307;
assign n9932 = n23762 & n2053;
assign n2086 = ~n3849;
assign n4641 = n8125 & n2550;
assign n6430 = n6122 ^ n19196;
assign n24497 = n25028 & n10871;
assign n20403 = ~(n18470 ^ n10793);
assign n12757 = n692 | n1991;
assign n20389 = ~(n7803 ^ n21630);
assign n15279 = n10751 | n14466;
assign n17736 = n7517 | n1026;
assign n17989 = n6715 & n3159;
assign n4627 = n25043 | n17901;
assign n8124 = n23758 | n10361;
assign n2935 = ~n16051;
assign n2876 = n25306 & n8038;
assign n11643 = ~(n11597 | n12888);
assign n3677 = ~n921;
assign n9608 = ~(n10608 ^ n12587);
assign n11712 = ~(n16463 ^ n16258);
assign n16460 = ~(n16710 ^ n11801);
assign n21289 = n15820 & n21824;
assign n19564 = n13076 & n17492;
assign n17283 = n15928 | n8444;
assign n11885 = n4801 & n11970;
assign n399 = ~(n5128 | n22926);
assign n314 = ~(n22764 ^ n2416);
assign n15794 = ~(n23166 ^ n18105);
assign n15449 = n3503 | n1875;
assign n8997 = ~(n17294 ^ n335);
assign n20303 = ~(n2909 | n19312);
assign n5339 = n18938 & n19957;
assign n6823 = n3586 | n1285;
assign n4279 = n16514 & n21825;
assign n26375 = ~(n19434 ^ n26965);
assign n21309 = ~(n25960 ^ n1102);
assign n22249 = ~(n11229 ^ n17195);
assign n7847 = n4304 | n23876;
assign n15736 = n2268 & n19153;
assign n21458 = ~(n15478 ^ n7369);
assign n18506 = ~n19228;
assign n12366 = ~n18183;
assign n21395 = n14936 | n15233;
assign n175 = ~(n18772 ^ n17654);
assign n4244 = n26465 | n9758;
assign n9385 = n6438 | n6473;
assign n3315 = n12400 & n2966;
assign n2797 = n25778 & n3134;
assign n7580 = ~(n12351 ^ n14323);
assign n6512 = n8746 | n620;
assign n10746 = ~(n1978 ^ n22884);
assign n7053 = ~(n26299 ^ n25208);
assign n4234 = n690 | n13036;
assign n13838 = n26557 | n4670;
assign n6185 = ~(n25595 ^ n909);
assign n10118 = n25891 | n2312;
assign n23519 = n6253 | n20664;
assign n26135 = ~(n4465 ^ n10271);
assign n338 = n5211 | n21832;
assign n12990 = ~n11589;
assign n13123 = ~(n12436 ^ n19475);
assign n23986 = ~(n16044 ^ n8113);
assign n1262 = ~n21832;
assign n13471 = n9027 | n22112;
assign n1032 = n22151 | n10960;
assign n9729 = n8713 | n6071;
assign n2261 = ~n23285;
assign n20606 = n3937 | n1243;
assign n3248 = ~(n1946 | n6648);
assign n17806 = ~n13452;
assign n5570 = n20453 & n1361;
assign n8839 = n1829 | n15371;
assign n10494 = ~(n2145 | n22021);
assign n179 = n24050 | n25737;
assign n7131 = ~(n3374 ^ n27101);
assign n25127 = n9623 & n3262;
assign n25726 = ~n5072;
assign n3686 = ~(n6261 ^ n19685);
assign n25121 = n19358 & n25302;
assign n18266 = n15827 & n15073;
assign n16510 = n5730 & n4825;
assign n6931 = n2577 & n4421;
assign n22291 = ~(n12396 | n20064);
assign n20805 = n2187 | n2161;
assign n12253 = n21886 | n2983;
assign n14244 = ~n7833;
assign n20757 = ~(n25345 ^ n9967);
assign n18788 = ~(n15636 | n18255);
assign n3816 = n16497 | n6848;
assign n2957 = ~(n7755 | n21097);
assign n10802 = ~n13468;
assign n784 = n14218 & n7737;
assign n5747 = n17041 & n25626;
assign n6937 = n23623 | n5412;
assign n1368 = n20983 & n18082;
assign n13800 = n20527 & n2525;
assign n21446 = ~(n25205 ^ n20356);
assign n9152 = ~(n10314 ^ n10242);
assign n21441 = n26912 ^ n13038;
assign n12290 = n16355 | n11371;
assign n19602 = ~(n24168 ^ n8271);
assign n1134 = n20826 | n14532;
assign n9785 = n7914 | n17767;
assign n19944 = ~n26979;
assign n6833 = ~n23039;
assign n25831 = ~(n13492 ^ n16536);
assign n20853 = ~(n23990 | n16960);
assign n21122 = n3145 & n10453;
assign n275 = ~(n23408 | n22660);
assign n17107 = n1540 | n13424;
assign n1523 = ~(n4576 ^ n17302);
assign n18591 = ~(n570 | n16211);
assign n16187 = n7065 | n18480;
assign n22825 = n26890 | n24117;
assign n19865 = ~(n3823 | n12262);
assign n12915 = n25204 | n19309;
assign n692 = ~(n4422 ^ n10442);
assign n5295 = ~(n20228 | n8717);
assign n11563 = n14736 | n21226;
assign n8674 = ~(n5122 ^ n19976);
assign n1071 = n18957 & n21660;
assign n4673 = ~n11810;
assign n12347 = n9295 & n15786;
assign n10986 = ~n3651;
assign n13181 = n22216 | n539;
assign n24397 = ~(n7756 | n20683);
assign n3782 = n5169 | n2085;
assign n2098 = n21649 & n17846;
assign n13131 = ~(n19701 | n7437);
assign n6544 = ~(n23529 ^ n10739);
assign n11520 = n12609 | n6954;
assign n23440 = n6834 | n5165;
assign n19859 = n22419 & n20390;
assign n14944 = ~(n3133 ^ n4379);
assign n7815 = n15541 & n16043;
assign n17441 = n13588 | n16318;
assign n8243 = n18355 | n21822;
assign n1895 = ~(n26716 ^ n16301);
assign n16366 = ~(n11654 ^ n8006);
assign n18318 = ~n3471;
assign n14109 = n16968 & n27189;
assign n22716 = ~(n13896 ^ n4661);
assign n19786 = n23015 | n24754;
assign n7336 = n25369 | n21329;
assign n20056 = ~n4877;
assign n15824 = n1558 | n5050;
assign n20154 = n21792 | n1478;
assign n10826 = n5226 & n11223;
assign n3351 = ~(n9076 | n24805);
assign n5994 = n3568 | n18202;
assign n18812 = ~(n18918 ^ n11787);
assign n16313 = ~n23833;
assign n3313 = n8568 | n1600;
assign n15933 = n11554 | n25521;
assign n9871 = n7728 & n1699;
assign n10862 = n21868 | n7892;
assign n7512 = n1762 | n711;
assign n19632 = ~n18314;
assign n15600 = n11503 | n18151;
assign n26508 = ~n15761;
assign n12718 = ~(n13650 | n14025);
assign n19156 = n22426 | n12543;
assign n8130 = ~(n3328 ^ n14970);
assign n8627 = n21777 | n4685;
assign n7523 = ~(n23556 ^ n27089);
assign n16780 = n13953 | n17511;
assign n4241 = ~(n2453 | n22492);
assign n16850 = n1492 & n6077;
assign n19124 = n25273 | n25777;
assign n3725 = ~(n9902 ^ n10913);
assign n19731 = n23104;
assign n21472 = ~(n19810 ^ n12273);
assign n26361 = n14518 | n18806;
assign n8007 = n16364 | n15495;
assign n7322 = n8094 | n5580;
assign n6476 = ~(n69 ^ n11593);
assign n8003 = ~n15643;
assign n22114 = n17013 & n7799;
assign n19209 = ~(n12009 | n10259);
assign n13771 = n5077 | n13914;
assign n7342 = n12513 & n8162;
assign n20007 = n18894 | n5186;
assign n27108 = ~(n161 ^ n12780);
assign n19834 = ~(n19236 ^ n21930);
assign n14588 = n744 | n9363;
assign n18238 = ~(n4394 ^ n672);
assign n15334 = ~(n4201 | n3045);
assign n3555 = ~(n22966 ^ n24722);
assign n17600 = ~(n16069 ^ n21673);
assign n10313 = n407 & n9717;
assign n14901 = n4034 & n15208;
assign n10424 = ~n665;
assign n26575 = n3309 & n23177;
assign n8335 = ~(n6731 ^ n7347);
assign n23459 = n4177 & n19482;
assign n17795 = n15318 & n7758;
assign n26747 = ~n21687;
assign n1098 = n4132 | n24301;
assign n25015 = ~n18125;
assign n12482 = n16743 | n5194;
assign n1638 = n9165 | n11319;
assign n9925 = ~(n22472 | n9125);
assign n1115 = n8333 & n7908;
assign n15799 = ~(n3681 | n18383);
assign n9188 = n17512 & n9606;
assign n7518 = ~(n5374 ^ n23002);
assign n26423 = ~(n17663 | n22862);
assign n25638 = n26845 | n3790;
assign n22152 = n1462 & n20007;
assign n13162 = n9378 & n10833;
assign n13462 = n13531 & n9745;
assign n17563 = ~(n10467 ^ n593);
assign n12022 = ~n19646;
assign n2648 = n6305 | n9197;
assign n18754 = ~n15910;
assign n10873 = ~(n11726 ^ n8401);
assign n14117 = ~(n2915 | n8363);
assign n20302 = ~(n19327 ^ n21934);
assign n18219 = n10156 & n26782;
assign n18084 = n838 & n10676;
assign n877 = n13103 | n14321;
assign n13455 = ~(n11988 ^ n17880);
assign n19790 = n26875 | n18487;
assign n10355 = ~(n13693 ^ n12650);
assign n13013 = n4278 & n15074;
assign n13600 = n22365 | n15359;
assign n11513 = ~(n21317 | n19196);
assign n18867 = ~n16078;
assign n25704 = ~n23653;
assign n20513 = ~n19540;
assign n15621 = n1356 | n13341;
assign n551 = ~(n13231 ^ n27115);
assign n9186 = n5113 | n5283;
assign n4323 = n19304 | n15497;
assign n3331 = n12534 | n3004;
assign n20260 = ~n80;
assign n20458 = ~(n11958 ^ n11483);
assign n10571 = ~n23213;
assign n10883 = n21471 | n19357;
assign n8135 = ~(n9092 ^ n13877);
assign n7600 = n25946 & n12512;
assign n22803 = n24200 | n14648;
assign n18541 = n7600 & n16757;
assign n24951 = ~(n26995 ^ n11658);
assign n11166 = ~(n16294 | n2160);
assign n3932 = ~(n11660 ^ n11512);
assign n17803 = ~n19691;
assign n4541 = n846 | n8407;
assign n23522 = n22083 | n1304;
assign n26389 = n3510 | n21523;
assign n24616 = ~(n4635 ^ n857);
assign n14644 = n22763 | n26865;
assign n9882 = n23063 | n11486;
assign n22241 = ~(n26919 ^ n11322);
assign n20238 = n17644 & n8924;
assign n7032 = ~(n12629 ^ n23212);
assign n5972 = n5512 | n27071;
assign n522 = ~(n20937 | n424);
assign n9192 = ~(n22254 ^ n22699);
assign n12090 = ~n6819;
assign n23905 = ~n23318;
assign n12620 = ~(n16151 ^ n18898);
assign n18886 = ~(n7723 ^ n25892);
assign n9656 = n20077 | n6794;
assign n1918 = ~(n9680 | n7364);
assign n13083 = n12789 | n23218;
assign n20876 = n6018 & n10099;
assign n18692 = ~(n330 ^ n5668);
assign n24298 = ~(n6224 ^ n11696);
assign n12728 = ~(n2308 | n2489);
assign n24537 = ~(n2381 ^ n22377);
assign n26923 = ~(n20834 ^ n16273);
assign n4581 = n26053 | n25461;
assign n12873 = ~(n18233 ^ n15535);
assign n24364 = ~n27146;
assign n2106 = ~(n25877 | n10057);
assign n21387 = n5363 | n9328;
assign n86 = ~(n3094 | n2191);
assign n23367 = n24273 | n14630;
assign n3395 = n14718 | n23705;
assign n15230 = ~(n13286 ^ n8514);
assign n20973 = ~(n5179 ^ n129);
assign n26736 = n16135 | n9168;
assign n7666 = ~(n25240 | n20707);
assign n9706 = n328 & n19387;
assign n12927 = n17522 & n9410;
assign n3449 = n1432 | n12040;
assign n27016 = n20952 | n20262;
assign n8916 = n8677 | n15146;
assign n26358 = ~(n910 | n12891);
assign n25776 = n18861 | n693;
assign n11834 = ~n22437;
assign n18764 = n21016 | n23956;
assign n3864 = n16565 | n11982;
assign n19812 = n16452 | n26840;
assign n21529 = ~(n21798 ^ n23969);
assign n5779 = ~(n4062 ^ n16499);
assign n13037 = n10908;
assign n15810 = n12602 & n24775;
assign n18088 = ~(n22660 | n24774);
assign n8264 = n18309 & n7433;
assign n3689 = n26530 & n25465;
assign n22564 = n20702 | n17774;
assign n15798 = n17402 & n5691;
assign n18940 = ~(n22532 ^ n15548);
assign n26738 = ~(n12650 | n13693);
assign n8728 = ~(n22410 ^ n15610);
assign n12163 = n4730 & n14030;
assign n9021 = ~(n11578 ^ n7335);
assign n17514 = n20728 & n1036;
assign n19697 = n22652 | n6267;
assign n10159 = ~n604;
assign n21257 = ~(n21784 | n18163);
assign n16804 = n5219 & n24454;
assign n487 = ~(n18869 | n10741);
assign n7813 = n22023 & n1017;
assign n3700 = n8189 & n24994;
assign n24906 = n7496 | n12151;
assign n9067 = ~n16965;
assign n18746 = ~n5098;
assign n8837 = ~(n18947 ^ n26797);
assign n7201 = n17578 | n8653;
assign n5167 = ~(n26747 ^ n9380);
assign n21392 = ~n11640;
assign n2407 = ~n16803;
assign n27067 = ~(n19110 ^ n10522);
assign n17074 = ~(n13734 ^ n6019);
assign n17774 = ~(n5919 | n3653);
assign n2909 = n27117 & n13836;
assign n25650 = ~n13851;
assign n10377 = n9286 & n7629;
assign n20198 = ~(n16009 ^ n6397);
assign n20029 = ~(n19249 ^ n12884);
assign n22284 = n18651 & n25307;
assign n6529 = n26227 & n23101;
assign n9634 = n20329 | n25464;
assign n16208 = ~(n6502 | n1630);
assign n19678 = n4581 & n3928;
assign n12864 = ~(n2716 ^ n18657);
assign n10969 = ~n755;
assign n19522 = n8373 & n18819;
assign n1495 = n9528 & n13055;
assign n8184 = ~(n14872 ^ n11903);
assign n25919 = ~(n977 ^ n2858);
assign n6031 = ~(n9524 ^ n2788);
assign n12833 = n23099 | n7402;
assign n5670 = n22912 | n7484;
assign n9519 = n13152 & n2688;
assign n23897 = ~(n5555 ^ n17323);
assign n14907 = n4515 & n19136;
assign n21234 = ~(n25701 ^ n1204);
assign n8416 = ~(n14696 ^ n19552);
assign n24791 = ~(n12664 ^ n24196);
assign n14093 = n17103 | n17795;
assign n23592 = ~n14130;
assign n10122 = n9735 & n2595;
assign n25612 = ~n11701;
assign n2846 = ~(n12929 | n16971);
assign n12079 = n21273 & n4302;
assign n2044 = ~n8728;
assign n16699 = n8414 | n24617;
assign n1259 = ~(n24620 | n22327);
assign n13628 = ~(n21322 ^ n19531);
assign n8774 = ~(n5133 ^ n2421);
assign n9676 = n18591 | n15726;
assign n24938 = n21247 | n24458;
assign n11578 = ~(n3171 ^ n3425);
assign n9282 = ~(n19360 | n12964);
assign n1971 = ~(n26295 ^ n16824);
assign n11574 = n25600 & n24123;
assign n8046 = ~(n7460 ^ n22068);
assign n9149 = n7377 & n21125;
assign n2045 = ~n5226;
assign n27002 = ~n2951;
assign n22692 = ~(n25419 ^ n17061);
assign n15777 = n14672 & n2258;
assign n113 = ~(n2980 | n12514);
assign n20842 = ~(n21597 | n22722);
assign n26431 = ~(n14509 ^ n825);
assign n21114 = ~n18395;
assign n7829 = ~(n5026 ^ n8581);
assign n13767 = ~n24429;
assign n7174 = ~(n6063 ^ n17862);
assign n3089 = ~(n27198 ^ n15469);
assign n14808 = n5724 & n2572;
assign n651 = n26043 | n6665;
assign n11618 = n24003 & n15472;
assign n3954 = n7757 | n16962;
assign n9273 = ~n231;
assign n23898 = ~n6819;
assign n26276 = n26329 | n4908;
assign n13694 = n17066 | n22325;
assign n1012 = ~(n23417 ^ n9513);
assign n3456 = ~(n10138 ^ n25054);
assign n23190 = ~n14256;
assign n15359 = ~(n14673 ^ n126);
assign n26740 = ~(n6501 ^ n20274);
assign n11038 = n1195 | n21412;
assign n7647 = ~(n2983 ^ n17519);
assign n4384 = ~(n19048 ^ n9536);
assign n2174 = ~n13460;
assign n20582 = ~(n19563 ^ n3189);
assign n11924 = ~n8847;
assign n26101 = n2376 | n6644;
assign n8436 = ~n13660;
assign n8682 = ~n1998;
assign n7092 = ~n5296;
assign n2526 = n12166 & n8346;
assign n17166 = ~(n17107 ^ n9228);
assign n14395 = ~n10917;
assign n13730 = n14965 | n25465;
assign n7375 = n19944 | n24366;
assign n17762 = ~(n13481 ^ n454);
assign n8293 = ~(n1777 ^ n16029);
assign n19891 = n9846 | n18099;
assign n1144 = n25113 | n24839;
assign n9367 = n4710 | n4526;
assign n22701 = n9464 & n5294;
assign n569 = n24786 | n1574;
assign n855 = n10715 & n12517;
assign n25089 = n16585 & n2751;
assign n18098 = ~(n8745 | n7532);
assign n7105 = n3923 & n12486;
assign n26928 = n13264 & n17982;
assign n301 = n23611 & n6512;
assign n7962 = ~(n13137 ^ n1288);
assign n4165 = ~(n5642 ^ n8731);
assign n16629 = n20975 | n18817;
assign n3566 = n10716 | n19132;
assign n23118 = ~n14921;
assign n4462 = ~(n17909 | n9172);
assign n23335 = n13591 | n3164;
assign n26355 = n4027 & n19065;
assign n24384 = n24850 | n12921;
assign n11323 = n26824 & n25761;
assign n18118 = n23084 & n3870;
assign n1427 = ~(n9957 | n6435);
assign n15842 = ~n3405;
assign n17319 = n8331 | n20176;
assign n20535 = ~n22057;
assign n18854 = ~(n11451 ^ n19770);
assign n10564 = ~(n105 ^ n2920);
assign n21039 = n10192 | n20335;
assign n2366 = ~(n22276 ^ n1113);
assign n23292 = ~(n6442 ^ n8959);
assign n1474 = n2377 | n12246;
assign n23442 = n465 & n24985;
assign n14924 = n23880 | n15166;
assign n17908 = ~(n5990 | n7326);
assign n1761 = n5237 & n7443;
assign n3383 = ~n22294;
assign n26063 = n26307 | n23799;
assign n9359 = ~(n2664 ^ n11301);
assign n18476 = n12016 | n23118;
assign n7 = ~(n11943 ^ n3369);
assign n10482 = ~(n11203 ^ n16978);
assign n26885 = ~(n6025 ^ n24788);
assign n10084 = ~(n5043 | n24726);
assign n7042 = n8784 | n17350;
assign n17781 = n11495 & n17275;
assign n23067 = ~(n13957 ^ n23392);
assign n22126 = ~(n3209 ^ n26685);
assign n16257 = ~n5255;
assign n20061 = ~(n20843 ^ n9879);
assign n20018 = n16766 & n25174;
assign n1325 = ~n15532;
assign n15584 = n4318 | n5562;
assign n17252 = ~(n20429 | n26054);
assign n2726 = ~(n6222 | n990);
assign n25954 = ~n5260;
assign n8850 = ~(n6681 ^ n10538);
assign n5708 = ~n25813;
assign n6896 = n20127 ^ n23842;
assign n5791 = n17251 | n7473;
assign n23512 = ~n23900;
assign n2760 = ~(n25602 ^ n15884);
assign n17503 = n24302 | n5238;
assign n4104 = n18907 | n18951;
assign n9144 = n5203 | n8297;
assign n10976 = n19680 & n18341;
assign n9672 = ~(n16473 ^ n22597);
assign n5809 = n641 & n14460;
assign n21355 = ~(n20290 ^ n9934);
assign n10686 = ~(n10075 ^ n15959);
assign n24009 = ~(n20823 ^ n5764);
assign n2031 = n13508 & n7400;
assign n19685 = ~(n23807 ^ n26443);
assign n12773 = ~(n15633 ^ n8097);
assign n2287 = ~(n11926 | n2090);
assign n633 = n1248 & n18222;
assign n24206 = n2216 & n22873;
assign n17726 = ~(n18724 | n138);
assign n16541 = ~(n16715 ^ n13255);
assign n25353 = n16521 | n7139;
assign n5788 = ~(n21104 ^ n6315);
assign n10760 = ~n1446;
assign n4878 = ~n26901;
assign n2665 = ~(n1618 ^ n17926);
assign n5510 = n16167 & n173;
assign n10339 = n7237 | n15087;
assign n8188 = n12337 | n18388;
assign n21603 = ~(n16687 ^ n20906);
assign n6675 = n10301 | n7001;
assign n5720 = n26920 | n3913;
assign n16047 = n12147 & n9485;
assign n16254 = ~(n2906 | n14187);
assign n2274 = ~n20570;
assign n2596 = ~(n10577 ^ n24196);
assign n4629 = n21783 & n26863;
assign n22138 = ~(n537 ^ n21221);
assign n4599 = ~n830;
assign n8054 = n17268 & n20636;
assign n12822 = ~(n8182 | n4659);
assign n26666 = n10574 | n16266;
assign n8520 = ~n7856;
assign n20374 = n8676 | n4672;
assign n21378 = ~(n26223 ^ n10950);
assign n18566 = n14638 & n11071;
assign n7290 = n21867 & n19155;
assign n22518 = ~(n9827 | n25799);
assign n9412 = ~(n22071 | n18452);
assign n5689 = n27142 & n2410;
assign n23266 = n26217 | n3698;
assign n25843 = n26972 | n9668;
assign n13922 = ~(n10951 ^ n15254);
assign n19765 = n2780 & n24212;
assign n28 = ~(n12754 | n2167);
assign n644 = ~(n2053 ^ n1503);
assign n6628 = ~(n14312 ^ n14451);
assign n20800 = n22301 & n14183;
assign n21021 = ~(n6972 ^ n3161);
assign n17659 = n19962 | n23793;
assign n1593 = ~(n2776 ^ n4853);
assign n12425 = n26704 | n3358;
assign n2519 = ~(n13378 | n2071);
assign n15723 = ~(n19154 ^ n13095);
assign n5920 = n9818 | n7530;
assign n13791 = n17099 | n15124;
assign n3915 = ~(n1897 ^ n7464);
assign n4309 = ~(n3554 | n167);
assign n12774 = ~n19737;
assign n14273 = ~n14381;
assign n11167 = n21565 | n6911;
assign n11170 = n17862 & n6063;
assign n8960 = n20820 & n16058;
assign n15149 = ~(n20896 | n6435);
assign n24202 = ~(n22521 ^ n26913);
assign n5893 = n469 & n25686;
assign n3929 = n19945 & n26190;
assign n21256 = ~(n23084 ^ n3870);
assign n20450 = ~(n20038 ^ n20947);
assign n5401 = n14899 | n10408;
assign n25012 = n22801 & n21033;
assign n23689 = n20078 & n6676;
assign n21739 = ~n3217;
assign n2336 = ~n11184;
assign n7164 = n5393 & n7986;
assign n1376 = ~(n12513 ^ n8162);
assign n20135 = n11906 & n14611;
assign n20425 = ~(n1221 ^ n16597);
assign n4264 = n22606 | n21381;
assign n17177 = n18200 | n19127;
assign n10012 = ~(n4326 ^ n12593);
assign n19987 = n5267 | n14038;
assign n6321 = ~n10017;
assign n23966 = ~n21538;
assign n11360 = n6638 | n6301;
assign n8484 = ~(n17090 ^ n20986);
assign n22694 = n10152 | n1700;
assign n11589 = ~(n3195 ^ n12998);
assign n24576 = ~(n13528 ^ n17274);
assign n23572 = ~n25540;
assign n16270 = n11586 | n3214;
assign n1366 = n5882 | n17064;
assign n1921 = n14204 | n14783;
assign n13618 = n2312 & n25891;
assign n15022 = n10158 & n25004;
assign n10779 = ~(n3840 ^ n8925);
assign n5552 = ~(n26486 ^ n2858);
assign n4975 = ~(n11499 ^ n16458);
assign n12126 = ~(n17570 ^ n11239);
assign n2307 = n12269 | n10069;
assign n24070 = n23211 | n17758;
assign n3784 = n18477 & n2060;
assign n3592 = n12427 | n23523;
assign n10842 = n1888 | n6817;
assign n26496 = n25950 & n16706;
assign n22381 = ~(n24226 ^ n17412);
assign n18091 = n3882 | n4112;
assign n17566 = n15980 & n5083;
assign n6684 = ~(n20337 ^ n16925);
assign n10030 = n13633 | n2675;
assign n11692 = n15675 | n6956;
assign n3978 = ~(n15539 ^ n17664);
assign n19533 = ~(n23724 ^ n17854);
assign n11242 = ~(n8713 ^ n20417);
assign n6100 = n25632 | n24399;
assign n12181 = n9872 | n2801;
assign n5758 = ~(n1630 | n11121);
assign n11994 = n2831 & n16409;
assign n25496 = n14640 | n15904;
assign n24685 = n12506 & n9819;
assign n15946 = ~(n4964 ^ n8259);
assign n579 = ~(n14158 ^ n11381);
assign n6095 = ~(n25757 ^ n26201);
assign n17411 = ~(n13692 ^ n12617);
assign n24280 = ~n11221;
assign n24680 = n6259 & n24152;
assign n19744 = n10542 | n10014;
assign n6002 = n1108 | n22075;
assign n2237 = n12153 | n10148;
assign n16845 = ~n20189;
assign n9177 = ~(n15932 | n2385);
assign n16109 = n12394 & n25034;
assign n18436 = n14551 | n16677;
assign n10961 = ~(n16001 ^ n1049);
assign n21140 = ~(n26328 ^ n4746);
assign n18784 = n25664 & n3008;
assign n16388 = n997 | n21480;
assign n7765 = ~(n25165 ^ n20308);
assign n26240 = ~(n14340 ^ n20302);
assign n95 = n24738 & n17546;
assign n18617 = ~n3118;
assign n2436 = ~(n17764 ^ n25858);
assign n4001 = n12791 & n16018;
assign n24120 = n20170 | n1827;
assign n4138 = n16777 & n13694;
assign n17979 = ~n11566;
assign n25292 = n3575 | n12936;
assign n24309 = ~(n3568 ^ n6071);
assign n18903 = ~(n13319 ^ n15490);
assign n13108 = ~n27078;
assign n18568 = n20606 & n5807;
assign n20590 = ~(n6266 ^ n447);
assign n2395 = n8770 | n2286;
assign n16115 = n12473 | n12681;
assign n5306 = n12354 | n8581;
assign n15843 = n23445 | n13733;
assign n8329 = ~(n22793 ^ n15077);
assign n26774 = n13391 & n21626;
assign n3722 = ~(n337 ^ n16507);
assign n23174 = ~(n109 ^ n592);
assign n15438 = ~(n7234 ^ n21146);
assign n10913 = ~(n26894 ^ n16573);
assign n24305 = ~n21489;
assign n12191 = ~(n56 ^ n20506);
assign n25184 = ~n9817;
assign n15869 = ~(n17289 ^ n9858);
assign n19421 = n14621 | n26581;
assign n20158 = ~(n3981 | n23805);
assign n17245 = n16324 | n10075;
assign n14587 = ~(n9789 ^ n2764);
assign n16057 = ~(n1171 | n3407);
assign n20758 = n1618 | n9218;
assign n4329 = n20743 | n25019;
assign n7328 = n12991 & n24700;
assign n27206 = n23449 & n5382;
assign n19573 = n3464 | n4217;
assign n26812 = n6602 | n24465;
assign n26791 = n14049 & n11360;
assign n23135 = n25072 & n16458;
assign n13659 = ~(n6580 | n16608);
assign n26664 = n18493 & n15356;
assign n2483 = ~(n8303 ^ n1733);
assign n14103 = n4556 & n254;
assign n25258 = ~n15447;
assign n12013 = ~(n2163 ^ n10346);
assign n16619 = n24327 | n23185;
assign n2133 = ~(n2281 ^ n6814);
assign n10696 = n16009 & n12910;
assign n3544 = ~(n4748 ^ n11486);
assign n23729 = n9050 & n11789;
assign n16392 = ~(n636 ^ n24256);
assign n17167 = n2190 & n17786;
assign n25434 = n11011 & n10217;
assign n5190 = n17254 | n14313;
assign n4564 = ~(n14256 ^ n25751);
assign n12289 = ~(n26661 ^ n26808);
assign n25017 = ~(n24143 ^ n13183);
assign n25713 = ~n24281;
assign n6220 = n6598 & n749;
assign n12352 = ~(n402 ^ n24815);
assign n15034 = ~(n5302 | n3694);
assign n19824 = n26678 | n12532;
assign n16506 = ~(n717 ^ n10927);
assign n15455 = n1735 | n20618;
assign n13601 = n22031 | n20824;
assign n13658 = ~(n9096 ^ n25937);
assign n20074 = ~n429;
assign n8113 = ~(n6030 ^ n2350);
assign n24988 = ~(n10955 ^ n12630);
assign n19302 = n4099 | n13717;
assign n12401 = n2689 | n21965;
assign n20043 = ~n11377;
assign n9497 = n20102 & n14269;
assign n16359 = ~(n7694 ^ n7650);
assign n25115 = ~(n10845 ^ n21705);
assign n10706 = n8964 | n18126;
assign n3173 = ~(n22180 ^ n8855);
assign n13743 = ~(n10074 ^ n1410);
assign n7332 = n22893 & n8481;
assign n5145 = n618;
assign n13785 = n24635 | n24162;
assign n3077 = ~(n2666 ^ n932);
assign n10311 = ~(n24443 ^ n9422);
assign n21852 = n1422 & n24246;
assign n25136 = n24209 | n7671;
assign n20930 = n1229 & n25410;
assign n18921 = ~n1618;
assign n26450 = ~n15182;
assign n26404 = ~(n5172 | n26124);
assign n6221 = ~(n12702 | n12507);
assign n9024 = ~(n20259 ^ n22043);
assign n9300 = ~n25192;
assign n10487 = ~(n22695 | n1278);
assign n25278 = n17422 & n9330;
assign n25518 = ~(n10609 ^ n466);
assign n26989 = ~(n20077 ^ n3952);
assign n14750 = ~n18734;
assign n20958 = n14297 & n18911;
assign n13457 = n9649 | n19613;
assign n14350 = ~(n15921 ^ n7691);
assign n20891 = ~(n18812 ^ n1222);
assign n5183 = ~(n16605 ^ n5804);
assign n23 = n8222 | n3435;
assign n14511 = ~(n2918 ^ n8305);
assign n12735 = ~n11467;
assign n13575 = ~(n8930 | n22772);
assign n4128 = n17740 & n25951;
assign n17915 = n3411 | n24824;
assign n7076 = n22441 & n21776;
assign n13201 = n9251 & n24851;
assign n22314 = n24227 | n22561;
assign n1491 = n13279 & n695;
assign n5874 = ~(n3341 ^ n16858);
assign n20867 = n15246 & n26338;
assign n8064 = ~n1002;
assign n25900 = ~n23688;
assign n15448 = n6357 | n16752;
assign n22695 = ~(n18630 ^ n8581);
assign n24197 = n24084 & n23458;
assign n21146 = n11897 | n4480;
assign n11276 = ~(n11018 ^ n1525);
assign n10026 = ~(n1380 | n10843);
assign n9356 = ~(n25038 | n22626);
assign n5639 = n20281 & n12193;
assign n21336 = n7775 | n24734;
assign n19551 = ~(n9411 ^ n12546);
assign n532 = n3518 | n935;
assign n23455 = n16029 & n25674;
assign n8308 = ~n26964;
assign n6653 = ~(n15127 | n13562);
assign n7200 = n3702 & n15634;
assign n8105 = ~(n27114 | n17727);
assign n16008 = n10448 | n6471;
assign n20736 = n17501 | n25991;
assign n26864 = ~(n9595 | n27066);
assign n25854 = n5140 & n6705;
assign n7115 = n13174 & n14263;
assign n16059 = n26036 & n1505;
assign n15381 = n9991 | n24061;
assign n20605 = ~(n13489 | n20575);
assign n821 = ~n22626;
assign n14407 = n22844 & n1836;
assign n8615 = ~(n20169 ^ n4426);
assign n22293 = n11610 & n9965;
assign n3627 = n15109 | n10125;
assign n1899 = n10548 | n9333;
assign n21762 = ~(n19084 ^ n9598);
assign n6159 = n26682 & n17964;
assign n17461 = ~(n19926 ^ n2193);
assign n18869 = ~n2657;
assign n24081 = ~n5882;
assign n13358 = n10568 | n8309;
assign n3762 = n24991 | n4321;
assign n5765 = ~(n9079 ^ n24632);
assign n2832 = ~(n13231 ^ n9003);
assign n18388 = n12954 & n21087;
assign n11401 = ~(n11924 ^ n3993);
assign n8631 = n20327 | n9538;
assign n16084 = ~n24170;
assign n12716 = n19109 | n5114;
assign n11432 = n5547 & n6625;
assign n12619 = n6750 | n11670;
assign n10637 = ~(n12944 | n3448);
assign n19041 = n20446 & n24606;
assign n12669 = n12872 | n8318;
assign n18670 = n18600 | n13723;
assign n2725 = ~(n7691 | n15921);
assign n13843 = ~n5357;
assign n11076 = n1706 | n13032;
assign n25896 = ~(n23849 | n16274);
assign n4479 = ~n692;
assign n10322 = ~(n10920 ^ n18537);
assign n21899 = n14641 | n11031;
assign n26929 = ~(n4372 ^ n5350);
assign n19689 = n26961 | n1639;
assign n16473 = ~(n17419 ^ n21134);
assign n21577 = ~(n3992 ^ n11882);
assign n21452 = n11232 | n15518;
assign n2939 = ~n23990;
assign n15549 = n21509 | n25608;
assign n21410 = ~(n15732 | n16058);
assign n9749 = ~(n7177 ^ n13393);
assign n554 = ~(n24332 ^ n13504);
assign n18780 = ~(n1384 ^ n17715);
assign n3086 = ~n3581;
assign n9606 = n22445 | n18492;
assign n16973 = ~(n19941 ^ n10577);
assign n13136 = ~n23885;
assign n18647 = ~(n18907 ^ n18901);
assign n2156 = ~n7305;
assign n6183 = ~(n23812 ^ n22099);
assign n5932 = n3050 | n7684;
assign n26220 = ~(n24809 ^ n434);
assign n12167 = ~(n19888 | n24188);
assign n22905 = ~(n20478 | n1204);
assign n8822 = n19789 | n4978;
assign n26069 = ~(n21493 ^ n15746);
assign n19418 = n15687 & n22048;
assign n25675 = n20191 | n20799;
assign n7575 = ~(n3194 ^ n7147);
assign n17124 = n3116 & n24980;
assign n10643 = ~(n1079 ^ n15411);
assign n16760 = ~(n15182 | n20065);
assign n13555 = ~(n527 ^ n6369);
assign n20628 = ~n22226;
assign n683 = n3225 | n9619;
assign n8389 = ~n2878;
assign n4739 = ~(n25797 ^ n10611);
assign n26896 = ~(n5633 ^ n13580);
assign n25983 = ~(n16261 ^ n15158);
assign n2674 = n4028 | n25870;
assign n7589 = n3100 | n5551;
assign n7991 = n22069 | n6943;
assign n13337 = ~(n11393 | n2409);
assign n17439 = ~(n13023 | n9548);
assign n4460 = n10949 | n22095;
assign n20208 = ~(n2252 | n18495);
assign n7405 = n17368 | n3019;
assign n8467 = ~(n1222 | n22021);
assign n24637 = n26949 | n4641;
assign n11550 = ~n7917;
assign n11646 = ~n16446;
assign n3387 = ~(n13463 ^ n25475);
assign n3496 = ~n6847;
assign n20098 = n6206 & n232;
assign n558 = n3896 & n5502;
assign n2155 = ~n3051;
assign n12896 = n11776 | n19629;
assign n14499 = ~(n4361 ^ n25514);
assign n1880 = ~(n13863 | n23160);
assign n14631 = ~(n1340 | n18742);
assign n11474 = ~(n11944 ^ n15167);
assign n14285 = n456 | n8437;
assign n3431 = ~(n3019 ^ n15241);
assign n8491 = ~(n181 ^ n15766);
assign n15523 = n22360 | n24776;
assign n11582 = ~n19147;
assign n3447 = n26747 | n24666;
assign n15515 = ~(n16524 ^ n987);
assign n1623 = n13519 & n10226;
assign n812 = ~n16562;
assign n12972 = n6795 & n21439;
assign n25447 = n8948 | n16474;
assign n14280 = ~(n8933 ^ n11321);
assign n18060 = ~(n11711 | n17308);
assign n14752 = n14104 | n10079;
assign n21362 = ~n11815;
assign n2618 = ~n4435;
assign n13955 = n2870 & n14667;
assign n8043 = n8840 | n25853;
assign n216 = ~n21751;
assign n8488 = ~(n23760 ^ n14528);
assign n6886 = n24183 | n12605;
assign n14665 = ~(n6494 | n8832);
assign n2768 = ~n2161;
assign n21065 = n9428 & n7851;
assign n3671 = ~(n1232 ^ n19913);
assign n26571 = n18409 & n4940;
assign n17204 = ~(n20547 ^ n26511);
assign n10736 = n26077 & n16751;
assign n23916 = n21623 | n20597;
assign n5717 = n4531 | n21833;
assign n16585 = n9910 | n7319;
assign n7783 = ~(n19888 ^ n20734);
assign n6963 = ~(n7614 ^ n4954);
assign n26332 = ~(n26587 ^ n25406);
assign n13682 = n19149 | n13133;
assign n22942 = ~(n11559 | n6351);
assign n538 = ~(n9373 ^ n24510);
assign n596 = n10469 | n11499;
assign n4668 = n2671 & n26183;
assign n25608 = ~(n13432 ^ n23174);
assign n14759 = n8736 | n5914;
assign n6954 = n26534 & n21199;
assign n15091 = n9540 | n12825;
assign n20568 = n7319 | n23488;
assign n8470 = n4328 | n25298;
assign n3239 = ~n1946;
assign n20559 = n16893 | n19779;
assign n17044 = ~(n17929 | n21923);
assign n21219 = ~n15333;
assign n6434 = n20567 | n6849;
assign n10859 = ~(n16458 ^ n20907);
assign n26775 = ~(n25750 ^ n6875);
assign n10350 = ~(n11467 ^ n26015);
assign n26192 = ~(n11929 ^ n26744);
assign n1416 = ~(n2705 ^ n535);
assign n7581 = ~(n5706 | n24821);
assign n17622 = n4217 | n18055;
assign n12248 = n7410 & n8458;
assign n14214 = n26971 | n10613;
assign n279 = ~n15872;
assign n22380 = ~(n2893 ^ n7039);
assign n10759 = n14964 | n12803;
assign n8354 = ~(n9632 | n197);
assign n20280 = n5583 & n26631;
assign n24020 = ~(n6877 ^ n874);
assign n22416 = ~(n16106 ^ n15000);
assign n7556 = n15837 | n14844;
assign n25295 = n25113 | n9881;
assign n12862 = n12258 | n8964;
assign n14934 = n5388 | n19341;
assign n17448 = ~(n26295 | n16896);
assign n15866 = ~(n7059 | n6202);
assign n8291 = n5071 | n3200;
assign n16072 = ~(n21232 ^ n22744);
assign n10775 = ~(n24591 ^ n20767);
assign n26225 = ~(n15894 ^ n18899);
assign n20307 = n20396 & n11332;
assign n7303 = n1437 | n12488;
assign n13760 = ~n16626;
assign n20965 = ~(n20153 | n2964);
assign n19820 = n19298 | n1173;
assign n18115 = ~n7524;
assign n19928 = n14143 & n18605;
assign n7394 = ~n26831;
assign n18197 = n18245 & n22965;
assign n15551 = n11963 | n6203;
assign n18885 = n1289 | n7813;
assign n26453 = n15668 & n13482;
assign n3719 = ~n1792;
assign n4609 = n1137 & n12290;
assign n14453 = n21334 & n15273;
assign n3179 = ~(n1878 ^ n9335);
assign n5667 = n5004 | n27171;
assign n6707 = ~(n383 ^ n16940);
assign n25557 = n6929 | n22008;
assign n11317 = ~n16360;
assign n11627 = ~n25317;
assign n11442 = ~n15024;
assign n5109 = ~(n22404 | n7324);
assign n18600 = ~(n25426 | n1532);
assign n12717 = n5268 | n16095;
assign n22927 = n6617 | n18941;
assign n11364 = ~(n24237 | n19592);
assign n14043 = n6987 & n18501;
assign n6798 = ~(n14661 ^ n25322);
assign n2903 = ~n3582;
assign n21211 = n971 | n1926;
assign n23772 = n12567 & n12279;
assign n2991 = n22905 | n26587;
assign n489 = ~(n5958 | n22349);
assign n22003 = ~n18496;
assign n24843 = n14802 & n5281;
assign n14677 = ~n4886;
assign n19328 = ~n21860;
assign n24055 = n1039 | n11110;
assign n7102 = ~(n25167 ^ n1104);
assign n24706 = ~(n3837 ^ n24374);
assign n2258 = n18594 | n20907;
assign n12016 = ~(n22783 ^ n18578);
assign n22736 = ~n9881;
assign n17704 = ~(n3203 ^ n2935);
assign n3730 = ~(n22229 ^ n7583);
assign n14845 = ~(n9163 ^ n11508);
assign n26359 = ~(n10509 ^ n9244);
assign n6378 = n26496 | n25800;
assign n14137 = n3239 | n14649;
assign n4874 = ~n17575;
assign n15388 = n9549 | n7489;
assign n25161 = ~(n25381 | n14573);
assign n9048 = ~(n22170 | n16848);
assign n15491 = n23746 & n7269;
assign n20676 = n5255 & n6446;
assign n12135 = n22595 | n15421;
assign n20080 = ~(n6823 ^ n2491);
assign n17807 = n22887 | n4700;
assign n26230 = n5055 & n1318;
assign n18038 = n12400 | n2966;
assign n7399 = ~n19568;
assign n16106 = ~n18137;
assign n13397 = n6042 | n5051;
assign n19640 = ~(n10683 | n21134);
assign n14335 = n17260 & n5457;
assign n862 = ~(n852 | n11848);
assign n23609 = ~(n22379 | n9967);
assign n18557 = ~n18263;
assign n3193 = ~(n16793 ^ n7692);
assign n24513 = n22558 | n16548;
assign n22369 = n2498 | n947;
assign n8752 = n1669 | n16639;
assign n9360 = n4234 & n18650;
assign n20665 = n5005 & n2654;
assign n26990 = ~(n2230 | n13842);
assign n19967 = ~(n6352 | n13435);
assign n5827 = ~(n16822 ^ n14580);
assign n17163 = ~(n4874 ^ n11708);
assign n5647 = n15861 | n4887;
assign n2460 = ~n11106;
assign n26698 = ~(n8956 ^ n8089);
assign n19990 = n17714 & n453;
assign n25382 = n6750 & n11670;
assign n10242 = ~(n14688 ^ n9084);
assign n22054 = ~(n11989 | n14087);
assign n2928 = ~(n22363 | n27065);
assign n20240 = n4527 & n5797;
assign n10911 = ~n7727;
assign n26656 = ~(n15385 ^ n24568);
assign n26106 = n5842 | n3590;
assign n1737 = n16958 & n18270;
assign n23446 = n9884 & n20093;
assign n4340 = ~(n20440 ^ n21731);
assign n9416 = ~(n7949 | n16609);
assign n1261 = ~(n27042 ^ n25415);
assign n25199 = ~(n18434 | n20051);
assign n3225 = n21915 & n2509;
assign n14259 = n782 | n27042;
assign n26862 = n21829 | n22465;
assign n16701 = ~(n17824 ^ n5860);
assign n17466 = ~(n17797 ^ n27021);
assign n15891 = ~n12297;
assign n25908 = ~(n5852 ^ n16963);
assign n24312 = n1749 & n15514;
assign n16470 = ~n23366;
assign n13590 = ~n25119;
assign n21659 = n1682 & n3318;
assign n8387 = n12634 & n16920;
assign n22481 = ~(n8456 ^ n26744);
assign n3016 = ~(n13114 ^ n16641);
assign n26566 = ~(n24560 ^ n27139);
assign n20002 = ~(n9747 ^ n17089);
assign n8923 = n17630 | n18557;
assign n22788 = n2799 | n2271;
assign n6703 = ~(n19120 ^ n5129);
assign n19714 = ~(n2281 ^ n18755);
assign n2895 = ~(n1345 ^ n9106);
assign n12250 = ~(n17380 | n10962);
assign n14487 = n26032 & n23171;
assign n9920 = ~(n8100 | n2481);
assign n22362 = n18971 | n1446;
assign n17693 = ~(n15456 ^ n25365);
assign n14506 = ~(n23285 ^ n25704);
assign n23940 = ~(n20043 | n23264);
assign n19785 = ~(n3802 ^ n8778);
assign n9885 = n20625 & n21453;
assign n24581 = n19668 | n21223;
assign n15992 = ~(n2139 ^ n3710);
assign n672 = ~(n17411 ^ n22727);
assign n21080 = n16154 & n6101;
assign n8621 = n9310 | n4119;
assign n9333 = n19991 & n16651;
assign n1888 = ~(n11186 | n12821);
assign n14009 = ~(n10053 ^ n15539);
assign n4176 = ~(n19498 ^ n8246);
assign n10296 = ~n5091;
assign n26462 = n11113 & n24272;
assign n9055 = n18714 | n729;
assign n25291 = ~n9873;
assign n11768 = n4986 | n21840;
assign n26888 = ~(n15796 ^ n8528);
assign n10592 = ~(n2897 ^ n22358);
assign n1298 = n21551 & n27013;
assign n12596 = ~(n20042 | n24466);
assign n7959 = ~(n22702 ^ n14074);
assign n9099 = ~n1040;
assign n20488 = ~n20489;
assign n18977 = ~(n5923 ^ n17481);
assign n25836 = n27172 | n20075;
assign n16843 = ~n161;
assign n1607 = n26125 & n26321;
assign n16901 = ~(n3740 | n21784);
assign n12373 = ~n17274;
assign n6769 = n5183 & n4448;
assign n6597 = ~(n20630 | n25312);
assign n24816 = ~(n16609 ^ n12906);
assign n2790 = ~n21981;
assign n24182 = n12757 & n3507;
assign n907 = n573 & n19345;
assign n10270 = n11399 | n15483;
assign n9436 = n18506 | n5226;
assign n9218 = ~(n9876 ^ n3330);
assign n1746 = n26133 | n16570;
assign n12569 = ~(n5600 ^ n8022);
assign n7463 = n16366 | n18203;
assign n15814 = ~(n24392 ^ n21779);
assign n1310 = ~(n15722 | n1184);
assign n17323 = ~n18950;
assign n23862 = ~(n2803 ^ n9645);
assign n24588 = n18754 | n24499;
assign n26795 = ~(n10418 ^ n3593);
assign n9906 = n4934 | n14061;
assign n17950 = n24267 | n5897;
assign n2181 = n17665 & n1496;
assign n20327 = ~n20770;
assign n26320 = n631 | n12734;
assign n24112 = ~(n9100 ^ n26264);
assign n13377 = ~(n16707 | n20120);
assign n11806 = ~n5408;
assign n25109 = n15396 & n25578;
assign n11301 = ~(n21839 ^ n16544);
assign n621 = ~(n23235 | n8253);
assign n1436 = n15740 | n2243;
assign n10156 = ~n7657;
assign n22097 = n19608 | n2730;
assign n2860 = ~(n1393 ^ n8936);
assign n18542 = n12554 & n20711;
assign n25748 = ~(n22609 ^ n22829);
assign n4949 = n26762 | n21555;
assign n26140 = n8117 & n3280;
assign n3076 = ~(n13502 ^ n27069);
assign n17520 = n4386 & n10583;
assign n13825 = ~(n12658 ^ n8232);
assign n26922 = n4915 | n5052;
assign n11864 = n4627 & n13334;
assign n1648 = ~(n1970 ^ n22043);
assign n8444 = n13087 & n13433;
assign n14781 = ~(n26363 | n21596);
assign n8724 = ~(n15657 ^ n14124);
assign n26688 = ~n25751;
assign n5304 = ~n8001;
assign n3117 = ~(n8745 ^ n24278);
assign n4132 = ~n9655;
assign n17354 = ~(n11751 | n3245);
assign n23809 = n16476 & n15008;
assign n17706 = ~n19508;
assign n24487 = n8704 & n18665;
assign n26416 = n22703 | n10299;
assign n8654 = n1819 | n15521;
assign n13696 = ~n19804;
assign n18735 = ~n26239;
assign n18968 = n18823 | n20147;
assign n20786 = ~(n17141 ^ n3299);
assign n24784 = ~(n26664 ^ n17538);
assign n12283 = n12316 | n19168;
assign n4218 = ~(n21632 | n26510);
assign n2722 = ~(n461 | n22387);
assign n8061 = n8643 | n26769;
assign n22950 = n6215 | n4636;
assign n15848 = n22676 & n11588;
assign n11252 = ~(n25221 ^ n22507);
assign n18265 = ~(n11454 ^ n8458);
assign n14374 = ~(n19941 | n10577);
assign n21223 = n25388 & n16288;
assign n22583 = ~(n6034 ^ n21934);
assign n24740 = n21653 & n21617;
assign n12035 = n446 | n11045;
assign n17797 = n9738 | n6048;
assign n9034 = n15433 | n24875;
assign n6444 = ~(n8783 ^ n7979);
assign n18071 = ~(n20910 ^ n6155);
assign n21962 = n5960 & n17830;
assign n2804 = ~(n25339 ^ n12700);
assign n26491 = n9365 | n9095;
assign n1594 = ~n13503;
assign n19076 = ~n1690;
assign n9847 = ~(n2113 ^ n14345);
assign n8098 = ~(n19219 | n25251);
assign n23126 = ~n26512;
assign n21571 = n20812 | n3135;
assign n18267 = n9400 & n11154;
assign n19970 = ~(n5103 | n21565);
assign n16543 = ~(n15561 ^ n19708);
assign n5369 = n13713 | n20001;
assign n12132 = ~(n10146 | n11152);
assign n25824 = n1725 | n39;
assign n15120 = ~(n2111 ^ n16473);
assign n8502 = n20531 & n7645;
assign n11570 = n4277 | n13685;
assign n3504 = n1654 | n2425;
assign n8709 = n4722 & n14323;
assign n15493 = n13912 | n11980;
assign n3803 = ~(n685 ^ n25586);
assign n11191 = ~(n11209 | n5495);
assign n13111 = n13751 | n3128;
assign n22949 = n17293 | n12298;
assign n18671 = n18003 | n26058;
assign n3165 = n26361 & n18470;
assign n6994 = n727 | n15637;
assign n10044 = ~(n13494 | n23983);
assign n19351 = n26797 & n16221;
assign n25446 = ~(n9817 ^ n13189);
assign n3547 = ~n26522;
assign n5950 = ~(n2336 | n19366);
assign n8249 = ~(n23657 ^ n23035);
assign n17367 = ~(n19971 ^ n6685);
assign n8927 = n8858 | n23602;
assign n14057 = n6868 & n5087;
assign n16235 = n884 & n4617;
assign n18551 = n240 | n3113;
assign n15696 = ~n17056;
assign n15993 = n26828 | n16070;
assign n10566 = n20362 | n3548;
assign n9364 = ~(n13121 ^ n5049);
assign n14271 = ~(n16945 ^ n15758);
assign n25580 = n25025 | n8356;
assign n14724 = n4040 | n18006;
assign n5583 = n22723 | n7006;
assign n3379 = ~(n23249 ^ n5077);
assign n18870 = n16294 | n2944;
assign n23594 = ~(n23983 ^ n13494);
assign n15402 = n25452 | n507;
assign n20521 = ~(n22517 ^ n9226);
assign n23239 = ~(n6595 | n6199);
assign n19360 = ~(n17283 ^ n9429);
assign n14378 = ~n1596;
assign n2499 = ~(n19856 ^ n21687);
assign n21468 = n9670 | n2873;
assign n25560 = n20064 & n215;
assign n19589 = ~(n24781 ^ n21426);
assign n20467 = n25095 & n7078;
assign n16071 = ~(n19361 ^ n15918);
assign n26650 = ~n20863;
assign n16300 = n1748 & n11353;
assign n25653 = ~(n5159 ^ n16734);
assign n10599 = ~(n10500 ^ n12493);
assign n23322 = n7237 & n4873;
assign n2108 = n12546 | n14614;
assign n16037 = ~n21080;
assign n15286 = ~(n17184 ^ n24487);
assign n25943 = n25441 | n21620;
assign n23478 = ~(n18227 | n17397);
assign n14250 = n5818 | n7365;
assign n9069 = ~(n4093 ^ n752);
assign n3992 = n4962 & n23214;
assign n19682 = ~(n23706 ^ n5984);
assign n23705 = ~n25331;
assign n21967 = ~(n23708 ^ n26808);
assign n3831 = ~(n25194 | n6935);
assign n13986 = n14140 | n20009;
assign n20966 = ~(n19016 ^ n12039);
assign n9169 = n16780 & n8188;
assign n17041 = n15415 | n12119;
assign n17842 = ~(n22716 ^ n23912);
assign n20644 = n16508 & n6976;
assign n16289 = n20681 | n15754;
assign n23371 = ~(n13733 ^ n16072);
assign n2916 = ~(n6356 | n8418);
assign n25065 = n8766 & n10690;
assign n25255 = n23281 & n20557;
assign n15185 = ~n2382;
assign n3913 = n5543 & n22409;
assign n15840 = n5123 & n15482;
assign n1022 = n19477 | n2114;
assign n2093 = ~(n22417 ^ n3595);
assign n8616 = n23001 & n5293;
assign n26653 = n17092 | n10543;
assign n6968 = n17509 & n9307;
assign n574 = n12508 | n25942;
assign n19704 = ~(n20296 | n20862);
assign n6565 = ~(n5211 | n15910);
assign n18055 = ~n22683;
assign n9888 = ~(n8263 ^ n2904);
assign n10245 = ~(n3149 ^ n5400);
assign n24945 = ~n25186;
assign n4002 = n3024 & n4949;
assign n17185 = ~(n24890 | n10411);
assign n15417 = ~n21833;
assign n13427 = n13028 | n11579;
assign n3177 = n15685 | n5477;
assign n21438 = ~(n4213 ^ n19454);
assign n19191 = ~(n27144 ^ n23980);
assign n7321 = n23841 & n556;
assign n27192 = n18758 ^ n20259;
assign n15457 = n2825 & n15948;
assign n13226 = n5533 & n12080;
assign n15138 = ~n25523;
assign n21563 = ~(n7991 | n3133);
assign n24900 = ~(n4492 ^ n23002);
assign n3381 = n14595 & n18367;
assign n26049 = n8932 | n7795;
assign n8422 = ~(n1737 ^ n15607);
assign n12522 = n18137;
assign n3380 = ~n13884;
assign n2489 = n26491 ^ n7894;
assign n12236 = ~(n10844 ^ n8615);
assign n2036 = ~n3014;
assign n17944 = ~(n19303 | n15313);
assign n9710 = n16033 | n15852;
assign n22505 = n11153 & n14639;
assign n7517 = ~n2013;
assign n6922 = n3904 | n1653;
assign n6541 = ~(n23197 ^ n11276);
assign n22832 = ~(n11459 ^ n1837);
assign n13721 = n450 | n16028;
assign n18405 = ~(n5545 ^ n4953);
assign n18167 = n12245 | n19666;
assign n24617 = ~n3002;
assign n14258 = n3320 | n7879;
assign n5681 = n1751 | n12008;
assign n25327 = ~n21216;
assign n15980 = n8858 | n5886;
assign n14264 = n1745 & n4135;
assign n13361 = n1587 & n1685;
assign n6012 = ~(n26242 ^ n24147);
assign n7599 = n18062 & n8478;
assign n25427 = ~(n22972 ^ n8003);
assign n4201 = ~(n14582 ^ n8946);
assign n11496 = ~(n26967 ^ n12203);
assign n23803 = ~(n23999 ^ n13190);
assign n4391 = n8996 | n9955;
assign n4682 = ~(n5555 ^ n21649);
assign n26249 = n5778 & n4965;
assign n8787 = ~(n8931 | n1003);
assign n5660 = ~(n7536 ^ n19200);
assign n19936 = n8727 & n21075;
assign n24980 = n26064 & n9095;
assign n9204 = ~(n26490 ^ n11168);
assign n23631 = ~n12375;
assign n24654 = ~(n1347 ^ n7962);
assign n16625 = ~(n12971 | n17953);
assign n10055 = ~(n13330 ^ n12256);
assign n17231 = n26514 | n23176;
assign n20688 = n6770 & n1175;
assign n14833 = n3416 | n3167;
assign n9028 = n10125 | n8522;
assign n2660 = ~(n331 ^ n24616);
assign n4608 = n4296 & n11019;
assign n10640 = n842 | n1543;
assign n2690 = ~(n12541 ^ n26901);
assign n3249 = ~(n7455 | n17255);
assign n21800 = ~(n3580 ^ n24724);
assign n18828 = n642 | n4127;
assign n20491 = n5304 & n15437;
assign n1207 = ~(n21627 | n5415);
assign n12945 = ~(n3009 | n6011);
assign n14594 = n5518 | n3194;
assign n6622 = ~(n11953 | n13896);
assign n14579 = n23813 & n3912;
assign n18054 = ~n4576;
assign n7197 = n5657 & n14395;
assign n16984 = ~(n24774 ^ n3460);
assign n128 = ~(n13329 ^ n15884);
assign n1597 = ~(n4957 | n7421);
assign n22177 = ~(n12686 | n5642);
assign n19726 = n17184 & n24487;
assign n4989 = ~(n27142 ^ n9312);
assign n20052 = n2594 & n21991;
assign n1561 = n8597 | n8194;
assign n13002 = n14942 | n3497;
assign n21101 = ~(n20711 ^ n16396);
assign n4366 = ~(n17213 ^ n11302);
assign n14186 = n1458 & n21372;
assign n299 = ~(n19357 ^ n21649);
assign n14204 = ~n6232;
assign n16339 = ~(n8471 ^ n21402);
assign n3006 = ~n7044;
assign n17766 = n15453 | n26012;
assign n23797 = ~(n9222 | n25054);
assign n25578 = n1797 | n1837;
assign n26291 = n24825 & n8009;
assign n4090 = n12056 & n9892;
assign n16349 = ~n14790;
assign n12523 = n2202 | n19072;
assign n20206 = ~n5140;
assign n10741 = ~n10482;
assign n22895 = ~(n10440 ^ n385);
assign n9238 = ~(n16507 ^ n23250);
assign n20337 = n22054 | n5473;
assign n18624 = ~n25278;
assign n24956 = ~(n13104 ^ n26420);
assign n16686 = n18835 & n26416;
assign n12469 = ~(n12781 ^ n9989);
assign n25462 = ~(n24004 ^ n12900);
assign n12067 = ~(n10470 | n4062);
assign n9381 = n18730 | n17753;
assign n16528 = ~(n11143 | n10709);
assign n14571 = n25624 | n9653;
assign n22268 = n10024 | n26141;
assign n13311 = n23835 & n10947;
assign n25360 = ~(n23881 ^ n5615);
assign n20236 = n11785 | n19713;
assign n19147 = n9927 & n19635;
assign n18993 = ~(n2498 ^ n26013);
assign n22741 = ~(n11578 | n2261);
assign n21239 = ~(n15539 ^ n24278);
assign n9504 = ~(n20039 ^ n8694);
assign n9528 = n6508 | n21710;
assign n26150 = ~(n13846 ^ n17090);
assign n4995 = ~n23185;
assign n22207 = ~n18953;
assign n7470 = ~n13567;
assign n3099 = ~(n13899 | n15242);
assign n16800 = ~(n11273 | n23086);
assign n20545 = n1264 | n26635;
assign n3267 = n4803 | n20408;
assign n20097 = n19894 | n22517;
assign n12500 = ~(n9373 | n7677);
assign n22654 = ~(n16518 ^ n23649);
assign n20150 = ~n5929;
assign n27001 = ~(n9274 | n9814);
assign n15795 = ~n7656;
assign n251 = ~n26915;
assign n402 = ~n22375;
assign n4857 = n15427 & n10168;
assign n20024 = n12976 | n18007;
assign n2362 = n9343 & n15656;
assign n20365 = ~n12950;
assign n10791 = ~n13119;
assign n13365 = ~(n20089 | n21216);
assign n7796 = n23757 | n8195;
assign n155 = n3791 | n26876;
assign n7275 = n4380 | n2998;
assign n26788 = ~(n22619 | n22043);
assign n5745 = ~n12152;
assign n26614 = n17996 | n4597;
assign n12510 = n15756 | n6484;
assign n2256 = n131 | n23542;
assign n11342 = n2780 | n2000;
assign n15050 = ~(n4603 | n26536);
assign n4488 = n3185 | n21996;
assign n454 = ~(n1136 ^ n11667);
assign n15882 = n14739 | n15458;
assign n18057 = ~(n20376 | n6202);
assign n24014 = ~(n12699 | n8688);
assign n10500 = ~n25685;
assign n18831 = ~(n1216 ^ n18680);
assign n21660 = n6140 | n22352;
assign n15431 = n22336 | n15724;
assign n2149 = ~(n24517 ^ n26327);
assign n19628 = n14519 & n14208;
assign n20657 = n18912 | n18198;
assign n24284 = ~(n26580 ^ n18768);
assign n2751 = n20178 | n20508;
assign n24161 = ~(n5897 ^ n12886);
assign n2280 = ~(n25471 ^ n23842);
assign n23618 = n14502 | n18230;
assign n23909 = n21580 | n16229;
assign n17180 = ~(n210 ^ n15873);
assign n20157 = n17793 | n20114;
assign n16833 = ~(n22392 ^ n8920);
assign n12910 = ~(n1381 ^ n19070);
assign n22805 = n3318 | n1682;
assign n27126 = n14017 | n19750;
assign n26821 = n9155 & n19490;
assign n9247 = ~(n17275 ^ n13014);
assign n493 = n18046 & n1025;
assign n19049 = n21141 | n26165;
assign n920 = ~(n4360 | n17368);
assign n971 = n21623 & n6503;
assign n11229 = ~n14078;
assign n5628 = n15398 | n21752;
assign n9508 = ~(n15868 ^ n7988);
assign n3896 = n24623 | n26638;
assign n24883 = ~n15254;
assign n20196 = ~n14394;
assign n11555 = n6588 & n2988;
assign n17840 = n16992 & n451;
assign n9516 = n8700 | n24884;
assign n11988 = ~n3323;
assign n10623 = ~(n2342 | n20245);
assign n6760 = ~n14510;
assign n759 = ~(n11901 | n10201);
assign n19931 = n15200 | n8783;
assign n16480 = n15284 & n26819;
assign n13888 = ~(n14288 | n20039);
assign n23762 = n11898 | n25063;
assign n17615 = ~(n1281 | n13169);
assign n12581 = n22540 | n21041;
assign n12491 = n19918 & n7404;
assign n15031 = n359 | n22710;
assign n24912 = n16540 | n9288;
assign n26691 = ~n24786;
assign n8024 = ~n19649;
assign n9127 = n25144 | n5972;
assign n8360 = n21678 & n684;
assign n20731 = ~(n12308 ^ n9145);
assign n20523 = ~(n13567 ^ n1730);
assign n2610 = n19657 & n17772;
assign n13167 = n13378 & n10444;
assign n4161 = n8078 | n15143;
assign n22567 = n8344 | n13913;
assign n1213 = n6721 | n7857;
assign n16219 = ~(n10914 ^ n1481);
assign n24660 = ~n18585;
assign n26002 = n15168 | n26720;
assign n7979 = ~(n26660 ^ n25643);
assign n24846 = n19864 & n12581;
assign n2520 = ~(n15884 | n2412);
assign n2449 = n8382 | n7644;
assign n13188 = ~(n26691 | n8661);
assign n207 = n13460 & n10008;
assign n2504 = n21118 | n2331;
assign n11078 = ~(n7219 ^ n21834);
assign n17744 = ~n20724;
assign n10568 = ~n10411;
assign n22014 = n18737 | n6109;
assign n10472 = n13708 | n23085;
assign n16170 = n5922 | n6624;
assign n9299 = n14 | n16897;
assign n25747 = n6164 | n25942;
assign n15001 = ~(n11220 ^ n2944);
assign n7246 = n25896 | n21184;
assign n15272 = ~(n10586 | n15253);
assign n18731 = n5753 & n5632;
assign n24351 = ~n12917;
assign n9313 = ~(n7565 ^ n22390);
assign n9222 = ~(n24046 ^ n10929);
assign n10987 = ~(n5785 | n16353);
assign n5230 = ~(n2057 | n21930);
assign n26903 = ~(n25872 ^ n19618);
assign n8695 = ~n23727;
assign n2503 = n3069 & n11654;
assign n26984 = n11384 | n16812;
assign n5046 = ~(n14591 ^ n14986);
assign n27196 = n13873 | n24355;
assign n12039 = ~(n17351 ^ n16507);
assign n26159 = ~(n10921 ^ n21357);
assign n24283 = ~(n16709 ^ n12272);
assign n17486 = n7935 | n11552;
assign n23973 = n10430 & n18575;
assign n10940 = n25157 & n26281;
assign n14518 = ~(n1944 ^ n897);
assign n11633 = n10311 & n14713;
assign n7397 = n24588 & n5102;
assign n7300 = n1757 | n11970;
assign n23920 = ~n677;
assign n24495 = ~n14448;
assign n18983 = ~n26304;
assign n26728 = n26956 & n7021;
assign n13109 = ~n21900;
assign n4841 = n11756 | n21175;
assign n19392 = ~n638;
assign n24724 = ~(n13539 ^ n20532);
assign n1621 = ~(n1704 ^ n3356);
assign n12941 = ~(n17327 ^ n10360);
assign n16044 = n14655 | n79;
assign n22514 = ~(n8869 ^ n8381);
assign n21632 = ~n1112;
assign n10578 = n27139 & n24560;
assign n20299 = ~n8864;
assign n16791 = n3937 & n1243;
assign n24189 = n4147 & n20862;
assign n19281 = n4431 & n11925;
assign n5731 = ~(n166 ^ n4376);
assign n15650 = ~n5125;
assign n21432 = n2731 & n16210;
assign n10689 = ~n14453;
assign n21775 = n9053 | n23488;
assign n25606 = ~(n8106 ^ n13262);
assign n6600 = n22298 & n19751;
assign n13793 = ~(n21412 ^ n9821);
assign n3470 = n26997 & n19059;
assign n8303 = n12597 & n19099;
assign n11684 = n26275 & n16434;
assign n22580 = n7741 | n3123;
assign n25192 = ~(n12032 ^ n2083);
assign n1428 = ~(n11273 ^ n7949);
assign n9031 = n5225 | n21652;
assign n19222 = ~(n25352 ^ n26823);
assign n79 = ~n22970;
assign n12575 = ~(n26673 | n15539);
assign n5490 = n18391 | n16421;
assign n26811 = n572 | n21076;
assign n16732 = n15608 | n24423;
assign n13926 = ~(n11954 ^ n9593);
assign n26936 = n26990 | n25012;
assign n15116 = n11707 | n15214;
assign n23606 = n4696 & n8515;
assign n6705 = ~n8079;
assign n16443 = ~n6154;
assign n21986 = ~(n11932 ^ n20720);
assign n22279 = n18914 | n4629;
assign n19356 = ~(n15500 ^ n16784);
assign n22497 = ~(n15007 ^ n14387);
assign n7685 = ~n23180;
assign n5350 = ~(n14265 ^ n2938);
assign n9955 = n3821 & n24781;
assign n21040 = n237 & n13688;
assign n19513 = ~(n4868 | n25345);
assign n2384 = n2146 & n212;
assign n8793 = n10357 | n20621;
assign n3596 = ~(n14130 ^ n23463);
assign n1338 = n2522 | n15764;
assign n25625 = n6764 | n5328;
assign n14427 = n25400 | n25975;
assign n24580 = ~n25739;
assign n597 = ~(n16513 ^ n6999);
assign n26603 = ~(n9983 | n16173);
assign n5030 = ~n9559;
assign n24126 = n5075 & n682;
assign n25753 = n23818 | n9360;
assign n25488 = n16943 | n22264;
assign n17843 = ~(n13944 ^ n7759);
assign n11792 = ~(n11789 ^ n26107);
assign n8081 = n2341 | n24620;
assign n3972 = ~(n9402 | n2439);
assign n14880 = ~(n3578 ^ n18181);
assign n21092 = ~(n19639 | n11207);
assign n713 = ~n17235;
assign n2072 = ~(n24921 ^ n6714);
assign n5134 = n348 | n6679;
assign n7188 = n15545 & n16461;
assign n21621 = ~(n27037 | n17605);
assign n24399 = ~(n15046 ^ n1156);
assign n9963 = ~(n10306 ^ n3710);
assign n13823 = n3136 | n5752;
assign n23979 = ~(n15023 | n10446);
assign n1691 = ~(n12453 ^ n14762);
assign n5137 = n1426 | n10105;
assign n21451 = ~(n24544 ^ n657);
assign n24881 = ~(n12751 ^ n7798);
assign n3664 = ~(n19025 | n16482);
assign n7924 = ~(n21791 ^ n22262);
assign n15962 = n8740 | n19638;
assign n18686 = ~(n15405 ^ n2223);
assign n3776 = ~n22399;
assign n13175 = n12642 | n5508;
assign n19760 = ~(n6492 | n9523);
assign n20760 = n16091 | n3012;
assign n19791 = ~(n1584 ^ n2743);
assign n24333 = n1658 | n384;
assign n22992 = n5854 & n24066;
assign n9659 = ~(n27149 | n15414);
assign n16469 = ~(n15182 ^ n17351);
assign n13189 = ~(n4563 ^ n23295);
assign n20518 = ~(n9934 | n2272);
assign n13722 = ~(n4827 ^ n15316);
assign n15505 = n23457 | n11006;
assign n6623 = ~(n24919 | n25261);
assign n23282 = n3942 | n26328;
assign n23785 = n13635 | n13067;
assign n25801 = n1326 | n2854;
assign n587 = n7801 & n8548;
assign n6878 = n2628 | n22554;
assign n17057 = n26895 | n2387;
assign n1363 = n20365 | n22571;
assign n7707 = n12289 | n552;
assign n22117 = n21609 | n20763;
assign n20947 = ~(n22363 ^ n27065);
assign n16785 = n19659 & n6646;
assign n1419 = ~(n2842 ^ n23678);
assign n14667 = n26314 | n14443;
assign n14433 = n22413 | n23302;
assign n23349 = n23129 | n9577;
assign n6316 = n9794 & n8503;
assign n17165 = n23164 | n16771;
assign n10056 = n3324 | n8612;
assign n16774 = ~n26077;
assign n7944 = ~(n12040 ^ n21085);
assign n3817 = ~(n17423 | n8614);
assign n12828 = n2805 | n1524;
assign n20874 = n5696 & n7871;
assign n23952 = n21054 & n21808;
assign n7168 = ~n18745;
assign n5497 = n8347 | n9019;
assign n847 = ~(n5421 ^ n13021);
assign n9495 = n12973 | n15867;
assign n24448 = n13084 & n14212;
assign n3754 = n25305 & n16749;
assign n17662 = ~(n24818 ^ n3981);
assign n26016 = ~(n16778 ^ n18691);
assign n25008 = ~(n13577 ^ n11374);
assign n11119 = ~(n15696 ^ n2109);
assign n13853 = ~(n25727 ^ n4253);
assign n19537 = n3114 | n20347;
assign n14548 = ~(n1682 ^ n18157);
assign n361 = ~(n13490 | n15769);
assign n24328 = n1163 | n5668;
assign n5806 = ~n5787;
assign n15414 = n952 & n3647;
assign n1110 = ~(n2858 | n977);
assign n4158 = ~(n3861 ^ n2809);
assign n15825 = n25021 | n20137;
assign n653 = n20964 | n18345;
assign n26743 = ~(n4435 ^ n274);
assign n9952 = ~(n11830 ^ n13775);
assign n24931 = n14260 | n4268;
assign n12286 = n19100 & n12074;
assign n12317 = ~n3186;
assign n24008 = ~n8255;
assign n17096 = n27183 | n23939;
assign n18992 = ~(n11901 | n4938);
assign n25542 = n21117 | n1112;
assign n14871 = n5654 & n17482;
assign n4645 = ~(n16949 | n3919);
assign n22216 = ~(n23285 | n25704);
assign n18838 = ~n15058;
assign n14324 = ~(n19128 ^ n7440);
assign n26897 = ~(n12962 | n1960);
assign n6860 = n8101 | n21912;
assign n12632 = ~(n196 ^ n9460);
assign n25282 = ~n3279;
assign n24548 = n24603 | n13022;
assign n7843 = n24059 | n2741;
assign n26734 = n1635 | n1592;
assign n22689 = n11847 | n1247;
assign n25112 = n21593 & n7787;
assign n19717 = ~(n24072 | n14312);
assign n12889 = ~n4956;
assign n22140 = n2251 | n20549;
assign n1364 = ~n17815;
assign n944 = ~n17940;
assign n5221 = ~(n16590 | n26090);
assign n1196 = ~(n8725 ^ n4077);
assign n5165 = ~n24298;
assign n17838 = ~(n16840 | n8302);
assign n21943 = ~(n2157 ^ n26136);
assign n6274 = n19531 | n21322;
assign n13407 = ~(n15330 ^ n16595);
assign n4144 = n15636 & n18255;
assign n12887 = ~n24677;
assign n8748 = n15100 & n11793;
assign n2105 = ~(n5632 ^ n16895);
assign n16258 = ~(n10749 ^ n7066);
assign n3041 = ~(n18504 ^ n11630);
assign n22160 = ~(n24700 ^ n26180);
assign n23991 = n13571 | n26028;
assign n10282 = n24150 | n7919;
assign n3484 = ~(n21424 ^ n14767);
assign n20316 = ~n11497;
assign n1806 = ~(n16166 | n10407);
assign n2977 = n18673 | n20953;
assign n7061 = ~(n12681 ^ n577);
assign n14503 = n15504 | n5441;
assign n4310 = n286 ^ n6294;
assign n11908 = n10935 & n1711;
assign n19782 = n1198 | n8593;
assign n5633 = ~(n21600 ^ n14261);
assign n19178 = n18444 | n17028;
assign n6674 = n2031 | n21369;
assign n24021 = ~n27082;
assign n4948 = n24605 | n10524;
assign n17067 = ~n20528;
assign n9761 = ~(n25093 ^ n10315);
assign n23843 = ~n15723;
assign n1866 = ~(n24327 | n663);
assign n4101 = n23281 | n20557;
assign n7455 = ~n22895;
assign n10780 = ~(n6305 ^ n1691);
assign n23012 = ~n10082;
assign n7072 = ~(n6181 ^ n4590);
assign n6038 = ~(n25623 ^ n145);
assign n2901 = ~(n8087 ^ n2041);
assign n24663 = n12932 & n22930;
assign n24062 = n3915 & n17411;
assign n23790 = ~(n1350 ^ n13368);
assign n21486 = ~(n14226 | n1255);
assign n23660 = ~(n4642 ^ n17658);
assign n14381 = ~(n10722 ^ n3893);
assign n16353 = ~(n9911 ^ n4120);
assign n8594 = ~(n16016 ^ n21797);
assign n4612 = n2180 | n20848;
assign n22430 = n27089 | n12657;
assign n21038 = ~n13714;
assign n1652 = ~n12646;
assign n14294 = ~(n3021 ^ n973);
assign n16483 = ~n7802;
assign n23922 = n25663 | n647;
assign n12268 = n21632 | n7751;
assign n19462 = ~(n24044 | n12657);
assign n27057 = ~n7991;
assign n5329 = ~(n18303 ^ n18558);
assign n18984 = n17717 | n21953;
assign n4122 = n3984 | n18251;
assign n13591 = ~n268;
assign n10025 = ~n21140;
assign n8895 = ~n8455;
assign n11960 = ~(n3349 ^ n6397);
assign n14854 = n10365 | n2951;
assign n21018 = n11434 & n5322;
assign n15922 = ~(n22852 ^ n5236);
assign n22000 = ~(n2421 | n5337);
assign n18491 = n23426 | n25885;
assign n6943 = ~n16212;
assign n24406 = n6708 & n16416;
assign n15751 = n24804 | n7809;
assign n11499 = ~n5599;
assign n18691 = ~(n13907 ^ n2858);
assign n16755 = ~n1222;
assign n13772 = n1490 | n9253;
assign n6270 = ~n19836;
assign n21901 = n12392 & n20648;
assign n22937 = n20389 | n2864;
assign n7795 = n7103 & n17849;
assign n5634 = ~(n467 ^ n27108);
assign n12073 = n306 | n26307;
assign n17447 = ~n15972;
assign n10870 = n12306 | n26545;
assign n503 = n6753 | n23529;
assign n652 = ~(n5 ^ n8255);
assign n2339 = ~(n17098 | n14273);
assign n19581 = n14088 & n23826;
assign n12890 = ~(n26528 ^ n12888);
assign n7039 = ~(n16465 ^ n5449);
assign n22491 = ~n23650;
assign n24607 = ~(n18537 | n24617);
assign n272 = n17822 & n10607;
assign n20502 = n12702 & n348;
assign n18104 = n10606 | n24743;
assign n18955 = n9233 | n15108;
assign n18207 = n8782 & n18643;
assign n3490 = ~(n25270 | n1339);
assign n7459 = n15422 | n2908;
assign n24331 = n21129 & n15159;
assign n8700 = ~(n4518 | n12990);
assign n9559 = ~(n9437 ^ n17720);
assign n26333 = ~(n14601 | n25297);
assign n443 = n14569 | n12004;
assign n15358 = ~(n4181 | n2633);
assign n17379 = ~n8402;
assign n6345 = ~(n16038 ^ n23901);
assign n7617 = n2175 & n4484;
assign n20133 = ~n4119;
assign n16260 = n10401 | n17437;
assign n14647 = ~n24679;
assign n21769 = n16813 | n11894;
assign n12451 = ~(n18649 | n3984);
assign n6515 = ~n26017;
assign n4788 = n22612 | n12360;
assign n486 = n22315 | n23877;
assign n8994 = ~(n14791 ^ n9557);
assign n7374 = ~n3213;
assign n6437 = ~(n2905 ^ n6807);
assign n25782 = n16884 | n5250;
assign n4422 = n20398 & n1517;
assign n24614 = n21824 & n11877;
assign n12977 = n4977 | n11320;
assign n17316 = ~n10124;
assign n8591 = n13302 & n11202;
assign n26121 = n15269 | n19377;
assign n7282 = n17020 & n17034;
assign n26998 = n16203 | n17816;
assign n22628 = n12233 & n25392;
assign n3797 = n10622 | n24166;
assign n13850 = ~(n23761 ^ n19040);
assign n1973 = ~n26545;
assign n19838 = ~(n16351 | n13549);
assign n25688 = ~(n22836 ^ n15636);
assign n25737 = ~n10667;
assign n9787 = ~(n17978 ^ n10650);
assign n4697 = ~(n12386 | n2696);
assign n20397 = ~(n20044 ^ n7421);
assign n4149 = ~n22492;
assign n10519 = n8492 | n20528;
assign n26299 = ~n15970;
assign n10935 = n10832 | n8352;
assign n24779 = n2277 & n26037;
assign n9046 = ~(n11820 ^ n11277);
assign n26529 = ~(n23689 ^ n24198);
assign n10037 = ~n1293;
assign n15639 = ~n4467;
assign n11246 = ~(n24799 ^ n22492);
assign n23301 = n24962 | n5644;
assign n6304 = ~(n13677 | n26752);
assign n21003 = n1781 | n26045;
assign n20503 = n26000 | n12137;
assign n16034 = ~(n23122 ^ n12587);
assign n15462 = ~(n7086 ^ n20462);
assign n9866 = n8198 | n11150;
assign n6712 = n218 | n4605;
assign n19723 = n16799 | n25148;
assign n10081 = n4993 & n9994;
assign n17965 = n7254 | n9599;
assign n12606 = ~(n9105 ^ n4449);
assign n7398 = n3029 | n16348;
assign n6477 = ~(n19581 ^ n12848);
assign n14145 = ~n1689;
assign n25716 = ~(n26162 | n21386);
assign n11244 = ~(n7168 | n17547);
assign n18656 = n3137 & n2838;
assign n6166 = n5460 | n7668;
assign n12924 = ~n3843;
assign n21893 = ~(n23862 ^ n4854);
assign n22513 = ~(n18008 ^ n14230);
assign n3822 = n16359 | n13257;
assign n24234 = n405 | n26109;
assign n18932 = n6910 | n25563;
assign n20384 = ~(n24422 ^ n4319);
assign n24019 = ~(n21272 | n3203);
assign n22405 = n21227 & n19813;
assign n25573 = n23288 | n3055;
assign n18437 = ~(n23780 ^ n25033);
assign n16957 = ~(n7652 ^ n16559);
assign n14625 = ~n16608;
assign n5558 = n22310 & n19209;
assign n17637 = ~(n3015 ^ n21272);
assign n5338 = ~n13941;
assign n21004 = ~n22413;
assign n7869 = n21282 & n19246;
assign n14092 = ~(n9942 ^ n2210);
assign n13488 = ~(n7693 | n3909);
assign n17229 = ~(n5886 ^ n1839);
assign n11101 = ~(n13211 ^ n16809);
assign n17267 = n20527 | n2525;
assign n15790 = ~(n19429 | n23519);
assign n27021 = ~(n18283 ^ n6924);
assign n11958 = ~n12081;
assign n20560 = n26660 & n17826;
assign n16372 = n2967 | n18907;
assign n18708 = ~(n13213 ^ n16011);
assign n18905 = ~(n12502 ^ n4320);
assign n20271 = ~n17166;
assign n9900 = ~(n835 ^ n20826);
assign n20398 = n24305 | n8823;
assign n26164 = n17911 | n17674;
assign n15649 = ~(n20470 ^ n4590);
assign n20864 = ~(n16928 | n19940);
assign n9733 = ~n22795;
assign n8084 = ~(n26950 ^ n1945);
assign n10620 = ~n3319;
assign n7633 = n13298 | n25231;
assign n3895 = ~(n966 ^ n12446);
assign n27167 = ~(n25139 | n15636);
assign n10416 = ~(n25724 | n24503);
assign n11027 = n26107 & n21636;
assign n12081 = ~(n9109 ^ n21354);
assign n8157 = n24005 | n15528;
assign n8737 = n26660 | n26810;
assign n26930 = ~(n14890 ^ n16375);
assign n10737 = ~(n22290 ^ n12562);
assign n26409 = n8571 & n10872;
assign n16835 = n4917 | n13841;
assign n25554 = n13750 & n20024;
assign n2279 = ~(n2123 ^ n1996);
assign n14027 = n12815 | n8441;
assign n9341 = ~(n19514 ^ n19228);
assign n13711 = n3460 & n16667;
assign n3257 = ~n14163;
assign n23503 = ~(n7010 ^ n13851);
assign n22751 = n9514 & n17204;
assign n8587 = ~(n26992 ^ n7437);
assign n22457 = ~(n9200 ^ n18758);
assign n6376 = n18850 | n15153;
assign n17195 = ~n4583;
assign n297 = n4592 & n24502;
assign n5744 = ~(n11579 ^ n8067);
assign n9443 = n22363 | n17291;
assign n11955 = ~(n24135 ^ n20291);
assign n15130 = n11997 | n18798;
assign n20732 = ~(n16573 | n26894);
assign n20508 = ~n14417;
assign n12678 = n6306 | n25396;
assign n27190 = ~(n23559 | n12048);
assign n7501 = ~(n18451 | n13081);
assign n20386 = n20226 & n21136;
assign n3396 = ~(n3668 | n2246);
assign n10950 = ~(n2570 ^ n10250);
assign n22576 = ~(n15332 | n8753);
assign n26880 = n1514 & n6922;
assign n12680 = ~(n4400 ^ n17739);
assign n22162 = ~(n2884 ^ n20455);
assign n26045 = n3991 & n13431;
assign n23467 = ~(n20645 ^ n21180);
assign n22239 = n21073 | n502;
assign n22772 = ~(n21564 ^ n11412);
assign n12177 = ~(n4970 ^ n2454);
assign n23989 = ~(n22602 | n12257);
assign n11900 = ~(n15204 ^ n12956);
assign n20940 = n2930 | n12885;
assign n23857 = ~(n17664 ^ n5115);
assign n4389 = n26833 | n22875;
assign n22288 = ~(n12068 | n18535);
assign n14299 = n26347 & n12393;
assign n7646 = n17245 & n8506;
assign n15447 = ~(n4474 ^ n23215);
assign n20509 = ~n26174;
assign n8437 = ~(n373 ^ n737);
assign n23211 = ~n7876;
assign n23273 = ~n18924;
assign n4408 = ~(n2432 ^ n11137);
assign n4821 = n8737 & n7699;
assign n796 = ~(n24612 | n9770);
assign n24741 = n16008 & n24287;
assign n15234 = ~(n26629 ^ n18690);
assign n25575 = ~(n23357 ^ n26958);
assign n14853 = n7198 | n16439;
assign n14979 = ~n25797;
assign n21699 = n25926 | n20385;
assign n18456 = n17458 | n17265;
assign n10694 = ~(n17309 ^ n2096);
assign n26014 = n7670 | n8227;
assign n14201 = ~(n13960 ^ n10405);
assign n21780 = ~n12744;
assign n19214 = ~(n22194 | n6104);
assign n18126 = ~n14504;
assign n6507 = n23365 | n12770;
assign n8392 = n13092 | n19237;
assign n18699 = n10810 | n17575;
assign n26615 = n23514 & n15132;
assign n20652 = ~(n15109 | n8677);
assign n14838 = n19788 & n1468;
assign n21251 = n3914 | n1717;
assign n4822 = ~(n4914 ^ n19338);
assign n8365 = n14213 & n14847;
assign n11552 = ~n24080;
assign n17121 = ~(n17973 | n26009);
assign n6066 = n15905 | n27118;
assign n18358 = n1790 | n20660;
assign n12375 = n22573 & n8400;
assign n8112 = ~(n20955 | n24322);
assign n17261 = ~n3786;
assign n13965 = ~(n17415 ^ n7593);
assign n24894 = n3180 | n10249;
assign n18748 = n7825 | n8511;
assign n23764 = n11659 | n4928;
assign n16992 = n7769 | n15245;
assign n24118 = n5167 & n4170;
assign n21293 = ~(n23136 ^ n15779);
assign n23944 = n8642 | n12172;
assign n22007 = ~(n16830 | n25688);
assign n5855 = ~n25069;
assign n17313 = n9434 & n5563;
assign n26842 = n21988 | n8380;
assign n10095 = ~(n18262 ^ n22588);
assign n16935 = n14145 | n20036;
assign n5970 = ~n17085;
assign n14955 = ~n3056;
assign n23338 = n2212 | n21393;
assign n10905 = ~(n4999 ^ n27017);
assign n12961 = ~n16846;
assign n1617 = n17789 & n1731;
assign n12228 = ~(n24986 ^ n9);
assign n9303 = ~n781;
assign n2110 = ~n7476;
assign n4211 = n9081 | n19597;
assign n24011 = n13771 & n14911;
assign n7257 = ~(n3591 ^ n647);
assign n26251 = ~(n16033 ^ n15946);
assign n9737 = ~(n24787 ^ n906);
assign n9420 = ~(n4856 ^ n23323);
assign n9636 = ~(n3049 ^ n25094);
assign n2233 = ~(n22195 ^ n1865);
assign n8651 = n10092 | n11477;
assign n2521 = n1740 & n4997;
assign n10068 = n13038 | n11306;
assign n19 = ~n8745;
assign n12241 = n9964 | n4880;
assign n7184 = n2894 & n22783;
assign n14308 = n6664 | n4114;
assign n18298 = ~n16263;
assign n24928 = ~(n3389 ^ n4148);
assign n17632 = ~(n26107 | n4376);
assign n22534 = n10471 & n8600;
assign n14355 = ~(n788 ^ n21780);
assign n1861 = n18704 | n5317;
assign n4375 = ~(n23734 ^ n25927);
assign n23685 = ~(n1894 ^ n3921);
assign n26466 = n19776 & n18932;
assign n5685 = ~n22340;
assign n26286 = n11601 & n4546;
assign n13019 = n13325 & n7176;
assign n26859 = n6206 | n17409;
assign n26537 = n17230 | n10792;
assign n1116 = ~(n10023 | n22715);
assign n2099 = ~(n21757 ^ n21239);
assign n7054 = n22750 | n13728;
assign n3999 = n6212 | n23375;
assign n20984 = n15259 | n7833;
assign n12439 = n8631 & n607;
assign n15246 = n21117 | n22332;
assign n8707 = n18737 & n15268;
assign n21848 = n17400 & n21196;
assign n25531 = n6812 | n14866;
assign n1727 = n319 & n23032;
assign n17112 = ~(n11098 ^ n15175);
assign n144 = ~n23529;
assign n16853 = ~(n27015 | n22993);
assign n9334 = n18633 | n24647;
assign n16132 = n6950 | n23275;
assign n15153 = ~(n4157 ^ n16503);
assign n1015 = n25524 | n2562;
assign n20566 = ~(n7060 | n19976);
assign n24209 = n4508 | n13843;
assign n17008 = n22348 & n7482;
assign n20998 = ~n11056;
assign n17282 = n14642 | n23417;
assign n2802 = ~(n23493 ^ n1222);
assign n17793 = n12083 & n7989;
assign n2052 = n19553 & n24195;
assign n8742 = n6635 & n121;
assign n24737 = n1404 | n18262;
assign n11763 = n12767 | n1658;
assign n17545 = n4621 & n10748;
assign n4920 = n21527 & n20509;
assign n21024 = ~(n10454 ^ n102);
assign n13830 = ~(n24170 ^ n18537);
assign n2414 = n17069 | n19446;
assign n15495 = ~(n21434 ^ n2715);
assign n13020 = n4510 | n24741;
assign n22482 = ~(n23609 | n14335);
assign n26114 = n7480 | n8122;
assign n2394 = n14100 | n2284;
assign n14325 = n10051 | n11047;
assign n19989 = ~n16097;
assign n7294 = n15 | n26706;
assign n18526 = ~(n1028 ^ n1994);
assign n7560 = ~(n12930 | n22084);
assign n16036 = n8886 | n2898;
assign n12123 = ~n19893;
assign n19491 = n13042 & n12721;
assign n9502 = n75;
assign n14905 = ~(n7561 ^ n3443);
assign n5933 = n4957 & n22688;
assign n25386 = n3419 | n25554;
assign n22095 = ~n17690;
assign n17194 = n24522 & n4450;
assign n17728 = ~n12964;
assign n14005 = ~(n4307 ^ n10964);
assign n3453 = n17789 | n1731;
assign n1174 = n15799 | n12496;
assign n23707 = ~n8497;
assign n21955 = n17535 & n6552;
assign n17502 = ~n19477;
assign n14980 = ~n24169;
assign n12060 = ~(n11118 ^ n4199);
assign n11779 = ~(n13960 ^ n12990);
assign n9016 = n17708 | n2769;
assign n17440 = ~(n24584 | n13802);
assign n10924 = ~(n18703 ^ n22530);
assign n5789 = ~(n9307 ^ n21963);
assign n24219 = ~(n22729 ^ n18744);
assign n10040 = n4856 | n14455;
assign n6425 = n2613 | n20851;
assign n8901 = ~(n8518 ^ n17677);
assign n4423 = n6385 | n8844;
assign n2292 = n9298 | n17339;
assign n20646 = n6801 & n16395;
assign n1760 = ~(n20980 ^ n4516);
assign n25118 = n8899 & n20873;
assign n4556 = n3014 | n23630;
assign n5622 = n23592 | n23463;
assign n13394 = n22658 | n4006;
assign n12826 = ~(n14365 ^ n11993);
assign n20012 = ~(n26822 ^ n22404);
assign n12672 = n24434 & n20585;
assign n12164 = n333 | n4798;
assign n9623 = n22206 | n9559;
assign n24110 = n17348 | n15335;
assign n730 = ~(n12385 | n4749);
assign n19973 = n24209 & n7671;
assign n18329 = n3409 | n2310;
assign n15568 = n26390 & n1489;
assign n10146 = ~n25643;
assign n17088 = ~n23660;
assign n25910 = n24850 | n16083;
assign n10533 = ~n18434;
assign n22368 = n6905 | n11587;
assign n23278 = n767 | n8806;
assign n9265 = n18966 | n19796;
assign n736 = ~(n23030 | n20829);
assign n24063 = n26393 & n13267;
assign n23029 = n21749 & n11676;
assign n1356 = ~(n19033 | n17037);
assign n2805 = ~(n1406 | n1978);
assign n388 = n16014 & n262;
assign n24138 = ~(n6847 ^ n12070);
assign n6508 = ~n14388;
assign n3736 = n8553 & n15502;
assign n4991 = n3169 | n8729;
assign n20401 = n18883 & n25146;
assign n4216 = n15189 | n24320;
assign n23774 = n9598 | n21570;
assign n7619 = ~n6185;
assign n18424 = n9099 & n19067;
assign n15797 = n22374 & n5118;
assign n10307 = ~(n21540 | n18768);
assign n7818 = ~n5077;
assign n24090 = ~n8009;
assign n2383 = ~(n25453 ^ n18743);
assign n8547 = n6847 & n2051;
assign n21026 = n13711 | n26586;
assign n9061 = n5907 | n24407;
assign n8489 = ~(n25410 ^ n21000);
assign n4923 = ~(n19628 ^ n2999);
assign n18648 = n17616 & n21391;
assign n8595 = n11961 & n22863;
assign n17362 = ~(n21287 ^ n25331);
assign n17748 = n10430 | n18575;
assign n18902 = ~(n4695 | n17371);
assign n16647 = n25274 & n3888;
assign n2150 = ~(n17989 ^ n20706);
assign n10348 = n14311 | n6335;
assign n19554 = n12390 | n9747;
assign n8993 = ~(n1598 ^ n12041);
assign n1233 = n25443 & n26761;
assign n5403 = ~(n22005 ^ n19854);
assign n23249 = ~n12739;
assign n26032 = n9479 | n3506;
assign n23364 = ~(n8472 ^ n23905);
assign n1392 = n16952 | n14756;
assign n21164 = ~(n9410 ^ n8762);
assign n7363 = ~(n5138 ^ n14669);
assign n26554 = n4363 & n13097;
assign n4295 = ~(n17935 ^ n8111);
assign n2130 = ~(n1876 | n5675);
assign n19241 = ~n5868;
assign n7821 = n20265 | n23297;
assign n9488 = ~(n12288 | n7932);
assign n313 = n11754 | n19885;
assign n17024 = n23500 | n4831;
assign n19373 = ~n21417;
assign n10253 = n23064 | n25818;
assign n3622 = ~n14957;
assign n1960 = ~n11980;
assign n18588 = n11753 | n19928;
assign n12536 = n1649 & n165;
assign n696 = ~(n1080 ^ n16356);
assign n617 = ~n12751;
assign n960 = ~(n8386 ^ n7641);
assign n6866 = n22767 | n7022;
assign n4628 = n22626 | n18765;
assign n9734 = n22935 | n12881;
assign n16169 = n16029 | n12088;
assign n309 = n11569 | n4921;
assign n6881 = ~(n26939 ^ n10057);
assign n11352 = ~(n1124 ^ n25999);
assign n6516 = n12097 | n9000;
assign n1232 = ~n23019;
assign n11508 = ~(n24529 ^ n18171);
assign n10743 = ~n12204;
assign n494 = ~(n15112 ^ n26035);
assign n1423 = ~(n11901 | n17911);
assign n14718 = ~n17911;
assign n11085 = n705 & n20047;
assign n8039 = n5335 | n5143;
assign n22529 = n11605 | n24399;
assign n24630 = ~n25556;
assign n22755 = ~n3169;
assign n4245 = n25556 & n12169;
assign n19937 = n26723 | n2205;
assign n9309 = ~(n11580 | n1799);
assign n16488 = n8553 | n15502;
assign n5262 = ~(n990 | n19097);
assign n11063 = ~(n19773 ^ n2885);
assign n5879 = n14830 | n6468;
assign n15074 = ~n18687;
assign n12261 = n6094 & n12877;
assign n18344 = ~(n17233 ^ n8160);
assign n24228 = ~(n15656 ^ n27177);
assign n1042 = n16927 & n16652;
assign n3407 = ~n10199;
assign n21119 = ~(n6883 | n14681);
assign n25918 = ~(n24123 ^ n9377);
assign n17336 = n18496 | n20201;
assign n727 = ~(n17295 | n14289);
assign n23197 = n25545 & n9585;
assign n3319 = ~(n11142 ^ n20703);
assign n2141 = ~n4100;
assign n25623 = n17331 | n11291;
assign n11507 = ~(n586 ^ n7566);
assign n23915 = ~(n22715 ^ n25900);
assign n10357 = ~n3623;
assign n698 = ~n20840;
assign n8013 = ~n9135;
assign n22759 = n2262 & n11735;
assign n171 = n15974 | n2593;
assign n2170 = n15652 | n8151;
assign n13317 = ~(n4896 ^ n2146);
assign n4278 = ~(n903 ^ n996);
assign n3120 = ~(n12504 ^ n24975);
assign n5357 = ~(n1349 ^ n23065);
assign n12995 = n3695 & n10953;
assign n381 = ~(n528 | n25471);
assign n2914 = ~n6381;
assign n25880 = n1058 | n2521;
assign n7097 = ~(n5245 ^ n26893);
assign n2843 = n17887 | n18417;
assign n22218 = n3450 & n10293;
assign n6532 = ~(n20700 ^ n26510);
assign n562 = n5931 | n25711;
assign n3140 = ~(n2036 | n12391);
assign n2474 = n6717 & n24912;
assign n17432 = ~(n38 ^ n19098);
assign n20927 = ~(n18624 ^ n21505);
assign n11754 = n9598 & n21570;
assign n6903 = ~(n23160 ^ n8067);
assign n24751 = n24381 | n40;
assign n7438 = ~(n4108 ^ n26689);
assign n13998 = ~(n19797 ^ n3903);
assign n24854 = n22617 & n19091;
assign n6656 = n3538 | n23515;
assign n25293 = ~(n4226 ^ n4548);
assign n24610 = ~(n4490 | n21846);
assign n14442 = ~(n6309 | n17572);
assign n12267 = ~n16949;
assign n19389 = ~(n19809 ^ n25223);
assign n22164 = n5719 | n17911;
assign n18967 = ~(n13460 ^ n11455);
assign n26464 = n6452 | n8475;
assign n5613 = n26450 | n23109;
assign n6882 = ~(n22736 | n12741);
assign n10124 = ~(n26283 ^ n16847);
assign n20913 = ~(n1587 | n16524);
assign n8570 = ~(n16024 ^ n8355);
assign n8970 = n1611 | n6718;
assign n26925 = ~n10481;
assign n14839 = ~(n4538 ^ n8776);
assign n21154 = ~(n1610 ^ n18685);
assign n20702 = n22422 & n18648;
assign n8783 = n12601 & n591;
assign n12137 = n8045 & n13779;
assign n17551 = n25974 & n6963;
assign n6918 = ~(n10169 ^ n19132);
assign n13475 = n15871 & n10572;
assign n19761 = ~(n8614 | n25972);
assign n2134 = n5089 & n6059;
assign n13363 = n15854 | n4821;
assign n20265 = n17251 & n23967;
assign n27150 = ~n13041;
assign n4141 = ~(n15087 ^ n15147);
assign n6883 = ~(n21288 | n26522);
assign n14172 = ~(n7374 ^ n13613);
assign n12772 = ~(n23467 ^ n6030);
assign n11979 = n26356 & n3838;
assign n12726 = n965 & n7483;
assign n5215 = n19239 | n4513;
assign n5385 = ~(n18710 ^ n5621);
assign n23630 = ~(n22785 ^ n3638);
assign n15633 = ~n7285;
assign n26015 = ~n11986;
assign n20729 = n17116 | n7717;
assign n15287 = ~n16581;
assign n1019 = ~(n4639 ^ n7506);
assign n27044 = ~(n19352 ^ n12593);
assign n5831 = ~(n13789 | n6971);
assign n12823 = n658 | n2723;
assign n9311 = n17126 & n18112;
assign n10912 = n12853 & n4535;
assign n9898 = ~(n20564 ^ n8721);
assign n21907 = ~(n7316 ^ n25068);
assign n15816 = ~(n18476 ^ n12144);
assign n11720 = ~(n8431 ^ n8244);
assign n4510 = n10448 & n6471;
assign n4749 = ~n13022;
assign n3928 = n86 | n11543;
assign n18182 = n4722 | n14323;
assign n25177 = n18924 | n12701;
assign n9447 = n17668 & n11167;
assign n2931 = ~(n27144 ^ n6774);
assign n5615 = ~(n9069 ^ n20470);
assign n25767 = n24659 | n590;
assign n22149 = ~(n4360 | n25923);
assign n2226 = ~(n19962 ^ n7139);
assign n6989 = n7263 & n24968;
assign n7947 = n20332 & n20987;
assign n10730 = n1877 & n7265;
assign n14349 = n7831 | n6005;
assign n26481 = n17002 | n18274;
assign n12652 = ~n5607;
assign n10235 = ~(n22700 ^ n9655);
assign n21923 = n21346 & n19548;
assign n18920 = ~n15161;
assign n9257 = n12702 & n11144;
assign n8147 = n21652 | n21600;
assign n13024 = n954 | n6208;
assign n2837 = n17554 & n11203;
assign n25004 = ~n9507;
assign n9978 = n1611 & n6718;
assign n23605 = ~(n7858 ^ n21294);
assign n14957 = ~(n6942 ^ n24953);
assign n17089 = n12390 ^ n6948;
assign n6621 = n7437 | n26992;
assign n21467 = ~(n23678 | n2842);
assign n14688 = n9950 | n16332;
assign n26914 = ~n3730;
assign n15964 = ~(n2978 ^ n20040);
assign n6026 = ~(n16210 | n166);
assign n13905 = n9639 & n22580;
assign n14886 = ~(n27152 ^ n15794);
assign n24500 = n14680 & n8948;
assign n18891 = n17266 & n25239;
assign n952 = n26688 | n16727;
assign n5160 = ~n14919;
assign n9732 = n3018 & n16366;
assign n14238 = n8559 & n9579;
assign n10761 = ~(n16826 ^ n6636);
assign n721 = ~(n12149 ^ n1952);
assign n11911 = ~(n12246 ^ n25204);
assign n24805 = ~n964;
assign n21537 = ~(n24390 ^ n13426);
assign n6006 = ~(n17379 ^ n16353);
assign n5129 = n8759 | n20456;
assign n12473 = ~(n22289 | n2509);
assign n16683 = ~(n3224 ^ n7873);
assign n7130 = n16541;
assign n19223 = ~(n23204 ^ n7474);
assign n700 = n24905 | n6033;
assign n25344 = ~(n23936 | n1386);
assign n17356 = n8324 | n5574;
assign n18673 = ~(n8540 | n2399);
assign n1566 = n24695 | n2088;
assign n16912 = n17115 | n5675;
assign n19857 = ~(n11302 ^ n2146);
assign n22191 = ~(n19206 ^ n11556);
assign n8507 = ~(n8515 ^ n14599);
assign n17994 = ~n16295;
assign n15118 = ~(n18087 ^ n10350);
assign n23109 = ~(n209 ^ n1288);
assign n2433 = ~(n11580 ^ n24620);
assign n18682 = n10399 & n13322;
assign n21704 = n12464 & n25352;
assign n23182 = ~(n4022 | n9569);
assign n15377 = n26358 | n1986;
assign n26576 = n13646 | n16137;
assign n24782 = ~(n5112 ^ n5417);
assign n25956 = ~(n7466 ^ n6659);
assign n990 = ~n7949;
assign n22316 = n7841 | n9445;
assign n17438 = n17470 & n25998;
assign n24929 = ~n24990;
assign n4011 = n3541 | n9219;
assign n13348 = ~n10046;
assign n23318 = ~(n10172 ^ n11104);
assign n25227 = ~(n10632 | n1824);
assign n18850 = ~n2666;
assign n5320 = ~n8025;
assign n2898 = n3406 & n19126;
assign n8692 = ~(n643 ^ n22635);
assign n19250 = n5887 | n10541;
assign n7840 = ~(n26422 ^ n21747);
assign n16311 = ~n26520;
assign n5191 = ~(n16496 ^ n22456);
assign n11851 = n24083 | n7409;
assign n8159 = ~(n1491 ^ n794);
assign n6262 = ~n11525;
assign n18464 = n23737 | n6361;
assign n6174 = ~(n12811 ^ n3260);
assign n2159 = n24170 | n23460;
assign n18249 = n13731 | n24630;
assign n9809 = ~(n7197 ^ n14609);
assign n9611 = n13414 & n25233;
assign n8750 = ~(n14008 ^ n3785);
assign n16378 = ~(n14740 | n14698);
assign n26426 = n4265 | n12995;
assign n8394 = n16561 | n18139;
assign n13536 = n9978 | n5598;
assign n3292 = n4594 | n21348;
assign n18636 = ~(n6917 ^ n2323);
assign n22913 = n11959 | n15312;
assign n17623 = ~(n2210 ^ n16608);
assign n8620 = ~(n4106 ^ n4943);
assign n1141 = ~n17488;
assign n10651 = ~(n2838 ^ n2438);
assign n3623 = ~(n1824 ^ n1457);
assign n2734 = ~(n12236 ^ n19785);
assign n24743 = n22504 & n2907;
assign n9 = ~(n20517 ^ n18735);
assign n15929 = ~(n26030 ^ n20478);
assign n390 = ~(n5678 ^ n2678);
assign n12799 = n22911 & n11396;
assign n11719 = n11473 | n15506;
assign n14537 = n8358 | n24344;
assign n5710 = n22492 | n9372;
assign n4043 = n19677 & n2554;
assign n19297 = ~n18024;
assign n9620 = ~(n14361 ^ n3120);
assign n10639 = ~(n13603 ^ n6756);
assign n12356 = ~n1055;
assign n15201 = n24164 | n14937;
assign n8101 = ~n15241;
assign n16154 = n6809 | n6847;
assign n11718 = n4220 & n22869;
assign n8490 = ~(n5927 ^ n17160);
assign n24403 = ~n19177;
assign n20388 = ~(n15351 ^ n10216);
assign n15742 = ~(n632 | n25827);
assign n25538 = ~(n2066 ^ n20478);
assign n24603 = ~n24015;
assign n566 = ~(n17784 | n24085);
assign n24446 = ~(n9096 ^ n485);
assign n923 = ~(n15808 ^ n4160);
assign n5991 = ~(n16994 ^ n16521);
assign n11425 = ~n23697;
assign n3769 = n18140 & n7085;
assign n22166 = n8382 & n7644;
assign n15925 = ~(n15271 | n12161);
assign n14384 = ~(n6712 ^ n5332);
assign n8205 = ~(n6259 ^ n14838);
assign n2694 = n3584;
assign n27069 = ~n11224;
assign n2927 = ~(n3086 | n18213);
assign n16864 = n2323 | n6917;
assign n23746 = ~n4325;
assign n3107 = n2612 | n27193;
assign n3008 = n4102 | n20744;
assign n22685 = n3283 & n25746;
assign n4621 = n12002 | n11918;
assign n11139 = n2542 & n17057;
assign n23178 = n8155 | n20920;
assign n16364 = ~n24599;
assign n20016 = ~(n1040 | n12152);
assign n8642 = ~(n11533 | n11095);
assign n6358 = n26787 & n13792;
assign n23162 = ~n21235;
assign n912 = ~n11719;
assign n22885 = ~(n8910 ^ n9246);
assign n6249 = ~(n9514 ^ n3939);
assign n7951 = n14133 | n7524;
assign n23756 = n15581 | n5407;
assign n10216 = ~(n17901 ^ n8430);
assign n18766 = n26478 | n19721;
assign n10868 = ~n21890;
assign n11636 = n5181 | n11282;
assign n16884 = ~(n8328 | n24601);
assign n9869 = ~(n13062 | n5341);
assign n11544 = ~n19282;
assign n12901 = n17983 & n10458;
assign n11140 = ~(n16029 ^ n19228);
assign n9398 = ~n15495;
assign n8020 = ~(n2415 ^ n172);
assign n22915 = n18828 & n23904;
assign n3804 = n18675 & n22423;
assign n14131 = ~n15220;
assign n26037 = n16717 | n1817;
assign n22907 = ~(n15306 ^ n6098);
assign n22765 = ~n24935;
assign n10045 = ~(n2964 ^ n11554);
assign n2562 = ~n6513;
assign n19198 = n7362 & n16143;
assign n16374 = ~(n4128 ^ n20891);
assign n18672 = n22212 | n12510;
assign n12455 = ~(n19081 | n6283);
assign n6308 = ~(n21616 ^ n12852);
assign n19518 = ~(n17108 | n4008);
assign n26716 = n12156 & n22242;
assign n2434 = ~(n7657 | n25316);
assign n26875 = ~n12960;
assign n9405 = n15315 | n10419;
assign n6459 = n18216 | n19259;
assign n349 = ~n9897;
assign n1674 = ~(n21848 ^ n7207);
assign n12929 = ~n19144;
assign n12108 = ~(n26914 ^ n8497);
assign n12058 = ~(n7486 | n15787);
assign n10898 = n17333 | n14783;
assign n23491 = n1672 & n16765;
assign n141 = ~n6064;
assign n22804 = ~n12663;
assign n26825 = n19327 | n25624;
assign n13183 = n8153 | n16333;
assign n5494 = ~(n1896 | n8381);
assign n19776 = n23089 | n12877;
assign n23652 = ~(n20201 ^ n18496);
assign n4271 = ~(n22182 ^ n22427);
assign n26204 = n2323 & n6917;
assign n6965 = ~(n5777 ^ n18010);
assign n5926 = n27199 | n20151;
assign n4072 = n9893 | n22104;
assign n15318 = n13451 | n949;
assign n26824 = n25004 | n7375;
assign n25384 = n17290 & n2034;
assign n12739 = n15546 | n24922;
assign n7090 = n1432 & n12040;
assign n7193 = ~(n20259 ^ n3925);
assign n18149 = n23477 | n7913;
assign n7763 = n4277 | n23843;
assign n8831 = n4486 | n19980;
assign n17288 = ~(n21824 ^ n11877);
assign n7475 = n11102 | n20454;
assign n9197 = n12453 & n2908;
assign n15823 = n1091 | n15079;
assign n9767 = ~(n6337 ^ n6128);
assign n1443 = ~(n778 | n16291);
assign n4405 = ~(n18421 ^ n19163);
assign n3122 = ~(n14345 ^ n14702);
assign n6725 = n5131 | n11719;
assign n15648 = n6912 | n25656;
assign n27156 = ~n17045;
assign n20180 = n14431 | n25739;
assign n3037 = ~(n11517 ^ n20484);
assign n15844 = n836 | n14696;
assign n10947 = ~n2950;
assign n25591 = n13117 | n18833;
assign n25050 = ~n12386;
assign n9713 = ~(n2293 ^ n6716);
assign n22311 = ~(n15934 ^ n10864);
assign n8948 = ~n5031;
assign n13517 = n9934 & n20290;
assign n22133 = ~(n251 | n8438);
assign n22383 = ~(n4870 ^ n1350);
assign n23612 = ~(n5824 ^ n17984);
assign n12072 = ~(n3008 ^ n22902);
assign n15963 = ~(n22047 ^ n6352);
assign n25247 = n98 & n4830;
assign n19775 = ~(n25521 ^ n11554);
assign n2039 = ~(n2146 ^ n6785);
assign n16669 = ~(n12049 | n10464);
assign n14766 = ~(n20639 | n24125);
assign n3074 = ~(n24081 | n14255);
assign n21109 = n4056 | n11555;
assign n21476 = ~(n9546 | n14758);
assign n13865 = ~(n24358 | n13781);
assign n24736 = ~(n2759 ^ n8052);
assign n769 = n8970 & n13536;
assign n26280 = ~(n24465 ^ n6602);
assign n24664 = ~n4183;
assign n4532 = ~(n14032 ^ n19152);
assign n26703 = ~(n12533 ^ n24927);
assign n4456 = n23997 | n15215;
assign n19993 = n24199 & n14020;
assign n1024 = n15157 & n8828;
assign n25041 = ~n26660;
assign n18651 = ~n14576;
assign n23379 = n11643 | n14590;
assign n4545 = n3349 & n10501;
assign n4980 = n13847 & n18206;
assign n14753 = n20105 & n9589;
assign n15576 = ~n8386;
assign n18112 = n8955 | n5741;
assign n16265 = n20569 & n3597;
assign n7622 = n20784 & n2897;
assign n9068 = ~n6971;
assign n12509 = ~n23789;
assign n21242 = n8430 | n11701;
assign n9965 = n22954 | n190;
assign n934 = n11418 & n14582;
assign n22593 = n22980 & n13363;
assign n2997 = ~n17171;
assign n481 = ~n2944;
assign n4968 = n26146 | n23891;
assign n1380 = n1917;
assign n20619 = n21291 & n14828;
assign n22151 = n15490 & n328;
assign n190 = n17011 & n23501;
assign n23045 = n14829 ^ n1165;
assign n19390 = n26546;
assign n10015 = n4507 & n9389;
assign n14248 = n13535 | n1047;
assign n9040 = ~(n11473 ^ n15506);
assign n19825 = ~(n21137 ^ n14130);
assign n22673 = ~(n1403 | n5284);
assign n14773 = ~(n24727 ^ n905);
assign n19182 = n9634 & n5190;
assign n22874 = n2972 & n8639;
assign n15881 = ~(n14965 ^ n10389);
assign n23568 = ~(n15212 ^ n8174);
assign n20407 = ~(n14444 | n5616);
assign n11032 = ~(n9242 ^ n25240);
assign n12966 = ~(n13137 ^ n7674);
assign n12567 = ~(n14179 ^ n19455);
assign n12704 = ~(n16683 | n16882);
assign n16245 = n3392 & n19582;
assign n4915 = ~(n9832 | n6513);
assign n1422 = n16856 | n21081;
assign n4850 = ~(n21597 ^ n440);
assign n11278 = ~n5374;
assign n1127 = ~(n5440 | n2724);
assign n10563 = ~(n14603 ^ n15053);
assign n12264 = n18994 | n7787;
assign n15813 = n2740 & n20949;
assign n8824 = ~(n192 ^ n26884);
assign n17872 = ~(n2267 ^ n6099);
assign n20533 = n10218 & n3523;
assign n4598 = n12126 | n7023;
assign n26790 = ~(n4663 | n19390);
assign n14114 = ~n4275;
assign n26074 = n12511 | n19196;
assign n11122 = ~(n7524 | n19680);
assign n22302 = ~n12015;
assign n12519 = n5549 | n8302;
assign n15792 = ~n23279;
assign n12664 = n24325 & n10937;
assign n2415 = ~(n12984 ^ n3468);
assign n1497 = n16833 & n20592;
assign n22732 = ~(n15182 | n12090);
assign n7091 = ~(n10501 ^ n3349);
assign n21671 = ~n16136;
assign n5479 = ~n14461;
assign n7362 = n1118 | n6477;
assign n17335 = n22770 | n14029;
assign n3304 = n2351 & n8377;
assign n11195 = ~n6501;
assign n25677 = n8927 & n17574;
assign n870 = ~(n21825 ^ n16514);
assign n21634 = ~n12821;
assign n975 = n23806 & n17629;
assign n25042 = n10837 & n1576;
assign n5784 = ~(n26660 ^ n1163);
assign n4625 = ~(n24982 ^ n20268);
assign n790 = ~(n4591 ^ n26562);
assign n6902 = ~(n15447 ^ n24951);
assign n8952 = ~n20707;
assign n8772 = ~(n22946 ^ n25053);
assign n6365 = n18030 & n4612;
assign n25811 = n15178 | n16263;
assign n21789 = ~(n1396 ^ n15967);
assign n22033 = n16120 & n19937;
assign n24401 = n4819 | n210;
assign n9094 = ~(n17995 | n462);
assign n25156 = n20413;
assign n10144 = n17083 | n17989;
assign n14202 = ~(n5739 ^ n16386);
assign n395 = ~n4822;
assign n12677 = n11563 & n24232;
assign n22084 = n5088 & n26110;
assign n25171 = ~n12322;
assign n10474 = n8580 | n587;
assign n3774 = n9617 | n10268;
assign n22948 = ~(n10470 | n11775);
assign n19898 = ~n2858;
assign n5545 = n25341 & n5173;
assign n7537 = n643 & n17804;
assign n10087 = n19950 | n24011;
assign n21326 = n19794 | n23810;
assign n23438 = n13117 | n20084;
assign n2684 = n7759 | n725;
assign n23156 = n10077 & n9285;
assign n3223 = ~(n17167 ^ n2546);
assign n15920 = n23592 | n14440;
assign n21996 = n11874 & n6994;
assign n7333 = n16067 & n6937;
assign n1894 = ~(n17139 ^ n25198);
assign n18027 = ~n26119;
assign n12926 = n24943 & n21027;
assign n1050 = n16102 & n3922;
assign n21917 = n616 | n13579;
assign n13270 = ~(n10515 ^ n16849);
assign n8792 = ~n10777;
assign n25710 = n1953 | n13585;
assign n22898 = n7901 & n13864;
assign n26368 = n10619 | n23675;
assign n1936 = n6675 & n12895;
assign n17948 = ~(n2909 ^ n9426);
assign n11657 = ~n11476;
assign n11819 = n16664 & n2848;
assign n2727 = n22275 | n17680;
assign n12004 = ~n18;
assign n21876 = n12650 & n14765;
assign n720 = n21068 & n11190;
assign n15389 = ~n8144;
assign n11705 = n6803 | n1509;
assign n26351 = ~n10560;
assign n20645 = n7676 & n12512;
assign n21964 = ~(n4022 ^ n14565);
assign n18988 = n8572 | n5939;
assign n324 = ~(n14684 ^ n22588);
assign n26473 = n16547 | n15;
assign n16744 = ~(n2558 ^ n14691);
assign n10584 = n4863 & n23622;
assign n26293 = ~n25885;
assign n11426 = ~(n10220 ^ n15901);
assign n2883 = n12002 & n27102;
assign n17182 = n8685 | n21283;
assign n17306 = ~(n9655 ^ n20946);
assign n21877 = n26588 & n4573;
assign n961 = ~(n24410 | n11662);
assign n19153 = n744 | n21038;
assign n23004 = n20049 & n13806;
assign n17942 = n11676 | n13037;
assign n23545 = n13411 | n4090;
assign n19894 = ~(n16171 ^ n5786);
assign n9817 = ~(n17330 ^ n5414);
assign n25163 = n337 | n16507;
assign n17264 = n24263 | n3608;
assign n18721 = ~(n22013 ^ n17681);
assign n12759 = n1938 | n25790;
assign n10673 = n4533 | n6340;
assign n21417 = ~(n5704 ^ n12315);
assign n19743 = n1183 | n8582;
assign n3370 = ~(n24620 ^ n7099);
assign n2961 = ~(n25290 ^ n10783);
assign n11927 = n1864 | n17035;
assign n18313 = ~(n2389 ^ n3007);
assign n7116 = n2589 & n3087;
assign n12467 = ~(n25186 ^ n1516);
assign n11833 = ~n24182;
assign n10875 = n12317 & n10394;
assign n1734 = ~(n11830 | n18006);
assign n23487 = ~n25074;
assign n3968 = ~(n8742 ^ n21789);
assign n26059 = ~(n1405 | n9067);
assign n20698 = n7915 | n5231;
assign n11415 = ~(n17734 ^ n10639);
assign n24778 = ~n4193;
assign n24367 = ~n7221;
assign n8598 = ~(n9332 ^ n5145);
assign n5004 = ~(n13898 | n14275);
assign n21606 = n7005 & n26820;
assign n13518 = n13833 ^ n1168;
assign n6577 = n7899 | n22388;
assign n7973 = ~n20382;
assign n22760 = ~(n11542 | n15079);
assign n13500 = ~(n9819 ^ n14960);
assign n4457 = n3520 & n19235;
assign n14765 = ~(n5234 ^ n12702);
assign n21182 = ~(n25428 ^ n16522);
assign n9705 = n20478 & n26030;
assign n16983 = ~(n25316 ^ n20385);
assign n18792 = ~(n7591 ^ n23680);
assign n4252 = n8958 | n21014;
assign n5852 = ~n1138;
assign n13883 = n23526 | n25081;
assign n26003 = n4446 | n4734;
assign n19345 = n15317 | n21568;
assign n25619 = ~(n5281 ^ n13176);
assign n16411 = n25287 & n23538;
assign n15426 = ~n26913;
assign n26465 = ~(n5402 | n7361);
assign n19869 = ~n1913;
assign n1182 = ~n3506;
assign n8702 = n16153 & n25116;
assign n21549 = ~(n8506 ^ n11584);
assign n17263 = ~(n3569 ^ n21013);
assign n22108 = ~n8583;
assign n21871 = ~n25494;
assign n9631 = ~n2331;
assign n4970 = ~n21082;
assign n16435 = n25255 | n17321;
assign n374 = n15823 & n15606;
assign n27204 = n21716 | n4457;
assign n16948 = ~(n15484 ^ n24964);
assign n17145 = n18740 & n20283;
assign n11368 = n22510 | n14306;
assign n4535 = n19718 | n16956;
assign n16232 = ~(n1653 ^ n8913);
assign n27050 = n6029 | n758;
assign n4548 = ~(n12944 ^ n2439);
assign n22882 = n7809 & n15038;
assign n8727 = n2416 | n16455;
assign n14414 = ~(n14213 ^ n18252);
assign n5632 = n7040 | n12799;
assign n24177 = ~(n20851 ^ n5385);
assign n20117 = ~n196;
assign n19113 = ~n26879;
assign n24152 = ~n9358;
assign n7889 = n24136 | n18806;
assign n24847 = ~(n27126 ^ n26068);
assign n25228 = ~n9192;
assign n24811 = n8077 | n10843;
assign n24810 = ~(n4626 | n21509);
assign n11601 = n27122 | n17251;
assign n6895 = ~n13858;
assign n6158 = n5735 & n9132;
assign n26166 = n9196 | n12354;
assign n20911 = n14823 | n12753;
assign n26367 = ~n14878;
assign n5897 = n12951 & n9704;
assign n13420 = ~n5673;
assign n12534 = ~(n10023 | n6670);
assign n23985 = n19293 & n659;
assign n9843 = n4236 & n8239;
assign n10142 = n4711 | n715;
assign n20092 = ~(n4032 ^ n17898);
assign n12531 = ~(n15308 ^ n3202);
assign n18811 = n16420 | n2233;
assign n6389 = n17655 & n10144;
assign n8813 = ~(n4469 | n23545);
assign n11795 = n5578 | n1493;
assign n10237 = n9291 | n1413;
assign n13947 = ~(n26942 ^ n9498);
assign n24237 = ~n25250;
assign n7914 = n3739 & n15892;
assign n24468 = ~n17792;
assign n12382 = n13105 & n1551;
assign n3549 = ~n10422;
assign n235 = ~(n5845 ^ n9566);
assign n1965 = n24330 & n5320;
assign n2218 = ~n16314;
assign n17431 = ~n10706;
assign n10267 = ~(n5322 ^ n21488);
assign n16314 = ~(n6455 ^ n25467);
assign n1846 = n20385 & n23932;
assign n2278 = n14557 | n16982;
assign n19399 = ~(n5307 ^ n22646);
assign n14528 = n12367;
assign n4547 = ~(n2732 | n21085);
assign n5888 = n26168 | n19660;
assign n2466 = n14309 | n9611;
assign n23125 = n6729 | n1106;
assign n1355 = n20945 | n22953;
assign n3881 = n12856 & n24703;
assign n22209 = ~(n19313 | n20444);
assign n5549 = ~(n23622 ^ n20199);
assign n7919 = ~(n1493 ^ n12585);
assign n3266 = ~(n7593 | n17415);
assign n9413 = ~(n12805 ^ n12350);
assign n23610 = ~(n8491 ^ n25586);
assign n13580 = n24442 & n4541;
assign n25061 = ~(n16276 ^ n24374);
assign n8999 = ~(n4665 | n7823);
assign n26033 = n20277 | n17460;
assign n21873 = ~(n22597 | n18901);
assign n9717 = ~n24842;
assign n1863 = ~(n1040 ^ n12152);
assign n21590 = ~(n13291 ^ n2443);
assign n13689 = n8838 & n1987;
assign n15585 = n2915 & n10625;
assign n5388 = ~(n12078 | n3354);
assign n24256 = ~(n19058 ^ n9445);
assign n11820 = n26574 | n5664;
assign n13977 = n6400 | n18554;
assign n7722 = ~(n5358 ^ n20726);
assign n2650 = ~(n20051 ^ n4901);
assign n6074 = n19934 & n24224;
assign n26956 = n23705 | n21287;
assign n14951 = n2254 & n13458;
assign n18021 = n24716 | n20875;
assign n14451 = ~(n2566 ^ n23677);
assign n5254 = n1459 & n8193;
assign n26080 = n8230 & n20653;
assign n23207 = ~(n18834 ^ n14231);
assign n1559 = ~(n26957 | n14130);
assign n26217 = n2886 & n16609;
assign n13529 = ~n27175;
assign n13557 = ~(n26951 ^ n22477);
assign n17636 = ~(n3116 ^ n24980);
assign n11673 = n8255 | n5;
assign n24797 = n8539 | n14610;
assign n21630 = ~(n13968 ^ n18649);
assign n14434 = n4780 | n15258;
assign n17890 = n16528 | n4503;
assign n17320 = ~(n25755 ^ n7358);
assign n19306 = n14156 | n11552;
assign n18075 = ~(n24323 ^ n1681);
assign n10148 = ~n8508;
assign n601 = ~(n19464 | n5108);
assign n13885 = ~(n26000 ^ n2394);
assign n10713 = ~(n12076 ^ n8856);
assign n4908 = n24564 & n15962;
assign n12988 = ~(n21520 | n19615);
assign n15957 = n20964 & n6762;
assign n4649 = ~(n9402 ^ n6864);
assign n8973 = ~(n20213 ^ n26725);
assign n20589 = ~(n19914 | n24551);
assign n23482 = n18546 | n25834;
assign n1501 = ~(n17616 ^ n959);
assign n21827 = ~(n1339 ^ n21842);
assign n18400 = ~(n12962 ^ n26662);
assign n988 = n146 | n16889;
assign n24606 = ~(n22810 ^ n22120);
assign n11723 = n7288 & n19064;
assign n20137 = ~n7437;
assign n7488 = n24574 | n16228;
assign n22061 = ~n18425;
assign n17292 = ~(n15087 | n3257);
assign n15145 = ~(n25894 ^ n8205);
assign n2379 = n20586 & n7299;
assign n7255 = n1418 | n2878;
assign n5256 = ~(n12270 ^ n15963);
assign n15253 = n26710 & n15418;
assign n12912 = n20463 & n13687;
assign n3552 = ~(n291 ^ n5117);
assign n6817 = n12221 & n19049;
assign n15888 = n25004 & n7375;
assign n19465 = n26312 & n26993;
assign n19324 = n15027 & n8030;
assign n2020 = n22161 & n19931;
assign n23473 = ~(n16313 ^ n15164);
assign n9121 = n13737 | n16907;
assign n26433 = ~n11670;
assign n12070 = ~(n25729 ^ n3279);
assign n11641 = n2317 | n5109;
assign n20916 = n5535 & n23137;
assign n21847 = ~(n11566 | n12198);
assign n4522 = ~(n6692 | n15661);
assign n4799 = ~(n24736 | n8713);
assign n12156 = n10037 | n19196;
assign n23105 = n16232 | n22294;
assign n21887 = n16830 | n18295;
assign n26028 = ~(n19820 ^ n1057);
assign n1107 = n7421 & n20044;
assign n4602 = n12318 & n25955;
assign n20664 = n2543 & n19810;
assign n14118 = ~n16260;
assign n16641 = n13357 & n11077;
assign n4906 = n8854 & n19145;
assign n16246 = ~(n1553 | n3547);
assign n24398 = n4615 | n26233;
assign n5229 = ~(n1839 | n5886);
assign n2857 = ~n9110;
assign n9715 = n12356 | n1545;
assign n4097 = n504 & n26135;
assign n212 = ~n6785;
assign n22509 = ~(n20470 ^ n3366);
assign n17279 = ~(n5260 ^ n16130);
assign n20078 = n17002 | n7731;
assign n7276 = ~(n12163 ^ n10139);
assign n4236 = ~n14258;
assign n9433 = ~(n11580 | n19230);
assign n24867 = n9143 & n16697;
assign n2954 = ~(n13288 ^ n18874);
assign n20379 = ~(n8722 | n10791);
assign n6726 = ~(n19824 ^ n22406);
assign n25346 = ~(n17926 ^ n17598);
assign n21089 = ~(n22742 ^ n26903);
assign n25939 = ~n5231;
assign n19676 = n13842 | n13708;
assign n3360 = n8610 & n4689;
assign n14894 = n5540 & n14179;
assign n23636 = ~(n802 ^ n21629);
assign n10506 = ~(n9576 ^ n21599);
assign n17708 = ~(n26222 | n12565);
assign n24242 = ~(n21907 ^ n26054);
assign n19134 = ~n6915;
assign n22337 = n6996 | n8570;
assign n10366 = n25054 & n10138;
assign n11298 = ~(n13081 ^ n18729);
assign n2157 = n8086 & n26948;
assign n24739 = ~(n22203 ^ n20259);
assign n18974 = ~(n6118 ^ n1521);
assign n4417 = n3061 | n2808;
assign n17912 = ~(n6353 ^ n12242);
assign n22512 = n17794 | n22551;
assign n20899 = n6010 | n22989;
assign n10418 = n4679 & n19102;
assign n2497 = n23467 | n10772;
assign n7436 = ~(n13458 ^ n25793);
assign n5050 = ~(n10308 ^ n7163);
assign n22860 = n24170 | n24085;
assign n22352 = n3005 & n9348;
assign n20660 = ~(n20088 | n5086);
assign n25460 = ~(n14744 ^ n691);
assign n3150 = ~(n316 ^ n24210);
assign n11378 = n17568 & n3171;
assign n27140 = ~(n11714 | n10861);
assign n19741 = ~(n2215 ^ n8706);
assign n5035 = n736 | n9148;
assign n16532 = ~n4787;
assign n4730 = n4132 | n2005;
assign n7359 = ~n12610;
assign n16263 = n5879 & n20806;
assign n1893 = ~(n7846 ^ n9609);
assign n15538 = n400 | n19478;
assign n22618 = ~(n7619 ^ n11044);
assign n25197 = n26766 | n21664;
assign n22648 = n15102 & n8237;
assign n1793 = ~(n26882 | n106);
assign n20346 = n24972 | n5429;
assign n5396 = n11205 | n19975;
assign n21886 = n379 & n20671;
assign n22408 = ~n1441;
assign n9842 = n1290 & n22657;
assign n3905 = n22116 | n15605;
assign n8926 = n21969 | n19284;
assign n18363 = ~n15392;
assign n4947 = ~(n19096 ^ n19063);
assign n17046 = n18643 | n14314;
assign n24827 = ~(n21037 | n13899);
assign n23206 = n21961 | n16121;
assign n10890 = n21947 & n16525;
assign n8266 = ~n690;
assign n20512 = ~(n27184 ^ n4812);
assign n7642 = ~(n11457 | n6385);
assign n15641 = n7921 | n1065;
assign n41 = n2773 | n12927;
assign n12713 = n19672 & n19987;
assign n15605 = n1189 & n15195;
assign n603 = n9598 | n7759;
assign n6501 = ~(n21656 ^ n20519);
assign n5774 = ~n6229;
assign n23708 = ~n15960;
assign n1081 = ~(n10224 ^ n11481);
assign n2721 = ~n13549;
assign n20524 = n13577 | n23587;
assign n17301 = ~n8957;
assign n4377 = n21229 | n7036;
assign n17758 = ~(n5704 ^ n22309);
assign n47 = n21359 | n23384;
assign n13506 = ~(n24803 ^ n227);
assign n1756 = n8804 & n12729;
assign n2924 = n5705 & n3227;
assign n15409 = ~(n27104 | n19005);
assign n8481 = n23072 | n26384;
assign n25941 = ~n15586;
assign n10255 = ~n17142;
assign n4106 = ~(n13372 ^ n1681);
assign n3340 = ~(n23172 ^ n20578);
assign n10594 = n17022 | n150;
assign n5687 = ~(n24550 ^ n4791);
assign n21121 = n9102 | n19180;
assign n18943 = ~(n9204 ^ n7359);
assign n2581 = n1868 | n26791;
assign n15221 = ~n9003;
assign n4554 = ~(n5304 ^ n20516);
assign n12740 = ~(n4292 ^ n14454);
assign n14101 = n20753 & n14581;
assign n8366 = ~(n14255 ^ n5882);
assign n3477 = ~(n22382 ^ n23326);
assign n11001 = n10075 | n8225;
assign n14749 = ~(n10286 ^ n25044);
assign n17221 = n1595 & n12820;
assign n25903 = n15809 & n181;
assign n26268 = n12044 & n11231;
assign n18428 = ~(n25806 ^ n9445);
assign n25348 = n2436 | n11714;
assign n5588 = n4415 | n23859;
assign n14992 = ~n2416;
assign n12257 = n20501 & n14476;
assign n5664 = n21059 & n10921;
assign n7756 = ~(n12343 | n25568);
assign n13441 = n4413 & n23116;
assign n16595 = ~(n10760 ^ n10882);
assign n2699 = ~(n7497 ^ n22863);
assign n15000 = ~n12674;
assign n16336 = n15404 & n10610;
assign n20368 = n25716 | n25708;
assign n22453 = n23617 | n21493;
assign n25097 = ~(n25911 ^ n1724);
assign n3851 = ~(n2510 ^ n7678);
assign n5537 = n17841 & n19096;
assign n19075 = n503 & n25056;
assign n22501 = ~n25855;
assign n20673 = ~(n3734 ^ n25984);
assign n1105 = ~n1834;
assign n10180 = n15918 | n21021;
assign n5868 = ~(n5993 ^ n1185);
assign n1468 = n784 | n21692;
assign n24101 = ~n2551;
assign n18236 = ~(n6753 | n2453);
assign n13513 = ~(n21247 | n1631);
assign n1669 = ~(n6831 | n7546);
assign n11567 = ~(n6502 ^ n1630);
assign n18895 = ~(n14735 ^ n16812);
assign n22798 = n11796 & n21464;
assign n17699 = n16789 & n10962;
assign n3987 = ~(n23974 ^ n8309);
assign n19670 = ~(n1630 ^ n11121);
assign n12694 = n20990 & n13344;
assign n7262 = n13488 | n6520;
assign n18352 = ~(n7170 | n19186);
assign n3100 = ~(n10146 | n329);
assign n12993 = n3643 & n24883;
assign n14037 = n8801 | n5889;
assign n8239 = ~n22846;
assign n20879 = ~(n13509 ^ n4861);
assign n6275 = ~(n3832 | n20006);
assign n24802 = ~n8170;
assign n13315 = n5576 & n1763;
assign n22388 = n25472 & n1966;
assign n2840 = n20112 | n2161;
assign n15658 = ~(n7297 | n304);
assign n15446 = n24480 & n14634;
assign n24794 = n14440 | n7523;
assign n19562 = ~(n13677 ^ n26752);
assign n2444 = ~(n4336 ^ n24967);
assign n20373 = n8117 | n3280;
assign n26313 = ~(n15659 ^ n5213);
assign n24681 = ~(n4685 ^ n21213);
assign n20707 = ~(n7562 ^ n5584);
assign n14212 = n23322 | n12185;
assign n9738 = n18511 & n14361;
assign n513 = n14192 ^ n3320;
assign n25521 = ~n24188;
assign n13748 = ~n5288;
assign n5655 = n5207 | n21284;
assign n956 = ~(n11623 ^ n19938);
assign n20111 = ~(n5400 ^ n9512);
assign n17132 = ~(n6755 ^ n13988);
assign n8379 = ~(n683 ^ n21299);
assign n20428 = n18053 & n2844;
assign n8590 = n11964 | n12345;
assign n22275 = n1099 & n3379;
assign n10213 = n11947 | n23271;
assign n8536 = n25439 | n14782;
assign n3303 = n944 | n22738;
assign n17940 = ~(n21878 ^ n17743);
assign n2595 = n9638 | n18631;
assign n2772 = n11170 | n8260;
assign n20355 = ~(n11784 ^ n70);
assign n5168 = ~(n8392 ^ n27153);
assign n348 = ~(n16704 ^ n5981);
assign n18243 = ~(n19153 ^ n27044);
assign n5429 = ~n11611;
assign n8759 = ~(n17056 | n23545);
assign n6928 = ~(n23464 ^ n9877);
assign n7989 = n9206 | n6597;
assign n17412 = ~(n15471 ^ n17712);
assign n26687 = n18950 | n17846;
assign n23850 = n24054 | n14032;
assign n26954 = ~(n25068 ^ n8324);
assign n23263 = n25340 | n15744;
assign n23863 = ~n14345;
assign n10488 = ~(n8472 | n6150);
assign n10380 = n19297 | n23754;
assign n21541 = n9294 | n18880;
assign n12499 = n19546 | n5130;
assign n20795 = ~(n14016 ^ n21106);
assign n15021 = n24325 | n21353;
assign n13558 = ~(n22205 ^ n26288);
assign n24967 = ~(n23161 ^ n22237);
assign n16823 = ~(n9928 ^ n6785);
assign n16403 = n20931 & n6144;
assign n16570 = n1873 & n10814;
assign n24901 = n17164 & n18726;
assign n14138 = ~n1599;
assign n24378 = ~(n22567 ^ n4532);
assign n23911 = ~(n2944 ^ n13951);
assign n21498 = n13108 ^ n5026;
assign n6643 = n16335 & n23893;
assign n11502 = ~n502;
assign n274 = ~(n14208 ^ n2547);
assign n11918 = ~(n13313 ^ n18959);
assign n17162 = n24025 & n20951;
assign n24210 = ~(n7436 ^ n5098);
assign n11007 = n17066 | n22773;
assign n24960 = ~n8551;
assign n11431 = ~(n19594 ^ n6235);
assign n9677 = n7361 | n14885;
assign n2054 = ~(n16393 ^ n11653);
assign n1129 = ~(n19227 ^ n19005);
assign n11324 = n25957 & n19247;
assign n1176 = ~n3136;
assign n26290 = ~(n19797 ^ n24620);
assign n2486 = ~(n10660 | n8897);
assign n9191 = ~(n5725 ^ n1499);
assign n6552 = n225 | n26181;
assign n21470 = n14851 & n3036;
assign n2817 = ~(n20700 ^ n12875);
assign n4994 = n7569 | n1779;
assign n9981 = ~(n21841 ^ n12693);
assign n406 = n20155 & n24424;
assign n12247 = n2230 | n18295;
assign n4986 = ~(n9133 | n393);
assign n9997 = n23561 & n10364;
assign n20848 = n11778 & n21121;
assign n19414 = ~(n13181 ^ n16447);
assign n24595 = ~(n13419 | n23475);
assign n14567 = n23614 & n17611;
assign n25858 = ~(n4119 ^ n1525);
assign n8905 = n21061 & n22956;
assign n12200 = n7487 | n16571;
assign n25215 = ~(n12368 ^ n2881);
assign n20176 = ~(n23642 ^ n24309);
assign n24365 = ~(n15884 ^ n5213);
assign n5733 = ~(n19643 ^ n9694);
assign n21819 = n10013 | n25971;
assign n2381 = n9119 | n9929;
assign n12327 = ~(n21334 | n18399);
assign n2794 = ~(n25394 ^ n8964);
assign n13713 = ~(n21489 | n11151);
assign n2993 = ~(n2731 ^ n4812);
assign n11174 = ~(n15090 ^ n20608);
assign n11638 = n20336 & n23233;
assign n1466 = n3782 & n8474;
assign n7649 = n22670 | n21050;
assign n7548 = n20948 & n5946;
assign n6849 = n5663 & n4945;
assign n3862 = ~n3554;
assign n6380 = n13275 & n14427;
assign n22683 = ~(n18351 ^ n9024);
assign n20062 = ~(n9600 | n3791);
assign n22223 = ~(n22009 | n24839);
assign n1784 = ~(n15284 ^ n8772);
assign n17927 = ~(n24303 ^ n1027);
assign n26086 = ~n16971;
assign n24667 = n19763 | n4922;
assign n21520 = ~n19955;
assign n17663 = ~(n23149 ^ n7240);
assign n15890 = ~(n20415 | n14852);
assign n5287 = n18098 | n13530;
assign n19184 = ~(n16671 ^ n20690);
assign n16600 = ~(n23063 | n19494);
assign n21565 = ~n75;
assign n2947 = n26621 & n5136;
assign n22414 = ~(n5468 ^ n16801);
assign n14058 = n26246 & n20778;
assign n12233 = n9675 | n11723;
assign n11497 = ~(n24027 ^ n24956);
assign n2259 = n16162 & n693;
assign n15574 = ~(n10625 ^ n19454);
assign n20697 = n9232 & n11042;
assign n6134 = ~(n11740 | n19941);
assign n10501 = ~n9550;
assign n4397 = n1398 & n20548;
assign n1332 = ~(n26570 ^ n15105);
assign n10479 = ~(n12139 ^ n17891);
assign n15147 = ~n14163;
assign n229 = n3525 | n17935;
assign n25826 = ~(n9414 ^ n538);
assign n18420 = ~(n14336 | n20077);
assign n26685 = n17494 | n15450;
assign n26957 = ~n14440;
assign n6840 = n5846 | n21950;
assign n4212 = n16003 | n489;
assign n13396 = n13643 | n6466;
assign n24927 = ~(n10158 ^ n1136);
assign n13485 = ~n3716;
assign n7100 = ~(n25034 ^ n7975);
assign n530 = ~n21267;
assign n23208 = ~n24736;
assign n22224 = ~(n6355 | n8589);
assign n3361 = n19621 & n27204;
assign n20459 = n11655 | n4644;
assign n17208 = ~(n8492 | n25739);
assign n17946 = n20562 | n13109;
assign n20840 = ~(n4406 ^ n8810);
assign n7598 = ~(n14712 ^ n10714);
assign n20888 = n6641 | n17952;
assign n21303 = n20645 | n21475;
assign n5492 = n12129 | n26173;
assign n18874 = ~(n13158 ^ n8309);
assign n15038 = ~n25100;
assign n4685 = ~(n26004 ^ n26896);
assign n10520 = ~(n22671 ^ n17975);
assign n191 = ~(n14637 | n11210);
assign n22002 = ~(n24677 ^ n10866);
assign n15772 = n9642 & n6331;
assign n10709 = ~(n13140 ^ n4158);
assign n16828 = ~(n16455 ^ n2416);
assign n1494 = n12096 | n9488;
assign n23964 = ~(n22671 ^ n22017);
assign n14970 = ~(n6141 ^ n5028);
assign n21099 = n12435 | n16281;
assign n26089 = n15188 & n24725;
assign n14679 = ~(n16662 ^ n7769);
assign n13578 = ~(n15451 ^ n1949);
assign n14551 = ~(n5342 | n17559);
assign n16343 = n18266 | n11814;
assign n25533 = ~n5110;
assign n21104 = ~n5017;
assign n23876 = ~(n11197 ^ n25878);
assign n6217 = n14406 | n19643;
assign n12742 = ~(n2830 ^ n22394);
assign n9590 = n11286 | n7392;
assign n14577 = ~(n11486 ^ n20235);
assign n5962 = n20059 | n17671;
assign n21175 = ~(n17868 ^ n4141);
assign n11204 = n17745 & n15843;
assign n14127 = ~n15914;
assign n24536 = ~(n26338 ^ n18166);
assign n3917 = n25149 & n12948;
assign n13238 = n25099 | n20455;
assign n12406 = ~(n12691 ^ n25080);
assign n7419 = ~(n19869 | n676);
assign n5364 = ~(n905 | n24727);
assign n15663 = ~(n21 ^ n20923);
assign n5266 = ~n24745;
assign n6676 = n15311 | n7574;
assign n22490 = n17214 & n15907;
assign n3821 = n22764 | n2360;
assign n21205 = ~(n10070 ^ n26483);
assign n3137 = n17035 | n2680;
assign n9747 = n12955 & n7353;
assign n10681 = ~n25001;
assign n7001 = ~(n14873 ^ n9452);
assign n20051 = ~n24117;
assign n18412 = n11459 & n18781;
assign n1170 = ~(n20427 ^ n24860);
assign n17504 = ~(n2360 ^ n17458);
assign n16177 = n24765 | n23447;
assign n15855 = n23806 | n17629;
assign n10963 = n1978 | n17055;
assign n15293 = ~(n18506 | n19514);
assign n9015 = ~n16981;
assign n2856 = ~(n19514 | n2415);
assign n25359 = ~(n14122 ^ n22300);
assign n1520 = n1110 | n9553;
assign n4712 = ~(n6033 ^ n21658);
assign n20131 = ~n26557;
assign n605 = ~(n13301 | n23313);
assign n4287 = n14790 | n342;
assign n4324 = n20212 & n6472;
assign n27147 = ~n24194;
assign n7075 = n12303 | n2406;
assign n1903 = n17595 & n14134;
assign n18494 = n18848 & n20038;
assign n17216 = n5312 & n7800;
assign n15483 = n6040 & n26812;
assign n21321 = ~n4008;
assign n12802 = ~n15009;
assign n23935 = ~(n19436 ^ n9792);
assign n16574 = ~(n13053 ^ n24150);
assign n17684 = ~(n13949 ^ n5128);
assign n24918 = n13434 & n390;
assign n18166 = ~(n26510 ^ n22332);
assign n17532 = ~n11667;
assign n26713 = ~(n15125 ^ n9130);
assign n7895 = n23877 | n25918;
assign n11541 = n11788 | n5301;
assign n26227 = ~n4199;
assign n4601 = ~(n1452 ^ n14236);
assign n9053 = ~n3740;
assign n4373 = n14948 & n6973;
assign n5606 = n13188 | n5738;
assign n24071 = n20964 | n20946;
assign n2243 = n7228 & n2991;
assign n11304 = ~(n6168 ^ n7555);
assign n3824 = n18990 | n673;
assign n11735 = n21307 | n25103;
assign n12636 = ~(n9204 | n12251);
assign n18606 = ~n669;
assign n2656 = ~n1708;
assign n2269 = ~(n8647 | n24343);
assign n23187 = n16889 & n8278;
assign n12951 = n20737 | n919;
assign n18773 = ~(n15433 | n15539);
assign n3110 = n18318 | n20171;
assign n4914 = n3095 & n22199;
assign n23939 = ~(n11782 ^ n5591);
assign n21857 = ~(n12685 ^ n11274);
assign n1253 = ~(n15271 ^ n5822);
assign n19332 = ~(n8732 | n15914);
assign n6534 = n7952 | n3952;
assign n19217 = ~(n16765 ^ n26999);
assign n17893 = n12215 & n4979;
assign n24800 = n5104 & n3997;
assign n16639 = n24676 & n19407;
assign n25712 = ~(n24026 ^ n5780);
assign n23733 = n4876 | n11819;
assign n4521 = n2428 | n4280;
assign n21646 = n17862 | n6063;
assign n17518 = ~(n17390 ^ n21247);
assign n24670 = n17993 | n23145;
assign n20540 = n24007 | n22028;
assign n332 = ~(n9953 ^ n9487);
assign n23257 = ~(n24745 ^ n3724);
assign n11413 = ~(n821 | n8856);
assign n129 = ~(n8856 ^ n22442);
assign n13437 = n4236 | n21476;
assign n12381 = ~n7946;
assign n11406 = n25910 & n13009;
assign n9940 = ~(n21962 ^ n13074);
assign n25944 = ~(n3337 ^ n709);
assign n12071 = n14736 & n3529;
assign n12635 = n9663 | n1526;
assign n15717 = ~(n3284 | n8003);
assign n16680 = ~(n20032 | n7149);
assign n11262 = ~(n26425 ^ n2151);
assign n10816 = ~(n9909 | n1694);
assign n12642 = ~(n5131 | n19674);
assign n23718 = ~(n12875 | n12652);
assign n23643 = ~(n16971 ^ n19144);
assign n21302 = ~(n16751 ^ n24021);
assign n27039 = ~(n13897 | n13159);
assign n10281 = ~n26645;
assign n22838 = n15375 | n22483;
assign n26883 = ~n3260;
assign n25205 = n17588 | n5155;
assign n16597 = ~(n9026 ^ n11273);
assign n9524 = n26411 | n3965;
assign n7994 = ~(n3976 | n16882);
assign n5466 = ~n2909;
assign n26781 = n20250 | n1682;
assign n1156 = ~(n26594 ^ n18880);
assign n2251 = ~(n1662 | n26962);
assign n8347 = ~(n4692 | n26023);
assign n19021 = n4412 | n22109;
assign n8588 = n19862 | n16223;
assign n13928 = ~(n21841 ^ n17994);
assign n16690 = ~(n5077 ^ n13851);
assign n16498 = n16374 | n23181;
assign n2980 = ~n17558;
assign n20282 = n18901 | n638;
assign n7900 = n7264 & n21515;
assign n17882 = ~(n25568 ^ n16880);
assign n9973 = n4229 & n26973;
assign n24260 = ~(n20937 ^ n7810);
assign n178 = n26271 | n25152;
assign n9663 = ~(n23487 | n26658);
assign n12685 = n21983 & n25557;
assign n8931 = ~n434;
assign n22547 = n6393 | n2028;
assign n22342 = ~n8660;
assign n10821 = ~n19312;
assign n3326 = ~(n13995 | n21981);
assign n25030 = n7541 & n20632;
assign n13643 = ~n3743;
assign n24142 = n5675 | n5424;
assign n25368 = ~n8933;
assign n3884 = ~(n12090 ^ n8487);
assign n826 = ~(n21095 ^ n11192);
assign n19658 = ~n26226;
assign n8120 = n5912 & n14990;
assign n5463 = n21190 & n18458;
assign n22847 = n17722 & n6792;
assign n9357 = n26367 | n8930;
assign n7159 = n21926 | n19468;
assign n13144 = ~(n18306 ^ n3726);
assign n26239 = ~(n5086 ^ n20670);
assign n10076 = ~(n21923 ^ n5637);
assign n18393 = ~n18944;
assign n9327 = n17828 & n11361;
assign n23079 = n20782 | n4702;
assign n24253 = n24772 | n24207;
assign n14311 = ~n11414;
assign n5268 = n15189 & n24320;
assign n4689 = n16636 | n20877;
assign n1435 = ~(n8732 ^ n14127);
assign n11799 = ~(n6356 ^ n4665);
assign n21072 = n2032 & n19782;
assign n2673 = n12857 | n1931;
assign n19216 = ~(n26298 ^ n26625);
assign n20525 = ~n9342;
assign n25584 = n619 & n14880;
assign n706 = ~(n10499 | n9512);
assign n22286 = n7437 & n26992;
assign n1030 = n20417 & n3568;
assign n14303 = n18738 | n9457;
assign n6818 = n17336 & n19812;
assign n7977 = n19012 & n25456;
assign n13679 = n19446 & n3931;
assign n13216 = ~(n9962 ^ n24028);
assign n6403 = ~(n7651 ^ n581);
assign n12955 = ~n7139;
assign n23288 = ~(n22351 | n24093);
assign n25091 = n1280 | n24787;
assign n14392 = n15009 | n12733;
assign n22070 = n10338 & n425;
assign n26794 = ~(n12231 ^ n26821);
assign n5319 = ~n6449;
assign n16081 = n25941 | n9269;
assign n17258 = n9869 | n16066;
assign n17280 = n16227 | n6513;
assign n9771 = ~(n22852 ^ n18229);
assign n23228 = ~(n26189 | n24180);
assign n4299 = ~n1917;
assign n15961 = ~(n21041 ^ n7838);
assign n25366 = n8429 & n16039;
assign n10373 = n15258 & n2420;
assign n21945 = ~(n20525 ^ n12806);
assign n26760 = ~(n5965 | n9200);
assign n7507 = ~(n16131 ^ n2922);
assign n21286 = n5539 & n23019;
assign n22398 = ~n21967;
assign n21908 = n13490 | n6333;
assign n9239 = ~(n9875 | n25562);
assign n15548 = ~(n11010 ^ n17183);
assign n20633 = ~(n12595 ^ n4682);
assign n22720 = n14809 | n21736;
assign n14525 = n18496 & n20201;
assign n13053 = ~n7919;
assign n24684 = ~(n12193 ^ n10174);
assign n1425 = n3499 | n14315;
assign n4904 = ~(n16476 | n15539);
assign n8862 = ~(n22277 ^ n3628);
assign n6050 = n24417 | n10027;
assign n22041 = n7130 | n3075;
assign n23590 = n1329 | n5512;
assign n22022 = n17736 & n15951;
assign n10300 = n7355 & n18273;
assign n20256 = n329 | n6541;
assign n10801 = n23478 | n12684;
assign n14920 = ~(n11452 | n23068);
assign n13286 = ~n6299;
assign n21492 = n16750 | n9015;
assign n4005 = ~(n2009 ^ n7767);
assign n14154 = ~(n13206 ^ n17035);
assign n5930 = n20742 & n26861;
assign n22585 = ~n17090;
assign n7717 = n7283 & n24915;
assign n25821 = n14366 | n8477;
assign n24439 = ~(n23819 ^ n22861);
assign n22900 = n773 | n12798;
assign n24979 = ~(n7657 ^ n25316);
assign n7319 = ~n8526;
assign n1582 = n13210 & n14890;
assign n8554 = n18552 & n1315;
assign n24424 = n18424 | n3837;
assign n21805 = n9793 | n22361;
assign n6132 = n17339 ^ n6502;
assign n15127 = ~(n14903 ^ n9302);
assign n20226 = n2766 | n18248;
assign n19310 = ~(n10201 | n24043);
assign n18741 = ~n15865;
assign n19453 = ~n24171;
assign n6998 = ~(n14906 ^ n23565);
assign n20571 = n23722 | n5324;
assign n12129 = ~(n14902 | n4288);
assign n19231 = n26027 | n19198;
assign n14097 = ~(n2035 ^ n12821);
assign n11365 = ~n14749;
assign n13736 = ~(n5629 ^ n7377);
assign n4671 = n20429 | n22909;
assign n24455 = ~n25653;
assign n6152 = ~(n15769 ^ n13190);
assign n23998 = n8820 | n13197;
assign n5918 = ~n13951;
assign n21618 = n18776 | n1770;
assign n12554 = ~n16396;
assign n24016 = ~(n6068 ^ n18745);
assign n20125 = ~n10204;
assign n12155 = n9816 & n11;
assign n8058 = n25283 | n13193;
assign n18604 = n19949 | n11285;
assign n25208 = ~(n10079 ^ n1820);
assign n14732 = n19133 & n19014;
assign n6028 = ~n25302;
assign n8479 = n15636 | n9656;
assign n802 = n20089 | n5998;
assign n24290 = ~(n26875 | n5530);
assign n9907 = n5149 | n26703;
assign n21991 = n24282 | n23712;
assign n20538 = ~n1530;
assign n24991 = n26213 & n24773;
assign n714 = n14870 | n8888;
assign n27030 = ~n22388;
assign n16087 = n24338 | n20110;
assign n23936 = ~n5818;
assign n5045 = ~n21427;
assign n6155 = ~(n20338 ^ n9531);
assign n22230 = ~n23763;
assign n21617 = n18073 | n6767;
assign n8246 = ~(n19940 ^ n14705);
assign n26996 = n18921 | n1028;
assign n26780 = ~(n8752 ^ n23796);
assign n2204 = ~n24225;
assign n26686 = n22597 | n16473;
assign n8685 = ~(n11503 ^ n18151);
assign n20583 = n14431 & n22587;
assign n11809 = n22590 & n19053;
assign n25818 = ~n17591;
assign n3897 = ~(n1336 ^ n6265);
assign n17557 = ~(n12042 ^ n11514);
assign n548 = ~(n15067 ^ n11079);
assign n13930 = n1252 & n23427;
assign n12339 = n8048 & n13942;
assign n12490 = n20737 | n20036;
assign n26679 = n26532 | n526;
assign n21968 = ~(n15787 ^ n11408);
assign n3708 = ~(n18584 ^ n19803);
assign n11388 = n4665 | n24278;
assign n5725 = n15840 | n8364;
assign n21244 = ~(n8779 ^ n18290);
assign n11957 = ~(n12639 | n26986);
assign n24842 = ~(n19983 ^ n18433);
assign n22632 = ~(n21517 ^ n8582);
assign n8267 = ~(n26040 ^ n17228);
assign n17827 = ~(n26536 ^ n4603);
assign n13597 = n22337 & n19290;
assign n3595 = ~(n7829 ^ n12593);
assign n17491 = n26007 | n15126;
assign n18050 = ~(n26870 ^ n25864);
assign n5249 = n21760 | n11589;
assign n19804 = ~(n18590 ^ n25225);
assign n22526 = n16730 | n11066;
assign n7019 = n173 | n18008;
assign n10109 = ~n11630;
assign n19779 = n26398 & n17886;
assign n10951 = ~n1200;
assign n16695 = n2235 & n3556;
assign n2535 = ~(n6384 ^ n21788);
assign n20717 = ~(n14777 | n3236);
assign n21194 = ~n12430;
assign n23283 = ~(n12709 | n19989);
assign n17296 = n17995 & n4222;
assign n9201 = n21186 & n2215;
assign n8971 = ~(n20656 ^ n9845);
assign n23925 = n17414 | n19478;
assign n25731 = ~(n16468 ^ n17351);
assign n20311 = ~(n14139 | n14838);
assign n3753 = ~(n8068 | n1128);
assign n10927 = ~(n23383 ^ n771);
assign n23664 = ~n2249;
assign n5678 = ~n15245;
assign n21641 = n9557 | n16158;
assign n23132 = n16268 & n1647;
assign n16159 = n11745 & n18249;
assign n4966 = ~(n19101 ^ n11797);
assign n2788 = ~(n15808 ^ n16713);
assign n17868 = n27190 | n2531;
assign n7955 = n18960 | n14982;
assign n9254 = n11016 & n9883;
assign n24255 = n11089 | n972;
assign n21911 = ~(n24509 ^ n18065);
assign n1201 = n9652 & n901;
assign n3536 = n23497 & n22413;
assign n2219 = ~n1536;
assign n10343 = ~n24992;
assign n21304 = n18097 & n20354;
assign n22321 = ~(n7800 ^ n5626);
assign n20647 = ~(n1654 ^ n21997);
assign n7021 = n14613 | n6777;
assign n5379 = n22851 | n17610;
assign n20887 = n22019 & n13064;
assign n27103 = n10769 & n1174;
assign n17168 = ~(n9348 ^ n24712);
assign n20301 = ~(n7806 ^ n19933);
assign n1173 = ~n14044;
assign n15876 = n23894 | n4851;
assign n10386 = ~(n27114 ^ n4569);
assign n3501 = n2459 | n24838;
assign n15450 = n4971 & n9306;
assign n167 = ~n10392;
assign n8546 = ~(n17664 | n21253);
assign n8337 = n7841 | n8952;
assign n20219 = ~(n24746 ^ n4119);
assign n5904 = ~(n2800 ^ n8584);
assign n25003 = n25903 | n20697;
assign n9234 = n6726 & n18202;
assign n21692 = n25308 & n17777;
assign n10813 = n14928 & n1614;
assign n6543 = ~(n16539 ^ n15362);
assign n8074 = n5898 | n24182;
assign n18742 = ~n19117;
assign n5524 = ~(n9674 ^ n24585);
assign n2854 = n15068 & n5630;
assign n23134 = n26984 & n24720;
assign n6719 = n5016 | n12839;
assign n22873 = n13593 | n13845;
assign n25 = n11919 | n19037;
assign n8021 = n15768 & n16592;
assign n11035 = n2713 | n20479;
assign n8944 = ~(n19825 ^ n10117);
assign n25727 = n20511 & n11272;
assign n1305 = n15162 | n19936;
assign n14898 = n20498 | n15486;
assign n24932 = ~(n20280 ^ n515);
assign n6289 = ~(n13596 ^ n7805);
assign n3330 = ~(n23822 ^ n1637);
assign n19108 = ~(n6053 ^ n1907);
assign n23317 = ~n25178;
assign n4899 = n5451 | n17858;
assign n25374 = n21708 | n13604;
assign n24313 = n26986 & n12639;
assign n7552 = n25121 | n14161;
assign n22251 = ~(n9135 ^ n27147);
assign n10509 = ~n17115;
assign n20413 = ~(n11979 ^ n6822);
assign n15443 = n3996 | n20916;
assign n22551 = n5941 & n7964;
assign n9017 = ~n15821;
assign n20419 = n1768 | n19069;
assign n18755 = ~n17343;
assign n827 = ~(n11151 ^ n4295);
assign n9513 = ~(n8264 ^ n15765);
assign n26597 = n11743 & n13301;
assign n18783 = n12175 | n12949;
assign n10099 = n4857 | n7193;
assign n18365 = n15824 & n18490;
assign n5723 = n6498 | n20906;
assign n20449 = n23549 & n764;
assign n26598 = ~(n9743 ^ n17806);
assign n25847 = n3589 | n18223;
assign n3899 = n5466 | n10821;
assign n10338 = n8991 | n20755;
assign n11766 = n2579 | n3468;
assign n25131 = ~(n22631 ^ n2117);
assign n11399 = n6602 & n24465;
assign n4889 = n14963 | n3570;
assign n26546 = ~(n2028 ^ n17853);
assign n23788 = n22554 & n1414;
assign n8359 = n3204 | n12626;
assign n25025 = ~(n19042 | n19360);
assign n17206 = ~(n8266 ^ n13495);
assign n23999 = ~(n17634 ^ n8687);
assign n7719 = ~(n9957 ^ n2659);
assign n23509 = ~(n11895 ^ n5451);
assign n17540 = n13384 | n4459;
assign n1360 = ~(n24473 | n3614);
assign n6899 = n10 | n23407;
assign n11761 = n528 | n13627;
assign n13030 = n15369 | n12580;
assign n21926 = n7722 & n154;
assign n1237 = ~(n3938 ^ n6481);
assign n20333 = ~(n8377 ^ n13155);
assign n6708 = ~n25807;
assign n24006 = n18425 | n7970;
assign n21366 = n2026 & n14906;
assign n17039 = n25904 & n20657;
assign n1919 = n5594 & n15708;
assign n4952 = n10736 | n4663;
assign n15393 = ~(n11151 ^ n21489);
assign n8072 = ~(n10622 ^ n265);
assign n14107 = ~(n9979 ^ n15805);
assign n1789 = n15660 | n24814;
assign n2372 = n2454 & n4970;
assign n9812 = ~(n2804 | n18129);
assign n602 = ~n1138;
assign n3643 = ~(n20089 ^ n16502);
assign n9038 = n860 | n14330;
assign n6102 = n2278 & n7093;
assign n23995 = ~n25689;
assign n5437 = ~(n7693 | n19472);
assign n24624 = ~n2525;
assign n19495 = ~(n20604 ^ n21735);
assign n23744 = ~(n2816 | n26486);
assign n16064 = ~n25520;
assign n6408 = ~(n2562 | n8244);
assign n20483 = ~(n21400 ^ n19081);
assign n7745 = ~n22495;
assign n3976 = ~(n23975 ^ n16645);
assign n18479 = n9655 | n21908;
assign n14740 = ~(n6613 | n6703);
assign n13729 = ~n9172;
assign n23972 = n16836 & n10798;
assign n11670 = ~(n26352 ^ n22679);
assign n20651 = ~(n26962 ^ n3730);
assign n1583 = n12354 | n19321;
assign n23461 = n19139 | n211;
assign n12082 = n11038 & n10058;
assign n17923 = ~n26291;
assign n22691 = ~(n10451 ^ n17741);
assign n2425 = n13783 | n26394;
assign n1929 = ~(n19476 | n2325);
assign n21527 = ~(n20899 ^ n11960);
assign n16139 = n18981 | n11381;
assign n22372 = ~(n9569 ^ n21317);
assign n4364 = n13307 & n14784;
assign n24793 = ~(n24990 ^ n19502);
assign n4192 = n21841 | n16295;
assign n16189 = n23436 | n9003;
assign n5541 = ~(n21764 ^ n23529);
assign n18383 = ~n6861;
assign n17317 = ~(n13108 ^ n11174);
assign n3219 = ~(n23396 ^ n1121);
assign n14772 = ~(n19879 ^ n2282);
assign n11656 = n7948 & n1583;
assign n17982 = ~(n1967 ^ n26989);
assign n23560 = ~(n24116 | n20929);
assign n2028 = n19082 | n24630;
assign n20405 = n4242 & n17388;
assign n24635 = n1365 | n25924;
assign n3450 = n15905 | n2510;
assign n25660 = ~(n24902 ^ n8623);
assign n26388 = n23539 | n14488;
assign n12957 = n7722 | n154;
assign n2696 = ~(n15605 ^ n22575);
assign n12239 = ~n13734;
assign n3938 = n4142 & n19504;
assign n19886 = ~(n10615 ^ n6078);
assign n22148 = n23216 | n15093;
assign n26428 = ~(n1181 | n11428);
assign n14612 = ~n1949;
assign n24180 = ~n8358;
assign n15141 = n26372 & n8080;
assign n14796 = ~(n2218 ^ n18483);
assign n6996 = ~(n11869 ^ n20198);
assign n2803 = n4258 | n25922;
assign n14522 = n26858 & n17327;
assign n20474 = ~(n25972 | n21378);
assign n23119 = ~(n14744 | n17936);
assign n1094 = n16625 | n15032;
assign n23080 = n15595 & n20781;
assign n26514 = ~(n4040 | n3349);
assign n21225 = ~(n16122 ^ n4115);
assign n8670 = n20622 & n25880;
assign n15726 = n1588 & n22229;
assign n12280 = n20613 | n14138;
assign n7286 = ~(n1406 | n4940);
assign n2432 = ~n10116;
assign n8252 = ~(n18290 | n25160);
assign n3765 = n11187 | n547;
assign n422 = ~(n651 ^ n11845);
assign n27203 = n866 | n9449;
assign n1065 = n14420 & n15664;
assign n1533 = ~n8724;
assign n15134 = ~(n9679 | n22442);
assign n88 = ~n25164;
assign n248 = ~(n20569 ^ n14120);
assign n18530 = n7566 & n22640;
assign n18820 = ~(n19946 ^ n12627);
assign n23351 = ~(n15058 | n1532);
assign n6461 = n603 & n16505;
assign n4977 = ~(n4003 | n22507);
assign n14531 = ~(n2242 ^ n12810);
assign n2672 = n16575 | n2379;
assign n12667 = ~(n19090 ^ n20271);
assign n26580 = ~n21540;
assign n9085 = ~(n3228 ^ n22470);
assign n3432 = n17014 | n17646;
assign n26637 = n20318 & n13345;
assign n3587 = ~n24399;
assign n7913 = ~(n19234 ^ n21398);
assign n12359 = n19731 & n23993;
assign n13217 = ~(n4708 ^ n19216);
assign n20099 = ~n9219;
assign n24845 = ~(n12481 | n9227);
assign n11485 = ~n26708;
assign n6261 = n22919 | n23044;
assign n742 = ~(n25465 ^ n26530);
assign n14269 = ~n2969;
assign n20743 = n4854 & n23862;
assign n16495 = n4574 | n25715;
assign n16103 = ~(n18995 | n17143);
assign n13122 = ~(n7483 ^ n10774);
assign n20922 = n13154 | n3918;
assign n24317 = n8352 | n22960;
assign n15598 = ~(n18547 ^ n26504);
assign n6103 = n5122 | n6483;
assign n881 = ~(n8814 ^ n21158);
assign n20123 = n5924 | n16201;
assign n7217 = n18300 & n9411;
assign n5851 = ~(n17626 ^ n2246);
assign n8375 = ~(n10152 ^ n7981);
assign n5352 = n5025 | n23162;
assign n11959 = n6908 & n9098;
assign n4208 = ~(n25036 | n11016);
assign n21169 = n417 | n4499;
assign n14825 = n13367 | n13074;
assign n6329 = ~(n6492 ^ n20835);
assign n26964 = ~(n6827 ^ n6055);
assign n24934 = ~(n25340 ^ n76);
assign n18512 = ~(n1505 ^ n26036);
assign n17993 = ~(n19182 ^ n22563);
assign n4184 = ~(n10784 ^ n6881);
assign n14312 = n10985 | n24122;
assign n13542 = n13224 | n21089;
assign n1568 = ~(n24355 | n1267);
assign n18415 = n11315 | n24918;
assign n21203 = ~(n25060 ^ n14832);
assign n2033 = n13184 | n13962;
assign n1552 = ~(n7442 ^ n8767);
assign n20680 = ~(n8987 | n14245);
assign n4938 = ~n23463;
assign n12754 = ~(n7073 ^ n13010);
assign n5742 = ~(n15329 ^ n13135);
assign n25469 = n6877 | n9108;
assign n11190 = n19732 | n14296;
assign n1820 = ~(n1163 ^ n18901);
assign n15711 = ~(n15905 | n23168);
assign n17219 = ~(n25148 ^ n21521);
assign n322 = n21083 | n7520;
assign n6783 = ~(n9485 ^ n12147);
assign n11620 = n16056 | n13540;
assign n3311 = ~(n413 ^ n5409);
assign n8421 = n14306 | n2599;
assign n24195 = n12582 | n6681;
assign n14595 = n23141 | n22981;
assign n8946 = ~(n8399 ^ n8052);
assign n17660 = ~n1512;
assign n868 = ~n4775;
assign n5286 = ~(n20040 ^ n9396);
assign n13963 = ~(n25558 ^ n18904);
assign n1518 = ~(n18127 ^ n2402);
assign n13989 = ~n19494;
assign n76 = ~(n15447 ^ n6838);
assign n4204 = ~(n3926 ^ n492);
assign n25308 = n19383 | n10422;
assign n24704 = ~(n1485 ^ n24518);
assign n18189 = ~n4626;
assign n15368 = ~(n18419 | n22005);
assign n13124 = ~n16392;
assign n7210 = ~(n17156 ^ n4872);
assign n21421 = ~(n19634 | n2731);
assign n710 = ~(n17894 ^ n1982);
assign n17707 = n18649 | n11278;
assign n6924 = ~(n15731 ^ n12300);
assign n8095 = n10002 | n21861;
assign n8933 = ~(n19120 ^ n16027);
assign n25539 = ~(n15755 ^ n14468);
assign n16838 = n4709 | n16088;
assign n21528 = n18926 | n2705;
assign n24774 = ~n2059;
assign n18402 = n6007 & n24641;
assign n26281 = n25190 | n24281;
assign n7227 = n18415 & n19369;
assign n16165 = n11486 | n13781;
assign n24286 = n14083;
assign n21684 = n24670 & n2182;
assign n21107 = ~n9274;
assign n25317 = n337 | n5340;
assign n8331 = ~(n11661 ^ n324);
assign n2260 = n23537 & n11010;
assign n2373 = n22487 | n13645;
assign n11525 = ~(n11608 ^ n17693);
assign n18544 = ~(n21276 ^ n18157);
assign n19312 = ~(n17659 ^ n3833);
assign n23672 = n24845 | n9641;
assign n3563 = ~(n14235 ^ n9796);
assign n20620 = ~n3830;
assign n20294 = n23320 | n19564;
assign n20920 = n18953;
assign n13353 = ~n5834;
assign n7921 = ~(n14612 | n20169);
assign n5225 = n10395 & n15476;
assign n25951 = n22994 | n9025;
assign n9780 = ~n9749;
assign n15090 = ~(n19023 ^ n8330);
assign n22090 = ~(n188 ^ n25551);
assign n7448 = ~n13257;
assign n12175 = n22820 & n19137;
assign n5871 = n4544 | n23701;
assign n21502 = ~(n8287 ^ n12483);
assign n19432 = ~(n5318 ^ n3943);
assign n12537 = n12673 | n21529;
assign n573 = n21701 | n21547;
assign n9980 = ~(n4570 ^ n17458);
assign n11577 = ~n18729;
assign n13382 = n8068 | n11192;
assign n6808 = n10575 & n7246;
assign n16943 = n6859 & n17600;
assign n17818 = n17675 & n26412;
assign n19983 = n26976 & n22947;
assign n1627 = n5883 | n20764;
assign n15093 = ~(n1787 ^ n10618);
assign n6320 = ~(n12204 | n22478);
assign n23425 = ~(n14967 | n20013);
assign n15035 = n23464 | n25966;
assign n26847 = ~(n5676 ^ n22381);
assign n17158 = n22749 | n5468;
assign n11530 = n6051 | n593;
assign n18528 = n5349 & n3990;
assign n19194 = ~n25383;
assign n20711 = n13898 & n7311;
assign n12083 = n11941 | n1890;
assign n24108 = n888 | n25977;
assign n15525 = n23631 | n24935;
assign n15205 = ~(n16686 ^ n14047);
assign n2871 = n832 | n11938;
assign n14969 = ~n6891;
assign n722 = ~(n3045 ^ n4201);
assign n6089 = ~n9168;
assign n18014 = ~(n19085 | n24592);
assign n3023 = n113 | n2604;
assign n3101 = n7046 & n7853;
assign n9331 = n10646 & n12106;
assign n26410 = n20237 & n13111;
assign n9544 = n1427 | n25497;
assign n18089 = ~(n9942 ^ n10739);
assign n6063 = ~n2443;
assign n224 = ~(n1928 ^ n21256);
assign n9560 = n14710 | n2219;
assign n4337 = n23852 | n17430;
assign n26895 = ~n6794;
assign n24303 = n6813 | n14347;
assign n20101 = n5727 | n3477;
assign n22340 = ~(n5681 ^ n9461);
assign n9194 = ~(n11099 ^ n915);
assign n23888 = ~(n4147 ^ n6700);
assign n18717 = ~(n2155 | n7097);
assign n14106 = ~(n19772 ^ n2571);
assign n20739 = n18749 | n4156;
assign n12830 = n15447 | n24951;
assign n14136 = ~(n16198 ^ n8184);
assign n5546 = n16534 | n5070;
assign n6118 = n26052 | n8054;
assign n12689 = n26555 & n18795;
assign n25892 = ~(n22260 ^ n10964);
assign n23728 = ~(n6502 | n19494);
assign n25107 = n9894 & n14793;
assign n7243 = n10247 & n14253;
assign n18013 = n6369 & n527;
assign n22823 = n7377 | n21125;
assign n20341 = n4502 | n25536;
assign n13078 = n4022 | n13110;
assign n20175 = ~n4122;
assign n21533 = ~(n6713 ^ n14528);
assign n7816 = n22996 & n163;
assign n11400 = n6239 | n25685;
assign n3262 = n13223 | n5545;
assign n13609 = n27157 & n16802;
assign n9810 = n20466 | n23323;
assign n26542 = n10743 | n26584;
assign n24463 = n4727 | n11207;
assign n21173 = ~(n12721 ^ n24095);
assign n24258 = ~(n2317 ^ n25385);
assign n8417 = ~(n17146 ^ n12207);
assign n26714 = n24240 & n4406;
assign n25975 = n6735 & n6045;
assign n19929 = n3074 | n2220;
assign n13911 = n26481 & n16976;
assign n20070 = ~(n2187 | n9572);
assign n14102 = ~(n90 ^ n23994);
assign n2807 = ~(n305 | n2610);
assign n8601 = n18742 | n14319;
assign n24289 = ~(n25039 ^ n5279);
assign n18395 = ~(n11197 ^ n17766);
assign n26154 = n22985 & n3156;
assign n10463 = n23216 & n15093;
assign n4221 = ~(n3774 ^ n7754);
assign n6043 = ~(n13322 ^ n18698);
assign n27205 = n23091 | n18735;
assign n4733 = n13452 & n9743;
assign n10486 = ~n6279;
assign n947 = ~(n11628 ^ n17325);
assign n2761 = ~(n21452 ^ n9467);
assign n4497 = ~n10185;
assign n24393 = ~(n1380 ^ n3324);
assign n7858 = n7003 | n2480;
assign n5612 = ~(n1346 | n442);
assign n21199 = n12178 | n7116;
assign n11972 = n6154 | n23996;
assign n9948 = ~(n25265 | n23773);
assign n12597 = n25331 | n2189;
assign n24343 = ~n26733;
assign n1829 = ~(n18855 | n20925);
assign n10277 = ~n18006;
assign n23226 = n22176 | n120;
assign n2275 = ~(n21520 ^ n19615);
assign n19330 = n8305 & n2918;
assign n19656 = n23306 | n9201;
assign n20956 = ~(n27008 | n21194);
assign n10748 = n20200 | n9156;
assign n2223 = ~n881;
assign n26671 = n15842 | n12606;
assign n25882 = ~(n3018 | n2731);
assign n24815 = ~n14380;
assign n26620 = ~(n6385 ^ n18171);
assign n25202 = ~(n14596 ^ n23635);
assign n3118 = ~(n520 ^ n6593);
assign n2919 = ~n25355;
assign n773 = ~(n23095 | n1112);
assign n2139 = n26318 | n15860;
assign n7938 = ~n22378;
assign n24502 = n4113 | n21278;
assign n8863 = ~(n12878 ^ n14539);
assign n10157 = ~n19335;
assign n2320 = ~(n17695 ^ n7692);
assign n2491 = ~(n23098 ^ n4434);
assign n21501 = n17035 | n1872;
assign n18164 = n9539 | n12255;
assign n1579 = n20912 & n2245;
assign n5737 = ~(n9621 ^ n17367);
assign n606 = n14242 & n12595;
assign n21770 = n14529 & n9477;
assign n22400 = ~(n25073 ^ n12152);
assign n13812 = ~(n12232 ^ n3740);
assign n10948 = ~n16945;
assign n9984 = ~(n4469 ^ n960);
assign n25141 = n20890 & n24952;
assign n17415 = ~(n20797 ^ n2978);
assign n20529 = n18278 & n19932;
assign n12357 = ~(n1639 ^ n5128);
assign n16965 = ~(n5450 ^ n5469);
assign n3048 = n18026 & n6188;
assign n21810 = n8440 & n2304;
assign n3029 = ~(n2698 | n16961);
assign n8174 = ~(n12612 ^ n20794);
assign n21324 = ~(n24751 ^ n8604);
assign n12660 = ~(n6812 ^ n2614);
assign n26639 = ~(n7331 ^ n12171);
assign n10139 = ~(n21322 ^ n25345);
assign n4525 = n7378 | n634;
assign n6661 = ~(n2926 ^ n12586);
assign n6357 = ~n24788;
assign n17451 = n9832 | n11831;
assign n7941 = ~(n8813 | n10770);
assign n1676 = n7590 | n16413;
assign n10830 = n22257 | n22287;
assign n5245 = n17188 | n24408;
assign n14711 = n48 | n1309;
assign n1200 = ~(n24323 ^ n6775);
assign n22508 = ~(n2976 ^ n13262);
assign n8447 = ~(n17718 | n7020);
assign n4611 = n418 & n16726;
assign n15847 = ~(n10116 | n15017);
assign n4151 = ~(n19994 ^ n6329);
assign n6224 = n26469 | n3867;
assign n14592 = n12261 | n22221;
assign n14530 = n544 | n8170;
assign n17437 = n12759 & n18156;
assign n22676 = n8875 | n259;
assign n14121 = ~(n13272 ^ n25346);
assign n10677 = ~(n20369 | n19034);
assign n9597 = ~n7241;
assign n6079 = ~n19660;
assign n4361 = ~n6335;
assign n5139 = ~(n19273 ^ n18347);
assign n540 = ~(n17679 | n8414);
assign n14291 = n288 | n2144;
assign n1441 = n6510 | n20482;
assign n14653 = n26895 | n6611;
assign n17 = n6274 & n3277;
assign n1390 = n6892 | n14428;
assign n12021 = ~(n3241 | n13944);
assign n12690 = n5553 | n18716;
assign n26237 = ~(n20762 ^ n2468);
assign n11872 = n17698 & n10450;
assign n9579 = n18056 | n2474;
assign n4974 = n18794 & n16038;
assign n16294 = ~n11220;
assign n18208 = ~(n6385 ^ n8869);
assign n15244 = ~(n17664 | n7532);
assign n27056 = n6061 | n12685;
assign n14480 = ~(n2538 ^ n19857);
assign n7109 = ~(n25779 | n26161);
assign n13205 = ~n10792;
assign n3655 = n11481 | n23493;
assign n9134 = n5149 & n26703;
assign n27077 = n3784 | n13121;
assign n25286 = n6485 | n18676;
assign n4305 = n3519 | n7687;
assign n403 = n6811 | n10860;
assign n24809 = n3213 & n8143;
assign n22226 = n10568 & n5848;
assign n22661 = n27000 & n6292;
assign n18408 = ~(n10324 | n9779);
assign n2377 = ~n25204;
assign n19870 = n13629 | n3693;
assign n4258 = n4086 & n1533;
assign n22060 = n21857 | n10861;
assign n13022 = ~(n7969 ^ n21827);
assign n21731 = ~(n21113 ^ n16019);
assign n13390 = ~(n25376 | n1752);
assign n12048 = ~n2055;
assign n15089 = n7360 | n18598;
assign n9709 = ~(n2586 ^ n11743);
assign n22227 = ~n2244;
assign n5144 = ~(n26703 | n7615);
assign n25935 = n15018 & n8426;
assign n4597 = n11200 & n8723;
assign n8567 = ~(n4301 | n16330);
assign n694 = n22958 | n19157;
assign n1852 = n24811 & n11500;
assign n15820 = ~(n10351 ^ n26318);
assign n201 = n5467 & n19110;
assign n16902 = ~(n24952 ^ n22371);
assign n22378 = ~(n26166 ^ n4124);
assign n9025 = n13254 & n24570;
assign n1786 = ~n9605;
assign n8608 = ~(n17340 ^ n15303);
assign n16635 = ~(n19610 | n18539);
assign n8725 = ~(n1577 ^ n14405);
assign n20577 = n17789 | n15337;
assign n19258 = ~n8943;
assign n25116 = n8301 | n20449;
assign n5568 = ~(n24850 ^ n22706);
assign n2585 = ~(n3740 | n2545);
assign n23280 = n16628 & n7028;
assign n8771 = ~n10104;
assign n16262 = ~(n20289 ^ n9300);
assign n8426 = n14479 | n17060;
assign n26601 = ~n13471;
assign n23423 = ~(n17483 ^ n18504);
assign n24104 = n26494 & n365;
assign n1548 = n22443 | n23938;
assign n22864 = n5084 | n8011;
assign n4734 = ~(n22350 ^ n2747);
assign n20974 = n12932 | n22370;
assign n6372 = n6724 | n11329;
assign n3606 = ~(n4074 ^ n15593);
assign n5973 = n3487 & n20889;
assign n11256 = ~(n22723 | n20923);
assign n26157 = n25721 | n24067;
assign n17192 = ~(n18909 | n18203);
assign n13891 = n576 & n13969;
assign n5305 = n2840 & n19079;
assign n8088 = ~(n13046 ^ n15216);
assign n3858 = n13659 | n14932;
assign n14777 = ~n22079;
assign n2295 = ~(n24403 ^ n26768);
assign n7058 = ~n24860;
assign n26741 = ~(n290 ^ n24086);
assign n497 = n7242 ^ n3311;
assign n18138 = n17120 | n7751;
assign n5003 = n446 | n25318;
assign n2929 = ~(n929 ^ n1376);
assign n21381 = n1407 & n7655;
assign n8898 = ~(n14417 ^ n3054);
assign n23396 = n8931 | n24809;
assign n6342 = ~(n12068 ^ n18535);
assign n8519 = ~(n4508 ^ n5357);
assign n3081 = n14080 | n24494;
assign n10782 = n22081 & n21382;
assign n8539 = ~n21073;
assign n4836 = ~(n11985 ^ n18116);
assign n5296 = ~(n14348 ^ n22393);
assign n15321 = n963 | n13071;
assign n23855 = ~(n1844 ^ n21300);
assign n10692 = ~(n9891 ^ n14461);
assign n1967 = n26895 | n5512;
assign n9859 = ~n22325;
assign n6022 = ~(n4488 ^ n15803);
assign n2063 = ~(n6685 | n19971);
assign n12345 = ~n16150;
assign n15367 = n25099 | n4442;
assign n9782 = ~(n12161 | n106);
assign n5955 = n11424 & n12692;
assign n6135 = ~(n14045 ^ n9936);
assign n8541 = n18008 | n17869;
assign n7350 = ~n1910;
assign n17651 = ~(n1837 ^ n9961);
assign n26102 = ~(n26997 ^ n19059);
assign n7863 = n25747 & n17661;
assign n20865 = ~(n20284 | n3779);
assign n16466 = ~n19845;
assign n27073 = n10604 & n17424;
assign n21157 = ~(n12711 ^ n3436);
assign n11377 = n10164 ^ n12983;
assign n3802 = n8556 & n18259;
assign n20096 = ~(n22614 ^ n8234);
assign n21611 = n580 | n3053;
assign n19992 = n3150 | n24929;
assign n24972 = ~(n21112 ^ n8309);
assign n10323 = ~(n14695 | n10125);
assign n9873 = ~(n508 ^ n12518);
assign n1322 = n8101 & n21912;
assign n23401 = ~(n5118 ^ n25944);
assign n3625 = ~n19478;
assign n16934 = n19440 & n27198;
assign n13564 = n8851 & n15212;
assign n16926 = n10097 | n18002;
assign n17417 = ~(n21912 ^ n15241);
assign n9211 = n18136 & n24976;
assign n5412 = n4919 & n17222;
assign n5021 = n24383 | n6403;
assign n2478 = ~(n1777 ^ n21832);
assign n383 = n14930 | n4002;
assign n11395 = ~(n17295 ^ n14289);
assign n24239 = ~n6095;
assign n22562 = ~n9986;
assign n16216 = ~(n5112 | n5417);
assign n12617 = ~(n20365 ^ n22571);
assign n7886 = n19110 ^ n2470;
assign n10852 = n22123 | n82;
assign n24214 = n1338 & n27180;
assign n8028 = ~(n21291 ^ n218);
assign n8189 = n4514 | n5111;
assign n6294 = n5558 | n23280;
assign n24226 = ~(n19871 ^ n25996);
assign n6771 = n5499 | n17773;
assign n13247 = ~(n25074 ^ n10053);
assign n7561 = ~n48;
assign n23874 = ~(n1817 ^ n159);
assign n26789 = ~(n14317 ^ n25797);
assign n8868 = ~(n4699 | n16946);
assign n17286 = ~n24768;
assign n12316 = n596 & n22790;
assign n22326 = ~(n25855 ^ n26461);
assign n8649 = ~(n8652 ^ n16973);
assign n26968 = ~(n20794 ^ n23333);
assign n25433 = n102 | n15192;
assign n7012 = n21134 & n4930;
assign n6235 = ~n7100;
assign n26349 = n4942 | n13147;
assign n3946 = ~n1714;
assign n22074 = n6218 & n9296;
assign n895 = n14519 | n3164;
assign n10547 = ~(n9942 ^ n23923);
assign n19444 = ~n23258;
assign n25405 = ~n25251;
assign n24122 = n4655 & n16629;
assign n8982 = ~(n21657 ^ n22241);
assign n9082 = n8032 | n14394;
assign n23523 = n8667 & n16977;
assign n22500 = n2997 | n6445;
assign n24859 = ~(n17090 ^ n22173);
assign n15851 = n10641 & n3469;
assign n15486 = n158 & n21053;
assign n18315 = ~(n9557 ^ n24170);
assign n16089 = n16606 & n5896;
assign n10665 = ~(n22274 ^ n22591);
assign n11892 = n16147 | n11367;
assign n18103 = ~n7249;
assign n4223 = n6734 & n3;
assign n19003 = ~n6082;
assign n3485 = ~n450;
assign n4215 = ~(n18930 ^ n9126);
assign n14946 = ~(n6492 ^ n17718);
assign n13621 = ~(n13252 ^ n9463);
assign n25841 = n20425 & n12332;
assign n19526 = n14724 & n9555;
assign n25832 = n12014 | n1222;
assign n15173 = n21261 & n18204;
assign n19751 = ~(n2876 ^ n19193);
assign n18619 = ~(n11670 ^ n16439);
assign n15346 = n24624 ^ n21095;
assign n22176 = ~n6773;
assign n6254 = ~(n4065 ^ n7479);
assign n20224 = n20470 & n14052;
assign n6894 = ~(n7311 ^ n13781);
assign n22203 = ~(n22619 ^ n6775);
assign n16012 = n528 & n17556;
assign n927 = n1319 | n3448;
assign n3705 = n14091 | n6693;
assign n19527 = ~n24049;
assign n21842 = ~n10392;
assign n6133 = ~(n23486 ^ n16663);
assign n3473 = ~(n15883 | n11096);
assign n9091 = n12508 & n25942;
assign n17834 = n22290 | n12562;
assign n14437 = ~(n23447 ^ n11225);
assign n2284 = n20503 & n5153;
assign n17614 = n21954 & n21548;
assign n5875 = ~n15119;
assign n11108 = ~(n8436 ^ n16167);
assign n22928 = ~(n8381 ^ n18295);
assign n16129 = ~n20040;
assign n21878 = n24780 & n16134;
assign n26142 = n18035 | n92;
assign n2116 = ~(n7892 ^ n15734);
assign n3811 = ~(n26508 | n61);
assign n21437 = n12657 & n10092;
assign n16014 = n10124 | n18734;
assign n15066 = ~(n26093 | n5745);
assign n12285 = n24594 & n15912;
assign n5641 = n20489 & n21693;
assign n10512 = n12962 & n26662;
assign n10526 = n26790 | n13366;
assign n12526 = ~(n1299 | n19411);
assign n3021 = n21102 & n8005;
assign n14627 = ~(n16294 | n12507);
assign n25369 = ~(n15580 | n9050);
assign n9437 = n5249 & n9516;
assign n9556 = ~(n15688 ^ n11169);
assign n4946 = n25639 | n12648;
assign n9585 = n4582 | n19993;
assign n10344 = n18186 & n1664;
assign n6279 = ~(n12382 ^ n26754);
assign n19154 = n14726 & n18695;
assign n1968 = n27188 | n8890;
assign n6484 = ~(n2585 | n7179);
assign n16950 = n1775 | n21170;
assign n1539 = ~(n11159 ^ n9477);
assign n13376 = ~n26191;
assign n1482 = ~(n7935 ^ n11552);
assign n4400 = ~n18500;
assign n11183 = n23304 | n17069;
assign n3082 = ~(n18806 ^ n24136);
assign n2380 = ~(n3257 | n3677);
assign n25507 = ~(n19327 | n21934);
assign n24658 = ~n21473;
assign n7848 = n5277 | n19123;
assign n11257 = ~n10631;
assign n17493 = ~(n23147 ^ n6536);
assign n6581 = ~(n16257 | n4119);
assign n16709 = ~n15291;
assign n2365 = ~(n24786 ^ n20036);
assign n2575 = n16622 & n23946;
assign n25596 = ~(n557 | n16006);
assign n5971 = n586 | n21825;
assign n6694 = n7661 | n459;
assign n11029 = ~(n14323 ^ n14071);
assign n7338 = ~(n20230 ^ n18034);
assign n5969 = ~(n23212 ^ n2728);
assign n7156 = n2341 & n2503;
assign n21734 = ~n25568;
assign n17783 = n23055 | n3696;
assign n12291 = ~(n26635 ^ n12399);
assign n16152 = n8672 & n5296;
assign n3208 = ~(n23902 ^ n7132);
assign n25848 = n17357 & n20419;
assign n14047 = ~(n9110 ^ n13282);
assign n10922 = n12520 & n26933;
assign n9693 = ~n15062;
assign n14151 = ~n8418;
assign n2144 = ~(n17370 | n11061);
assign n19133 = n14133 | n4024;
assign n5328 = ~n12169;
assign n506 = ~n24326;
assign n23950 = ~(n3887 ^ n327);
assign n12297 = ~(n8336 ^ n2985);
assign n23821 = n20446 | n24606;
assign n17455 = ~(n2812 ^ n5736);
assign n15437 = ~(n26360 ^ n110);
assign n12145 = ~(n2256 ^ n20694);
assign n24769 = n16002 | n3945;
assign n25453 = n2846 | n23087;
assign n22715 = ~n16324;
assign n12189 = ~(n21247 | n17390);
assign n19226 = n3958 & n10746;
assign n17318 = n17834 & n22663;
assign n21912 = ~(n1286 ^ n15645);
assign n9969 = ~n19940;
assign n14370 = n13131 | n5528;
assign n23976 = ~(n13037 | n13129);
assign n12303 = ~(n25119 | n21934);
assign n632 = n19267 | n4177;
assign n1543 = n21241 & n10060;
assign n10162 = n7051 | n6749;
assign n19766 = n15517 | n8120;
assign n10542 = n5802 & n19368;
assign n19605 = ~n10884;
assign n25342 = ~(n19673 | n5462);
assign n15559 = n26451 | n26155;
assign n7852 = n13162 | n23346;
assign n14762 = ~(n15431 ^ n25310);
assign n16452 = n26224 & n8672;
assign n15342 = ~(n22654 ^ n21915);
assign n11132 = ~(n3808 ^ n923);
assign n2714 = n10078 | n4373;
assign n11354 = ~(n26324 ^ n12262);
assign n7044 = n11324 | n20168;
assign n2288 = n4304 ^ n21114;
assign n22463 = ~(n27118 ^ n7678);
assign n13657 = n22879 & n12616;
assign n26436 = n21489 | n4085;
assign n498 = ~(n20296 ^ n17338);
assign n10259 = ~(n12046 | n6072);
assign n11612 = n1509 | n16913;
assign n15014 = ~(n5140 ^ n6105);
assign n14298 = ~(n11305 ^ n3001);
assign n11943 = n15983 | n23117;
assign n3781 = ~(n6969 ^ n22339);
assign n7415 = n7844 & n9541;
assign n1512 = ~(n15288 ^ n12361);
assign n5760 = ~n8151;
assign n843 = n20373 & n1375;
assign n21312 = n8322 | n19081;
assign n26878 = ~(n24116 | n11580);
assign n16126 = ~(n16234 ^ n4673);
assign n23468 = n2396 & n432;
assign n23955 = ~(n23290 ^ n10709);
assign n18883 = ~(n15652 ^ n4939);
assign n18128 = n19375 | n9278;
assign n24608 = ~(n4750 ^ n7859);
assign n17097 = n23359 | n11898;
assign n2305 = ~(n4941 ^ n9780);
assign n46 = n8561 & n4470;
assign n2635 = n10366 | n16814;
assign n19292 = n11429 | n12969;
assign n16767 = ~(n10773 | n22470);
assign n4048 = n21686 | n17191;
assign n16233 = ~(n8596 ^ n15508);
assign n8969 = n12264 & n27137;
assign n15750 = n10044 | n24999;
assign n20809 = ~(n25953 | n24460);
assign n1223 = ~(n24043 ^ n10201);
assign n8265 = n2421 & n11243;
assign n15634 = n24555 | n5985;
assign n4582 = ~(n16988 | n20442);
assign n14960 = ~(n13492 ^ n23763);
assign n7824 = ~(n10667 ^ n19636);
assign n1821 = ~(n10477 ^ n6548);
assign n24136 = ~(n13854 ^ n18503);
assign n25024 = ~(n21547 | n6003);
assign n11068 = n6482 & n8710;
assign n14191 = n17065 | n11124;
assign n12712 = ~(n10053 | n5329);
assign n23682 = n6833 | n24615;
assign n6088 = ~(n15572 ^ n2989);
assign n4102 = n11089 & n972;
assign n16731 = ~n13284;
assign n25553 = ~(n12900 | n1255);
assign n2936 = n5244 | n16373;
assign n12055 = ~n24714;
assign n2367 = ~(n1308 ^ n7734);
assign n3531 = ~(n4075 | n12120);
assign n7766 = n1742 | n14251;
assign n3221 = n12305 | n24817;
assign n5496 = ~(n24519 ^ n12161);
assign n3028 = n24792 & n18299;
assign n26381 = n25940 | n22325;
assign n15110 = n27071 | n18595;
assign n8673 = n19949 | n11136;
assign n17790 = ~n17311;
assign n17814 = ~(n4304 | n19413);
assign n1162 = ~(n12103 ^ n9448);
assign n2447 = n12914 | n6846;
assign n16414 = n24414 | n22434;
assign n11182 = ~(n11977 ^ n10059);
assign n994 = n7094 | n21163;
assign n6283 = ~(n15730 ^ n2331);
assign n15514 = ~n19431;
assign n7778 = ~(n1279 | n14875);
assign n20288 = ~(n9711 ^ n19064);
assign n19303 = ~(n18913 ^ n15352);
assign n10492 = ~(n1594 | n16602);
assign n23968 = ~(n16781 | n15777);
assign n25708 = n22430 & n9676;
assign n12188 = ~(n23779 ^ n11615);
assign n393 = ~n1924;
assign n6870 = ~(n15743 | n2809);
assign n4903 = n9296 | n25915;
assign n4885 = ~(n17390 ^ n22736);
assign n26908 = n21937 | n25355;
assign n12069 = n7716 | n22654;
assign n15956 = ~(n3209 ^ n9306);
assign n615 = n26222 & n12565;
assign n11697 = ~n15108;
assign n20750 = ~(n10557 | n18113);
assign n14731 = ~(n22861 ^ n4426);
assign n7272 = ~(n20620 ^ n14575);
assign n8579 = ~(n14996 | n10357);
assign n13821 = ~n6483;
assign n14044 = ~(n13731 ^ n13714);
assign n15259 = ~n16705;
assign n4650 = ~(n19842 | n7258);
assign n5340 = n3228 | n20189;
assign n23483 = n649 | n26065;
assign n4502 = ~(n25718 ^ n4634);
assign n15988 = n21395 & n10856;
assign n17129 = ~(n16751 | n25018);
assign n5914 = n8280;
assign n24366 = ~n1152;
assign n6423 = ~(n21471 ^ n19357);
assign n8767 = ~(n9399 ^ n9507);
assign n10668 = n11976 & n11437;
assign n1618 = ~(n22354 ^ n5744);
assign n6811 = n11485 & n11582;
assign n6912 = ~(n18881 ^ n25016);
assign n3268 = n26797 | n16221;
assign n10904 = ~n13262;
assign n16040 = ~(n17184 ^ n18587);
assign n10805 = n6239 | n8319;
assign n12066 = ~n20013;
assign n14541 = ~(n15650 ^ n15691);
assign n544 = ~n9359;
assign n345 = ~(n6908 ^ n26972);
assign n3287 = n2241 & n16418;
assign n11362 = n26122 | n26306;
assign n19249 = n4698 & n14623;
assign n16642 = ~n3217;
assign n4276 = n19746 & n22693;
assign n13798 = ~(n10471 ^ n13403);
assign n15049 = ~n19039;
assign n16142 = ~(n24661 ^ n15462);
assign n7155 = ~(n8708 | n9402);
assign n12965 = ~(n19460 | n16064);
assign n9320 = n13861 & n4021;
assign n5676 = n25206 & n10502;
assign n6720 = n7099 | n18888;
assign n7880 = ~(n23039 | n4590);
assign n13662 = n2314 | n25643;
assign n11881 = ~(n24557 | n15630);
assign n3713 = ~(n1082 ^ n10277);
assign n19185 = n9351 | n16360;
assign n1500 = n7822 & n24543;
assign n5886 = ~n10024;
assign n4811 = ~(n16075 ^ n9370);
assign n24765 = ~(n776 | n13494);
assign n22996 = n21078 | n13725;
assign n11954 = n12140 | n8791;
assign n6875 = ~(n17333 ^ n14783);
assign n8633 = n9493 | n12297;
assign n169 = n16853 | n8768;
assign n24015 = ~(n11061 ^ n1971);
assign n7049 = ~(n21882 ^ n26694);
assign n9837 = n844 | n3103;
assign n21487 = ~(n23262 ^ n12931);
assign n25522 = n14052 | n18925;
assign n2329 = ~(n23582 | n16738);
assign n8170 = ~(n19159 ^ n23399);
assign n22461 = n18581 | n12567;
assign n25272 = n11996 | n7430;
assign n13970 = n25408 | n15781;
assign n6073 = n5395 & n11991;
assign n5512 = ~n12315;
assign n315 = n17978 | n3134;
assign n9791 = n1792 & n19521;
assign n10173 = n7461 & n26464;
assign n20068 = ~(n10602 ^ n22395);
assign n26992 = ~(n22142 ^ n26081);
assign n24461 = ~(n25980 ^ n15182);
assign n20769 = n3453 & n6487;
assign n14316 = n1341 & n7821;
assign n12518 = ~(n2312 ^ n10378);
assign n17567 = n13078 & n19183;
assign n12914 = n21101 & n17779;
assign n25478 = n2482 | n19104;
assign n10135 = ~(n15490 ^ n18);
assign n20210 = ~(n6489 ^ n16743);
assign n20231 = ~(n6049 ^ n23816);
assign n16897 = n4392 & n14834;
assign n27135 = ~(n18742 ^ n14319);
assign n12169 = ~(n5816 ^ n5438);
assign n9379 = n15571 & n16838;
assign n3465 = ~(n2843 ^ n25232);
assign n26234 = ~(n7963 ^ n6590);
assign n8802 = ~(n6523 | n24479);
assign n26052 = n10333 & n2100;
assign n27099 = ~n24444;
assign n8193 = n11862 | n23070;
assign n2611 = ~(n17607 ^ n23366);
assign n12641 = ~(n26991 | n23330);
assign n17337 = ~(n24895 ^ n21970);
assign n20293 = ~(n6937 ^ n17843);
assign n22258 = n7165 | n23239;
assign n23268 = ~(n9895 ^ n15537);
assign n2724 = ~n14275;
assign n24787 = n6958 & n2912;
assign n10134 = n14619 | n26251;
assign n16450 = n14566 & n11895;
assign n7410 = ~n11454;
assign n19398 = ~(n8119 | n26135);
assign n24828 = ~(n5679 ^ n20839);
assign n15665 = n17630 & n18557;
assign n10866 = ~(n17250 ^ n11044);
assign n12112 = ~n21620;
assign n17654 = n11834 & n5788;
assign n24590 = ~n6492;
assign n19858 = ~(n16271 ^ n3117);
assign n495 = n8981 | n22593;
assign n4029 = ~n2530;
assign n4 = n2159 & n5056;
assign n23256 = n17707 & n27133;
assign n4260 = ~(n17250 ^ n15241);
assign n4477 = ~(n17517 ^ n23099);
assign n18621 = ~n5034;
assign n751 = ~(n5031 | n6510);
assign n18804 = n11972 & n19507;
assign n17281 = n25671 | n17040;
assign n16952 = ~(n25365 | n15456);
assign n11050 = n21992 & n13289;
assign n23838 = n5410 | n8358;
assign n19123 = n16341 & n11218;
assign n1741 = ~(n8720 ^ n3803);
assign n9146 = ~(n15310 ^ n5844);
assign n11921 = ~n23216;
assign n9297 = ~(n26170 | n23664);
assign n1585 = n21821 | n25530;
assign n2040 = n22851 & n5988;
assign n508 = ~n14199;
assign n8958 = ~(n3704 ^ n9021);
assign n12905 = ~(n23704 ^ n2659);
assign n19917 = n20814 | n22936;
assign n13675 = n12567 | n12279;
assign n5433 = ~n16411;
assign n6948 = ~n477;
assign n18900 = n27199 | n12964;
assign n7730 = n26634 | n7314;
assign n14015 = ~(n6895 ^ n20462);
assign n2038 = ~(n26190 ^ n12355);
assign n16397 = ~(n11533 ^ n14398);
assign n25045 = ~(n3136 ^ n5752);
assign n17407 = ~(n24656 | n13583);
assign n11586 = n19568 & n162;
assign n12030 = ~(n27053 | n12544);
assign n11340 = n18709 & n27016;
assign n9347 = n212 & n9928;
assign n12971 = ~n2608;
assign n26296 = n14510 & n8994;
assign n19402 = ~(n2036 ^ n2891);
assign n6651 = n23537 | n11010;
assign n13822 = ~n22793;
assign n6761 = n17319 & n9511;
assign n6735 = n25650 | n5077;
assign n23315 = ~n6387;
assign n17571 = n11966 & n6722;
assign n15416 = n15576 | n21739;
assign n17561 = n8690 & n9363;
assign n20499 = n23949 & n17093;
assign n13343 = ~n6372;
assign n12056 = n5918 | n2944;
assign n16297 = n7632 | n14384;
assign n17117 = ~(n8083 ^ n18705);
assign n4116 = ~n25995;
assign n2644 = n7146 | n3549;
assign n5786 = ~(n17959 ^ n6861);
assign n20473 = n22256 | n16220;
assign n13280 = ~n3480;
assign n22486 = n1831 | n10022;
assign n1210 = n11700 & n13398;
assign n5096 = ~(n23709 ^ n19282);
assign n11854 = ~(n12464 | n18907);
assign n20185 = n21597 & n22722;
assign n24314 = ~(n1432 | n2852);
assign n25787 = ~n17694;
assign n14945 = n14128 & n2256;
assign n19885 = n23774 & n24751;
assign n17179 = n26191 | n13284;
assign n26622 = n16402 & n24944;
assign n6140 = n22439 & n26235;
assign n3628 = ~(n13539 ^ n20973);
assign n5362 = n7951 & n15443;
assign n18139 = ~(n6208 ^ n10177);
assign n21400 = ~n13963;
assign n2314 = ~n329;
assign n18305 = ~(n8428 | n25961);
assign n5015 = n21856 | n24163;
assign n6829 = ~(n1118 ^ n10053);
assign n3647 = n4686 | n21836;
assign n1948 = n34 | n13625;
assign n8482 = ~(n24488 ^ n23250);
assign n22857 = ~(n3346 ^ n8044);
assign n21401 = n19129 & n20855;
assign n10105 = ~n12419;
assign n23943 = ~(n23798 | n12217);
assign n25620 = n5101 & n17423;
assign n26606 = n10156 | n12416;
assign n14119 = ~n6590;
assign n16613 = n11580 | n2035;
assign n5978 = ~(n22640 ^ n7566);
assign n22185 = ~(n1209 | n13599);
assign n68 = ~(n6731 | n7347);
assign n17801 = n23315 | n14463;
assign n9340 = ~n15458;
assign n19393 = ~(n3732 ^ n23196);
assign n4069 = n2631 & n7559;
assign n17065 = ~(n20151 | n5852);
assign n22704 = ~(n7407 ^ n9625);
assign n7412 = n1259 | n44;
assign n665 = ~(n12077 ^ n3596);
assign n25566 = ~n18213;
assign n26563 = n8895 | n13727;
assign n26755 = n10273 | n24648;
assign n3559 = ~(n27188 ^ n4326);
assign n2819 = ~(n12771 ^ n5025);
assign n17894 = n2877 | n20457;
assign n18108 = ~(n16070 ^ n20008);
assign n6841 = ~n7330;
assign n17598 = ~(n12677 ^ n10974);
assign n23114 = ~n10751;
assign n11005 = ~(n19407 ^ n25398);
assign n22397 = ~n14057;
assign n16632 = n14401 | n26306;
assign n14914 = n8200 & n21192;
assign n15084 = n23477 | n1365;
assign n21227 = n12702 | n13672;
assign n10879 = n3775 & n23221;
assign n23725 = ~n11933;
assign n238 = n2445 | n7511;
assign n6869 = ~(n13957 | n13343);
assign n21475 = ~(n27120 | n23264);
assign n5550 = n12578 & n16671;
assign n611 = n23396 & n17790;
assign n23997 = n6464 & n7351;
assign n21931 = n5345 & n17363;
assign n26478 = ~(n12258 | n14774);
assign n7331 = ~n6038;
assign n23390 = n22198 & n24493;
assign n6237 = ~(n5465 ^ n17505);
assign n14971 = ~(n1765 ^ n25119);
assign n17032 = ~(n20845 | n26848);
assign n12458 = ~(n5288 | n24923);
assign n8468 = n16034 | n10451;
assign n15595 = n25021 | n26495;
assign n23958 = ~(n22098 ^ n7174);
assign n1010 = n16767 | n23606;
assign n21814 = ~n4062;
assign n20025 = ~(n25974 ^ n19005);
assign n10328 = n3970 | n4059;
assign n25113 = ~(n3572 ^ n3148);
assign n3638 = ~(n21652 ^ n5225);
assign n2169 = ~n19531;
assign n14379 = n13601 & n20540;
assign n6172 = ~(n19875 ^ n9737);
assign n17585 = ~(n20794 ^ n25471);
assign n21281 = ~(n12343 | n14106);
assign n11840 = ~n323;
assign n17010 = ~n17530;
assign n2201 = ~(n1112 ^ n7751);
assign n23427 = n20536 & n2749;
assign n1057 = ~(n2093 ^ n22173);
assign n24344 = ~(n2924 ^ n13669);
assign n828 = n4967 | n18559;
assign n24731 = ~n6135;
assign n4086 = ~(n14210 ^ n21078);
assign n2053 = n25791 | n15088;
assign n17584 = ~n26986;
assign n16520 = ~(n8443 ^ n5170);
assign n13458 = n11179 | n6668;
assign n8575 = n7827 | n23203;
assign n20534 = n20798 & n9878;
assign n7089 = ~(n10937 ^ n16376);
assign n18150 = n21260 | n24121;
assign n130 = n13800 | n25766;
assign n4686 = ~(n25751 | n21850);
assign n19896 = ~(n3393 ^ n1465);
assign n4345 = ~(n13502 ^ n21055);
assign n2507 = ~(n14148 ^ n14275);
assign n8395 = ~n14102;
assign n18912 = ~(n9877 | n23464);
assign n21657 = n23584 & n26020;
assign n10408 = ~(n23740 ^ n2858);
assign n25853 = n11859 & n15770;
assign n2440 = ~(n5656 ^ n21005);
assign n20982 = ~n12696;
assign n17138 = ~(n15849 ^ n7278);
assign n22752 = n2842 | n20933;
assign n1463 = n19469 | n13989;
assign n13180 = n16221 | n21444;
assign n21139 = n25588 | n25613;
assign n24425 = ~(n18983 ^ n4487);
assign n2682 = n21380 | n15659;
assign n20166 = n20589 | n26021;
assign n26693 = ~(n14633 ^ n2886);
assign n24587 = n6996 & n8570;
assign n3982 = n2230 | n19227;
assign n1263 = n17077 & n14620;
assign n5577 = n24607 | n7903;
assign n20701 = n19541 | n25749;
assign n3338 = n5141 & n24637;
assign n10974 = ~(n19042 ^ n23586);
assign n20801 = ~(n26450 | n17351);
assign n26285 = ~(n8163 ^ n2688);
assign n10155 = ~n18171;
assign n22600 = ~n25115;
assign n11290 = n15044 | n12377;
assign n26216 = ~(n4985 ^ n11242);
assign n2332 = ~(n8003 | n22972);
assign n23356 = n6871 | n18328;
assign n26943 = ~(n25732 ^ n11565);
assign n23960 = ~(n11337 ^ n11893);
assign n18722 = n21280 | n7002;
assign n8060 = n14778 | n13510;
assign n26578 = n20978 | n25243;
assign n8207 = n9147 & n24597;
assign n26360 = n20504 & n14896;
assign n23662 = n21879 | n8853;
assign n19754 = n21956 & n17700;
assign n21375 = n24461 & n26095;
assign n16347 = ~(n9107 | n18360);
assign n5826 = ~n6265;
assign n19083 = ~(n839 | n6139);
assign n18137 = ~(n13219 ^ n19376);
assign n3799 = ~(n7242 ^ n880);
assign n18185 = n26069 | n23277;
assign n24808 = n8435 & n9580;
assign n15398 = n20076 & n4970;
assign n1387 = ~n10699;
assign n15229 = ~n20014;
assign n22886 = ~(n20127 | n19927);
assign n9070 = n4149 | n12875;
assign n12018 = ~n11671;
assign n15835 = ~(n3045 ^ n9376);
assign n20184 = ~(n4326 | n3952);
assign n2571 = n7124 | n16510;
assign n7698 = ~(n14729 ^ n1976);
assign n10921 = n438 | n18784;
assign n9580 = n3422 | n22525;
assign n12196 = ~(n24237 | n4017);
assign n19095 = n5329 & n2694;
assign n10846 = ~(n16882 ^ n3976);
assign n21688 = n25068 | n23535;
assign n7440 = n6869 | n1159;
assign n20818 = n26092 | n24930;
assign n16067 = n7759 | n10479;
assign n7988 = ~(n22772 ^ n8930);
assign n6839 = n17856 | n18790;
assign n20433 = ~n17824;
assign n26942 = ~(n24308 ^ n13075);
assign n5781 = n2058 & n10112;
assign n15037 = n15154 | n19445;
assign n8643 = n17371 & n4695;
assign n8647 = ~n271;
assign n26675 = ~(n5370 ^ n9685);
assign n2084 = ~(n23913 | n3710);
assign n21485 = ~n15190;
assign n3709 = n18994 & n7787;
assign n18269 = ~n10057;
assign n4859 = ~n10250;
assign n15828 = ~(n19701 ^ n7437);
assign n18440 = n7602 & n4475;
assign n13163 = ~(n905 | n4706);
assign n17378 = ~(n6270 | n27121);
assign n19344 = n24890 | n4665;
assign n15716 = ~(n720 ^ n6888);
assign n18509 = ~(n5459 ^ n6467);
assign n19926 = ~n23776;
assign n12361 = ~(n18255 ^ n15636);
assign n16055 = n7161 | n16411;
assign n2286 = n8921 & n26734;
assign n6200 = ~n4184;
assign n9030 = n11980 | n19446;
assign n25448 = n8021 | n25309;
assign n6844 = n21613 | n8974;
assign n16021 = n18244 & n4107;
assign n9373 = ~n24928;
assign n14492 = ~(n10758 | n13562);
assign n22862 = ~n11295;
assign n2835 = n23428 | n8649;
assign n20519 = ~(n13945 ^ n12341);
assign n22384 = n18114 | n1;
assign n15690 = n18761 | n5665;
assign n19708 = ~(n8006 ^ n5211);
assign n9992 = ~(n13891 ^ n11140);
assign n13316 = n1414 | n4005;
assign n18703 = n2789 & n13640;
assign n5502 = n22318 | n1162;
assign n3486 = n375 & n25771;
assign n5086 = n22299 & n13294;
assign n174 = n22737 | n3767;
assign n23585 = ~(n3467 ^ n19456);
assign n11538 = ~(n156 ^ n22058);
assign n5818 = ~(n212 ^ n17150);
assign n14574 = n21777 | n15392;
assign n18010 = ~(n4230 ^ n8378);
assign n14158 = ~n24219;
assign n26753 = n12505 | n24497;
assign n2389 = ~(n24436 ^ n21885);
assign n20926 = n7577 & n15731;
assign n14987 = n24540 | n14901;
assign n5142 = ~(n974 ^ n18668);
assign n15328 = ~(n22972 ^ n3945);
assign n5556 = ~(n7787 ^ n23722);
assign n13958 = ~(n7014 ^ n13611);
assign n21212 = ~(n24902 ^ n25572);
assign n9212 = ~n16814;
assign n4709 = n6204 & n23898;
assign n19434 = n25823 | n2018;
assign n1430 = n24532 & n18021;
assign n25541 = n19699 & n24526;
assign n3433 = n12787 & n2016;
assign n16318 = n25776 & n628;
assign n19404 = ~(n15924 ^ n2680);
assign n1795 = n19061 | n13436;
assign n16676 = n9471 | n6589;
assign n15627 = n17251 | n23967;
assign n2827 = ~(n23631 ^ n22765);
assign n7630 = ~(n25995 ^ n21115);
assign n22581 = ~(n12734 ^ n631);
assign n26282 = ~(n8722 ^ n13119);
assign n1145 = n1932 & n14526;
assign n12996 = ~n18145;
assign n8283 = ~(n7805 ^ n7657);
assign n15763 = n7089 & n16793;
assign n22953 = ~(n18614 ^ n19420);
assign n24683 = n331 | n684;
assign n7045 = ~(n9655 ^ n13074);
assign n20415 = ~(n11883 ^ n14064);
assign n16549 = n3676 & n9224;
assign n15454 = ~n9554;
assign n11160 = n9070 & n10842;
assign n18593 = n2085 & n5169;
assign n9937 = ~(n6319 ^ n442);
assign n21252 = ~(n17734 ^ n23253);
assign n13266 = ~(n9535 ^ n2615);
assign n10518 = n23808 | n20887;
assign n22776 = ~(n9993 ^ n25926);
assign n19446 = ~(n19545 ^ n25749);
assign n11622 = ~(n8371 | n4410);
assign n10489 = ~(n11396 ^ n14797);
assign n3426 = ~(n11693 ^ n13375);
assign n19031 = n9913 | n20428;
assign n2637 = ~(n11363 | n14119);
assign n5271 = n5355 | n17659;
assign n22687 = ~(n9333 ^ n14666);
assign n19884 = ~n8635;
assign n12282 = ~(n25974 | n2355);
assign n21399 = ~(n23421 ^ n10846);
assign n18839 = n9262 | n16934;
assign n19981 = n4256 | n5713;
assign n9262 = n11089 & n4955;
assign n16085 = ~(n25324 | n1630);
assign n9037 = n26782 | n20089;
assign n915 = n7325 ^ n15232;
assign n20737 = ~n15167;
assign n9989 = ~(n10218 ^ n19547);
assign n21970 = ~(n20771 ^ n18639);
assign n20501 = n5304 | n13115;
assign n5805 = ~(n3785 ^ n21);
assign n15039 = ~(n18295 ^ n16223);
assign n18577 = ~(n11499 ^ n18570);
assign n19860 = n21360 & n2311;
assign n6655 = ~(n13067 ^ n25735);
assign n25416 = n7991 ^ n13323;
assign n22305 = n24737 & n25767;
assign n10865 = n176 | n1452;
assign n25878 = n5836 | n17788;
assign n24141 = ~(n5909 ^ n15401);
assign n23066 = n22011 & n17042;
assign n2921 = n6533 | n24685;
assign n4658 = ~n4869;
assign n1379 = n18274 | n24383;
assign n23793 = ~n15508;
assign n13151 = ~(n9717 ^ n407);
assign n12045 = n15699 & n25732;
assign n15335 = n10292 & n20559;
assign n26097 = n12471 | n23533;
assign n11671 = ~(n7415 ^ n8242);
assign n17241 = n21892 & n20779;
assign n5906 = n23304 | n1465;
assign n25779 = ~n3078;
assign n2573 = ~(n13806 ^ n20351);
assign n22611 = n23830 | n19342;
assign n25813 = ~(n24075 ^ n20941);
assign n147 = ~n11721;
assign n10660 = ~(n22951 ^ n14561);
assign n11037 = n7705 | n19016;
assign n18875 = ~(n16500 ^ n8678);
assign n804 = ~(n20051 ^ n18434);
assign n23302 = ~n18265;
assign n15360 = n19632 | n6085;
assign n5325 = ~(n20116 ^ n12054);
assign n9642 = n12562 | n12351;
assign n14803 = n15135 & n25712;
assign n2340 = ~(n26443 | n10017);
assign n10991 = n19954 & n9596;
assign n21082 = ~(n21345 ^ n9190);
assign n20653 = n4834 | n23823;
assign n19876 = n17090 | n6773;
assign n13169 = n5704 & n5512;
assign n15007 = ~n4513;
assign n7239 = n12434 & n11681;
assign n9616 = ~(n17146 ^ n4004);
assign n16798 = ~(n12332 ^ n20692);
assign n26585 = ~(n420 ^ n18219);
assign n7503 = ~n8622;
assign n27149 = ~(n25586 | n8491);
assign n1252 = ~n3795;
assign n12120 = n21539 & n6200;
assign n18523 = n2102 | n598;
assign n21264 = n18237 & n2847;
assign n10589 = n25763 | n13145;
assign n10864 = ~(n1705 ^ n9456);
assign n21440 = n16453 | n12033;
assign n5642 = n21383 & n13624;
assign n4744 = ~n766;
assign n2467 = ~n25718;
assign n13326 = ~(n18157 | n2698);
assign n21826 = ~(n7335 | n4319);
assign n7177 = ~n7010;
assign n25770 = ~(n5847 ^ n27188);
assign n12493 = n24425;
assign n20412 = n4341 | n5069;
assign n20020 = ~n3072;
assign n347 = n25 & n23382;
assign n14735 = ~n21688;
assign n3093 = ~n15421;
assign n13434 = n22644 | n8918;
assign n10822 = n12846 & n10968;
assign n9165 = n9821 & n11838;
assign n25214 = ~(n25967 ^ n4409);
assign n21944 = n3136 | n4423;
assign n23722 = ~(n16936 ^ n7515);
assign n3183 = ~(n4999 ^ n19196);
assign n7807 = ~(n21982 | n5760);
assign n3011 = ~(n1387 | n2782);
assign n21070 = ~n6549;
assign n16361 = n22362 & n26589;
assign n21248 = ~n20080;
assign n9883 = n21510;
assign n7259 = n12962 | n18322;
assign n935 = ~(n9347 | n3723);
assign n16083 = ~(n23930 ^ n14055);
assign n8630 = ~(n18371 | n7933);
assign n3277 = n9587 | n18816;
assign n3741 = ~(n26915 ^ n14598);
assign n152 = ~(n7498 ^ n14180);
assign n891 = n19588 | n8041;
assign n11828 = n19152 & n22567;
assign n12259 = n13781 & n10917;
assign n10900 = n18035 | n3279;
assign n5618 = n18383 | n17959;
assign n27106 = n3480 & n11393;
assign n6788 = ~(n19680 | n17360);
assign n10973 = ~(n17386 ^ n5073);
assign n4181 = ~n25628;
assign n2176 = n6851 & n2656;
assign n19200 = n19955;
assign n4901 = ~(n20193 ^ n16768);
assign n2715 = n4297 & n9171;
assign n27101 = ~(n17198 ^ n19170);
assign n21061 = n7930 | n20929;
assign n17568 = ~n3425;
assign n21176 = ~(n15181 ^ n9503);
assign n25193 = n16760 | n7415;
assign n9108 = ~n16874;
assign n19009 = n26606 & n16914;
assign n20553 = n14518 & n18806;
assign n25367 = n1226 & n26610;
assign n22964 = ~n2850;
assign n16097 = ~(n6089 ^ n25476);
assign n8372 = ~n1558;
assign n22944 = ~(n6397 | n10995);
assign n18889 = n22268 & n11931;
assign n26435 = n11363 | n12161;
assign n3825 = n25522 & n484;
assign n10283 = ~(n15766 ^ n6105);
assign n6561 = ~n10076;
assign n14768 = ~(n13846 ^ n26625);
assign n20934 = n8949 | n20469;
assign n14482 = ~(n6694 ^ n21707);
assign n5529 = n7954 & n4157;
assign n10384 = n14719 & n24215;
assign n1726 = ~n25843;
assign n26919 = ~n791;
assign n22370 = ~n21934;
assign n5979 = n14086 | n25077;
assign n3760 = ~(n509 ^ n403);
assign n11082 = n19074 | n15936;
assign n20668 = ~(n15417 ^ n24578);
assign n11477 = ~n26851;
assign n13206 = ~n22121;
assign n10167 = n23141 & n1370;
assign n13284 = ~(n19149 ^ n11409);
assign n2127 = n5479 & n9891;
assign n16514 = ~n3614;
assign n15343 = ~(n10660 ^ n8897);
assign n3693 = n10380 & n1548;
assign n16210 = ~n4376;
assign n21729 = n25376 & n2378;
assign n10884 = n10747 & n9578;
assign n13444 = ~(n22012 ^ n18883);
assign n2591 = n9706 | n24554;
assign n20806 = n15056 | n13572;
assign n8182 = ~(n19433 ^ n13951);
assign n9215 = ~(n8831 ^ n20539);
assign n19286 = n26029 & n17582;
assign n17668 = n26760 | n25596;
assign n8704 = ~n6032;
assign n23083 = ~(n7799 ^ n24879);
assign n21834 = ~(n6471 ^ n15489);
assign n26 = n13332 | n6112;
assign n4498 = n16477 | n10767;
assign n13140 = n23793 | n8596;
assign n16776 = ~(n4199 | n6529);
assign n2853 = ~(n7732 ^ n4898);
assign n25377 = ~n11293;
assign n25645 = n12513 | n8395;
assign n23372 = ~(n20129 ^ n24035);
assign n6081 = n15049 | n5139;
assign n24889 = ~n2186;
assign n11175 = n6456 | n17978;
assign n11009 = ~(n6729 | n11192);
assign n6988 = ~(n12635 ^ n17791);
assign n9569 = ~n8251;
assign n9196 = ~n24323;
assign n6777 = n20095 & n6980;
assign n4882 = n1898 | n14395;
assign n3583 = n19035 & n3539;
assign n16803 = ~(n10730 ^ n14399);
assign n12433 = ~(n3284 ^ n15643);
assign n9684 = ~(n19609 | n19132);
assign n14903 = n3956 | n23167;
assign n22441 = n19460 | n17530;
assign n8967 = n17979 | n13578;
assign n3806 = ~(n162 ^ n26174);
assign n3735 = ~(n18975 ^ n8411);
assign n3771 = n19384 | n14041;
assign n18535 = ~n18488;
assign n22032 = n17817 | n19900;
assign n1922 = ~(n15769 ^ n13490);
assign n13929 = ~(n8185 | n18402);
assign n609 = ~n16840;
assign n3723 = n17608 & n2591;
assign n15015 = ~(n18031 | n21537);
assign n26444 = ~(n953 ^ n14501);
assign n25191 = n8181 & n15953;
assign n146 = ~n11898;
assign n22452 = ~(n5629 ^ n15546);
assign n11130 = n5215 & n14368;
assign n19977 = n1892 & n26277;
assign n5143 = ~n307;
assign n4740 = n26618 | n12658;
assign n17413 = n14289 | n17132;
assign n26827 = n8680 | n16611;
assign n8010 = ~(n20512 | n25726);
assign n3307 = ~(n21192 ^ n13003);
assign n23040 = n16993 | n3829;
assign n23761 = n19921 | n14238;
assign n17006 = ~(n18464 ^ n5548);
assign n12270 = n12722 & n20236;
assign n4810 = ~(n23350 ^ n2303);
assign n26735 = ~n6053;
assign n24651 = n20417 | n3568;
assign n19746 = n12380 | n4191;
assign n11449 = ~(n10481 | n3407);
assign n9286 = n26312 | n8079;
assign n26960 = n16041 | n5659;
assign n9494 = ~(n13160 ^ n12148);
assign n25528 = n10650 & n17978;
assign n2368 = n9210 | n2729;
assign n19673 = ~n7769;
assign n20105 = n472 | n23586;
assign n8333 = n15135 | n25712;
assign n17941 = n19268 | n20452;
assign n14420 = n13378 | n9323;
assign n1905 = ~n4201;
assign n12737 = n6424 & n15720;
assign n5122 = ~n7060;
assign n13886 = ~n24926;
assign n22525 = n12823 & n2674;
assign n24696 = ~(n3018 ^ n9557);
assign n3682 = ~(n10049 | n7621);
assign n15349 = n14129 | n18286;
assign n16371 = n23776 | n20556;
assign n22396 = ~(n15659 | n6988);
assign n23164 = ~(n17593 | n21376);
assign n2455 = n21934 | n18277;
assign n22863 = ~(n5785 ^ n6006);
assign n640 = ~(n11670 | n8266);
assign n1775 = ~(n15073 | n19814);
assign n14279 = n10492 | n13467;
assign n4777 = ~(n940 ^ n26763);
assign n24040 = ~n5789;
assign n26670 = ~(n5891 | n26100);
assign n5856 = ~(n23321 ^ n6300);
assign n19364 = ~(n16066 ^ n1712);
assign n12087 = n17425 | n4068;
assign n18744 = n5318 & n3943;
assign n13908 = n13138 & n2068;
assign n13324 = n2791 & n24027;
assign n2203 = n22131 | n24064;
assign n21794 = n2184 | n23109;
assign n5843 = n26646 & n4329;
assign n11894 = n24794 & n7826;
assign n11236 = ~(n12406 | n16203);
assign n13525 = n14510 & n7292;
assign n13125 = n11049 & n15097;
assign n8225 = ~(n15786 ^ n12177);
assign n26994 = n10136 & n19519;
assign n8131 = n2626 & n5821;
assign n6060 = n7405 & n3350;
assign n12687 = ~(n14335 ^ n7356);
assign n23108 = n8782 | n24561;
assign n26890 = ~n4901;
assign n7505 = ~(n15146 ^ n5532);
assign n20504 = n23208 | n26583;
assign n16440 = ~(n13416 ^ n20339);
assign n24604 = ~(n18819 ^ n18011);
assign n7356 = ~(n22379 ^ n9967);
assign n21364 = n23157 | n20016;
assign n1588 = n11841 | n17077;
assign n20599 = ~n18926;
assign n12263 = n7648 & n5289;
assign n7237 = ~n23272;
assign n14281 = n13894 | n10277;
assign n14847 = n27057 | n2408;
assign n4583 = ~(n312 ^ n799);
assign n13134 = n19759 | n23941;
assign n19027 = n5696 & n23463;
assign n18442 = n277 | n5112;
assign n1465 = ~(n20559 ^ n14657);
assign n5559 = ~(n10931 ^ n12615);
assign n998 = n22599 | n17897;
assign n5729 = ~(n19608 | n15378);
assign n23552 = n2770 & n2558;
assign n9326 = n8153 & n19355;
assign n21813 = n2987 | n13905;
assign n16344 = n11364 | n18654;
assign n7194 = n15167 & n25330;
assign n758 = n2624 & n23336;
assign n7312 = n2358 & n1208;
assign n17082 = ~(n16697 ^ n9143);
assign n13614 = ~(n9655 ^ n23849);
assign n2778 = n25668 | n18336;
assign n1051 = ~(n25524 | n16325);
assign n19343 = n23062 & n5166;
assign n25984 = ~(n1987 ^ n11161);
assign n21719 = ~(n17701 ^ n18092);
assign n4262 = n18296 | n14207;
assign n1336 = ~n23597;
assign n9537 = n19935 | n8195;
assign n1090 = ~(n19157 ^ n22878);
assign n4860 = n12719 & n22187;
assign n3511 = n4868 | n11425;
assign n992 = ~(n5346 ^ n19121);
assign n22158 = ~n16016;
assign n16228 = n4899 & n1256;
assign n24450 = n9444 & n12425;
assign n11036 = n8265 | n23462;
assign n14084 = n5658 & n15966;
assign n15198 = ~(n7743 | n13263);
assign n13043 = ~(n1173 ^ n91);
assign n8073 = n11057 & n10149;
assign n25652 = n21904 & n17057;
assign n22859 = ~n8352;
assign n4776 = ~(n21780 | n788);
assign n5042 = ~(n26240 ^ n20700);
assign n1409 = n7836 | n19343;
assign n21363 = ~(n3868 | n13259);
assign n5982 = n23726 & n7659;
assign n22161 = n10146 | n26660;
assign n13279 = n14955 | n13098;
assign n26068 = ~(n1658 ^ n19464);
assign n4044 = n24856 | n17724;
assign n25924 = n22128 & n5306;
assign n12023 = n24771 & n22046;
assign n4059 = n21815 & n11012;
assign n26626 = n25941 | n13958;
assign n9633 = ~(n5311 ^ n11717);
assign n23456 = ~n13133;
assign n26420 = ~(n5718 ^ n22643);
assign n53 = n18220 & n20634;
assign n3278 = n20505 | n11539;
assign n16024 = ~n886;
assign n24661 = ~n6102;
assign n13610 = ~(n4230 ^ n16290);
assign n3633 = ~(n3601 | n23894);
assign n5462 = n6400 | n17864;
assign n18631 = n17123 & n21026;
assign n11750 = ~(n25164 | n6285);
assign n1909 = ~n9289;
assign n20526 = n1015 & n26922;
assign n2559 = ~n22631;
assign n6203 = ~n9512;
assign n1492 = n24485 | n14356;
assign n7236 = ~(n14039 ^ n4396);
assign n17792 = ~(n10329 ^ n23222);
assign n17249 = n13721 & n16353;
assign n7251 = n6209 | n4326;
assign n16688 = ~(n10073 ^ n6683);
assign n22139 = ~n8997;
assign n6196 = ~(n23290 ^ n1939);
assign n8557 = n19082 | n8910;
assign n23240 = ~(n7750 ^ n7284);
assign n18536 = n23742 & n6425;
assign n24591 = n11790 | n8279;
assign n6387 = ~(n3060 ^ n3979);
assign n6169 = ~(n20322 ^ n19334);
assign n23543 = ~(n3018 ^ n18537);
assign n5911 = ~(n19537 ^ n26668);
assign n9697 = n23497 | n22413;
assign n23205 = n21681 | n15373;
assign n11747 = n25457 & n9949;
assign n8801 = ~(n10405 | n25370);
assign n25864 = ~(n10782 ^ n15150);
assign n5361 = n7877 & n21591;
assign n4507 = n24403 | n13667;
assign n12364 = ~(n15110 ^ n22940);
assign n25663 = ~n19941;
assign n17547 = ~n5510;
assign n3564 = ~(n12470 ^ n14750);
assign n25198 = ~(n61 ^ n15761);
assign n9230 = n11338 | n12633;
assign n19342 = n74 & n22984;
assign n27163 = ~(n3557 ^ n14985);
assign n4849 = ~(n16364 | n7680);
assign n14467 = n25126 | n22097;
assign n11240 = ~n1218;
assign n12308 = n11021 & n26507;
assign n15199 = n386 | n21758;
assign n23639 = ~n9179;
assign n13962 = n11072 | n18728;
assign n22914 = ~(n7054 ^ n3057);
assign n13980 = ~n21451;
assign n20955 = ~(n8520 | n17590);
assign n11688 = ~(n17043 ^ n23103);
assign n10522 = n4534 | n10654;
assign n6318 = n12530 | n23657;
assign n9056 = n5977 | n8894;
assign n26362 = n8209 | n19479;
assign n5147 = n17453 | n16903;
assign n6977 = n3452 | n555;
assign n26506 = ~n3483;
assign n18232 = ~(n23519 ^ n4092);
assign n25809 = n17021 & n1010;
assign n19996 = ~(n11459 | n18781);
assign n18311 = ~(n8513 ^ n8578);
assign n22991 = n2423 | n2197;
assign n22334 = n7571 | n21484;
assign n1013 = n10424 | n21206;
assign n1321 = n4669 & n7556;
assign n24269 = ~(n17705 ^ n22421);
assign n19555 = n21951 | n10383;
assign n22053 = ~(n22849 | n405);
assign n10978 = ~n22097;
assign n19691 = ~(n12576 ^ n18130);
assign n12192 = ~(n1194 ^ n7881);
assign n20418 = ~(n20444 ^ n12112);
assign n5205 = ~(n19739 ^ n25883);
assign n18210 = ~(n10514 ^ n6105);
assign n20636 = n13304 | n14416;
assign n15575 = n13189 | n18258;
assign n12992 = ~(n7159 ^ n21818);
assign n12695 = n12879 & n9338;
assign n9054 = ~(n11036 ^ n22618);
assign n23124 = ~(n26344 | n14754);
assign n21049 = ~(n15417 ^ n18792);
assign n10033 = ~(n23162 ^ n19241);
assign n8746 = ~(n6946 | n20124);
assign n17059 = n16648 | n13377;
assign n24870 = ~(n7823 ^ n1);
assign n20735 = n16415 | n8465;
assign n16467 = n21784 & n18163;
assign n12015 = n1582 | n17699;
assign n13510 = ~(n26749 | n2938);
assign n13556 = ~(n12758 ^ n8760);
assign n26596 = n24417 & n24907;
assign n7776 = ~n9809;
assign n24359 = ~n14080;
assign n16651 = n1423 | n5346;
assign n11386 = ~(n18458 ^ n5470);
assign n8327 = n20597 | n109;
assign n1996 = ~(n22492 ^ n25523);
assign n1969 = n8322 | n15659;
assign n21833 = ~(n380 ^ n824);
assign n14215 = ~(n24124 ^ n10838);
assign n4413 = n13137 | n3274;
assign n25081 = n23869 & n22127;
assign n19502 = ~n3150;
assign n20072 = ~(n13543 ^ n6794);
assign n6431 = ~(n23459 ^ n6196);
assign n26604 = ~(n19531 ^ n1999);
assign n21757 = n16454 | n10584;
assign n1702 = n15221 | n21853;
assign n15421 = n24652 & n26418;
assign n13985 = n5255 & n25289;
assign n14344 = ~n7593;
assign n23044 = n23470 & n9009;
assign n19946 = n25754 & n12294;
assign n14143 = n23002 | n13556;
assign n26387 = ~(n26968 ^ n25336);
assign n11382 = ~(n15523 ^ n7711);
assign n25933 = n17069 & n19446;
assign n6090 = n12973 | n19742;
assign n14341 = ~n2728;
assign n26946 = ~n15961;
assign n11637 = n8713 & n54;
assign n23088 = ~(n387 | n12293);
assign n15412 = n16216 | n18356;
assign n20898 = ~(n25376 ^ n2378);
assign n16979 = ~(n6670 ^ n10023);
assign n12582 = ~(n21998 | n25779);
assign n26547 = n20497 | n21997;
assign n21171 = n2628 | n15383;
assign n10230 = ~n5490;
assign n24054 = n13913 | n13843;
assign n3014 = n23386 | n15374;
assign n12019 = n4087 | n4667;
assign n6706 = ~(n558 ^ n2765);
assign n7727 = n24065 | n20307;
assign n25487 = ~(n8305 ^ n22253);
assign n27088 = n19192 | n15511;
assign n1088 = ~n7207;
assign n15616 = ~n26306;
assign n18051 = n22285 | n25998;
assign n1808 = ~(n9979 ^ n27007);
assign n521 = ~(n25495 ^ n9152);
assign n11269 = n1786 | n5408;
assign n15045 = n3568 & n18202;
assign n23688 = ~(n19995 ^ n1008);
assign n1556 = n22135 | n1609;
assign n19909 = ~(n13990 ^ n2307);
assign n17094 = n9318 | n1022;
assign n23171 = n13817 | n272;
assign n15352 = ~(n6691 ^ n21753);
assign n22578 = n20158 | n4538;
assign n17030 = n11592 | n14003;
assign n13313 = n22572 & n12752;
assign n26233 = n27166 & n10850;
assign n15553 = ~(n15164 | n16313);
assign n20689 = ~(n25231 ^ n11109);
assign n14397 = ~n18326;
assign n7160 = ~n4288;
assign n18124 = n22134 | n11940;
assign n23361 = ~(n10201 ^ n6814);
assign n8237 = n12579 | n14043;
assign n25519 = ~(n11066 ^ n1552);
assign n9120 = ~(n15787 ^ n7486);
assign n18734 = ~(n495 ^ n22999);
assign n14156 = ~(n9320 ^ n13614);
assign n18832 = n6584 | n4474;
assign n25839 = ~(n24686 ^ n25451);
assign n4198 = ~(n12477 ^ n18035);
assign n3243 = n13039 & n6043;
assign n5773 = n10302 & n2273;
assign n27133 = n23781 | n22904;
assign n21339 = n11914 & n17158;
assign n19672 = n20342 | n14826;
assign n18031 = ~n16744;
assign n15958 = ~(n6964 ^ n22064);
assign n9829 = ~(n11220 | n4299);
assign n7180 = ~(n19078 ^ n18039);
assign n12872 = ~(n18269 | n5026);
assign n24905 = ~(n6082 | n23097);
assign n9754 = n2995 | n17428;
assign n10999 = n19025 & n21962;
assign n25413 = ~(n9721 ^ n3916);
assign n5120 = ~(n4684 ^ n23220);
assign n20792 = n19081 | n26316;
assign n10166 = ~(n23168 | n3962);
assign n16852 = n24301 & n9669;
assign n26112 = n14936 | n6502;
assign n12279 = ~(n23394 ^ n2305);
assign n19468 = n14592 & n12957;
assign n22371 = ~(n22382 ^ n26471);
assign n26081 = ~(n26224 ^ n18483);
assign n5975 = n15083 | n22431;
assign n18275 = n1651 & n23350;
assign n3510 = n16604 & n23348;
assign n22571 = ~n949;
assign n22363 = ~n852;
assign n10193 = n16825 & n17703;
assign n22570 = n4849 | n26245;
assign n9543 = n24391 | n12704;
assign n8639 = n12250 | n24525;
assign n2851 = n3000 | n26385;
assign n6842 = ~n19366;
assign n10828 = n15943 | n19591;
assign n10059 = ~(n18710 ^ n21796);
assign n17272 = n19974 & n22440;
assign n10433 = n20956 | n6699;
assign n2750 = ~n15675;
assign n17747 = n9099 | n5745;
assign n22327 = ~(n17783 ^ n16337);
assign n2126 = ~n23591;
assign n20551 = n26782 | n11088;
assign n6845 = n14145 | n22436;
assign n8031 = n4645 | n7985;
assign n19077 = n2579 | n19081;
assign n1438 = n15884 | n5213;
assign n37 = n24316 & n12745;
assign n13918 = n23837 | n23242;
assign n18102 = ~(n17251 ^ n4913);
assign n19690 = n22155 | n11823;
assign n7634 = ~(n5528 ^ n15828);
assign n8972 = n8754 | n10344;
assign n8930 = n18429;
assign n8078 = ~(n20151 | n20429);
assign n2612 = ~(n10037 ^ n13148);
assign n24192 = n12513 | n8162;
assign n4955 = ~n6925;
assign n8929 = n13714 & n1329;
assign n7280 = ~(n18658 ^ n11928);
assign n21906 = n4882 & n12637;
assign n6702 = ~(n3498 | n14289);
assign n20344 = ~n25415;
assign n11928 = ~(n5949 ^ n21969);
assign n7686 = ~(n19091 ^ n2275);
assign n15591 = n3172 & n17238;
assign n21700 = n13677 & n10451;
assign n24521 = ~(n8367 | n726);
assign n10336 = n24142 & n10569;
assign n887 = ~(n1471 ^ n3152);
assign n6559 = ~(n25296 ^ n23717);
assign n26400 = n9216 | n25107;
assign n18179 = ~n8814;
assign n19213 = n21218 | n9815;
assign n9641 = n12953 & n22328;
assign n13765 = ~(n481 | n15474);
assign n1718 = n26789 | n11733;
assign n719 = n14358 & n6986;
assign n3153 = ~(n19482 | n4177);
assign n27112 = ~(n21130 ^ n18154);
assign n25603 = ~(n3954 ^ n18611);
assign n771 = ~(n26889 ^ n6961);
assign n4063 = ~(n16722 ^ n6385);
assign n25812 = ~(n23254 ^ n27008);
assign n11052 = ~n17784;
assign n5783 = ~n7670;
assign n19828 = ~n20819;
assign n18291 = ~(n14886 ^ n933);
assign n11263 = n2023 | n19489;
assign n17043 = n20985 | n25304;
assign n13761 = ~(n13436 ^ n25693);
assign n22386 = ~n16701;
assign n25155 = ~(n6989 ^ n23257);
assign n10888 = n22948 | n18165;
assign n25995 = n9874 | n6816;
assign n11307 = n8419 | n23727;
assign n10198 = n10473 & n25429;
assign n11831 = ~n16117;
assign n18045 = ~(n9237 ^ n24508);
assign n1274 = n13237 | n5568;
assign n2492 = ~n23346;
assign n10872 = n14695 & n15473;
assign n24798 = ~(n22626 ^ n3324);
assign n23693 = ~(n22314 ^ n22473);
assign n27128 = n707 | n21418;
assign n7901 = n1646 | n4191;
assign n24156 = ~(n24045 ^ n21433);
assign n4298 = ~n17705;
assign n26184 = ~(n5098 | n7436);
assign n5992 = n12583 | n25593;
assign n10116 = ~(n27014 ^ n10322);
assign n17462 = ~(n10001 ^ n21263);
assign n9159 = n21974 & n22284;
assign n15025 = ~(n6814 | n8084);
assign n223 = ~n21223;
assign n11897 = ~(n7234 | n15360);
assign n18862 = ~(n18247 ^ n2409);
assign n19264 = ~(n9359 | n24802);
assign n26341 = n162 & n20509;
assign n6115 = ~(n4504 ^ n14577);
assign n4008 = ~(n11621 ^ n23965);
assign n19534 = ~(n6631 ^ n24732);
assign n8842 = n26168 & n19660;
assign n4463 = n15415 | n4395;
assign n24841 = ~(n17874 ^ n20802);
assign n12935 = n5635 & n17153;
assign n22278 = ~n25632;
assign n5185 = ~n13719;
assign n19853 = n25407 | n20979;
assign n18074 = n15204 | n18478;
assign n3869 = ~(n21722 ^ n10504);
assign n25540 = ~(n405 ^ n4561);
assign n25793 = ~(n26452 ^ n2999);
assign n5590 = n18428 & n16793;
assign n24171 = ~(n3009 ^ n21729);
assign n13670 = n535 | n2705;
assign n7472 = ~(n23161 | n3383);
assign n25219 = n6097 & n11686;
assign n13428 = ~(n25900 | n22715);
assign n7284 = ~(n15788 ^ n12556);
assign n17110 = ~n3460;
assign n13449 = n23863 & n11114;
assign n10088 = ~(n9554 | n8176);
assign n11283 = ~(n6610 | n7752);
assign n6635 = n18100 | n16231;
assign n18120 = n25957 | n19247;
assign n15273 = ~(n5998 ^ n14352);
assign n25145 = n21883 | n15615;
assign n10820 = ~(n18333 ^ n11497);
assign n26178 = ~n1552;
assign n4706 = ~n19486;
assign n19872 = ~n21143;
assign n243 = ~(n25127 ^ n19734);
assign n19403 = ~(n4652 ^ n8521);
assign n21353 = ~(n25849 ^ n7167);
assign n23975 = n19088 | n17516;
assign n5703 = ~(n10072 ^ n21159);
assign n20730 = ~(n21334 | n15273);
assign n22135 = n18724 & n138;
assign n12684 = n9144 & n25236;
assign n1283 = n20292 | n15119;
assign n23262 = n20276 & n16292;
assign n9022 = ~(n23044 ^ n22201);
assign n12173 = n1597 | n26924;
assign n5525 = ~n6413;
assign n23784 = ~(n16471 ^ n12835);
assign n16120 = n20796 | n26444;
assign n2032 = n17626 | n25241;
assign n23305 = ~(n21569 ^ n13151);
assign n415 = ~(n25566 | n16233);
assign n21129 = n14718 | n14440;
assign n18866 = n6600 | n18910;
assign n19368 = ~(n7653 ^ n579);
assign n7742 = n4049 & n19529;
assign n17722 = n25931 | n1510;
assign n17936 = ~(n4028 ^ n17569);
assign n9403 = ~(n14220 ^ n10362);
assign n10073 = n17105 | n24819;
assign n9566 = ~(n25452 ^ n3673);
assign n2185 = ~(n5205 ^ n23586);
assign n15364 = ~(n13349 | n8856);
assign n9935 = ~n7131;
assign n13817 = ~(n1182 | n2743);
assign n23770 = n5590 | n18682;
assign n25069 = ~(n17442 ^ n15424);
assign n4518 = ~n21760;
assign n9435 = ~(n7512 ^ n6133);
assign n1218 = n16358 & n21331;
assign n13228 = n1219 & n3374;
assign n928 = n12369 & n15646;
assign n23948 = n15747 | n11994;
assign n22750 = n3188 & n9862;
assign n16645 = ~(n19282 ^ n2978);
assign n2430 = n21421 | n16647;
assign n17098 = ~n15883;
assign n1447 = ~(n8155 | n17287);
assign n25938 = ~(n21447 ^ n7779);
assign n13318 = n16824 | n25353;
assign n3733 = ~(n17952 ^ n22756);
assign n1054 = ~(n2914 | n13914);
assign n26595 = n17352 | n4043;
assign n7287 = n19157 | n12138;
assign n6453 = ~(n11211 ^ n26522);
assign n15243 = ~(n2160 ^ n19282);
assign n8955 = ~(n13425 | n22215);
assign n6646 = n1018 | n2616;
assign n24860 = ~(n24070 ^ n661);
assign n18310 = ~(n25961 ^ n15225);
assign n4551 = n10898 & n25750;
assign n24834 = ~(n25370 ^ n4426);
assign n3580 = n18407 & n18866;
assign n11092 = n8255 & n5;
assign n6428 = n26268 | n1258;
assign n25185 = n15876 & n22367;
assign n26786 = ~n26422;
assign n15565 = n586 ^ n21226;
assign n26995 = n13086 & n14303;
assign n7812 = n1654 | n24245;
assign n2347 = n17100 | n24390;
assign n13128 = n23230 | n20488;
assign n13622 = ~(n18371 ^ n21151);
assign n23666 = n18344 & n2965;
assign n3554 = ~(n15777 ^ n5857);
assign n1148 = n119 & n20459;
assign n11674 = ~(n550 ^ n7928);
assign n1265 = ~(n11382 | n17607);
assign n19215 = ~n20530;
assign n19142 = ~(n2944 ^ n22270);
assign n18242 = n15640 | n1221;
assign n19984 = n14856 | n11192;
assign n24347 = ~(n19124 ^ n6897);
assign n24858 = n25201 | n4057;
assign n181 = n11043 & n25117;
assign n6692 = n2324;
assign n1778 = ~(n4003 ^ n17959);
assign n10954 = n13670 & n17029;
assign n9322 = ~(n14265 ^ n25667);
assign n10316 = ~(n9003 ^ n13453);
assign n11811 = n8326 & n26456;
assign n13889 = ~(n8638 | n23018);
assign n11767 = ~n3535;
assign n5700 = ~(n6396 ^ n26740);
assign n27116 = n1672 | n16765;
assign n22426 = ~n14575;
assign n9178 = n12900 | n16547;
assign n25080 = ~(n7841 ^ n22918);
assign n168 = n12094 | n25724;
assign n3391 = ~n21626;
assign n5813 = ~(n17250 ^ n10125);
assign n19117 = ~(n23 ^ n20626);
assign n23071 = ~n18466;
assign n26008 = ~n19638;
assign n23419 = ~(n21937 | n11736);
assign n3327 = ~(n17739 | n4400);
assign n15261 = ~(n19960 ^ n16140);
assign n18473 = ~n2731;
assign n18520 = ~(n4245 ^ n18577);
assign n17741 = ~(n7217 ^ n8324);
assign n26707 = ~(n21662 ^ n14943);
assign n26472 = n9204 & n12251;
assign n1714 = ~(n12972 ^ n16719);
assign n6892 = n15628 & n21722;
assign n6757 = n26415 | n24088;
assign n15599 = ~(n8625 | n7291);
assign n26717 = ~n12161;
assign n26484 = ~(n6179 ^ n18345);
assign n11489 = ~(n14062 ^ n8837);
assign n7902 = ~n25864;
assign n379 = ~(n26009 ^ n7354);
assign n1248 = n3173 | n2841;
assign n26176 = n750 & n11520;
assign n3698 = ~(n18287 | n406);
assign n25515 = ~(n3434 ^ n2301);
assign n26809 = ~(n14113 | n8172);
assign n15583 = ~n18877;
assign n22563 = ~(n6204 ^ n3795);
assign n17116 = ~(n5213 | n24617);
assign n26997 = ~n11044;
assign n20227 = n15838 & n2398;
assign n24052 = ~(n10932 ^ n26764);
assign n5019 = ~(n2780 | n10411);
assign n25355 = ~(n16535 ^ n15908);
assign n21791 = n5704 & n24665;
assign n20057 = ~(n20970 ^ n13367);
assign n26255 = ~n21078;
assign n2199 = ~(n5990 ^ n21208);
assign n8784 = ~(n18492 ^ n12813);
assign n17254 = ~(n20536 | n3349);
assign n18836 = n9103 & n3342;
assign n11855 = ~(n12861 | n15064);
assign n3573 = ~(n2675 ^ n5139);
assign n6286 = n2836 & n18436;
assign n14923 = ~n19982;
assign n3567 = n1541 | n25495;
assign n26640 = ~(n20009 | n23980);
assign n15786 = n20251 | n10942;
assign n17831 = ~(n22222 | n7761);
assign n16674 = ~(n26010 ^ n6661);
assign n25149 = n7111 | n926;
assign n15319 = ~(n5451 ^ n3918);
assign n25040 = n4304 & n19413;
assign n6859 = ~(n22218 ^ n3431);
assign n24862 = ~n23612;
assign n7767 = ~(n21764 ^ n5483);
assign n10934 = ~n9504;
assign n13773 = n3468 | n15289;
assign n5895 = ~(n3582 | n21784);
assign n10666 = ~n5167;
assign n21423 = ~(n23352 | n25659);
assign n18327 = ~(n18338 | n18672);
assign n15055 = ~(n13783 | n22332);
assign n4335 = n25566 | n3581;
assign n12954 = n14486 | n18735;
assign n15875 = ~n2233;
assign n24902 = ~n16374;
assign n23267 = n6935 | n16808;
assign n6282 = n2812 | n8363;
assign n18697 = n14402 | n20785;
assign n21449 = ~(n25015 ^ n1850);
assign n5282 = n16872 | n25027;
assign n8904 = n21450 & n4870;
assign n11384 = ~n25923;
assign n25568 = ~(n19772 ^ n6866);
assign n15779 = ~(n10995 ^ n11736);
assign n14387 = ~(n986 ^ n3122);
assign n22896 = n20037 | n1207;
assign n8951 = n23125 & n15080;
assign n14685 = ~(n8512 ^ n2819);
assign n10909 = ~(n306 | n13936);
assign n8521 = ~(n9132 ^ n3611);
assign n4015 = ~(n20120 ^ n13129);
assign n15267 = ~n15475;
assign n21397 = ~(n790 ^ n5914);
assign n4750 = n18408 | n4283;
assign n22476 = ~(n21937 ^ n10706);
assign n26185 = ~(n21 ^ n23513);
assign n2799 = n19531 & n26872;
assign n1153 = n14173 & n9772;
assign n9195 = n15173 | n6415;
assign n27014 = n9956 | n24294;
assign n15193 = ~n24496;
assign n6326 = n26423 | n21530;
assign n5921 = n458 & n26101;
assign n13808 = ~(n25330 ^ n15167);
assign n10051 = ~(n2379 ^ n15319);
assign n4318 = n14899 & n10408;
assign n16740 = n12688 | n26249;
assign n13392 = ~(n20707 | n9780);
assign n9839 = n22273 | n9605;
assign n6449 = n21756 | n17178;
assign n2775 = ~n5236;
assign n4332 = n6120 | n23197;
assign n14560 = ~(n5990 | n21208);
assign n12415 = n13763 & n118;
assign n7519 = ~(n20376 ^ n6202);
assign n7527 = n23219 & n23764;
assign n25037 = n17741 & n10451;
assign n15653 = n23029 | n17840;
assign n25762 = ~(n8496 | n1574);
assign n5214 = ~(n18994 ^ n2100);
assign n17529 = ~(n662 ^ n18736);
assign n19391 = ~n3836;
assign n9154 = n3622 | n15764;
assign n24969 = ~(n2493 ^ n9442);
assign n23276 = ~(n14936 | n5740);
assign n10585 = ~(n21489 ^ n4085);
assign n16070 = n10580 & n12084;
assign n15959 = ~n7216;
assign n23027 = n13237 | n1066;
assign n23567 = ~(n26939 ^ n20259);
assign n13647 = n23912 | n22716;
assign n16434 = n22687 | n11734;
assign n20624 = ~(n4612 ^ n7118);
assign n12350 = ~(n14244 ^ n16705);
assign n17721 = ~(n24525 ^ n22267);
assign n15427 = ~n16994;
assign n5808 = n5942 | n7023;
assign n22023 = n3623 | n6444;
assign n15532 = n12161 | n24886;
assign n3495 = ~(n3460 | n19477);
assign n12149 = ~n22557;
assign n5835 = n11183 & n16891;
assign n192 = n23119 | n16591;
assign n6660 = ~n6371;
assign n22446 = n26512 | n4909;
assign n10034 = ~(n87 ^ n10129);
assign n13807 = ~(n6239 | n20209);
assign n14053 = n379 | n20671;
assign n10523 = n10916 | n5835;
assign n21029 = ~n18107;
assign n24329 = ~n21884;
assign n5807 = n16791 | n26967;
assign n14748 = n22751 | n6505;
assign n25692 = ~n14458;
assign n3933 = n16227 | n21226;
assign n2359 = n9034 & n19959;
assign n11642 = n3134 | n24135;
assign n11094 = ~(n23941 ^ n11196);
assign n23260 = n25571 | n7978;
assign n4828 = ~(n6200 ^ n14257);
assign n16993 = ~(n21503 ^ n20269);
assign n2892 = ~(n3199 ^ n22782);
assign n14891 = ~(n27203 ^ n25202);
assign n5472 = ~(n1321 ^ n2665);
assign n7196 = n16103 | n4990;
assign n7907 = ~(n20411 | n9512);
assign n24848 = n6613 & n8933;
assign n14429 = n13664 & n6197;
assign n20178 = ~(n25120 | n8526);
assign n14799 = ~(n1534 | n6201);
assign n8607 = ~n25455;
assign n1408 = n17782 | n16782;
assign n21639 = n14966 | n19370;
assign n23563 = n26782 | n11069;
assign n13754 = ~(n27034 ^ n11995);
assign n328 = ~n24032;
assign n26629 = ~n1183;
assign n7833 = ~(n25366 ^ n25949);
assign n17224 = n5714 & n26409;
assign n23566 = n10156 & n20551;
assign n7225 = n13935 | n11841;
assign n4763 = n3749 | n21342;
assign n9084 = ~(n21089 ^ n23086);
assign n1563 = ~(n25040 | n9060);
assign n6446 = ~n851;
assign n23540 = n23923 & n23874;
assign n19460 = n1092;
assign n15132 = ~(n25357 ^ n15499);
assign n17490 = n17177 & n18712;
assign n11769 = n4740 & n26614;
assign n16173 = n7340 | n24448;
assign n1061 = ~n23201;
assign n26826 = ~(n9814 ^ n9274);
assign n119 = n18256 | n14958;
assign n13251 = ~(n24624 ^ n17090);
assign n18663 = n2371 | n14713;
assign n1983 = n25788 & n8697;
assign n2625 = n21301 & n8912;
assign n8440 = n15796 | n4836;
assign n1696 = n15321 | n1652;
assign n20203 = n22030 | n3754;
assign n13880 = n1954 | n4575;
assign n14882 = ~(n13621 | n16130);
assign n11992 = n14570 | n1528;
assign n288 = n16824 & n26295;
assign n13631 = ~(n9940 ^ n8013);
assign n12839 = n6004 & n18567;
assign n6549 = n6195 | n20608;
assign n8730 = n2775 & n22852;
assign n4747 = n18902 | n8643;
assign n18644 = ~(n19472 ^ n21226);
assign n24880 = ~n10787;
assign n4370 = ~(n26810 ^ n26660);
assign n12306 = ~n7837;
assign n25429 = n8998 | n25378;
assign n3576 = n6701 | n7195;
assign n5787 = ~(n24118 ^ n13271);
assign n3406 = n23231 | n10114;
assign n16998 = n1630 | n16147;
assign n9116 = n5877 & n11626;
assign n1073 = n777 | n3433;
assign n264 = n12016 | n17756;
assign n27178 = ~(n7428 | n17169);
assign n11716 = n8118 | n14359;
assign n10484 = ~(n18160 ^ n687);
assign n17906 = ~n14265;
assign n11505 = n24646 | n4288;
assign n18859 = ~(n18468 ^ n11639);
assign n778 = ~n13044;
assign n19340 = ~n22358;
assign n612 = n25930 | n15940;
assign n18775 = n23912 & n22716;
assign n26218 = ~n7850;
assign n16978 = ~(n16468 ^ n12720);
assign n18218 = ~(n7070 ^ n21661);
assign n8150 = ~(n17266 | n9151);
assign n8386 = n14339 | n25705;
assign n17580 = n10914 | n25014;
assign n1555 = ~(n7041 ^ n393);
assign n16614 = n13443 | n13783;
assign n5547 = ~n9598;
assign n21999 = ~n15710;
assign n10628 = ~(n13937 ^ n10836);
assign n18743 = ~(n10411 ^ n8309);
assign n3026 = n7119 | n14544;
assign n21920 = n321 | n16577;
assign n16267 = ~n10843;
assign n863 = ~(n2610 ^ n9406);
assign n24599 = ~(n13240 ^ n18897);
assign n18543 = n4796 | n20828;
assign n234 = ~n15977;
assign n16161 = n22173 | n17932;
assign n1455 = n26909 & n17618;
assign n25705 = n2392 & n9061;
assign n18696 = n6723 & n5370;
assign n6374 = n171 & n15680;
assign n16137 = n12738 & n10615;
assign n12379 = ~(n25422 ^ n6388);
assign n17196 = ~(n18643 ^ n15313);
assign n12923 = ~n14704;
assign n6913 = n11280 & n6479;
assign n1009 = ~n19196;
assign n19274 = ~(n24051 ^ n18158);
assign n5036 = ~n14391;
assign n13752 = ~(n8110 ^ n23691);
assign n18919 = ~(n18567 ^ n2164);
assign n3656 = n6090 & n17429;
assign n11102 = ~(n19110 | n10522);
assign n12044 = n19152 | n22567;
assign n13952 = n11125 | n22203;
assign n23856 = n10084 | n4372;
assign n18914 = ~(n17056 | n2109);
assign n21840 = n9515 & n19559;
assign n13893 = ~n8753;
assign n1493 = n3064 & n22746;
assign n22421 = ~n16290;
assign n25572 = ~n649;
assign n17230 = ~n6729;
assign n8701 = ~(n20056 ^ n11135);
assign n9865 = n18344 | n2965;
assign n21137 = ~n1097;
assign n26393 = n20040 | n23983;
assign n22912 = ~n3606;
assign n745 = n26739 & n24046;
assign n14878 = ~(n24720 ^ n4175);
assign n24677 = n1880 | n25227;
assign n21792 = ~(n15077 | n24112);
assign n17017 = ~(n23854 | n25533);
assign n13064 = n24051 | n20989;
assign n21830 = n3738 & n20193;
assign n26905 = ~(n21296 ^ n23229);
assign n4922 = ~n13175;
assign n25628 = n146 & n6832;
assign n20104 = ~(n21619 ^ n22974);
assign n4259 = ~(n814 ^ n4121);
assign n14572 = ~(n19170 | n3608);
assign n18847 = ~n8119;
assign n1858 = n6267 | n18319;
assign n4038 = ~n16291;
assign n20723 = ~(n14388 ^ n19892);
assign n21977 = ~n19583;
assign n4584 = n6373 | n13567;
assign n17400 = n2903 | n22015;
assign n5706 = ~(n5047 ^ n9934);
assign n16673 = n26086 | n19144;
assign n5954 = ~(n22539 ^ n6798);
assign n17363 = n22403 | n22681;
assign n18371 = ~n13844;
assign n15460 = n3745 | n21074;
assign n16865 = n10854 | n21969;
assign n22801 = n8381 | n23775;
assign n18555 = n26691 & n7563;
assign n21867 = ~n20259;
assign n22449 = n18423 & n19029;
assign n10658 = n14899 | n23308;
assign n5037 = ~(n2242 | n6449);
assign n10513 = ~n18421;
assign n21334 = n23563 & n21699;
assign n12061 = n25690 | n7273;
assign n2441 = n26062 | n25068;
assign n7648 = n21107 | n4675;
assign n15465 = ~(n2204 ^ n20252);
assign n4007 = ~(n17752 ^ n8383);
assign n24176 = ~(n8771 ^ n7897);
assign n3678 = n13977 | n15006;
assign n24310 = ~(n3097 | n26667);
assign n26605 = ~(n14500 ^ n26784);
assign n19480 = n26701 & n4233;
assign n19508 = n5560 | n16944;
assign n26133 = ~(n20923 | n5288);
assign n16400 = ~n24485;
assign n25631 = ~(n4869 ^ n11317);
assign n6831 = ~n14282;
assign n10292 = n6104 | n19985;
assign n10562 = n19962 | n12955;
assign n9137 = n680 & n4948;
assign n5314 = n6352 | n21288;
assign n15338 = ~(n3570 | n575);
assign n21504 = ~(n3506 ^ n9934);
assign n8442 = n9396 | n11817;
assign n9944 = ~n25471;
assign n11456 = ~(n5495 | n9366);
assign n19506 = n3260 | n20512;
assign n25930 = ~n13190;
assign n10390 = ~(n19290 ^ n20872);
assign n27155 = n15489 & n6471;
assign n24509 = n23741 & n12977;
assign n14270 = n24276 | n578;
assign n4542 = n1238;
assign n21310 = n20032 | n19227;
assign n22978 = ~(n15534 | n25572);
assign n27017 = ~(n14183 ^ n11509);
assign n3967 = ~n15521;
assign n19848 = n16427 & n1807;
assign n11380 = ~(n17230 | n3447);
assign n9330 = n7581 | n16933;
assign n10848 = n3368 & n23531;
assign n12485 = ~(n9399 | n9507);
assign n16575 = ~(n5451 | n3918);
assign n13252 = n831 & n5871;
assign n17849 = n23603 | n9720;
assign n22623 = n3734 | n10487;
assign n20721 = n7457 & n32;
assign n2697 = ~(n725 ^ n7759);
assign n4068 = n20246 & n6017;
assign n26763 = n15380 | n22576;
assign n21724 = n3457 & n15181;
assign n5417 = ~n7376;
assign n12931 = ~(n1759 ^ n25331);
assign n3773 = n286 | n13379;
assign n4929 = ~(n26529 ^ n17204);
assign n6604 = n7561 | n2849;
assign n13052 = n24004 | n21081;
assign n4246 = n22297 & n1633;
assign n6239 = ~n24425;
assign n1869 = ~(n22281 ^ n8537);
assign n13473 = ~(n21288 ^ n25238);
assign n22539 = n15632 & n5278;
assign n5152 = n698 | n18404;
assign n2351 = n26056 | n9314;
assign n11551 = ~n20001;
assign n8214 = ~(n5506 ^ n20923);
assign n25275 = n25837 | n5481;
assign n5315 = n11144 | n12702;
assign n25662 = n4691 | n4988;
assign n12008 = n1795 & n10824;
assign n27107 = ~n22465;
assign n13946 = n25643 | n27141;
assign n24619 = n20914 & n4528;
assign n11161 = ~(n6825 ^ n21498);
assign n7381 = n11903 | n14872;
assign n9619 = n23702 & n1038;
assign n7216 = ~(n25537 ^ n14971);
assign n9959 = n17151 | n3572;
assign n7964 = n13862 | n23976;
assign n4078 = n3217 | n3746;
assign n27171 = n16188 & n1566;
assign n1766 = n12143 | n1351;
assign n15166 = n7936 & n2962;
assign n4790 = n16488 & n5725;
assign n14582 = n15022 | n13125;
assign n2090 = ~n18302;
assign n3273 = n5183 | n4448;
assign n12529 = ~(n19116 ^ n3945);
assign n6950 = n7935 & n11552;
assign n8165 = ~(n19194 ^ n14805);
assign n11114 = n26241 & n918;
assign n13351 = ~(n22358 | n9597);
assign n15470 = ~(n27123 ^ n6884);
assign n9740 = ~(n15405 | n2223);
assign n10251 = ~n693;
assign n21282 = n9779 | n20205;
assign n7391 = ~(n23193 ^ n14154);
assign n26376 = n8298 | n5124;
assign n12442 = ~(n9671 | n19042);
assign n81 = ~(n9246 ^ n7876);
assign n25583 = n21467 | n23870;
assign n19568 = ~(n24082 ^ n11447);
assign n4083 = ~n10320;
assign n10590 = ~(n15584 ^ n21030);
assign n25187 = n6764 | n8344;
assign n13546 = ~(n16016 | n14365);
assign n24371 = ~n2139;
assign n1359 = n16476 & n19;
assign n7961 = n6262 | n18975;
assign n6885 = ~(n13333 ^ n9512);
assign n22116 = ~(n2045 | n19228);
assign n9376 = ~(n23404 ^ n7753);
assign n1117 = ~(n25643 ^ n20604);
assign n8162 = ~n22282;
assign n24281 = ~(n17162 ^ n17147);
assign n19260 = ~(n18814 | n25471);
assign n17928 = ~(n27084 ^ n19696);
assign n24662 = ~(n5715 | n20554);
assign n19000 = ~(n27188 | n4326);
assign n18048 = n10889 & n6696;
assign n24853 = ~(n15609 ^ n1560);
assign n15978 = n16180 & n19463;
assign n26872 = ~(n204 ^ n14704);
assign n1517 = n21128 | n13252;
assign n2990 = ~(n22332 ^ n7751);
assign n5746 = ~n11932;
assign n5068 = ~(n11740 | n3591);
assign n26754 = ~(n21749 ^ n919);
assign n21328 = ~(n6734 ^ n19404);
assign n13913 = ~n5208;
assign n7628 = n22975 | n18144;
assign n8441 = ~(n26021 ^ n4984);
assign n14505 = n14604 & n2851;
assign n20393 = ~n14156;
assign n25173 = ~(n5708 ^ n1181);
assign n9501 = n6229 | n7212;
assign n15159 = n23198 | n10822;
assign n17499 = n12618 & n7595;
assign n145 = ~(n23509 ^ n7731);
assign n12262 = ~n6359;
assign n25134 = n2125 | n20829;
assign n11748 = n5512 | n18962;
assign n5360 = ~(n21200 ^ n18549);
assign n6395 = n17664 & n21253;
assign n8160 = n2917 & n3771;
assign n4016 = n2605 & n3683;
assign n23242 = ~n4391;
assign n13047 = n19513 | n22137;
assign n21469 = ~n7391;
assign n8345 = ~(n5043 | n18133);
assign n15561 = n902 | n19620;
assign n24552 = ~n13708;
assign n16757 = n11377 | n16611;
assign n2661 = n25981 | n27003;
assign n11154 = n14814 | n6419;
assign n1510 = ~(n516 ^ n10020);
assign n2568 = ~(n226 ^ n18544);
assign n8980 = ~n13250;
assign n25132 = n18765 & n4659;
assign n22145 = n16880 | n18357;
assign n6354 = ~(n13218 ^ n17472);
assign n488 = n25586 & n8491;
assign n15802 = n11449 | n26154;
assign n24989 = ~(n4086 ^ n8724);
assign n8572 = ~n4708;
assign n23007 = ~(n20979 ^ n10779);
assign n17326 = n7305 | n830;
assign n8364 = n16563 & n9334;
assign n15411 = ~(n4641 ^ n7746);
assign n24251 = n25078 & n3023;
assign n25468 = ~(n21011 ^ n16299);
assign n9248 = n8256 | n17815;
assign n4983 = n21 | n23513;
assign n7558 = ~(n20540 ^ n26126);
assign n593 = n13220;
assign n10441 = ~n5182;
assign n16921 = n20650 & n4968;
assign n26586 = n21581 & n14741;
assign n9979 = ~(n23333 ^ n16502);
assign n19255 = ~n25659;
assign n13720 = n25237 | n13336;
assign n23329 = ~n14661;
assign n11371 = n21583 & n16756;
assign n11128 = ~(n4613 ^ n10076);
assign n20122 = n26596 | n6399;
assign n13491 = ~(n13494 ^ n3425);
assign n24892 = ~(n21471 | n24612);
assign n19171 = n13026 & n13906;
assign n16075 = n27048 | n24530;
assign n2166 = n19097 & n5333;
assign n20987 = n10373 | n25082;
assign n27141 = n9557 | n21944;
assign n2534 = ~(n8195 ^ n19935);
assign n4591 = ~n3214;
assign n7573 = ~(n1705 ^ n5354);
assign n2471 = n1106 | n26770;
assign n20193 = n4996 | n26669;
assign n16518 = n22111 & n13971;
assign n16841 = ~(n7637 ^ n3377);
assign n20677 = n14171 | n16739;
assign n24613 = n23647 & n24465;
assign n19878 = n23773 | n9358;
assign n14888 = ~(n3606 ^ n7484);
assign n20543 = n8843 & n9071;
assign n8505 = ~(n8157 ^ n22899);
assign n15846 = ~(n24628 ^ n9322);
assign n14706 = ~(n16058 ^ n18532);
assign n2615 = ~(n26260 ^ n4139);
assign n11682 = ~(n11969 ^ n7302);
assign n16748 = n1009 & n4999;
assign n5671 = n20988 | n26955;
assign n3856 = ~(n7008 | n25810);
assign n10462 = n11311 & n12903;
assign n26593 = n13591 | n3909;
assign n14709 = n25326 | n17752;
assign n25166 = ~(n7670 ^ n3253);
assign n3401 = n19032 | n23802;
assign n19407 = n13408 | n2450;
assign n18529 = n14625 | n2210;
assign n22091 = ~(n13852 ^ n4009);
assign n20395 = n3315 | n6214;
assign n9626 = ~(n14021 ^ n14202);
assign n7458 = n22666 | n18148;
assign n15815 = ~(n2182 ^ n12814);
assign n9481 = n19624 | n14625;
assign n20967 = ~(n15266 ^ n3506);
assign n1990 = n7623 | n16736;
assign n12547 = ~n18905;
assign n22515 = ~n13220;
assign n15048 = n26757 & n12504;
assign n11666 = n1896 | n11457;
assign n10721 = n7496 & n12151;
assign n9023 = n8338 & n3967;
assign n10726 = n17836 | n9684;
assign n18387 = n26560 & n9272;
assign n11179 = ~(n401 | n14519);
assign n10274 = ~n23369;
assign n9452 = ~(n25739 ^ n26443);
assign n20241 = n17062 & n21906;
assign n16894 = n16261 | n23013;
assign n25902 = n19387 & n1395;
assign n6219 = ~(n19303 ^ n8782);
assign n26646 = n8416 | n101;
assign n11803 = ~(n16261 ^ n24188);
assign n19247 = ~(n9562 ^ n19409);
assign n26189 = ~(n215 ^ n14702);
assign n5125 = n24686 | n9889;
assign n5648 = n19197 & n26099;
assign n21515 = n22411 | n3951;
assign n1732 = n1242 | n21031;
assign n17645 = ~n5521;
assign n27197 = n25405 ^ n20406;
assign n4881 = n5767 | n23435;
assign n15073 = ~n20505;
assign n4998 = n21905 | n24481;
assign n7036 = n16655 & n3339;
assign n9001 = n19427 | n18500;
assign n25592 = ~(n13352 ^ n2233);
assign n5059 = n13782 & n9568;
assign n2048 = ~n7924;
assign n8817 = ~(n12125 ^ n25327);
assign n6107 = ~(n24851 ^ n12495);
assign n2172 = n12513 | n14106;
assign n21583 = n9180 | n2514;
assign n20816 = n23788 | n4249;
assign n17855 = ~(n1818 ^ n13557);
assign n11439 = ~(n3360 ^ n26006);
assign n24320 = ~(n11930 ^ n1277);
assign n2826 = ~(n5241 ^ n1177);
assign n2422 = ~(n14462 ^ n5784);
assign n12920 = ~(n25991 ^ n1840);
assign n25007 = ~n23187;
assign n2945 = n2099 | n21948;
assign n10749 = ~n9413;
assign n10750 = ~(n24645 ^ n13714);
assign n26498 = ~n5450;
assign n12686 = ~(n15693 | n21626);
assign n15974 = ~(n12068 | n4558);
assign n5111 = ~(n15414 ^ n23610);
assign n5331 = ~(n25007 | n19048);
assign n20796 = ~n8079;
assign n1045 = n17631 & n24068;
assign n5530 = ~n1344;
assign n17350 = ~n22456;
assign n6097 = n6613 | n8933;
assign n19219 = n13528 | n12373;
assign n7289 = n681 & n18491;
assign n4250 = n23438 & n7603;
assign n15864 = ~(n1536 | n21743);
assign n11453 = ~n23026;
assign n5087 = n22740 | n24169;
assign n890 = ~(n17605 ^ n25533);
assign n10605 = ~(n5934 ^ n7776);
assign n6822 = ~(n17716 ^ n14704);
assign n18628 = ~(n18452 ^ n1752);
assign n13202 = ~(n972 ^ n11155);
assign n4464 = ~(n13489 ^ n20575);
assign n22647 = n15075 & n19800;
assign n959 = ~n9966;
assign n23191 = n21801 & n15597;
assign n3998 = n13392 | n23394;
assign n26494 = n19277 | n13963;
assign n15181 = n18209 | n8047;
assign n15086 = n11069 | n6743;
assign n7304 = n17439 | n24966;
assign n19028 = ~n19786;
assign n21896 = ~n22634;
assign n3256 = ~(n3809 | n8406);
assign n16432 = n1715 & n19371;
assign n5927 = ~(n7153 ^ n15325);
assign n17105 = n9713 & n1471;
assign n13334 = n15900 | n15351;
assign n21726 = ~(n3184 ^ n7209);
assign n17483 = ~n7436;
assign n2733 = n20642 | n22932;
assign n6889 = n12453 | n2908;
assign n631 = ~(n8786 ^ n25381);
assign n8785 = n16998 & n10134;
assign n3015 = ~n5701;
assign n14421 = ~(n3861 ^ n6631);
assign n21629 = ~(n20043 ^ n20986);
assign n23946 = n740 | n14318;
assign n19070 = ~(n17605 ^ n4263);
assign n14068 = n16464 | n4844;
assign n12655 = ~(n3405 | n24165);
assign n1882 = ~n12754;
assign n4175 = ~(n16812 ^ n25923);
assign n4307 = ~n17159;
assign n18065 = ~(n16077 ^ n26300);
assign n8306 = ~(n12721 ^ n13465);
assign n5877 = n8773 | n11657;
assign n14361 = ~(n24246 ^ n14883);
assign n18036 = ~(n16993 ^ n24601);
assign n22089 = ~(n23849 | n19702);
assign n19439 = ~(n2995 | n15678);
assign n27070 = ~(n575 ^ n22198);
assign n18101 = ~(n11378 | n22110);
assign n25614 = ~(n11383 ^ n16859);
assign n15303 = ~(n21071 ^ n8945);
assign n11903 = ~(n10808 ^ n3077);
assign n15767 = n271;
assign n23050 = ~n4115;
assign n19609 = n10169 & n7133;
assign n6539 = n17005 | n12117;
assign n17791 = ~(n8006 ^ n19514);
assign n26083 = n10265 | n241;
assign n19396 = ~(n1336 ^ n3843);
assign n12982 = n10003 | n8929;
assign n9574 = ~n6658;
assign n117 = ~(n11209 ^ n5495);
assign n18700 = ~n26608;
assign n20910 = n14146 & n2437;
assign n20255 = n11357 & n10286;
assign n12218 = ~(n13190 | n9318);
assign n18308 = n6338 & n3070;
assign n11138 = ~(n264 ^ n1261);
assign n17998 = ~(n14159 ^ n5770);
assign n18909 = ~(n22226 ^ n23430);
assign n11540 = n7062 & n14349;
assign n5841 = ~(n24971 ^ n9687);
assign n27199 = ~n17959;
assign n12392 = n19297 | n24042;
assign n4026 = ~(n20196 ^ n26748);
assign n11033 = ~(n20032 | n25974);
assign n1515 = n6764 | n6611;
assign n9769 = n12122 | n19320;
assign n14332 = n12468 | n22224;
assign n16581 = n21019 & n10433;
assign n3483 = ~(n23729 ^ n22597);
assign n735 = ~(n5227 ^ n2140);
assign n21012 = n25334 | n18978;
assign n92 = n5077 | n12739;
assign n9755 = n18504 & n17483;
assign n397 = n13757 | n25654;
assign n10199 = ~(n23292 ^ n11423);
assign n4172 = ~(n7611 ^ n6342);
assign n23551 = ~(n2057 ^ n21930);
assign n11732 = ~(n7305 | n23061);
assign n15606 = n25897 | n17573;
assign n13794 = ~(n8285 ^ n20036);
assign n22391 = ~(n21450 ^ n24821);
assign n600 = n20393 | n26832;
assign n2548 = n26572 | n4029;
assign n7203 = n505 | n9748;
assign n463 = ~(n11437 ^ n13740);
assign n3949 = ~n1543;
assign n9002 = ~(n9940 ^ n11455);
assign n17972 = ~(n21824 ^ n15820);
assign n13732 = ~(n20365 ^ n14127);
assign n3298 = ~(n17005 ^ n25303);
assign n8226 = ~(n23032 ^ n22863);
assign n19381 = n5723 & n6324;
assign n20102 = ~(n7659 ^ n7031);
assign n2950 = ~(n2206 ^ n24412);
assign n23767 = ~(n20526 ^ n24139);
assign n17916 = n8943 | n9683;
assign n3636 = n24972 & n5429;
assign n13698 = ~(n24125 ^ n20639);
assign n18545 = ~(n14158 ^ n5140);
assign n22365 = ~n12587;
assign n19137 = ~(n4096 ^ n22778);
assign n7496 = ~(n11722 ^ n1316);
assign n492 = ~(n21420 ^ n9820);
assign n11603 = ~n863;
assign n202 = n17701 | n10531;
assign n6495 = ~(n23865 ^ n19200);
assign n17988 = n22074 | n15484;
assign n5132 = n17212 & n14634;
assign n19103 = ~(n17762 ^ n22433);
assign n8538 = ~(n22964 | n21060);
assign n11709 = n7328 | n20493;
assign n26344 = n24873;
assign n1769 = n25139 | n1794;
assign n4956 = ~(n8201 ^ n20317);
assign n2208 = ~n2221;
assign n25996 = ~(n21378 ^ n25972);
assign n21913 = n15782 & n14334;
assign n5393 = n26957 | n18662;
assign n24107 = n604 | n4626;
assign n4736 = ~(n22597 ^ n18901);
assign n19375 = n6750 & n13328;
assign n10335 = n6894 & n2894;
assign n3043 = n8568 & n13140;
assign n12176 = n3091 | n26031;
assign n9610 = n13225 & n10115;
assign n22545 = n2915 & n23559;
assign n19350 = n22626 & n25038;
assign n677 = ~(n9052 ^ n4982);
assign n16826 = n19944 | n1451;
assign n17405 = ~(n20077 ^ n22433);
assign n6164 = ~(n1093 ^ n3718);
assign n18216 = ~(n832 | n23506);
assign n4114 = n10005 & n12691;
assign n7636 = ~(n25089 ^ n11721);
assign n21305 = n19074 | n8581;
assign n16182 = ~(n3239 ^ n1464);
assign n9575 = ~(n24920 ^ n26806);
assign n20953 = n15674 & n17270;
assign n2913 = n3081 & n19512;
assign n4539 = ~(n22198 | n8774);
assign n14180 = ~(n8964 ^ n1293);
assign n2836 = n16874 | n18589;
assign n22845 = ~(n7149 | n22871);
assign n14031 = n25345 | n18479;
assign n15975 = ~(n4485 ^ n19906);
assign n4839 = n9050 | n16210;
assign n17878 = n23493 | n8405;
assign n10641 = n16822 | n23329;
assign n20249 = ~n23034;
assign n24911 = ~(n25171 ^ n3577);
assign n7414 = n9779 & n24663;
assign n24154 = ~(n20649 ^ n15565);
assign n3265 = ~(n22782 ^ n24455);
assign n22404 = ~(n16676 ^ n16612);
assign n26645 = n21674 | n5791;
assign n18987 = n7953 & n20908;
assign n17572 = ~n10897;
assign n17745 = n21232 | n7471;
assign n18645 = n18306 & n3303;
assign n19625 = ~(n18107 ^ n10859);
assign n16900 = ~(n14332 ^ n3662);
assign n27117 = ~(n19962 ^ n15508);
assign n3649 = ~(n11532 ^ n8375);
assign n3726 = ~(n111 ^ n17940);
assign n19201 = ~n9246;
assign n15069 = n12751 | n24847;
assign n22669 = ~(n9394 ^ n6039);
assign n7982 = n24130 | n16531;
assign n17679 = ~(n21007 ^ n3018);
assign n8156 = n9210 & n2729;
assign n22265 = ~(n14158 | n11381);
assign n20964 = ~n2289;
assign n2951 = n1650 & n3272;
assign n10268 = n21837 & n25845;
assign n17776 = n5025 | n12771;
assign n7906 = ~n17808;
assign n22069 = ~n11006;
assign n2324 = ~(n13867 ^ n1922);
assign n12943 = n11924 | n13072;
assign n24963 = ~(n11824 | n14152);
assign n22868 = ~(n26054 | n21907);
assign n18679 = ~(n18396 ^ n16923);
assign n18067 = ~(n626 | n21772);
assign n1070 = n16307 & n14742;
assign n639 = n3346 | n8044;
assign n25868 = ~(n755 | n23366);
assign n26012 = n5314 & n25878;
assign n18813 = n15489 | n6471;
assign n25064 = n11279 & n6336;
assign n16530 = n20998 | n22281;
assign n676 = ~n1741;
assign n10113 = n2219 & n8059;
assign n1489 = n14392 & n18164;
assign n14061 = n8780 & n3154;
assign n3436 = ~(n12049 ^ n10464);
assign n15475 = n18176 & n25847;
assign n298 = ~(n14912 ^ n4989);
assign n21185 = n24672 & n12748;
assign n13360 = ~n24969;
assign n14377 = n16787 | n7115;
assign n23878 = n8988;
assign n23576 = n17937 | n11253;
assign n17933 = n23895 & n8491;
assign n2343 = ~(n8397 ^ n23872);
assign n6112 = n11946 & n24033;
assign n23530 = ~(n1568 | n24571);
assign n16616 = n27084 & n11307;
assign n16671 = n14800 | n13824;
assign n12059 = ~(n5143 ^ n9040);
assign n3261 = ~(n24919 ^ n21915);
assign n20251 = n19488 & n18355;
assign n16557 = n4764 | n6043;
assign n5565 = n10067 | n12818;
assign n15644 = ~n5001;
assign n25551 = ~(n16246 | n21119);
assign n18253 = n10406 & n8947;
assign n18930 = ~n22070;
assign n24089 = ~(n3839 | n21774);
assign n3691 = n7625 & n17785;
assign n7755 = ~(n6777 ^ n17362);
assign n9891 = ~(n10951 ^ n8794);
assign n11211 = ~n14907;
assign n9157 = ~(n18345 | n25168);
assign n19026 = n2382 | n22169;
assign n8376 = ~(n5359 ^ n19912);
assign n9397 = n23925 & n16964;
assign n2753 = n17434 & n16737;
assign n8008 = ~n8679;
assign n6970 = ~(n7150 | n22062);
assign n6514 = ~(n10103 ^ n8274);
assign n27200 = ~n17845;
assign n26145 = ~(n5783 | n6682);
assign n5415 = n24550 & n22182;
assign n22031 = ~(n11625 ^ n13959);
assign n9153 = n24587 | n13597;
assign n16535 = n24710 & n16431;
assign n25696 = ~(n15143 ^ n6527);
assign n12894 = ~(n15153 | n9340);
assign n26236 = n14322 & n8726;
assign n16974 = n25863 | n23626;
assign n7536 = ~(n14144 ^ n17478);
assign n13100 = n25886 | n19005;
assign n19784 = n19651 & n6298;
assign n10477 = n10815 | n2655;
assign n8717 = ~(n16631 ^ n17395);
assign n40 = ~(n24211 | n8304);
assign n23131 = ~(n1654 ^ n16482);
assign n4792 = ~n17870;
assign n24096 = ~(n21484 ^ n26639);
assign n19004 = ~(n6200 | n6672);
assign n1475 = n1477 | n3957;
assign n25206 = n5471 | n2864;
assign n3414 = ~(n5801 ^ n1004);
assign n19815 = n20112 | n23746;
assign n16527 = ~(n18741 ^ n3265);
assign n22115 = n9180 | n18754;
assign n26915 = ~(n17057 ^ n27049);
assign n11047 = ~(n26697 ^ n24439);
assign n26843 = n26551 | n22035;
assign n9390 = n11450 & n3489;
assign n1318 = ~n14767;
assign n25668 = n14899 & n18496;
assign n10867 = ~(n25413 ^ n1293);
assign n11584 = ~(n22715 ^ n10023);
assign n2477 = ~n12541;
assign n1803 = ~n26405;
assign n12703 = n13453 | n4434;
assign n10399 = n18428 | n16793;
assign n22756 = ~(n14139 ^ n9358);
assign n6585 = ~(n2244 ^ n543);
assign n11528 = n11211 | n13774;
assign n25489 = ~(n15894 ^ n24378);
assign n5146 = ~(n17381 | n23731);
assign n25988 = n6647 | n9457;
assign n10036 = ~(n24578 | n15417);
assign n22040 = n9598 & n19084;
assign n19051 = ~n19625;
assign n25921 = n1262 & n1084;
assign n12116 = n13190 & n21632;
assign n8168 = n15533 & n18839;
assign n23121 = ~(n9832 | n3959);
assign n3475 = n5745 | n25073;
assign n5112 = ~n12211;
assign n24650 = ~n22597;
assign n10465 = n16225 & n4680;
assign n10629 = ~(n901 ^ n8258);
assign n2710 = n6202 | n2366;
assign n26446 = n475 | n10517;
assign n8047 = n1276 & n5311;
assign n12885 = n3517 & n15377;
assign n11568 = n21803 & n13768;
assign n14890 = n1006 | n6531;
assign n17535 = n6946 | n8485;
assign n1000 = ~n3903;
assign n13774 = ~(n24270 ^ n17958);
assign n22938 = n12167 | n13956;
assign n7175 = ~(n24208 | n2423);
assign n10271 = ~(n23097 ^ n14749);
assign n3105 = n280 | n16214;
assign n6314 = n17562 | n16804;
assign n23967 = ~(n8650 ^ n20826);
assign n7925 = ~n10460;
assign n18892 = ~(n8087 | n14795);
assign n26501 = ~n24592;
assign n26162 = ~n27089;
assign n13331 = n20435 | n10085;
assign n1825 = ~(n16257 | n6861);
assign n21168 = ~(n16220 ^ n4774);
assign n3509 = ~(n18358 ^ n14206);
assign n6335 = ~(n7371 ^ n7438);
assign n15302 = ~(n4659 | n1835);
assign n4800 = ~n15719;
assign n10066 = ~(n1236 | n23717);
assign n9800 = ~(n2341 | n6596);
assign n4783 = n21389 & n413;
assign n22698 = n24941 | n3961;
assign n22655 = ~n13387;
assign n12323 = ~(n17599 ^ n665);
assign n9792 = ~(n21948 ^ n26805);
assign n11237 = n644 | n12868;
assign n18613 = n24791 & n2291;
assign n24301 = ~n20946;
assign n25546 = n12154 & n12103;
assign n25595 = n23074 & n26395;
assign n24574 = n5451 & n1533;
assign n9004 = ~(n18968 ^ n18753);
assign n13374 = n22202 | n19983;
assign n11312 = ~n15268;
assign n14331 = n5852 & n16963;
assign n2030 = ~(n17578 ^ n4085);
assign n22175 = ~(n10833 ^ n9378);
assign n26004 = n26003 & n20166;
assign n16093 = ~(n8994 ^ n14510);
assign n9361 = n1293 & n15921;
assign n17019 = n540 | n9342;
assign n15383 = ~(n6977 ^ n23096);
assign n9897 = ~(n7009 ^ n4300);
assign n3545 = ~(n8964 | n22554);
assign n4022 = ~n21317;
assign n7620 = n13311 | n17332;
assign n19040 = ~(n9935 ^ n22841);
assign n15054 = ~(n12380 | n16638);
assign n4615 = ~(n13842 | n23670);
assign n17709 = n9275 & n25597;
assign n17123 = n13190 | n23999;
assign n12746 = ~(n13528 ^ n4417);
assign n3758 = ~(n5864 ^ n14587);
assign n19835 = ~(n7671 ^ n197);
assign n5762 = n14933 | n17386;
assign n21868 = ~n21912;
assign n18319 = ~(n2541 ^ n1722);
assign n20733 = ~n8439;
assign n25211 = ~(n22660 ^ n21753);
assign n10115 = n381 | n24356;
assign n13309 = ~n19911;
assign n26047 = ~n17200;
assign n17732 = n22895 | n17203;
assign n13018 = ~(n25042 ^ n7421);
assign n1052 = ~(n3780 ^ n5075);
assign n18552 = n5498 | n16544;
assign n3080 = ~(n16713 ^ n17497);
assign n20431 = ~(n3203 ^ n21272);
assign n26564 = ~(n19753 ^ n16369);
assign n11663 = n23328 | n11117;
assign n20242 = n3260 & n21832;
assign n11755 = ~n4485;
assign n21116 = n1902 & n15441;
assign n24493 = ~n7536;
assign n11311 = n3099 | n23418;
assign n1125 = n24544 & n21167;
assign n385 = ~(n20455 ^ n5376);
assign n17613 = ~n5817;
assign n10417 = n17004 & n24496;
assign n24772 = ~(n10773 | n13460);
assign n26952 = n8860 & n4313;
assign n23684 = ~(n19538 ^ n17227);
assign n13173 = n5790 | n14398;
assign n14737 = ~(n3132 ^ n21957);
assign n17924 = n15697 | n7104;
assign n7806 = n18316 & n15480;
assign n19036 = n13440 & n23944;
assign n14791 = ~n21944;
assign n6491 = ~(n1765 ^ n12875);
assign n23064 = n8898;
assign n14091 = ~(n18441 ^ n1117);
assign n20343 = n24761 & n13746;
assign n9432 = ~(n2850 | n19907);
assign n9542 = n25263 | n18387;
assign n22867 = ~(n6051 | n25276);
assign n7570 = ~(n18145 ^ n26191);
assign n23246 = n9131 & n15704;
assign n18655 = ~n5419;
assign n2001 = n16930 & n662;
assign n966 = ~n18720;
assign n27183 = ~n16449;
assign n3001 = ~(n7402 ^ n7305);
assign n20004 = ~(n22219 ^ n11553);
assign n1849 = n1116 | n7646;
assign n20886 = ~n14792;
assign n24233 = n5348 | n19226;
assign n24594 = n3393 | n1465;
assign n15541 = n18090 | n1252;
assign n22538 = ~(n17212 ^ n20411);
assign n4040 = ~n6397;
assign n13587 = ~(n9431 ^ n27076);
assign n2937 = ~(n2213 ^ n26269);
assign n18156 = n15125 | n11929;
assign n2620 = n24562 | n14018;
assign n19577 = ~(n5213 ^ n19081);
assign n20799 = n9470 & n15320;
assign n14628 = ~n20970;
assign n23428 = ~n18035;
assign n571 = ~(n17568 | n2978);
assign n5661 = n7841 | n19595;
assign n18505 = n16473 | n2111;
assign n24116 = ~n24620;
assign n25766 = n17267 & n23517;
assign n22665 = n11237 & n10091;
assign n15771 = n18118 | n1928;
assign n352 = n7123 & n6615;
assign n7346 = ~(n17001 ^ n1784);
assign n2027 = ~n9498;
assign n3718 = ~(n6319 ^ n19836);
assign n1472 = ~(n56 | n20506);
assign n19277 = ~n19081;
assign n23176 = n11208 & n20899;
assign n15759 = n11465 & n21109;
assign n7469 = n10593 | n1662;
assign n9419 = ~(n8357 ^ n17082);
assign n19151 = n14961 | n5520;
assign n22038 = ~(n2013 | n22640);
assign n14851 = n14760 | n6734;
assign n13706 = n20108 | n12411;
assign n20823 = n21781 | n25549;
assign n12598 = n7550 & n7858;
assign n22262 = ~(n18409 ^ n8259);
assign n7240 = ~(n23430 ^ n19081);
assign n23885 = ~(n4888 ^ n1572);
assign n25135 = n19805 | n5125;
assign n11999 = n840 | n19719;
assign n14389 = ~n26177;
assign n8087 = ~(n1206 ^ n4260);
assign n16479 = ~(n4217 ^ n22683);
assign n24920 = ~(n18338 ^ n12644);
assign n12421 = ~n25449;
assign n5616 = ~n12999;
assign n9374 = n3604 | n11815;
assign n14203 = ~(n14465 | n6356);
assign n4680 = n4312 | n21903;
assign n26324 = ~n3823;
assign n6177 = ~(n15633 | n8097);
assign n22688 = ~n12075;
assign n14073 = ~(n1939 | n13818);
assign n22946 = n6938 | n1201;
assign n10321 = ~(n10764 ^ n2253);
assign n25260 = ~n11230;
assign n8845 = ~(n14804 ^ n20579);
assign n27125 = n4614 | n15132;
assign n26945 = ~(n19172 | n7371);
assign n5697 = ~n8511;
assign n20022 = ~(n11550 | n13884);
assign n22180 = n14098 & n18124;
assign n24486 = ~(n17897 ^ n20278);
assign n5242 = n13902 & n3557;
assign n21258 = ~(n5752 ^ n14071);
assign n16807 = ~(n26026 ^ n4905);
assign n11087 = ~(n19005 | n12889);
assign n9680 = ~n2102;
assign n25062 = ~(n16950 ^ n11632);
assign n8703 = n8448 | n15892;
assign n20759 = ~(n4938 | n25345);
assign n18667 = ~(n9748 ^ n3037);
assign n7682 = ~n18409;
assign n8697 = n16326 | n7199;
assign n12180 = n3605 & n2748;
assign n10361 = n6108 & n20911;
assign n5891 = ~n9011;
assign n16102 = n24219 | n8792;
assign n22638 = n916 & n21211;
assign n14606 = ~(n14397 ^ n10125);
assign n23277 = ~(n9278 ^ n5561);
assign n16880 = n9140;
assign n1729 = n23115 & n1849;
assign n6637 = ~(n22084 ^ n4765);
assign n12525 = ~(n3124 | n24170);
assign n14585 = n3938 | n9853;
assign n1507 = n18212 | n15223;
assign n6837 = ~(n7693 ^ n3909);
assign n8 = ~(n26688 | n14256);
assign n12051 = n6218 & n7669;
assign n25959 = n992 & n19311;
assign n14745 = n19761 | n26684;
assign n12092 = n9970 & n24413;
assign n4188 = n19090 | n13085;
assign n8154 = ~(n14130 ^ n468);
assign n21804 = ~n21654;
assign n5294 = n3231 | n3533;
assign n11420 = ~(n8906 ^ n2420);
assign n5332 = ~(n24592 ^ n21291);
assign n15784 = ~(n25582 ^ n17035);
assign n17711 = ~(n11 ^ n20331);
assign n25362 = ~(n14915 ^ n9510);
assign n19774 = n13316 & n6266;
assign n21595 = n11672 | n6401;
assign n7355 = n468 | n22322;
assign n1946 = ~(n16282 ^ n20714);
assign n14018 = n23391 & n6763;
assign n13056 = ~(n11229 ^ n9741);
assign n12765 = ~(n13906 ^ n13026);
assign n9193 = n24552 | n24618;
assign n1744 = n26568 | n13767;
assign n15673 = n1946 | n1629;
assign n12208 = ~n13384;
assign n15030 = n688 | n7674;
assign n17963 = ~(n21747 ^ n25397);
assign n21098 = ~(n11394 ^ n17847);
assign n26545 = ~(n18314 ^ n20635);
assign n13066 = ~n23876;
assign n18165 = n14434 & n14869;
assign n8410 = ~(n12663 | n14974);
assign n26582 = ~(n19564 ^ n7918);
assign n20239 = ~(n26265 ^ n6485);
assign n4452 = n23245 | n3778;
assign n1923 = ~n6955;
assign n27009 = ~n6362;
assign n22824 = ~(n10998 ^ n22793);
assign n5070 = n15578 & n17991;
assign n26394 = n26660 | n3232;
assign n14865 = ~(n16319 ^ n23882);
assign n27114 = ~n18123;
assign n24028 = ~(n15681 ^ n13333);
assign n19272 = n7402 & n23099;
assign n3855 = n4499 | n16136;
assign n20172 = ~(n21710 ^ n6508);
assign n10475 = ~(n25962 | n17468);
assign n14619 = ~(n6209 | n12241);
assign n8171 = n134 | n17702;
assign n49 = ~(n5740 ^ n25770);
assign n14978 = n11452 | n3460;
assign n1637 = ~n8272;
assign n4317 = ~n4104;
assign n18005 = ~(n4479 ^ n23724);
assign n14550 = ~(n24184 ^ n25923);
assign n24738 = n1587 | n13303;
assign n25018 = ~(n19527 ^ n21993);
assign n4553 = ~(n21406 ^ n11165);
assign n9605 = ~(n19687 ^ n6219);
assign n21680 = ~(n16997 ^ n60);
assign n1631 = ~n10219;
assign n26745 = ~(n15907 ^ n24404);
assign n23363 = n25868 | n13200;
assign n9877 = ~n19284;
assign n5158 = ~(n18019 ^ n186);
assign n25577 = n3774 & n1613;
assign n22906 = ~n17636;
assign n24022 = n13897 | n22121;
assign n10596 = ~(n20131 ^ n10048);
assign n9825 = n6400 | n11069;
assign n4388 = n16614 & n4238;
assign n23422 = ~(n12567 ^ n11048);
assign n20107 = ~(n17108 ^ n4008);
assign n9431 = ~(n26286 ^ n16492);
assign n3557 = n12053 | n7527;
assign n17712 = ~(n2565 ^ n23261);
assign n2338 = n12389 & n23143;
assign n148 = ~(n5299 ^ n15546);
assign n13178 = n4623 & n373;
assign n17176 = ~(n21235 ^ n5025);
assign n18390 = n2712 & n26221;
assign n10876 = ~(n10587 | n9163);
assign n23354 = ~(n17672 ^ n2832);
assign n9392 = ~n9901;
assign n8254 = ~(n12971 | n13553);
assign n8346 = n19611 | n22582;
assign n10414 = ~(n17035 | n13206);
assign n20438 = ~n21585;
assign n21074 = n18276 & n17086;
assign n6522 = ~n9022;
assign n17029 = n228 | n9239;
assign n7348 = ~n274;
assign n17548 = n17966 & n5762;
assign n1848 = ~(n11044 | n4325);
assign n17811 = ~(n5673 ^ n16146);
assign n14624 = ~(n26748 | n20196);
assign n14356 = ~n24907;
assign n3 = ~(n16348 ^ n25321);
assign n3489 = n4547 | n7540;
assign n4501 = ~(n5194 ^ n12161);
assign n20360 = n8223 & n10678;
assign n4495 = n26519 | n6194;
assign n19570 = ~(n12782 ^ n17811);
assign n996 = ~(n10571 ^ n9431);
assign n21710 = ~(n1143 ^ n11709);
assign n24111 = ~n20234;
assign n23577 = n9432 | n24803;
assign n4450 = n8018 | n16700;
assign n5830 = n19011 & n22117;
assign n1653 = n23858 & n24702;
assign n18860 = n478 & n19421;
assign n14087 = ~n11047;
assign n575 = ~n6733;
assign n23398 = n12751 | n12696;
assign n21100 = ~(n15427 | n14337);
assign n26208 = ~(n11747 ^ n15161);
assign n8197 = ~n20887;
assign n4969 = ~(n4883 | n27076);
assign n17056 = n22366 | n5550;
assign n21094 = ~(n8438 ^ n3741);
assign n26852 = n17725 | n1562;
assign n21160 = ~(n5211 ^ n21832);
assign n23057 = ~(n7470 | n1730);
assign n19854 = ~(n12248 ^ n1696);
assign n22401 = n12891 | n9266;
assign n24694 = n9719 & n21639;
assign n6843 = ~(n12002 | n11056);
assign n2531 = n25311 & n380;
assign n15579 = n26450 | n6819;
assign n2621 = n992 | n19311;
assign n26405 = ~(n5714 ^ n26409);
assign n19583 = ~(n26979 ^ n18962);
assign n11644 = ~(n13261 ^ n22591);
assign n2019 = n19525 | n25862;
assign n20674 = ~(n26744 | n8456);
assign n18749 = ~n9971;
assign n3336 = n12698 | n18443;
assign n16769 = ~(n25494 ^ n1314);
assign n10003 = ~(n2268 | n4326);
assign n25685 = ~(n23080 ^ n2133);
assign n20610 = ~(n10405 ^ n23974);
assign n8688 = ~(n14869 ^ n24795);
assign n26468 = n16601 | n18580;
assign n359 = ~(n23024 | n10522);
assign n24184 = ~(n15472 ^ n22821);
assign n12299 = ~n11019;
assign n177 = n19437 & n18640;
assign n27087 = n3511 & n11602;
assign n5881 = n25015 | n4890;
assign n19546 = ~(n14431 | n25877);
assign n278 = n8654 & n1094;
assign n6229 = n24370 | n18868;
assign n25473 = n10166 | n26652;
assign n17785 = n15301 | n24789;
assign n6610 = ~n10083;
assign n1370 = ~(n12501 ^ n8067);
assign n12224 = ~(n23396 | n17790);
assign n19449 = n2694 | n7823;
assign n6497 = n26259 & n10016;
assign n16775 = n8155 | n15077;
assign n23034 = ~(n11762 ^ n20190);
assign n22247 = ~n25439;
assign n19737 = ~(n26979 ^ n5704);
assign n26099 = n21036 | n4118;
assign n1958 = n25068 & n17881;
assign n12848 = ~(n342 ^ n14570);
assign n12919 = n7731 | n19858;
assign n8432 = ~(n17429 ^ n22255);
assign n12119 = ~(n17542 ^ n19840);
assign n19715 = n23397 & n5398;
assign n24962 = n11151 & n4295;
assign n5170 = ~(n12317 ^ n1186);
assign n15857 = ~(n602 ^ n4858);
assign n2008 = n18335 | n16911;
assign n16025 = ~(n3925 ^ n12121);
assign n14609 = ~(n1552 ^ n27006);
assign n9336 = n27063 | n10203;
assign n14635 = ~(n21480 ^ n14225);
assign n24777 = n3329 | n23358;
assign n917 = ~(n15038 ^ n2217);
assign n20495 = ~(n4916 ^ n18346);
assign n19544 = n5147 & n20350;
assign n18790 = ~(n24218 ^ n4501);
assign n18945 = ~(n16660 ^ n25687);
assign n14940 = ~(n3161 | n11630);
assign n3512 = n1350 | n6637;
assign n14422 = n16477 & n10767;
assign n3975 = ~(n6895 | n20462);
assign n1072 = n21888 | n18044;
assign n4254 = ~(n21846 | n19608);
assign n7425 = n10391 & n10383;
assign n13917 = n19510 & n5175;
assign n4125 = ~n2114;
assign n820 = ~(n13772 ^ n14668);
assign n11527 = n6800 | n22152;
assign n1932 = n14936 | n25324;
assign n9083 = n275 | n12133;
assign n10975 = n10909 | n2541;
assign n208 = n18269 | n10784;
assign n27043 = n14818 & n16631;
assign n982 = ~(n2627 ^ n26489);
assign n5404 = ~(n9897 ^ n19132);
assign n24095 = n23137 & n13320;
assign n10682 = n5512 | n5067;
assign n21973 = ~n4118;
assign n13856 = ~(n139 | n914);
assign n4509 = ~(n25835 ^ n7519);
assign n24316 = n6760 | n21649;
assign n15578 = n18814 | n17090;
assign n12147 = ~(n18365 ^ n12850);
assign n20443 = ~(n24961 ^ n5243);
assign n14889 = n9813 | n953;
assign n10006 = n23343 | n21064;
assign n980 = ~(n14655 ^ n22970);
assign n1291 = ~(n3465 | n2244);
assign n11625 = n12136 | n15531;
assign n20322 = n7311 | n15780;
assign n15115 = n2519 | n8951;
assign n852 = ~(n2778 ^ n21504);
assign n9050 = ~n26107;
assign n19488 = ~(n7213 ^ n9172);
assign n21787 = n10881 | n17324;
assign n16866 = n5400 | n9512;
assign n19530 = n12996 | n13376;
assign n22969 = n20909 | n7397;
assign n6040 = n13080 | n12362;
assign n16227 = ~n8244;
assign n3109 = n11199 & n15757;
assign n8736 = ~n12406;
assign n14874 = ~(n23791 | n20925);
assign n24079 = n17899 | n9169;
assign n2252 = n17299;
assign n375 = n14580 | n14195;
assign n13640 = n20056 | n17692;
assign n6828 = ~n14838;
assign n7952 = ~n10158;
assign n20200 = n12002 & n11918;
assign n9457 = ~n7805;
assign n18168 = ~(n17690 ^ n713);
assign n14573 = ~n15383;
assign n11181 = ~(n8792 ^ n26334);
assign n11575 = n2940 & n2464;
assign n12010 = n1389 | n2677;
assign n23558 = ~(n21667 ^ n26387);
assign n22465 = n4903 & n20858;
assign n21778 = n15444 & n4072;
assign n13503 = ~(n20314 ^ n10046);
assign n576 = n25936 | n16712;
assign n26799 = n23804 | n10997;
assign n2298 = ~(n19597 ^ n21785);
assign n3356 = n1512;
assign n17974 = n150 & n17022;
assign n10452 = ~n16524;
assign n3325 = n11244 | n7587;
assign n8603 = n26580 | n3716;
assign n26346 = n2975 | n20938;
assign n5278 = n22319 | n17134;
assign n18429 = ~(n21026 ^ n23803);
assign n18477 = ~(n15898 ^ n11271);
assign n7749 = n21279 & n4389;
assign n9464 = n25954 | n25241;
assign n9953 = n2928 | n18494;
assign n5238 = ~n4410;
assign n26438 = ~(n15678 ^ n13475);
assign n5289 = n17939 | n24214;
assign n25213 = ~(n26724 ^ n5226);
assign n4737 = n9887 | n10630;
assign n228 = n23083 & n17858;
assign n22377 = ~(n2978 ^ n3425);
assign n12549 = n9078 & n10759;
assign n13678 = n7895 & n26349;
assign n13484 = ~(n24743 ^ n5191);
assign n2567 = n19949 | n15210;
assign n19130 = ~(n493 | n14969);
assign n16511 = n13109 & n24898;
assign n21695 = n23121 | n23395;
assign n20616 = ~(n27183 ^ n2150);
assign n22367 = n699 | n23661;
assign n10546 = n15110 | n16701;
assign n10470 = ~n15258;
assign n9849 = ~(n880 | n19328);
assign n26363 = ~n10795;
assign n7018 = ~(n13376 | n16731);
assign n17049 = n8781 | n21058;
assign n7995 = n10403 | n23956;
assign n22780 = ~(n21506 ^ n19911);
assign n10994 = n22739 & n13970;
assign n22356 = n8793 & n15804;
assign n8553 = ~(n6316 ^ n18647);
assign n6677 = ~(n26660 | n18907);
assign n21851 = n12202 | n12672;
assign n20670 = ~(n23693 ^ n10505);
assign n8738 = ~n19089;
assign n23675 = ~(n5449 | n9647);
assign n1984 = ~n354;
assign n1550 = n27060 & n25543;
assign n20817 = n10841 | n2386;
assign n12256 = ~(n4194 ^ n8795);
assign n13489 = ~(n6625 ^ n9598);
assign n26761 = n25866 | n14836;
assign n16062 = ~(n13259 ^ n12252);
assign n17175 = n20470 | n14052;
assign n24427 = ~(n13303 ^ n3785);
assign n12424 = ~(n27188 ^ n6502);
assign n15100 = n26925 | n9394;
assign n8624 = ~n10984;
assign n17655 = n7802 | n10785;
assign n17703 = ~(n17769 ^ n7638);
assign n18195 = n21312 & n13673;
assign n5539 = ~(n19465 | n2126);
assign n16821 = n6759 | n10755;
assign n13766 = ~n7272;
assign n2304 = n361 | n13867;
assign n10457 = ~n23375;
assign n25820 = n24638 | n19327;
assign n3574 = n7849 | n6123;
assign n22844 = n22442 | n22253;
assign n23987 = ~(n18585 ^ n25713);
assign n21311 = n16542 | n24655;
assign n6786 = ~(n20415 | n255);
assign n8456 = ~n23587;
assign n10286 = n3514 | n20867;
assign n5321 = n11737 & n14274;
assign n22236 = n20289 | n6184;
assign n11163 = n25584 | n18435;
assign n10496 = ~(n19110 | n26753);
assign n3738 = n24018 | n13074;
assign n14371 = n1673 | n14579;
assign n15808 = ~(n3339 ^ n15252);
assign n9087 = n25379 & n11625;
assign n2485 = n644 & n154;
assign n26163 = n16947 | n25899;
assign n7386 = n15992 | n6093;
assign n12654 = ~(n21492 ^ n10605);
assign n6966 = n14600 | n563;
assign n19017 = ~n13625;
assign n13613 = ~(n13569 ^ n17553);
assign n21499 = n2055 | n619;
assign n289 = n26459 | n21195;
assign n13442 = n25820 & n22032;
assign n25201 = ~(n22219 | n12514);
assign n3497 = n15987 & n9139;
assign n19078 = n13797 & n13496;
assign n19426 = n14825 & n10931;
assign n11010 = ~(n370 ^ n2228);
assign n17847 = ~n259;
assign n22985 = n15072 | n8748;
assign n3424 = ~(n3356 | n19758);
assign n10228 = ~(n2346 ^ n14768);
assign n19322 = ~(n11366 ^ n11669);
assign n25309 = ~(n16339 | n5569);
assign n20106 = n19042 & n18846;
assign n12450 = n20903 & n624;
assign n19125 = ~(n2452 ^ n16484);
assign n20811 = ~n24200;
assign n523 = n18383 | n5255;
assign n14964 = ~(n26252 | n7750);
assign n22897 = ~(n2977 ^ n325);
assign n22255 = ~(n26499 ^ n22083);
assign n18407 = n22298 | n19751;
assign n7538 = ~(n10811 ^ n8965);
assign n19045 = ~(n21542 ^ n1378);
assign n8286 = ~(n3587 ^ n22278);
assign n9184 = n18131 & n13724;
assign n23255 = n16906 | n16138;
assign n17143 = ~n2389;
assign n20671 = ~(n24197 ^ n10094);
assign n23435 = ~(n589 ^ n23293);
assign n21652 = ~n14261;
assign n16918 = n1282 & n9167;
assign n3476 = n8359 & n27040;
assign n2193 = n21865 | n12628;
assign n11162 = ~n17756;
assign n22997 = n6779 | n14463;
assign n25850 = ~(n18926 ^ n6513);
assign n425 = n3174 | n3006;
assign n16721 = n14293 & n26886;
assign n12222 = n3405 & n24165;
assign n26981 = n25542 & n26214;
assign n15106 = n5619 | n22541;
assign n21812 = n17579 | n4859;
assign n12849 = n4436 & n21406;
assign n12272 = ~(n14504 ^ n8964);
assign n9317 = ~(n9394 ^ n26925);
assign n11249 = ~n23717;
assign n5436 = ~n580;
assign n4784 = n5349 | n3990;
assign n23988 = n25832 & n2188;
assign n24597 = n16975 | n24470;
assign n1581 = ~(n19023 | n18375);
assign n14367 = n7678 | n11579;
assign n2189 = ~(n2882 ^ n17190);
assign n3104 = n12115 | n23256;
assign n8185 = ~(n19974 | n22440);
assign n15096 = n10554 & n330;
assign n24114 = ~(n12258 | n19116);
assign n25597 = n207 | n25030;
assign n11559 = ~n7731;
assign n6348 = n23789 | n25555;
assign n7003 = n10096 & n24511;
assign n4163 = ~(n17572 ^ n6692);
assign n10595 = ~(n18382 ^ n18142);
assign n25994 = ~(n9891 ^ n15872);
assign n23581 = ~n5674;
assign n18514 = ~n17351;
assign n17020 = n24768 | n1019;
assign n1102 = ~(n10710 ^ n26510);
assign n11758 = ~(n15557 ^ n18807);
assign n9609 = ~(n15113 ^ n26832);
assign n9858 = ~(n17004 ^ n15193);
assign n7930 = ~n6596;
assign n8843 = n19361 | n15918;
assign n22891 = ~(n19421 ^ n8217);
assign n26804 = ~(n11158 ^ n11566);
assign n21342 = ~(n6948 | n1911);
assign n20021 = ~(n12956 ^ n26913);
assign n22624 = ~(n5855 ^ n7693);
assign n25893 = ~(n6814 ^ n10763);
assign n20507 = n20563 | n21191;
assign n158 = n14431 | n22587;
assign n20681 = ~(n2768 | n5924);
assign n20436 = ~(n3969 ^ n18998);
assign n26904 = ~n2570;
assign n9886 = n2395 & n11259;
assign n15387 = n10941 | n12901;
assign n13956 = n15933 & n6153;
assign n25971 = ~(n4187 ^ n4225);
assign n8628 = n2939 | n2316;
assign n7136 = n15736 | n19352;
assign n823 = n24170 & n23460;
assign n19995 = n6066 & n7701;
assign n13835 = ~(n21990 ^ n17427);
assign n15604 = ~(n2750 | n25393);
assign n9583 = n12553 & n14872;
assign n14112 = n18170 & n3444;
assign n20270 = n26528 | n25017;
assign n18247 = ~n25057;
assign n18474 = ~n14845;
assign n15425 = n21520 | n24106;
assign n16045 = ~(n26241 | n2999);
assign n8117 = ~(n233 ^ n22583);
assign n13445 = ~(n17674 ^ n17911);
assign n13404 = n22585 | n26837;
assign n6904 = ~n21134;
assign n3005 = n22439 | n26235;
assign n21391 = n19155 | n25458;
assign n14436 = n1637 | n23822;
assign n8312 = n6408 | n14815;
assign n10304 = ~(n17069 ^ n16608);
assign n13673 = n24127 | n9207;
assign n3836 = ~(n7312 ^ n4180);
assign n618 = ~(n13240 ^ n21473);
assign n24306 = n10882 & n8719;
assign n180 = ~n25265;
assign n17564 = n25932 & n14771;
assign n14816 = ~(n16303 ^ n4481);
assign n7337 = ~(n17728 ^ n17959);
assign n7151 = ~(n23708 | n6013);
assign n16277 = ~(n11243 ^ n2421);
assign n25200 = ~(n5875 ^ n13473);
assign n2642 = ~(n5728 ^ n24704);
assign n15877 = ~(n15439 | n7248);
assign n26117 = ~(n8220 ^ n7361);
assign n4235 = n11695 | n2135;
assign n17796 = ~(n19247 ^ n25957);
assign n14373 = n7357 & n24332;
assign n2852 = ~(n13234 ^ n18737);
assign n23312 = ~n11747;
assign n18466 = ~(n1601 ^ n24151);
assign n13583 = n8655 & n11037;
assign n7827 = ~n19263;
assign n24121 = ~(n20018 ^ n10033);
assign n5594 = n2657 | n10482;
assign n4455 = n13361 | n8300;
assign n4380 = ~(n19138 | n24984);
assign n1809 = ~(n18027 ^ n25101);
assign n14021 = ~n17040;
assign n8126 = ~(n22824 ^ n8385);
assign n3152 = n21469 ^ n9713;
assign n2361 = ~(n25774 ^ n4885);
assign n14072 = n9094 | n22655;
assign n14459 = ~(n14514 ^ n24536);
assign n14818 = ~n1136;
assign n11944 = ~n17261;
assign n9778 = ~(n22689 ^ n2650);
assign n24125 = ~n24932;
assign n11662 = ~(n14588 ^ n10288);
assign n1862 = n13343 ^ n11784;
assign n12409 = n24850 | n15271;
assign n12545 = ~(n4210 ^ n10790);
assign n21238 = ~(n16629 ^ n1214);
assign n7543 = ~n6956;
assign n7202 = n898 | n10503;
assign n10247 = n3366 | n4753;
assign n11158 = ~n10973;
assign n6303 = ~n26371;
assign n876 = n26980 | n8387;
assign n1974 = n12247 & n15971;
assign n18597 = n17797 & n10789;
assign n20314 = ~n25089;
assign n22820 = n26119;
assign n6742 = n17251 | n26107;
assign n24158 = ~(n4371 | n11849);
assign n504 = ~(n22900 ^ n13142);
assign n9968 = ~(n1916 ^ n23749);
assign n5074 = ~(n7023 ^ n12126);
assign n11458 = ~(n23932 ^ n20385);
assign n26245 = n13634 & n16997;
assign n11623 = ~(n22608 ^ n2101);
assign n17463 = n23963 & n20807;
assign n7020 = ~n17703;
assign n7468 = ~(n4713 ^ n7805);
assign n9284 = ~(n4721 | n5140);
assign n4224 = ~(n1849 ^ n12034);
assign n21123 = ~(n18932 ^ n14243);
assign n8398 = ~(n18132 ^ n14527);
assign n9595 = ~n25515;
assign n11698 = ~(n4659 ^ n8182);
assign n19315 = ~(n14784 ^ n20058);
assign n15800 = n25710 & n18162;
assign n26649 = ~(n11186 | n7099);
assign n12670 = ~(n9446 ^ n17372);
assign n4428 = n16383 | n21742;
assign n9394 = ~(n23292 ^ n17533);
assign n21572 = n15751 & n20434;
assign n26103 = ~(n26510 ^ n1112);
assign n14516 = ~n8379;
assign n8300 = n25459 & n23282;
assign n8675 = ~n4967;
assign n19867 = n5785 & n16353;
assign n17487 = ~(n26872 ^ n19531);
assign n18928 = ~n7752;
assign n964 = ~(n2162 ^ n7941);
assign n20159 = ~(n12509 | n7761);
assign n9147 = n25540 | n14845;
assign n1347 = n13390 | n8053;
assign n17917 = n13542 & n14688;
assign n19131 = n16557 & n12934;
assign n23022 = n23921 | n5946;
assign n14458 = ~(n211 ^ n195);
assign n23826 = n16061 | n7614;
assign n23336 = n6192 | n20885;
assign n14584 = ~(n26684 ^ n9088);
assign n26815 = ~(n21966 ^ n24269);
assign n24836 = ~(n2829 | n23620);
assign n750 = n23746 | n13161;
assign n17212 = ~(n20074 ^ n20409);
assign n25829 = ~(n14172 | n611);
assign n26599 = ~(n1584 | n17690);
assign n26539 = n24484 | n23995;
assign n11724 = ~(n4535 ^ n17662);
assign n21245 = ~(n25345 | n21322);
assign n21966 = n24477 | n13091;
assign n19806 = ~n11738;
assign n15983 = ~(n12145 | n9814);
assign n13786 = n1541 & n25495;
assign n13395 = n9309 | n3119;
assign n11209 = ~(n10999 ^ n23463);
assign n22726 = n11316 | n10663;
assign n16386 = ~(n1056 ^ n16689);
assign n6029 = ~(n4426 | n13109);
assign n7390 = ~(n25702 ^ n6462);
assign n6973 = n23640 | n1083;
assign n9821 = ~(n18801 ^ n10130);
assign n21983 = n832 | n15424;
assign n21539 = n18963 | n19956;
assign n1405 = ~n6138;
assign n20857 = n14870 & n8888;
assign n4164 = n23666 | n26134;
assign n13000 = ~(n13480 | n11544);
assign n3634 = n3909 & n24200;
assign n23532 = n524 | n18027;
assign n6589 = n1805 & n14674;
assign n26337 = ~(n24839 ^ n22009);
assign n18467 = ~(n1579 ^ n22822);
assign n4066 = n1705 | n5354;
assign n7860 = ~n6710;
assign n13734 = n20787 | n13769;
assign n13476 = ~(n4203 ^ n20207);
assign n19387 = n15695 | n13502;
assign n5468 = n11594 & n1342;
assign n8483 = ~(n16012 | n20127);
assign n5627 = ~(n20043 ^ n16611);
assign n17497 = ~n7086;
assign n9429 = ~(n10712 ^ n23586);
assign n25442 = ~(n27161 ^ n21448);
assign n6046 = ~(n2410 ^ n23370);
assign n9064 = ~(n23144 | n1662);
assign n15301 = n13263 & n8979;
assign n20130 = n15149 | n21955;
assign n10800 = ~(n27089 ^ n8806);
assign n12223 = ~(n25541 ^ n1575);
assign n16790 = n24939 | n18416;
assign n9089 = ~(n5709 ^ n26834);
assign n23285 = ~(n24339 ^ n17176);
assign n681 = n3097 | n3764;
assign n6227 = n11516 | n4513;
assign n12583 = n4858 & n8224;
assign n12225 = ~(n12243 ^ n2642);
assign n19797 = ~n22327;
assign n19501 = ~(n20235 ^ n8259);
assign n24380 = n5391 & n7784;
assign n8132 = ~n20054;
assign n25034 = n15050 | n26700;
assign n13464 = n7814 & n1393;
assign n4360 = ~n16812;
assign n11066 = ~n17408;
assign n2352 = ~(n8351 ^ n25519);
assign n25691 = ~n26394;
assign n13756 = n7517 & n24318;
assign n20962 = n15899 & n18520;
assign n25058 = ~(n11044 | n7619);
assign n4694 = n13525 | n3691;
assign n26315 = n17954 | n23608;
assign n3645 = n5226 | n21205;
assign n9180 = ~n5211;
assign n14621 = ~(n13037 | n8295);
assign n24555 = ~(n2230 | n8869);
assign n5673 = ~(n17194 ^ n17417);
assign n13218 = n10291 | n5192;
assign n11788 = ~(n4410 | n9456);
assign n16301 = ~(n13775 ^ n6397);
assign n16704 = n9801 & n21574;
assign n21046 = ~(n10532 ^ n4782);
assign n2946 = ~(n24281 ^ n8492);
assign n2604 = n8866 & n26570;
assign n8355 = ~(n10501 ^ n5914);
assign n17108 = ~(n18033 ^ n10478);
assign n5694 = ~(n3186 ^ n23224);
assign n20191 = n13708 & n21083;
assign n18377 = ~(n21917 ^ n8585);
assign n22652 = ~n19360;
assign n7544 = ~(n10017 ^ n5026);
assign n24143 = ~n8313;
assign n8092 = ~(n3441 | n8959);
assign n18632 = ~(n25084 ^ n8366);
assign n15288 = n11227 & n16370;
assign n2378 = n4022 & n14565;
assign n5860 = ~(n10383 ^ n25336);
assign n2187 = ~n9054;
assign n15326 = ~(n10405 | n23974);
assign n10269 = n6688 & n1746;
assign n2550 = n20560 | n14462;
assign n2533 = ~(n25986 ^ n16959);
assign n26776 = ~(n182 ^ n17171);
assign n26288 = ~(n8869 ^ n1738);
assign n16065 = ~n8166;
assign n23683 = n2858 | n18727;
assign n4239 = n5935 & n13952;
assign n16825 = ~(n14671 ^ n9707);
assign n15827 = ~(n18805 ^ n8614);
assign n20527 = n5167 & n6458;
assign n13939 = n26200 & n13233;
assign n23163 = ~(n24015 | n4749);
assign n1308 = ~(n5089 ^ n17947);
assign n7768 = ~(n9180 | n18537);
assign n6109 = n14603 | n1141;
assign n19382 = n22476 | n25748;
assign n6099 = ~(n2412 ^ n15884);
assign n23360 = n9598 | n350;
assign n12468 = n19839 & n6518;
assign n4848 = n16189 & n7451;
assign n2508 = n12875 | n7751;
assign n13213 = n19518 | n15677;
assign n9947 = n17635 | n20080;
assign n13329 = ~n26001;
assign n17402 = n26658 | n18991;
assign n10301 = ~n15688;
assign n13544 = n11996 & n7430;
assign n26021 = n20270 & n23379;
assign n8796 = ~(n23369 | n22906);
assign n23800 = ~n7734;
assign n25798 = ~(n24348 | n8332);
assign n13863 = ~n2421;
assign n7643 = n22085 | n15368;
assign n5095 = ~n15775;
assign n7344 = ~(n528 | n1639);
assign n4719 = ~(n5667 ^ n26953);
assign n8975 = n21867 & n22248;
assign n2397 = n20577 & n6519;
assign n16056 = n3809 & n8406;
assign n21097 = ~n23829;
assign n26590 = ~(n358 ^ n19274);
assign n4440 = ~(n312 | n799);
assign n8602 = ~n6808;
assign n2348 = ~(n18649 | n3795);
assign n4207 = n9941 & n9868;
assign n20245 = ~n15289;
assign n26520 = ~(n1367 ^ n8296);
assign n11353 = n16293 | n5600;
assign n7990 = ~(n17599 ^ n9093);
assign n12085 = n6203 | n13333;
assign n5867 = ~(n25524 | n16117);
assign n8665 = ~(n21565 ^ n5103);
assign n17171 = ~(n24253 ^ n398);
assign n21640 = n18349 & n25703;
assign n22107 = ~(n25482 ^ n2901);
assign n6657 = n19332 | n4001;
assign n7557 = n3026 & n8752;
assign n15640 = ~(n11273 | n9026);
assign n14282 = ~(n10269 ^ n14135);
assign n4982 = ~n13573;
assign n10171 = n20842 | n5054;
assign n9298 = n19469 & n25625;
assign n24602 = ~(n10091 ^ n22376);
assign n365 = n24387 | n13507;
assign n25343 = n2296 | n13582;
assign n2097 = n17838 | n8954;
assign n23252 = n11616 & n981;
assign n19336 = n26658 | n1118;
assign n11871 = ~n3414;
assign n16869 = n23068 | n13171;
assign n12793 = n16244 | n19741;
assign n16446 = n11243 | n26497;
assign n6010 = ~(n1009 | n1742);
assign n22455 = n22173 | n583;
assign n25212 = n14974 | n12652;
assign n7851 = n3162 | n24878;
assign n7250 = n11008 | n12743;
assign n19166 = ~(n11479 | n679);
assign n11810 = n11566 | n13150;
assign n13792 = n16347 | n13261;
assign n15236 = ~n25359;
assign n26429 = ~(n8514 ^ n17189);
assign n9434 = n6485 | n26265;
assign n4076 = ~(n8539 | n7627);
assign n13132 = n10623 | n7613;
assign n19256 = n7917 | n3380;
assign n22575 = ~(n19228 ^ n5226);
assign n6533 = ~(n23763 | n13492);
assign n15329 = n14846 & n16297;
assign n24073 = n3635 | n22635;
assign n7645 = n9044 | n21183;
assign n20908 = n10037 & n13148;
assign n26384 = n27035 & n11163;
assign n12472 = ~(n22318 | n3391);
assign n1440 = n24252 | n10081;
assign n23658 = n24187 & n19331;
assign n16772 = n19 | n16476;
assign n25611 = ~(n4832 ^ n2534);
assign n15757 = n5781 | n14112;
assign n7777 = ~(n6115 | n7385);
assign n16802 = n3856 | n20834;
assign n3159 = n12819 | n23186;
assign n22722 = ~n20002;
assign n6877 = ~n866;
assign n233 = n20282 & n20294;
assign n6285 = ~n14447;
assign n1576 = n8568 & n23793;
assign n2122 = ~(n1627 ^ n14773);
assign n5741 = n18979 & n23138;
assign n10177 = ~(n1099 ^ n6381);
assign n16962 = ~(n14362 | n14240);
assign n7904 = n20686 & n20507;
assign n26270 = n26457 & n7063;
assign n3993 = ~n13072;
assign n26077 = ~(n5328 ^ n15780);
assign n14761 = ~(n22234 ^ n2175);
assign n5658 = n10668 | n13212;
assign n9828 = ~(n14704 | n17716);
assign n20497 = ~n5400;
assign n24488 = ~(n9553 ^ n25919);
assign n6014 = n9357 & n23155;
assign n22854 = n9718 | n5425;
assign n1143 = ~(n18314 ^ n12644);
assign n26321 = n7553 | n10879;
assign n22656 = n11030 & n6141;
assign n24211 = ~(n22290 | n13018);
assign n16000 = n5994 & n18348;
assign n21580 = ~(n17231 ^ n16354);
assign n1481 = ~(n4934 ^ n20658);
assign n25937 = ~(n24920 ^ n21639);
assign n10617 = ~(n24589 ^ n3588);
assign n16066 = n8790 & n7633;
assign n6670 = ~n8225;
assign n23365 = ~n16713;
assign n2494 = n17017 | n19418;
assign n1076 = n23804 | n21138;
assign n3250 = n3689 | n20135;
assign n15651 = n6485 & n18676;
assign n15909 = ~(n25941 ^ n17495);
assign n11194 = ~(n13494 ^ n4319);
assign n26854 = n16812 | n14397;
assign n20317 = ~(n18295 ^ n25974);
assign n16272 = n4729 | n10096;
assign n16356 = ~(n13529 ^ n5474);
assign n10186 = n23303 & n15067;
assign n10236 = ~(n22118 ^ n1170);
assign n4489 = ~(n17316 ^ n18734);
assign n22615 = ~n22303;
assign n16553 = n10213 & n14924;
assign n14182 = n6904 & n17419;
assign n14840 = ~(n19616 | n1118);
assign n5711 = n26552 & n3337;
assign n18364 = n23230 | n4665;
assign n8280 = ~(n2595 ^ n26484);
assign n2675 = ~n8988;
assign n26881 = n26659 & n16187;
assign n4130 = ~n7871;
assign n4020 = n10025 & n24456;
assign n14536 = ~n5443;
assign n18198 = n9181 & n8926;
assign n5925 = ~n20961;
assign n21555 = n1260 & n22555;
assign n13499 = ~(n20138 ^ n25073);
assign n15242 = n22792 | n1550;
assign n17036 = n21535 & n19787;
assign n23424 = ~(n111 ^ n5587);
assign n9491 = n16106 | n26964;
assign n20014 = ~(n4303 ^ n4387);
assign n23951 = ~(n1019 ^ n24768);
assign n1625 = n12260 & n25990;
assign n8123 = n11201 | n26340;
assign n25189 = n8060 & n9482;
assign n5631 = ~(n18191 | n18188);
assign n10606 = ~(n16496 | n17350);
assign n2522 = ~n985;
assign n5391 = n18601 | n19874;
assign n26724 = ~n9992;
assign n27012 = ~(n4100 | n24609);
assign n17172 = ~(n5329 ^ n10053);
assign n9148 = n26868 & n22205;
assign n16035 = n2746 | n4609;
assign n4798 = ~n22091;
assign n23087 = n16673 & n1408;
assign n3198 = n11736 | n18183;
assign n2357 = n19849 | n26585;
assign n9538 = ~n10468;
assign n21233 = ~(n24403 ^ n23175);
assign n14475 = ~(n5282 ^ n17837);
assign n6419 = n2866 & n19645;
assign n10608 = ~n15359;
assign n16041 = ~(n9570 | n6785);
assign n14829 = ~n15214;
assign n18375 = ~(n6631 | n7339);
assign n8858 = ~(n5135 ^ n7792);
assign n23199 = ~(n8371 ^ n6464);
assign n18681 = n4868 | n23820;
assign n11802 = ~n16910;
assign n14795 = ~n2041;
assign n26115 = n1029 | n19281;
assign n15026 = ~n4293;
assign n14334 = n2502 | n366;
assign n20432 = n18525 & n876;
assign n18225 = ~(n22755 ^ n310);
assign n3215 = n6027 | n7239;
assign n21383 = n14515 | n10735;
assign n10871 = n13163 | n6497;
assign n18339 = ~(n7671 ^ n4959);
assign n17322 = ~(n3837 ^ n7325);
assign n21016 = n8248 & n22917;
assign n19246 = n2207 | n22142;
assign n10212 = ~(n23460 ^ n24170);
assign n16369 = ~(n1742 ^ n19196);
assign n26130 = n5657 | n733;
assign n10819 = n2721 | n14826;
assign n1399 = n16607 | n1244;
assign n11542 = ~n2409;
assign n19289 = n22545 | n7875;
assign n16525 = n5426 | n8028;
assign n21243 = n5750 | n2249;
assign n11515 = ~(n19480 ^ n14787);
assign n5227 = ~n20432;
assign n2598 = ~(n13339 ^ n12562);
assign n23738 = n19653 & n18132;
assign n14313 = n11781 & n24396;
assign n26887 = ~(n10788 | n16900);
assign n26146 = ~(n3946 | n18318);
assign n7694 = n14722 | n13442;
assign n6864 = ~n15969;
assign n11993 = ~(n22591 ^ n26167);
assign n1480 = ~(n23064 ^ n3582);
assign n5375 = n874 | n12267;
assign n5574 = ~n2510;
assign n258 = ~n8799;
assign n10642 = n24823 | n13893;
assign n7041 = ~n9133;
assign n921 = ~(n15509 ^ n14304);
assign n6054 = ~(n4195 | n21671);
assign n25437 = n23162 | n5868;
assign n6297 = ~(n7096 ^ n7876);
assign n22535 = ~n6360;
assign n14423 = ~(n21071 ^ n7906);
assign n23747 = ~(n10117 ^ n3306);
assign n21429 = n15796 | n10739;
assign n16872 = n25237 & n21710;
assign n12465 = ~n16126;
assign n11547 = n2949 | n43;
assign n12227 = n15240 | n27185;
assign n26830 = ~n20687;
assign n3373 = n22176 | n21662;
assign n12991 = ~n7466;
assign n1915 = ~(n4261 ^ n117);
assign n27075 = ~n303;
assign n12502 = ~(n26541 ^ n4967);
assign n14674 = n6815 | n19505;
assign n12246 = ~(n27204 ^ n18545);
assign n1036 = ~n18438;
assign n3060 = n4654 | n25874;
assign n13502 = n9052 & n11082;
assign n15915 = n20513 | n12605;
assign n21581 = n3460 | n16667;
assign n20500 = ~(n3164 ^ n2547);
assign n22267 = ~(n17380 ^ n20927);
assign n70 = n18190 | n3084;
assign n19484 = n25738 | n11265;
assign n25009 = ~(n11503 ^ n12593);
assign n2600 = n14441 | n20240;
assign n11293 = n9942 | n13946;
assign n19409 = ~(n20284 ^ n3779);
assign n5823 = n20378 & n4677;
assign n25558 = ~n20923;
assign n11077 = n13376 & n4643;
assign n12605 = ~(n21474 ^ n11354);
assign n13430 = n18506 | n4812;
assign n8729 = ~(n6240 ^ n19497);
assign n23982 = ~(n1036 ^ n20728);
assign n2572 = n23043 | n26622;
assign n24494 = n22308 | n14407;
assign n16307 = n26460 | n19649;
assign n3064 = n19902 | n12535;
assign n16660 = ~n18063;
assign n11396 = n18352 | n2129;
assign n18039 = ~(n3018 ^ n2731);
assign n11680 = ~(n22077 | n21838);
assign n18852 = n3120 & n14361;
assign n26497 = ~n1434;
assign n22474 = ~(n2291 ^ n24791);
assign n19829 = n25643 | n20604;
assign n23980 = ~(n1755 ^ n24993);
assign n2523 = n741 & n7594;
assign n10531 = n20425 & n15498;
assign n17805 = ~(n2281 ^ n1047);
assign n6398 = ~(n840 | n11186);
assign n9535 = ~(n10223 ^ n17078);
assign n10010 = ~(n18588 ^ n3845);
assign n13652 = ~(n15696 ^ n13709);
assign n2069 = n9678 | n1484;
assign n14787 = ~(n23612 ^ n14488);
assign n23561 = n20554 | n19058;
assign n6307 = ~(n21993 ^ n14575);
assign n18975 = ~(n16838 ^ n20267);
assign n22986 = ~(n16561 ^ n23596);
assign n18066 = n20747 | n18540;
assign n21079 = n2403 | n25125;
assign n11554 = n8626;
assign n4659 = ~n3955;
assign n18094 = ~(n19005 ^ n7149);
assign n20257 = n11550 | n1626;
assign n14320 = ~(n2980 ^ n4781);
assign n19105 = n20880 | n376;
assign n23231 = ~n3668;
assign n7729 = ~(n27015 ^ n22993);
assign n8798 = ~(n5527 ^ n25218);
assign n1307 = ~(n6865 | n3727);
assign n22473 = ~(n8418 ^ n6356);
assign n21491 = n25480 | n16904;
assign n12134 = ~(n19340 | n234);
assign n19082 = ~n6775;
assign n25356 = ~(n25011 ^ n2943);
assign n22122 = ~(n4580 ^ n5057);
assign n1172 = ~(n26892 ^ n26047);
assign n17051 = ~(n2160 ^ n7335);
assign n9217 = ~(n12694 ^ n22450);
assign n26891 = ~(n11840 | n23059);
assign n17675 = n23800 | n1308;
assign n13551 = ~(n7552 ^ n26609);
assign n22808 = ~(n14041 ^ n10359);
assign n14424 = n20826 | n17326;
assign n10175 = n12454 | n16755;
assign n15260 = ~(n21540 | n13485);
assign n9470 = n21083 | n13708;
assign n10756 = ~(n5995 ^ n22627);
assign n3333 = ~n21727;
assign n8311 = n16937 | n14002;
assign n10931 = n14517 | n2839;
assign n24002 = ~(n8839 ^ n25852);
assign n1202 = ~(n8305 | n2918);
assign n15710 = n9196 | n6775;
assign n8757 = ~(n2017 | n650);
assign n14032 = ~(n8645 ^ n15635);
assign n4565 = n9401 | n22121;
assign n945 = ~n19569;
assign n23281 = ~n2696;
assign n20190 = ~(n2816 ^ n1222);
assign n12511 = ~n1742;
assign n15880 = ~(n8422 | n25627);
assign n6061 = ~(n18261 | n12398);
assign n555 = n12244 & n14673;
assign n5301 = n8421 & n4305;
assign n24069 = n989 | n22847;
assign n15013 = n22804 | n21309;
assign n18923 = n17446 | n11606;
assign n2584 = n16298 | n3819;
assign n4402 = n4704 | n14365;
assign n10630 = n4976 & n15694;
assign n19664 = ~(n2741 ^ n5581);
assign n18020 = ~(n21850 ^ n25751);
assign n17120 = ~n22332;
assign n26369 = n19574 & n13185;
assign n6298 = ~(n21070 ^ n17317);
assign n10896 = n8978 & n27123;
assign n2512 = ~(n20794 | n25471);
assign n12278 = ~(n4181 ^ n13879);
assign n2311 = n2668 | n12807;
assign n22440 = ~n23435;
assign n24582 = ~(n14692 | n14437);
assign n20860 = n19594 | n12749;
assign n11653 = ~(n25746 ^ n8973);
assign n22786 = n20 | n16907;
assign n17456 = ~(n18741 | n22782);
assign n18899 = ~(n5972 ^ n1823);
assign n2875 = ~n27126;
assign n526 = n16916 & n3624;
assign n15976 = n24806 | n5342;
assign n21105 = n7973 | n15179;
assign n24060 = n4132 | n13074;
assign n8173 = n4875 & n4209;
assign n26374 = ~(n16309 | n23873);
assign n6887 = ~n24984;
assign n26127 = n20945 & n22953;
assign n14538 = ~(n13207 ^ n24427);
assign n17837 = ~(n5669 ^ n21575);
assign n18191 = ~n1570;
assign n20404 = ~n25322;
assign n13236 = n24631 | n352;
assign n23771 = ~(n16249 | n14557);
assign n8155 = ~n22379;
assign n26445 = ~(n19144 | n5496);
assign n6087 = n303 | n25101;
assign n17922 = ~(n4749 ^ n24015);
assign n5964 = ~(n13236 ^ n3355);
assign n15689 = n25649 | n19581;
assign n22681 = n7222 & n19601;
assign n22699 = n22723 & n5692;
assign n15896 = n2334 | n12598;
assign n22811 = n20404 | n14661;
assign n21612 = n23753 | n3240;
assign n624 = n18465 | n3580;
assign n15292 = ~(n21599 | n9576);
assign n16454 = ~(n4844 | n8052);
assign n21821 = n26539 & n8476;
assign n17897 = n19815 & n2581;
assign n19155 = n8910 & n25018;
assign n23933 = n1291 | n4829;
assign n18044 = n12409 & n17934;
assign n3269 = n21871 | n6659;
assign n14132 = n1654 & n7893;
assign n10914 = ~(n12774 ^ n12121);
assign n2994 = ~n5568;
assign n12805 = n23082 & n9613;
assign n20883 = ~n12137;
assign n25825 = n17919 & n26773;
assign n18425 = ~(n13813 ^ n17496);
assign n6553 = ~(n962 ^ n9318);
assign n12292 = n10426 & n12635;
assign n14618 = n5407 | n20604;
assign n12217 = ~n1674;
assign n1337 = n18406 & n9959;
assign n22020 = ~(n20854 ^ n20352);
assign n18548 = n16252 & n17943;
assign n15914 = ~(n15798 ^ n20832);
assign n13256 = n18847 | n12110;
assign n5182 = ~(n11006 ^ n16212);
assign n21051 = n144 | n11919;
assign n6351 = ~n19858;
assign n12798 = n12268 & n5573;
assign n13784 = ~(n5988 ^ n13677);
assign n21041 = n6405 & n3765;
assign n23296 = n9671 & n5205;
assign n3950 = n26079 | n7863;
assign n24913 = ~(n21194 ^ n27008);
assign n27179 = ~(n7692 ^ n25464);
assign n6226 = ~n19678;
assign n24761 = n10514 | n10041;
assign n18414 = ~(n19536 ^ n1764);
assign n23069 = ~(n3239 | n1464);
assign n78 = ~(n18035 ^ n5834);
assign n25785 = n4411 & n14197;
assign n18518 = ~(n570 | n2479);
assign n12078 = ~(n21612 ^ n23825);
assign n2577 = n21749 | n2298;
assign n18223 = ~n13218;
assign n18615 = ~n19262;
assign n21368 = ~(n9076 ^ n704);
assign n13138 = n14684 | n1667;
assign n18519 = ~(n7920 ^ n20976);
assign n14171 = n16713 & n17497;
assign n13890 = n10514 & n10041;
assign n5482 = ~(n10135 ^ n2809);
assign n362 = ~(n20655 ^ n19951);
assign n25092 = n14520 & n21712;
assign n25098 = n27033 | n4207;
assign n13899 = ~n26208;
assign n5154 = ~(n15282 | n9859);
assign n25385 = ~(n5475 ^ n7324);
assign n6171 = ~(n14371 ^ n17997);
assign n1720 = ~n2747;
assign n20376 = ~n2719;
assign n7158 = n20994 & n12669;
assign n20421 = ~(n23993 ^ n19731);
assign n2976 = ~(n19286 ^ n10245);
assign n14607 = ~(n1522 ^ n1599);
assign n22159 = ~(n14974 ^ n12663);
assign n6338 = n21456 | n22537;
assign n17575 = n14224 & n11097;
assign n15524 = n173 | n16167;
assign n4846 = ~n5862;
assign n27124 = n14367 & n11142;
assign n15164 = ~n13558;
assign n18276 = n14337 | n24865;
assign n4707 = n13899 | n8233;
assign n16713 = ~(n21039 ^ n14694);
assign n18229 = ~(n24732 ^ n12892);
assign n9461 = ~(n1519 ^ n5263);
assign n8662 = ~(n13524 ^ n9225);
assign n19649 = ~(n12676 ^ n18791);
assign n23237 = ~(n9671 | n10712);
assign n14629 = n16747 | n15520;
assign n17312 = ~(n26564 ^ n22744);
assign n16508 = n14040 | n8477;
assign n1535 = n1989 & n18369;
assign n7539 = n17330 & n24140;
assign n24556 = n18447 & n24350;
assign n26932 = n341 & n21569;
assign n13477 = ~(n22737 ^ n17220);
assign n11083 = n10819 & n1813;
assign n6579 = n19448 & n21966;
assign n10049 = ~n25068;
assign n4174 = ~n7082;
assign n15476 = n18134 | n16539;
assign n5088 = n23877 | n20354;
assign n18586 = ~(n23800 ^ n5163);
assign n7701 = n6391 | n24800;
assign n11798 = n6456 & n17978;
assign n19614 = ~n18820;
assign n20951 = ~n13940;
assign n10060 = n26767 | n21470;
assign n4179 = n8509 | n17087;
assign n12346 = ~(n20003 ^ n15343);
assign n26555 = n19770 | n11451;
assign n8585 = ~(n7071 ^ n14848);
assign n6312 = n11011 | n1019;
assign n23139 = ~(n7143 ^ n10728);
assign n13983 = ~(n22083 | n26215);
assign n18367 = n22868 | n1153;
assign n11137 = ~n20485;
assign n1537 = ~(n18295 | n16223);
assign n11889 = ~n2337;
assign n760 = n5682 | n3862;
assign n11804 = n10792 & n17230;
assign n19066 = ~(n17203 | n17597);
assign n1303 = n3334 | n9998;
assign n19969 = n22518 | n14824;
assign n23238 = ~(n10459 ^ n12313);
assign n26619 = n16144 | n18107;
assign n17521 = n9829 | n22181;
assign n14006 = n25855 | n26461;
assign n11634 = n17037 | n21385;
assign n20596 = ~(n7656 | n669);
assign n14885 = ~(n1529 ^ n14786);
assign n16891 = n14001 | n20543;
assign n11595 = ~(n15586 | n17495);
assign n22331 = n14699 | n21300;
assign n747 = ~(n16687 | n5319);
assign n26046 = ~(n8607 ^ n25523);
assign n21841 = ~n23864;
assign n11023 = ~(n3787 ^ n22818);
assign n24415 = ~(n8021 ^ n10591);
assign n7288 = n17091 | n9711;
assign n21207 = ~n6691;
assign n6908 = ~(n5035 ^ n18531);
assign n25328 = ~(n20395 ^ n21746);
assign n336 = ~(n13424 ^ n23831);
assign n2215 = n15806 | n20300;
assign n19816 = n12301 | n560;
assign n3727 = ~n6703;
assign n3513 = ~(n1028 ^ n1618);
assign n3808 = n7192 & n11956;
assign n2956 = n14540 & n16023;
assign n10106 = ~n7883;
assign n19285 = n16796 & n10256;
assign n4336 = n9740 | n17850;
assign n15363 = n13967 | n20964;
assign n13747 = ~(n23508 ^ n22945);
assign n12266 = ~(n19926 ^ n1243);
assign n8981 = n13783 & n6341;
assign n12130 = ~(n2914 | n16376);
assign n19064 = ~(n1128 ^ n19948);
assign n14022 = n25817 & n23052;
assign n15178 = n22634 & n17816;
assign n14805 = ~(n650 ^ n9872);
assign n22815 = ~(n4461 ^ n17954);
assign n3568 = ~(n26234 ^ n18697);
assign n15560 = ~n20826;
assign n19818 = ~(n15415 | n25523);
assign n25639 = ~n4602;
assign n4064 = ~(n20751 ^ n16466);
assign n24698 = n15279 & n23817;
assign n24812 = ~(n14218 ^ n7737);
assign n10982 = ~(n26197 | n4555);
assign n7192 = n8689 | n21508;
assign n14876 = n8562 | n8941;
assign n3844 = ~(n150 ^ n24315);
assign n13408 = ~(n25604 | n26499);
assign n22468 = ~(n2017 | n11649);
assign n354 = ~(n4502 ^ n24901);
assign n103 = n10593 | n5817;
assign n7718 = n2883 | n4018;
assign n25422 = n25640 & n5702;
assign n21803 = n25049 | n20731;
assign n8533 = ~(n26373 ^ n25418);
assign n15803 = ~(n2566 ^ n4894);
assign n12570 = ~(n11006 ^ n10113);
assign n18622 = n15825 & n14370;
assign n9822 = ~(n8088 ^ n8624);
assign n14526 = n7074 | n19000;
assign n13909 = ~(n27037 | n23913);
assign n2011 = n2023 | n15675;
assign n11896 = ~(n20102 | n14269);
assign n12204 = ~(n14209 ^ n6162);
assign n10009 = ~(n12231 ^ n724);
assign n23141 = ~n26054;
assign n8815 = n12613 | n22680;
assign n2996 = ~n25980;
assign n14958 = ~n8272;
assign n557 = ~(n24863 ^ n5252);
assign n1771 = ~(n19227 | n24298);
assign n26530 = ~(n1761 ^ n2817);
assign n15632 = n8629 | n21352;
assign n7449 = n20315 | n11869;
assign n18359 = n6844 & n15040;
assign n24345 = ~(n11809 ^ n16957);
assign n26302 = ~n4786;
assign n9337 = n1333 & n19051;
assign n5104 = n1587 | n14008;
assign n20872 = ~(n8570 ^ n6996);
assign n2042 = ~(n10092 ^ n23644);
assign n21771 = ~n25031;
assign n13829 = n7367 & n15993;
assign n26342 = n12258 | n152;
assign n2541 = n18041 & n21012;
assign n22708 = n1896 | n25886;
assign n724 = ~(n1833 | n9834);
assign n18015 = n23771 | n907;
assign n25955 = n2239 | n23415;
assign n2442 = n17351 | n26528;
assign n21636 = ~(n21172 ^ n6369);
assign n4392 = n13384 | n16106;
assign n1330 = n25693 | n7131;
assign n16150 = n22243 | n2143;
assign n5231 = ~(n9724 ^ n17689);
assign n413 = n24382 | n24262;
assign n18752 = n3645 & n3747;
assign n24437 = ~(n22962 | n12209);
assign n14561 = ~(n27037 ^ n11736);
assign n18807 = ~(n1293 ^ n19196);
assign n589 = n17577 & n20341;
assign n24542 = ~(n18608 ^ n19899);
assign n20292 = ~(n21288 | n25238);
assign n11165 = ~n10034;
assign n12732 = n17970 | n3700;
assign n15009 = ~(n17453 ^ n26783);
assign n15626 = ~n19484;
assign n5370 = n4133 | n2335;
assign n16500 = ~(n7317 ^ n21471);
assign n26327 = ~n12939;
assign n16605 = n12021 | n7333;
assign n9914 = ~(n6255 ^ n21984);
assign n21031 = n8136 & n14371;
assign n18406 = n21853 | n17410;
assign n12727 = ~(n14616 ^ n10573);
assign n7122 = ~(n6915 ^ n18158);
assign n1158 = n26907 | n26152;
assign n6265 = ~(n4997 ^ n9864);
assign n25165 = n16650 & n4323;
assign n4892 = ~(n18798 | n9332);
assign n8221 = n276 & n15386;
assign n19069 = n3286 & n785;
assign n18448 = n3607 | n16463;
assign n21661 = ~(n13489 ^ n4913);
assign n21202 = n9064 | n23446;
assign n17269 = ~(n11210 ^ n14637);
assign n3135 = ~(n14545 | n18070);
assign n13345 = n3495 | n9525;
assign n21587 = ~n17016;
assign n16328 = n19178 & n21147;
assign n9555 = n22944 | n19249;
assign n7652 = ~(n7116 ^ n22569);
assign n26132 = ~(n23528 | n10852);
assign n3914 = ~(n15752 ^ n10506);
assign n24250 = n11116 | n2608;
assign n12818 = n2744 & n7626;
assign n5997 = ~(n26951 ^ n27054);
assign n7831 = ~(n16633 | n4622);
assign n6879 = ~(n3694 ^ n5302);
assign n12429 = n1727 | n8595;
assign n2358 = n16830 | n26741;
assign n9692 = ~(n19134 | n18158);
assign n7373 = ~(n18542 ^ n25074);
assign n18563 = ~(n4136 ^ n4826);
assign n4824 = n10762 & n26050;
assign n2629 = n11980 & n19446;
assign n23010 = n19494 & n1458;
assign n22797 = ~n4005;
assign n11848 = ~n17291;
assign n22510 = ~n7072;
assign n10806 = n85 | n10475;
assign n14474 = n8327 & n13432;
assign n15070 = n9076 | n25368;
assign n20108 = n12017 & n15807;
assign n13769 = n7926 & n27152;
assign n7764 = ~(n10622 ^ n12064);
assign n12106 = n1021 | n11009;
assign n4662 = n6356 | n4067;
assign n13148 = n20544 & n12071;
assign n4644 = n25175 & n18023;
assign n15997 = ~(n18676 ^ n24731);
assign n16004 = n21873 | n22690;
assign n25711 = n22564 & n18671;
assign n9225 = ~(n17010 ^ n19460);
assign n2593 = n15648 & n18160;
assign n2345 = ~(n6185 ^ n10125);
assign n4492 = ~n23950;
assign n8828 = n13388 | n19318;
assign n24030 = ~(n23321 ^ n20429);
assign n10288 = ~(n15258 ^ n2420);
assign n10093 = ~(n1190 ^ n17852);
assign n10667 = n6058 | n21056;
assign n21732 = ~(n19872 ^ n21462);
assign n3455 = ~(n12341 | n22515);
assign n8321 = ~(n23654 ^ n19225);
assign n12960 = ~(n14432 ^ n10283);
assign n10303 = ~(n16247 ^ n23541);
assign n14025 = ~(n10335 | n10141);
assign n5958 = n1205 & n7494;
assign n3608 = ~n757;
assign n1557 = ~(n25639 | n21337);
assign n24346 = n14624 | n5448;
assign n24109 = ~(n11270 ^ n10732);
assign n5179 = n217 & n22165;
assign n22778 = ~(n5855 ^ n14576);
assign n22961 = ~(n14532 | n17635);
assign n9643 = n19679 & n26379;
assign n21870 = n26238 | n10753;
assign n20844 = n17734 | n10639;
assign n4343 = n6619 & n12176;
assign n14589 = ~(n8176 ^ n8827);
assign n3833 = ~(n6640 ^ n25565);
assign n9418 = ~(n18415 ^ n2536);
assign n17510 = ~(n25276 | n6137);
assign n14430 = n19899 & n18608;
assign n17961 = n8410 | n22826;
assign n14010 = ~(n6206 ^ n17409);
assign n2114 = n11223 | n7710;
assign n10812 = n7649 & n5864;
assign n19457 = ~(n26214 ^ n26103);
assign n12229 = ~n7445;
assign n21676 = ~(n3030 | n7407);
assign n10768 = ~(n19177 | n26768);
assign n17103 = ~(n3483 | n19556);
assign n16116 = n9186 & n2716;
assign n19207 = n5816 | n15780;
assign n22402 = ~(n11195 | n20274);
assign n18897 = n17054 | n24063;
assign n11444 = n7748 & n26203;
assign n7218 = n15448 & n24034;
assign n19273 = n970 | n12292;
assign n5488 = n5440 & n24366;
assign n5239 = n5455 | n1530;
assign n20430 = n6786 | n11872;
assign n22739 = n3785 | n21;
assign n22339 = ~(n23354 ^ n2950);
assign n1064 = n18746 | n17483;
assign n3154 = n24049 | n16025;
assign n9189 = n17063 | n5843;
assign n15162 = n2416 & n16455;
assign n6432 = n468 & n22322;
assign n1972 = ~(n5520 ^ n24977);
assign n16125 = ~(n26135 ^ n504);
assign n26947 = ~n14048;
assign n23820 = ~(n11468 ^ n26604);
assign n2473 = n11016 & n25036;
assign n17496 = ~(n7669 ^ n6218);
assign n7464 = ~(n20512 ^ n3260);
assign n2266 = ~(n12465 ^ n19575);
assign n12662 = n25876 | n24541;
assign n726 = ~n22082;
assign n25051 = n20101 & n8705;
assign n8294 = n21222 | n277;
assign n18087 = n3033 | n22701;
assign n26079 = n8106 & n10904;
assign n26202 = ~n14467;
assign n14859 = n11938 | n7162;
assign n24240 = n14979 | n4957;
assign n18241 = ~(n9654 ^ n20523);
assign n5985 = n13787 & n20545;
assign n9700 = ~(n3691 ^ n10272);
assign n7182 = n15408 | n19111;
assign n16019 = ~n2792;
assign n19902 = ~n21749;
assign n21817 = n3367 & n16063;
assign n10091 = n19811 | n534;
assign n22263 = n14874 | n22661;
assign n19881 = n16576 | n10437;
assign n10218 = n3403 | n24778;
assign n6030 = ~n10772;
assign n18202 = ~n22934;
assign n3528 = ~(n10226 ^ n9547);
assign n7292 = ~n16988;
assign n22775 = ~(n18157 | n26030);
assign n12254 = n21270 | n19823;
assign n8391 = ~(n2040 ^ n23039);
assign n4127 = ~n19377;
assign n4339 = ~(n9108 | n8873);
assign n21548 = n3438 | n25848;
assign n14428 = n21524 & n18532;
assign n22112 = n2508 & n17127;
assign n6616 = n11525 | n19569;
assign n11899 = ~(n1176 | n7254);
assign n18237 = n4537 | n6446;
assign n12580 = n9895 & n760;
assign n25532 = ~(n5250 ^ n18036);
assign n6336 = n16995 | n25229;
assign n22333 = ~n20512;
assign n5208 = n8645 | n13365;
assign n23421 = n14508 | n13778;
assign n14241 = n19094 & n1197;
assign n10483 = ~(n17784 ^ n24085);
assign n24926 = ~(n21687 ^ n19922);
assign n5258 = ~(n9990 | n7134);
assign n17650 = n21245 | n12163;
assign n26845 = n18814 & n802;
assign n11346 = n26307 & n23799;
assign n18052 = n25498 & n8132;
assign n3282 = ~(n14195 ^ n14580);
assign n17469 = n2811 | n4239;
assign n7635 = ~(n16743 ^ n24485);
assign n561 = ~(n4940 | n7609);
assign n2829 = ~(n12608 ^ n25323);
assign n14982 = ~n12716;
assign n13007 = n9944 | n20986;
assign n12337 = ~(n23076 | n3509);
assign n9577 = n4806 & n11883;
assign n16243 = ~(n22141 ^ n10858);
assign n8289 = n23467 & n10772;
assign n16281 = n11570 & n21103;
assign n25088 = n19935 & n8195;
assign n16496 = ~(n10695 ^ n4794);
assign n1697 = ~(n16546 ^ n24283);
assign n4802 = n22254 | n6733;
assign n21856 = ~(n12593 ^ n13714);
assign n17515 = n23769 & n13747;
assign n9076 = ~n19499;
assign n4484 = ~(n7125 ^ n24418);
assign n13699 = n24279 & n6106;
assign n26335 = n5253 & n20146;
assign n4425 = n286 ^ n7234;
assign n5420 = n23837 & n4384;
assign n3571 = n5783 | n2043;
assign n16705 = ~(n7414 ^ n18496);
assign n4664 = ~n21638;
assign n23189 = ~(n18035 | n12477);
assign n19019 = n8454 | n1061;
assign n7030 = ~(n8616 ^ n3875);
assign n106 = ~n16083;
assign n14985 = ~(n19658 ^ n15767);
assign n5527 = ~(n23770 ^ n16082);
assign n1 = ~n3584;
assign n4480 = n24395 & n1303;
assign n27078 = n5596 ^ n9427;
assign n14164 = ~(n25624 ^ n9653);
assign n2735 = n16627 | n16393;
assign n24930 = n12378 & n1072;
assign n22743 = ~n26625;
assign n19679 = n5006 | n23529;
assign n4047 = n17403 | n13288;
assign n10163 = n7175 | n22621;
assign n12978 = ~(n656 ^ n1007);
assign n4496 = n24305 | n20231;
assign n6625 = n15114 & n25699;
assign n6232 = ~(n25182 ^ n25211);
assign n19887 = n25120 & n2903;
assign n16832 = n21287 | n19981;
assign n17190 = ~(n12900 ^ n1255);
assign n20352 = ~(n26876 ^ n21997);
assign n2190 = n20100 | n18720;
assign n806 = n23054 | n22630;
assign n8847 = ~(n14290 ^ n19562);
assign n23414 = ~(n25689 ^ n6852);
assign n636 = ~n6060;
assign n7490 = n26854 & n19206;
assign n20498 = n24417 & n10027;
assign n23020 = n16139 & n2225;
assign n22187 = n7296 | n3562;
assign n9036 = n15089 & n16740;
assign n15537 = ~(n5682 ^ n3554);
assign n8953 = n11249 | n25296;
assign n24907 = ~(n21139 ^ n2039);
assign n15818 = ~n367;
assign n14478 = ~(n14016 | n14102);
assign n23494 = n6281 | n8661;
assign n13717 = ~(n24314 | n9236);
assign n7206 = n12422 | n12999;
assign n9765 = ~n22986;
assign n18949 = n23124 | n2136;
assign n20058 = ~(n6734 ^ n3);
assign n3191 = n6959 | n19819;
assign n18461 = n5006 & n7156;
assign n4879 = n19027 | n12647;
assign n24679 = ~(n16968 ^ n21654);
assign n23221 = n16917 | n938;
assign n7784 = n3308 | n18623;
assign n22399 = ~(n12213 ^ n132);
assign n17200 = ~(n41 ^ n21718);
assign n25415 = ~(n17892 ^ n9915);
assign n11389 = n6603 | n21263;
assign n2129 = ~(n13040 | n23204);
assign n22306 = ~(n12301 | n26467);
assign n12903 = n11669 | n9561;
assign n15366 = ~(n14357 ^ n9714);
assign n11216 = n19833 & n18178;
assign n11814 = ~n10955;
assign n22713 = n3606 & n24643;
assign n13541 = n8074 & n22239;
assign n21624 = n11092 | n6642;
assign n24855 = ~n20646;
assign n20954 = ~n6603;
assign n5555 = ~(n22876 ^ n18312);
assign n7403 = ~(n25315 ^ n21323);
assign n14686 = n8270 | n5610;
assign n18657 = ~(n26667 ^ n3097);
assign n2636 = ~n17169;
assign n4748 = ~(n7311 ^ n9399);
assign n20115 = n25382 | n518;
assign n2376 = n16366 & n18203;
assign n19943 = n4236 | n6622;
assign n3098 = n22968 | n17186;
assign n4186 = ~(n2127 ^ n2285);
assign n17516 = n27059 & n23368;
assign n19097 = ~(n406 ^ n15297);
assign n12097 = n10546 & n6052;
assign n2216 = n8818 | n5171;
assign n8212 = n14198 & n12902;
assign n14193 = ~(n19177 | n23175);
assign n23486 = ~(n20817 ^ n27195);
assign n15655 = ~(n3460 | n24774);
assign n24059 = n22034 & n2110;
assign n18248 = n25478 & n22143;
assign n26617 = n19984 & n26978;
assign n7023 = ~(n14663 ^ n20247);
assign n17294 = n8707 | n2807;
assign n8683 = n3995 | n26333;
assign n17901 = ~(n11448 ^ n1391);
assign n7533 = n5276 | n16810;
assign n22076 = ~(n13589 ^ n12476);
assign n25457 = n16129 | n396;
assign n25564 = n6645 & n17379;
assign n1562 = ~n3245;
assign n9441 = ~(n8381 ^ n23775);
assign n21890 = n20429 | n14922;
assign n17627 = n12671 | n15196;
assign n12505 = ~(n21272 | n3015);
assign n14721 = ~n23568;
assign n20746 = n20821 | n7972;
assign n13077 = n14438 | n13265;
assign n2469 = ~(n24031 | n6204);
assign n26149 = ~n19104;
assign n14337 = ~n4964;
assign n22842 = n21088 | n11247;
assign n13012 = n7025 | n7706;
assign n21785 = ~(n1689 ^ n17095);
assign n7166 = n4854 | n23862;
assign n4438 = n22579 & n18834;
assign n3886 = n7605 | n13518;
assign n4042 = ~(n4447 ^ n16786);
assign n24868 = ~n8845;
assign n5402 = ~n2173;
assign n4759 = ~(n5270 ^ n610);
assign n22344 = n20406 & n24013;
assign n21508 = ~(n4428 ^ n17140);
assign n12501 = n20923 | n7983;
assign n23819 = ~(n14629 ^ n17244);
assign n9552 = ~(n1375 ^ n10447);
assign n11791 = ~(n13359 | n1);
assign n21866 = n8423 | n358;
assign n20719 = ~(n931 ^ n3792);
assign n16685 = n2008 & n21478;
assign n17921 = n11993 | n8541;
assign n15912 = n21236 | n23738;
assign n26987 = n20070 | n11222;
assign n8076 = ~n4923;
assign n13725 = ~n27102;
assign n20329 = ~n3349;
assign n25404 = n3098 & n21296;
assign n19098 = ~(n25178 ^ n25103);
assign n13844 = ~(n23037 ^ n21409);
assign n21197 = n21435 | n9643;
assign n24097 = ~(n14333 ^ n9532);
assign n11785 = ~(n18333 | n20316);
assign n2885 = ~(n5471 ^ n12679);
assign n12591 = ~(n22254 | n8067);
assign n16180 = n18514 | n25261;
assign n7774 = n4053 | n13846;
assign n7113 = n25109 | n7187;
assign n17900 = ~(n9010 ^ n5707);
assign n18933 = ~(n27111 ^ n24701);
assign n4294 = ~(n6515 ^ n3282);
assign n16478 = n5132 | n18146;
assign n12743 = ~(n11060 | n25249);
assign n16611 = ~n23264;
assign n13724 = n1265 | n18308;
assign n24174 = n21281 | n20656;
assign n1157 = n11393 | n5580;
assign n16183 = ~(n9799 ^ n414);
assign n9578 = n11968 | n20958;
assign n9751 = n24205 & n6069;
assign n9928 = ~(n26234 ^ n23033);
assign n16194 = n2707 & n6755;
assign n20785 = n10221 & n9052;
assign n936 = n12017 | n15807;
assign n24971 = n19915 | n21985;
assign n8477 = ~n19060;
assign n23219 = n21113 | n21945;
assign n25588 = ~(n22527 | n24032);
assign n3352 = ~(n4384 ^ n21778);
assign n7891 = ~(n24383 ^ n6403);
assign n23110 = n5620 & n23814;
assign n21357 = ~(n14040 ^ n24711);
assign n21190 = n12375 | n17003;
assign n26528 = ~(n6429 ^ n20757);
assign n15351 = n5670 & n1800;
assign n4214 = n8419 | n24580;
assign n22799 = n7019 | n17649;
assign n2178 = n19551 & n2705;
assign n16653 = n1776 & n17962;
assign n7997 = ~(n19184 | n14661);
assign n409 = ~(n22309 ^ n19107);
assign n7542 = n18517 | n15759;
assign n13820 = n871 & n7412;
assign n8666 = n8254 | n17874;
assign n26516 = n940 | n8462;
assign n12880 = ~(n14484 ^ n21617);
assign n815 = n11343 & n23618;
assign n17970 = n488 | n5121;
assign n13625 = ~(n25675 ^ n21477);
assign n11372 = n2737 & n24303;
assign n14707 = ~(n647 | n26408);
assign n1599 = ~(n6643 ^ n21252);
assign n19720 = ~(n19789 ^ n21226);
assign n5715 = ~n7841;
assign n2164 = ~(n12457 ^ n11758);
assign n14651 = ~n10093;
assign n12014 = ~n23493;
assign n8063 = n26272 & n3184;
assign n2060 = ~n10629;
assign n25179 = n23345 | n26788;
assign n12194 = ~(n1594 ^ n762);
assign n16421 = ~n16410;
assign n14662 = n17960 | n7418;
assign n14661 = ~(n24931 ^ n7890);
assign n3454 = ~n14466;
assign n410 = ~(n1510 ^ n24150);
assign n25879 = ~(n11743 | n13301);
assign n3888 = n19558 | n4648;
assign n9349 = n23477 | n1334;
assign n5041 = n1694 | n8206;
assign n6059 = n2146 | n20216;
assign n13674 = n21674 & n5090;
assign n11476 = ~(n8696 ^ n1593);
assign n23366 = ~(n23041 ^ n6172);
assign n15817 = ~(n18163 ^ n21784);
assign n8534 = n24452 & n13528;
assign n9339 = n370 & n23022;
assign n17513 = n23244 | n23842;
assign n6247 = ~(n15801 | n26047);
assign n18978 = n2237 & n20475;
assign n22271 = ~(n23207 | n15930);
assign n26772 = n23800 | n3445;
assign n15397 = ~(n7524 ^ n15967);
assign n19280 = n18844 & n17107;
assign n25676 = ~n25054;
assign n21008 = ~(n18855 ^ n20218);
assign n26893 = n8770 & n2286;
assign n13666 = n27046 | n24125;
assign n19313 = n6678;
assign n25379 = n22365 | n11356;
assign n26006 = ~(n3062 ^ n11185);
assign n12794 = n1220 | n13950;
assign n18257 = ~n3030;
assign n9813 = ~(n22729 | n21698);
assign n14828 = n6712 | n26501;
assign n5377 = ~(n17412 ^ n22562);
assign n23866 = ~(n9246 | n23120);
assign n10276 = n25246 & n24728;
assign n7864 = ~(n22571 ^ n11792);
assign n307 = ~(n18149 ^ n19103);
assign n15856 = ~(n17549 | n4095);
assign n10305 = ~(n21764 ^ n23900);
assign n3009 = ~n13137;
assign n20145 = ~n448;
assign n19712 = ~(n933 | n5378);
assign n21835 = n22759 | n19066;
assign n11919 = ~n20700;
assign n23587 = ~(n7429 ^ n9323);
assign n8872 = n10008 | n27025;
assign n18785 = ~n8207;
assign n5743 = ~n20176;
assign n19823 = n6889 & n2648;
assign n13992 = ~(n11583 | n17959);
assign n20603 = ~(n15918 ^ n21735);
assign n16362 = n19041 | n21006;
assign n20788 = ~(n14279 ^ n6921);
assign n14943 = ~n7568;
assign n18259 = n24877 | n26549;
assign n10412 = n22171 & n12283;
assign n24986 = n11852 & n15037;
assign n8292 = ~(n17924 ^ n27098);
assign n1673 = ~(n11408 | n15787);
assign n11376 = ~(n6262 ^ n945);
assign n25669 = ~(n7692 | n25464);
assign n10410 = ~n1050;
assign n24669 = n21702 | n7815;
assign n23377 = n7664 | n13678;
assign n12698 = ~(n27142 | n9312);
assign n26900 = ~(n12523 ^ n4454);
assign n17014 = ~(n3324 | n4299);
assign n5043 = n13977 & n14650;
assign n25790 = n10137 & n26298;
assign n24094 = n22138 | n10086;
assign n19034 = n12280 & n24520;
assign n15002 = ~(n24598 ^ n22326);
assign n12699 = ~n18052;
assign n24041 = ~(n20542 | n9575);
assign n18532 = ~(n6645 ^ n7050);
assign n2021 = ~(n22173 ^ n24032);
assign n8273 = n24171 | n11671;
assign n509 = n15973 | n21631;
assign n12940 = ~(n19025 | n9655);
assign n9062 = n14442 | n2634;
assign n634 = n18214 & n900;
assign n18789 = n12871 & n8888;
assign n9510 = ~(n455 ^ n3603);
assign n20576 = n18452 | n3118;
assign n18181 = ~(n10408 ^ n14899);
assign n2390 = ~(n21710 ^ n25237);
assign n9819 = n16236 | n20019;
assign n17904 = n25972 | n3707;
assign n6238 = n8782 & n24561;
assign n15299 = ~(n23114 ^ n3454);
assign n6891 = ~(n8000 ^ n22156);
assign n23847 = n2754 & n9195;
assign n9107 = ~n22591;
assign n2026 = n25156 | n2073;
assign n13846 = ~(n10792 ^ n19922);
assign n10767 = ~(n4617 ^ n24261);
assign n16890 = ~n1682;
assign n7673 = n12882 & n3325;
assign n18439 = ~(n4949 ^ n14170);
assign n20479 = ~n24612;
assign n9644 = n9172 | n10571;
assign n25788 = n27114 | n3247;
assign n1062 = ~n21906;
assign n10771 = ~(n23230 | n10053);
assign n9287 = ~(n3859 ^ n21603);
assign n4944 = n7912 & n18949;
assign n26860 = ~(n6064 ^ n4405);
assign n24612 = ~(n3994 ^ n19228);
assign n1229 = n24928 | n18187;
assign n3927 = ~(n3981 | n24818);
assign n26737 = n25188 | n1042;
assign n1874 = n9149 | n23564;
assign n15208 = n19804 | n13567;
assign n5887 = ~(n7693 | n9453);
assign n4300 = ~(n10158 ^ n3952);
assign n24568 = ~(n5925 ^ n9058);
assign n452 = n8192 | n26716;
assign n2915 = ~n11481;
assign n6271 = ~(n23439 ^ n7573);
assign n10440 = n19689 & n16384;
assign n2662 = n19797 | n21497;
assign n685 = ~(n1328 ^ n13987);
assign n4745 = ~(n8915 ^ n27067);
assign n9781 = n13838 & n3357;
assign n8038 = n9326 | n1466;
assign n6327 = ~n6283;
assign n2273 = n16588 | n27047;
assign n5663 = n23250 | n16856;
assign n6738 = n17748 & n47;
assign n20909 = ~(n22327 | n4559);
assign n407 = ~(n15720 ^ n18512);
assign n10752 = n22365 | n20429;
assign n10538 = ~(n21998 ^ n25779);
assign n9702 = ~(n19366 ^ n11184);
assign n2396 = n5794 | n12744;
assign n27172 = ~n14386;
assign n19321 = ~n12121;
assign n14192 = n11177 & n10254;
assign n24173 = n193 | n19415;
assign n12238 = ~(n1802 | n7331);
assign n17938 = ~n11688;
assign n9103 = n19161 | n7966;
assign n15661 = ~n7940;
assign n5721 = n2118 & n19960;
assign n5677 = ~(n10763 ^ n5696);
assign n22206 = ~n4714;
assign n21884 = n8601 & n23815;
assign n14824 = n15207 & n21787;
assign n10019 = ~(n22806 ^ n19972);
assign n12659 = ~(n12090 ^ n12018);
assign n20005 = ~(n7540 ^ n7944);
assign n1244 = n238 & n24333;
assign n26609 = ~(n18263 ^ n12475);
assign n25884 = ~(n8661 ^ n8496);
assign n17016 = n16551 | n19166;
assign n7494 = n12543 | n4934;
assign n17144 = n4490 | n1949;
assign n27031 = ~(n22564 ^ n772);
assign n16859 = ~(n23558 ^ n12421);
assign n5748 = n5434 | n10074;
assign n16168 = ~(n18173 | n5101);
assign n25942 = ~n22850;
assign n21153 = n19 | n26673;
assign n1911 = n24575 & n15232;
assign n8263 = n11256 | n745;
assign n4394 = n2413 | n10449;
assign n16696 = ~(n21058 ^ n9111);
assign n4818 = ~n21361;
assign n7145 = ~(n14016 ^ n14102);
assign n25536 = ~(n16626 | n1998);
assign n23640 = ~(n14089 | n15930);
assign n6526 = n4311 & n11660;
assign n1614 = n20476 | n6159;
assign n14523 = ~(n24475 | n14749);
assign n21481 = n442 & n6319;
assign n12588 = n2505 | n6969;
assign n24524 = ~(n16091 | n16602);
assign n2391 = ~n14091;
assign n5349 = ~(n5563 ^ n20239);
assign n13235 = ~(n21280 ^ n24364);
assign n11265 = n21471 | n22014;
assign n16005 = n11180 & n20510;
assign n24878 = n8499 & n8388;
assign n10258 = ~n7612;
assign n13796 = ~(n12014 | n8405);
assign n11225 = ~(n13494 ^ n18880);
assign n6128 = ~(n3686 ^ n21155);
assign n14836 = n675 & n14934;
assign n14804 = n16996 & n22025;
assign n7108 = ~(n22428 ^ n1269);
assign n11521 = ~(n6753 | n8779);
assign n7704 = n9679 | n13405;
assign n5232 = n4619 & n10901;
assign n12707 = ~(n8817 ^ n19583);
assign n23731 = ~(n22904 ^ n19571);
assign n8287 = n13600 & n14108;
assign n15361 = ~(n7785 | n8853);
assign n15597 = n18253 | n5756;
assign n18762 = n14344 | n6521;
assign n8143 = n14569 | n24049;
assign n9784 = ~(n9768 | n16276);
assign n3675 = ~n4723;
assign n27011 = ~(n24773 ^ n7492);
assign n14504 = n11583 & n14085;
assign n22037 = n20905 | n8670;
assign n17819 = n23528 & n10852;
assign n16703 = ~(n16722 ^ n13708);
assign n7748 = n21213 | n4685;
assign n1433 = ~n7002;
assign n16504 = n19881 & n11532;
assign n24248 = n8076 | n22031;
assign n14200 = ~(n5559 ^ n26036);
assign n6093 = ~n22435;
assign n24584 = ~n13085;
assign n1890 = ~n25312;
assign n4769 = ~(n21073 | n15975);
assign n13094 = ~(n6632 ^ n1831);
assign n21348 = n14123 & n2494;
assign n16485 = n26312 | n17453;
assign n2758 = ~(n26065 ^ n13136);
assign n8769 = ~(n8704 ^ n15596);
assign n9972 = ~(n16737 ^ n10342);
assign n10110 = n6709 | n24386;
assign n11030 = ~n5028;
assign n20298 = n23695 | n854;
assign n11410 = ~(n22688 | n3474);
assign n26557 = ~(n7336 ^ n11105);
assign n4365 = ~(n26408 | n12477);
assign n4415 = n4614 & n15132;
assign n24337 = n25749 | n22082;
assign n25598 = n18386 | n6689;
assign n11678 = n2688 | n8163;
assign n7434 = n16465 | n5709;
assign n14401 = ~n20104;
assign n1722 = ~(n13936 ^ n11201);
assign n21799 = n23835 | n10947;
assign n1128 = n23932 | n2606;
assign n13003 = ~(n20754 ^ n593);
assign n8071 = ~n13915;
assign n1195 = ~(n16966 ^ n14796);
assign n21411 = n15938 | n5747;
assign n14896 = n4799 | n11411;
assign n9288 = n3974 & n717;
assign n386 = n23281 & n5142;
assign n25231 = n24687 & n23301;
assign n24728 = ~(n10953 ^ n2734);
assign n20214 = ~(n1118 | n20489);
assign n8025 = ~(n22686 ^ n15464);
assign n14990 = n22536 | n22955;
assign n15207 = n13360 | n16724;
assign n15459 = n8532 | n22685;
assign n22754 = n14337 & n24865;
assign n21149 = n5968 | n5180;
assign n10443 = ~(n25119 | n12652);
assign n24577 = n15890 | n1384;
assign n11320 = n15235 & n10545;
assign n25700 = ~n7538;
assign n23346 = n11505 & n24352;
assign n3586 = n20044 & n11835;
assign n22483 = n4809 & n6114;
assign n17579 = ~n1831;
assign n4017 = ~n10873;
assign n17716 = ~n23820;
assign n25525 = ~(n8455 ^ n24835);
assign n23136 = n26342 & n26906;
assign n26697 = n10840 | n14914;
assign n6013 = ~(n20608 ^ n6195);
assign n13864 = n15054 | n25031;
assign n4032 = ~n10652;
assign n26570 = n9526 | n25349;
assign n17648 = n4200 & n19302;
assign n6641 = ~(n14139 | n24152);
assign n26347 = n10151 | n5324;
assign n19809 = n716 & n15543;
assign n26591 = n10090 | n16377;
assign n30 = n11058 & n14616;
assign n10671 = ~(n12375 | n22765);
assign n2781 = n8574 & n22188;
assign n8222 = n19327 & n25624;
assign n5940 = ~(n12821 ^ n5579);
assign n2443 = ~(n17964 ^ n20651);
assign n131 = ~(n1262 | n9557);
assign n7567 = ~(n6037 ^ n5376);
assign n6993 = n867 & n11341;
assign n16011 = ~(n11751 ^ n3245);
assign n13400 = ~(n22965 ^ n19791);
assign n9867 = ~(n24279 ^ n3296);
assign n25549 = n26091 & n17349;
assign n18370 = ~(n23686 | n8084);
assign n8826 = ~(n22480 ^ n7020);
assign n24516 = n24684 & n12880;
assign n17314 = ~(n14845 ^ n2274);
assign n14717 = ~(n13872 | n14279);
assign n26594 = ~(n24813 ^ n9396);
assign n2058 = ~(n3123 ^ n4393);
assign n26031 = n0 & n22796;
assign n5089 = n930 | n2638;
assign n8545 = ~(n11336 ^ n10201);
assign n811 = ~(n22375 | n5722);
assign n7625 = n8979 | n13263;
assign n22234 = ~n15384;
assign n20580 = n22889 & n24790;
assign n12975 = ~(n26056 ^ n27151);
assign n23696 = n13335 & n11547;
assign n6310 = n10964 | n17159;
assign n24916 = ~(n15456 ^ n18880);
assign n2374 = ~(n7908 ^ n12723);
assign n12854 = n24077 | n17615;
assign n7423 = ~(n2055 | n17938);
assign n12613 = n2415 & n8414;
assign n25241 = ~(n25753 ^ n26018);
assign n8271 = ~(n1731 ^ n16430);
assign n25561 = ~(n9881 ^ n12741);
assign n19733 = ~(n12153 | n9490);
assign n24649 = ~n19608;
assign n22285 = ~n12098;
assign n8758 = n25282 | n10577;
assign n27085 = n17892 | n3371;
assign n6170 = ~n2548;
assign n25602 = ~(n27156 ^ n3909);
assign n12416 = ~n25316;
assign n24518 = ~(n8439 ^ n3710);
assign n23692 = ~(n2823 ^ n3630);
assign n9237 = ~n9931;
assign n8278 = n9586 & n12778;
assign n12372 = n8797 | n23485;
assign n3280 = ~n2574;
assign n6149 = ~(n10217 ^ n11011);
assign n16584 = ~(n3023 ^ n14320);
assign n9708 = n10497 & n6656;
assign n17203 = ~n17255;
assign n11039 = ~n20389;
assign n13227 = ~(n10324 | n13719);
assign n10400 = n15367 & n8350;
assign n25323 = ~(n10593 ^ n1662);
assign n2101 = ~(n16496 ^ n17647);
assign n22987 = ~n655;
assign n13634 = n24599 | n12766;
assign n6949 = ~(n5606 ^ n1698);
assign n25634 = ~(n18788 | n15288);
assign n2493 = n10835 | n7490;
assign n13543 = ~(n14090 ^ n18962);
assign n19162 = ~(n7530 ^ n4189);
assign n7069 = ~(n23851 ^ n4100);
assign n21443 = n18537 | n10920;
assign n24747 = n19451 & n25828;
assign n20846 = n8467 | n4128;
assign n24893 = n7081 | n24213;
assign n16375 = ~(n10962 ^ n16789);
assign n22962 = ~n6631;
assign n16806 = ~(n20365 | n8083);
assign n22010 = n2590 | n21901;
assign n11951 = n682 | n5075;
assign n18756 = ~(n20719 ^ n22918);
assign n8698 = n20040 | n16555;
assign n22598 = n20324 | n810;
assign n18250 = n21977 & n8817;
assign n12033 = n22500 & n21601;
assign n17592 = ~(n6615 ^ n22493);
assign n2192 = ~(n11958 | n1036);
assign n20691 = ~(n23759 ^ n13984);
assign n18334 = n2976 & n10904;
assign n24074 = ~n10854;
assign n7520 = ~n6834;
assign n14539 = ~n14215;
assign n874 = ~n3919;
assign n7933 = ~n7516;
assign n23827 = n13153 & n9230;
assign n1431 = ~(n18974 ^ n26380);
assign n26805 = ~n2099;
assign n16726 = n12551 | n23442;
assign n11817 = n1999 | n766;
assign n12730 = ~(n23877 ^ n9830);
assign n64 = ~n18815;
assign n16707 = ~(n912 ^ n5131);
assign n13960 = ~n12236;
assign n24435 = ~(n10505 | n6925);
assign n10550 = n13229 & n18670;
assign n11915 = n20358 & n3960;
assign n10032 = ~(n16038 ^ n18794);
assign n24904 = ~(n15405 | n3940);
assign n10837 = ~n19680;
assign n25053 = ~(n12488 ^ n1437);
assign n10702 = n22547 & n10428;
assign n7504 = ~(n26458 | n6073);
assign n20708 = ~(n13915 | n23644);
assign n2346 = ~n5899;
assign n8448 = ~(n14291 ^ n20285);
assign n3263 = ~(n1554 ^ n21397);
assign n24480 = ~(n7860 ^ n13719);
assign n9272 = n2329 | n2753;
assign n14917 = ~(n3990 ^ n5349);
assign n10557 = n12322;
assign n5866 = ~(n20384 ^ n8008);
assign n4155 = ~n13502;
assign n7479 = ~(n19227 ^ n8381);
assign n21568 = n25836 & n23569;
assign n20067 = n24157 | n1910;
assign n19431 = n25234 & n9405;
assign n19880 = ~(n2156 | n5796);
assign n22850 = ~(n21851 ^ n20868);
assign n15861 = ~(n7339 ^ n26808);
assign n16923 = ~(n21678 ^ n24616);
assign n23058 = ~(n6126 ^ n1420);
assign n14153 = ~(n17876 ^ n17508);
assign n14563 = ~(n27104 | n13317);
assign n3518 = ~(n212 | n9928);
assign n5283 = ~n26667;
assign n18114 = ~n5976;
assign n7207 = n20568 & n9861;
assign n18553 = ~(n1798 ^ n8930);
assign n1930 = n16022 | n1519;
assign n755 = ~(n7574 ^ n16675);
assign n26198 = n21450 | n4870;
assign n6179 = ~(n5092 ^ n19270);
assign n10481 = n11798 | n7509;
assign n23151 = ~(n2481 ^ n9477);
assign n9527 = ~(n17022 ^ n9506);
assign n13654 = ~(n7752 ^ n12541);
assign n15109 = ~n15146;
assign n15350 = n446 | n13349;
assign n19801 = n20071 | n12026;
assign n17366 = ~n18790;
assign n17738 = ~(n5890 | n22838);
assign n26396 = n10417 | n8362;
assign n21385 = ~(n12474 ^ n15713);
assign n25443 = n20921 | n22552;
assign n12313 = ~(n23962 ^ n2274);
assign n25808 = ~(n21585 ^ n23146);
assign n12595 = n2354 | n8940;
assign n7890 = ~(n19282 ^ n26986);
assign n7601 = n3285 & n21463;
assign n3624 = n1665 | n19269;
assign n21093 = ~(n15800 ^ n3772);
assign n18490 = n7384 | n6931;
assign n24308 = n12708 | n9529;
assign n15754 = n14605 & n22010;
assign n12111 = ~n14382;
assign n17854 = ~(n2867 ^ n20756);
assign n9584 = ~n15910;
assign n23748 = ~(n8811 ^ n645);
assign n3653 = ~(n19155 ^ n27192);
assign n22429 = n2372 | n12347;
assign n198 = ~n9028;
assign n21189 = ~(n25160 ^ n18290);
assign n25400 = ~(n7818 | n13851);
assign n16166 = ~(n25403 ^ n22973);
assign n25509 = ~n4345;
assign n13550 = n11144 | n11640;
assign n7697 = ~n9527;
assign n14028 = n25348 & n7153;
assign n14116 = n17844 & n1962;
assign n18099 = ~(n8107 | n18363);
assign n15163 = n13901 | n4860;
assign n18841 = ~n26703;
assign n11451 = ~(n15626 ^ n5302);
assign n2439 = n4178 | n16763;
assign n15731 = n12276 | n22992;
assign n17820 = ~(n8034 ^ n19724);
assign n17259 = n9839 & n6754;
assign n5105 = ~(n4599 ^ n7305);
assign n14837 = n15643 | n3393;
assign n10968 = n14132 | n3338;
assign n13571 = n378 & n5779;
assign n18264 = n3840 & n24908;
assign n12750 = n21516 & n26336;
assign n15076 = n14323 & n12351;
assign n18100 = ~n13319;
assign n22017 = ~(n21116 ^ n1448);
assign n14637 = ~(n21725 ^ n19283);
assign n18306 = n9976 | n13702;
assign n14330 = ~(n13006 ^ n15092);
assign n4442 = ~n6037;
assign n24462 = ~(n11938 | n8244);
assign n10002 = ~(n24244 | n11577);
assign n15250 = n9826 | n26505;
assign n8910 = ~n3925;
assign n15117 = n7172 | n19806;
assign n12600 = n9910 | n20342;
assign n12868 = ~n4429;
assign n15504 = ~(n11303 | n23200);
assign n19639 = n19340 & n234;
assign n4288 = ~(n10328 ^ n7579);
assign n21637 = ~(n11206 ^ n6840);
assign n8338 = ~(n19929 ^ n23787);
assign n3087 = n18067 | n2333;
assign n15502 = ~n20391;
assign n24279 = n18852 | n20815;
assign n5351 = ~(n51 ^ n21513);
assign n18043 = ~(n19591 ^ n22667);
assign n8574 = n10159 | n14790;
assign n7311 = ~n2088;
assign n15419 = n11831 | n14777;
assign n20880 = ~n7721;
assign n23781 = n18649 & n11278;
assign n5944 = n21325 & n27069;
assign n7161 = n12143 & n20215;
assign n5896 = n12359 | n22528;
assign n17358 = n14027 & n23421;
assign n19146 = ~(n6170 ^ n5115);
assign n10101 = ~(n15510 ^ n22496);
assign n23549 = n25218 | n5527;
assign n883 = ~(n26951 | n27054);
assign n6051 = ~n12341;
assign n21948 = ~(n2720 ^ n21228);
assign n24012 = n10040 & n9810;
assign n17470 = ~(n24331 ^ n24798);
assign n21559 = ~(n21317 ^ n13110);
assign n14351 = n8976 & n2466;
assign n15947 = n2607 & n11687;
assign n21042 = n8694 | n6900;
assign n4431 = n13293 | n17388;
assign n20466 = ~(n22422 | n13521);
assign n16287 = ~(n5527 ^ n6551);
assign n15768 = n16873 | n6591;
assign n17980 = n16699 & n11621;
assign n27018 = ~n16058;
assign n5698 = n15695 | n18;
assign n18711 = ~(n9399 ^ n14275);
assign n6618 = n15101 | n3663;
assign n3288 = n23105 & n19637;
assign n22098 = n19777 | n17036;
assign n16961 = ~n10869;
assign n22237 = ~n4509;
assign n12902 = ~n7314;
assign n21987 = n2175 | n4484;
assign n24549 = ~(n11707 | n13643);
assign n436 = n16053 & n1807;
assign n4170 = ~n9489;
assign n14784 = n26082 | n5210;
assign n25946 = ~(n22176 ^ n23065);
assign n18072 = n19669 & n23933;
assign n20168 = n18120 & n11620;
assign n14231 = ~(n10593 ^ n19701);
assign n24817 = n2081 & n8693;
assign n24396 = n2692 | n21394;
assign n4524 = ~(n4897 ^ n8772);
assign n2855 = n26132 | n23184;
assign n15859 = ~(n3191 ^ n25831);
assign n8686 = n3927 | n10912;
assign n16384 = n11913 | n14109;
assign n9074 = n24277 | n20863;
assign n8257 = n4969 | n18390;
assign n5626 = ~(n10000 ^ n6790);
assign n22390 = ~(n21101 ^ n17779);
assign n3233 = ~(n5320 ^ n19663);
assign n23638 = ~(n8745 | n24278);
assign n20319 = n23833 | n13558;
assign n3859 = n17438 | n22490;
assign n24270 = n11440 | n25111;
assign n18282 = ~(n4217 ^ n25565);
assign n13321 = n8975 | n26939;
assign n7211 = ~(n2666 ^ n14739);
assign n12780 = ~n2197;
assign n16644 = n14646 | n22543;
assign n20694 = ~(n25643 ^ n21753);
assign n17202 = ~(n26527 ^ n18686);
assign n10200 = n20998 | n20250;
assign n26708 = n2570 | n17239;
assign n11774 = n12020 | n26447;
assign n26589 = n18646 | n1140;
assign n23099 = n7221;
assign n15675 = ~(n1931 ^ n9980);
assign n15088 = n24053 & n2727;
assign n19509 = n25277 & n21860;
assign n1609 = ~(n17726 | n14969);
assign n6743 = ~n11435;
assign n4731 = ~(n17148 ^ n9807);
assign n2676 = n23210 & n18127;
assign n20634 = n24305 & n2580;
assign n14879 = ~(n8255 | n5625);
assign n23026 = n13537 & n18285;
assign n3749 = ~(n24575 | n15232);
assign n840 = ~n11580;
assign n3296 = ~(n18283 ^ n13400);
assign n16558 = ~(n7364 ^ n2102);
assign n21457 = n9601 & n26070;
assign n24756 = n26167 & n18554;
assign n13133 = ~(n24090 ^ n13110);
assign n23873 = ~(n27040 ^ n3711);
assign n19777 = n15411 & n1079;
assign n22083 = n3429;
assign n9342 = n22384 & n26910;
assign n21561 = ~(n23670 ^ n23775);
assign n17920 = ~(n16427 ^ n1807);
assign n6108 = n24766 | n19529;
assign n14168 = ~n26572;
assign n15254 = ~(n23504 ^ n13940);
assign n2736 = n9752 & n4467;
assign n4316 = ~n9936;
assign n15745 = n8051 & n25573;
assign n10265 = ~(n4040 | n655);
assign n20375 = n11600 | n2423;
assign n24363 = ~(n22764 ^ n1536);
assign n1479 = ~(n15229 | n8050);
assign n22233 = n6901 & n23385;
assign n20063 = n22673 | n16265;
assign n16920 = n2957 | n19285;
assign n18498 = ~n9983;
assign n14963 = ~n8067;
assign n14642 = ~n3770;
assign n18809 = n26030 | n3752;
assign n15316 = ~(n17411 ^ n3915);
assign n18361 = ~(n14393 | n26239);
assign n4616 = ~(n5380 ^ n19296);
assign n1792 = ~(n8879 ^ n6544);
assign n24311 = ~(n3600 ^ n12836);
assign n12696 = ~(n20534 ^ n17131);
assign n23978 = ~(n23266 ^ n7580);
assign n10624 = ~(n12567 ^ n12279);
assign n20410 = ~(n16400 ^ n17561);
assign n10092 = ~(n9923 ^ n767);
assign n26916 = n26371 | n2418;
assign n2553 = ~(n16652 ^ n12141);
assign n26832 = ~(n511 ^ n703);
assign n18328 = ~(n11318 | n2615);
assign n12881 = n13237 & n1066;
assign n14997 = n21514 | n7947;
assign n10714 = ~(n14361 ^ n18511);
assign n16284 = n23828 & n26346;
assign n16425 = n23311 | n284;
assign n18858 = ~(n169 ^ n13934);
assign n23721 = n19358 | n25302;
assign n26543 = ~(n2160 | n7335);
assign n4261 = n24981 & n4091;
assign n23138 = n26067 | n6643;
assign n15540 = n20293 | n22006;
assign n17253 = ~(n12821 ^ n6596);
assign n24080 = ~(n262 ^ n4489);
assign n20877 = n15261 & n14630;
assign n17918 = n24130 | n4721;
assign n24541 = n8633 & n22810;
assign n25915 = ~n5703;
assign n5313 = ~n11737;
assign n2540 = ~(n25625 ^ n6132);
assign n18499 = ~(n5330 | n919);
assign n22643 = ~(n8856 ^ n8305);
assign n24027 = n525 | n2501;
assign n21623 = ~(n15257 ^ n604);
assign n12309 = n15202 | n25805;
assign n389 = ~(n13944 ^ n23871);
assign n10551 = ~(n26876 ^ n1662);
assign n4434 = ~(n13177 ^ n3164);
assign n9214 = n4237 & n4495;
assign n17533 = n13410 | n12564;
assign n26340 = ~n13936;
assign n3562 = n4378 & n23929;
assign n14739 = ~n15153;
assign n25153 = n25928 | n17109;
assign n12649 = ~(n19297 | n21248);
assign n19675 = n7974 | n23369;
assign n8419 = ~n15931;
assign n14463 = ~(n19065 ^ n26232);
assign n9329 = n14162 | n1947;
assign n25771 = n12183 | n26017;
assign n26062 = ~n6790;
assign n2325 = n7287 & n20154;
assign n6420 = n5884 & n26468;
assign n12692 = ~n12102;
assign n21885 = ~(n1777 ^ n4812);
assign n16972 = ~(n25830 ^ n23897);
assign n10798 = n3252 | n7637;
assign n26866 = ~(n13267 ^ n16310);
assign n24746 = ~(n9113 ^ n25643);
assign n9855 = ~(n23173 | n15046);
assign n8272 = ~(n2255 ^ n12558);
assign n4778 = n7089 | n16793;
assign n10294 = n4741 | n17818;
assign n21323 = ~(n1532 ^ n25426);
assign n17880 = ~(n9069 ^ n22169);
assign n20155 = n9099 | n19067;
assign n24527 = n15334 | n11084;
assign n3958 = n18205 | n18595;
assign n22469 = n17451 & n22343;
assign n19261 = ~(n20655 ^ n23170);
assign n26521 = ~n12717;
assign n26868 = n8869 | n1738;
assign n3128 = n12073 & n14234;
assign n25445 = n26186 & n19556;
assign n22186 = ~n12426;
assign n2917 = n7237 | n2813;
assign n4834 = ~(n1329 ^ n12315);
assign n17467 = ~n21353;
assign n19437 = n25171 | n7946;
assign n16589 = ~(n17025 ^ n14419);
assign n3716 = ~(n13175 ^ n9567);
assign n20925 = ~(n9548 ^ n1885);
assign n18175 = ~(n3612 | n21274);
assign n12551 = ~(n24862 | n24996);
assign n14218 = ~n2575;
assign n21644 = ~n25370;
assign n5812 = ~n19058;
assign n12816 = ~(n3331 ^ n1023);
assign n14295 = n333 | n19017;
assign n22821 = ~(n16812 ^ n1279);
assign n18255 = ~n18108;
assign n26048 = n10109 & n26742;
assign n24029 = n7155 | n805;
assign n445 = n24721 | n863;
assign n16241 = ~(n524 | n7566);
assign n25681 = n18825 & n21866;
assign n4095 = ~(n22405 ^ n24416);
assign n18817 = n17413 & n12340;
assign n21054 = n10274 | n18108;
assign n12006 = n26997 | n23746;
assign n24178 = n2368 & n9029;
assign n10543 = n5900 & n23079;
assign n17330 = n13031 & n9615;
assign n6047 = n10957 & n12758;
assign n25746 = n26897 | n5217;
assign n14967 = ~n7788;
assign n14630 = ~n16902;
assign n8789 = n6507 & n9524;
assign n24390 = n1274 & n17469;
assign n25110 = ~n17239;
assign n15494 = n14730 | n13308;
assign n15420 = n23073 | n8190;
assign n553 = ~n2583;
assign n23061 = ~n26332;
assign n18162 = n7297 | n24102;
assign n11837 = ~(n4353 ^ n17903);
assign n26764 = ~(n18344 ^ n2965);
assign n11604 = n13269 | n13022;
assign n3837 = ~(n15743 ^ n20658);
assign n21782 = n23914 | n16501;
assign n4817 = n13810 | n27024;
assign n5848 = ~n4578;
assign n5378 = ~n14886;
assign n9950 = ~(n22683 | n17553);
assign n27071 = ~n11429;
assign n5381 = ~(n22619 ^ n22043);
assign n24400 = n20372 & n6434;
assign n20461 = n22146 & n21709;
assign n13050 = ~(n4184 ^ n4075);
assign n4123 = ~(n10481 ^ n15802);
assign n22487 = ~(n5834 | n3186);
assign n622 = ~(n23114 ^ n27009);
assign n8754 = n19444 & n20689;
assign n20904 = n26038 | n8473;
assign n16868 = n69 & n8115;
assign n11780 = n17607 | n16470;
assign n1904 = ~n16183;
assign n12553 = ~(n1789 ^ n5246);
assign n4108 = ~(n7690 ^ n1428);
assign n13089 = ~(n4860 ^ n20248);
assign n4561 = n14337 & n23211;
assign n15770 = n9282 | n11962;
assign n290 = n15589 & n25531;
assign n431 = ~(n2603 ^ n14917);
assign n2889 = ~(n2813 ^ n1536);
assign n27007 = ~n25948;
assign n17058 = n26877 | n10440;
assign n24246 = n20857 | n4808;
assign n20783 = n14940 | n27029;
assign n21152 = n27139 | n24560;
assign n18729 = n11889 & n14249;
assign n10555 = ~(n10405 | n13960);
assign n26871 = n7935 & n18608;
assign n10833 = ~(n8291 ^ n14459);
assign n437 = n26689 & n12906;
assign n12959 = ~(n12208 ^ n27074);
assign n17618 = n24709 | n9997;
assign n25049 = ~n23048;
assign n23001 = n6393 | n25877;
assign n14157 = ~(n5727 ^ n6137);
assign n1642 = ~n3952;
assign n939 = n11902 & n10827;
assign n12578 = n20342 | n8526;
assign n24441 = ~(n2818 ^ n15536);
assign n24368 = ~(n16896 ^ n9303);
assign n9529 = n6627 & n4377;
assign n1657 = ~n18338;
assign n13799 = n10429 & n2627;
assign n11058 = n9797 | n6095;
assign n7267 = ~(n7193 ^ n16994);
assign n17197 = n7948 & n19321;
assign n5023 = n26320 & n6166;
assign n6867 = ~(n7202 ^ n11772);
assign n25425 = n21839 | n19282;
assign n8133 = ~(n6079 ^ n2483);
assign n19102 = n20243 | n10015;
assign n11976 = ~n25607;
assign n27121 = ~n3835;
assign n13342 = n26123 | n7456;
assign n27086 = n2453 | n1765;
assign n13671 = ~n22359;
assign n5133 = n17539 & n6377;
assign n16418 = n13564 | n12612;
assign n7758 = n18908 | n848;
assign n23596 = n5203 & n26048;
assign n19290 = n7582 | n15797;
assign n80 = ~(n22272 ^ n21654);
assign n21267 = ~(n10377 ^ n19731);
assign n10368 = n18678 & n12372;
assign n1774 = n7140 | n8641;
assign n20978 = ~n22607;
assign n26489 = ~(n4338 ^ n25106);
assign n13707 = n21269 | n5789;
assign n380 = n640 | n20227;
assign n16285 = n19872 & n360;
assign n21178 = n9143 | n16697;
assign n12515 = ~(n23332 ^ n2199);
assign n9682 = n12227 & n26558;
assign n5241 = n12537 & n283;
assign n20440 = n20066 & n24295;
assign n24036 = n296 | n16686;
assign n18702 = n24044 | n8937;
assign n4009 = ~(n18558 ^ n10411);
assign n183 = n8243 & n22190;
assign n18800 = ~n23545;
assign n21822 = ~(n9071 ^ n16071);
assign n3448 = ~n2439;
assign n16906 = n481 & n18111;
assign n9261 = ~(n12097 ^ n14810);
assign n25781 = n2235 & n22812;
assign n9753 = ~(n1003 ^ n23233);
assign n16237 = n14465 | n15204;
assign n18927 = n26315 & n9982;
assign n16735 = n22601 | n25727;
assign n10458 = n24500 | n10208;
assign n17011 = n14603 | n15053;
assign n18623 = n23909 & n3812;
assign n22742 = n22178 | n25783;
assign n763 = ~(n8507 ^ n15602);
assign n17155 = n13011 & n3104;
assign n25969 = n7373 | n13069;
assign n6673 = ~(n2587 ^ n21859);
assign n23745 = ~(n27169 ^ n26940);
assign n2220 = n1366 & n25084;
assign n6435 = n25947;
assign n15122 = ~(n16400 | n24907);
assign n3115 = ~n4743;
assign n19054 = n10086 | n20176;
assign n139 = ~(n25946 ^ n9380);
assign n20326 = ~n8292;
assign n5508 = ~(n20534 | n13146);
assign n25803 = n2663 | n7911;
assign n24948 = ~(n14555 ^ n23912);
assign n7931 = ~(n18749 ^ n4156);
assign n6609 = n21487 | n10749;
assign n11126 = n3906 | n16856;
assign n22830 = n9693 & n10767;
assign n1082 = ~(n24747 ^ n14737);
assign n14326 = ~(n9169 ^ n11304);
assign n2313 = ~(n20822 ^ n14692);
assign n16990 = n24844 | n16224;
assign n11308 = ~(n1600 ^ n5482);
assign n11518 = ~(n1578 | n20254);
assign n17157 = ~(n2852 ^ n1432);
assign n7842 = n26963 & n22828;
assign n8900 = ~(n1352 | n10844);
assign n14150 = ~(n2156 | n7402);
assign n20803 = ~(n19413 ^ n2288);
assign n10856 = n11909 | n12660;
assign n22943 = ~(n5938 | n25071);
assign n974 = n11342 & n4047;
assign n15941 = n23679 & n1569;
assign n26531 = n13227 | n21503;
assign n15756 = n3740 & n2545;
assign n27115 = ~n20618;
assign n564 = ~(n16166 ^ n14705);
assign n24682 = ~(n13 | n23792);
assign n11523 = ~(n23428 | n5834);
assign n11482 = ~(n17646 ^ n24393);
assign n8604 = ~(n21570 ^ n9598);
assign n7661 = ~(n23819 | n22861);
assign n11875 = ~(n14904 | n11575);
assign n9757 = ~(n4473 | n3798);
assign n24626 = ~(n14043 ^ n2076);
assign n7040 = n17122 & n23383;
assign n13507 = ~n5038;
assign n6555 = ~(n16755 ^ n367);
assign n4087 = ~n23333;
assign n9106 = ~(n18537 ^ n5211);
assign n7043 = n6164 & n25942;
assign n438 = n21517 & n16972;
assign n16424 = ~(n2854 ^ n2660);
assign n20825 = n21582 & n24553;
assign n13813 = n23472 & n20736;
assign n18848 = n852 | n13476;
assign n4315 = ~n19116;
assign n9905 = n2219 | n2813;
assign n24024 = ~n5737;
assign n24099 = n14626 & n20843;
assign n14613 = n21287 & n23705;
assign n9104 = ~(n24653 ^ n26602);
assign n5293 = n21869 | n21999;
assign n23723 = n2369 | n18899;
assign n21396 = ~(n13192 ^ n18050);
assign n21921 = n14958 | n5800;
assign n4785 = ~(n11934 ^ n2094);
assign n25968 = n6222 | n19378;
assign n22351 = ~n8194;
assign n18503 = ~(n1364 ^ n8256);
assign n11536 = n12147 | n9485;
assign n13533 = ~(n2225 ^ n11181);
assign n19170 = ~n2923;
assign n2297 = n16833 & n21910;
assign n4990 = n6236 & n13160;
assign n17753 = ~(n16197 | n24936);
assign n16291 = ~(n6143 ^ n1689);
assign n4071 = ~(n11247 ^ n19919);
assign n20128 = ~(n21378 | n14584);
assign n23052 = n3900 | n16202;
assign n6205 = n26087 | n7243;
assign n19326 = n27205 & n6858;
assign n17629 = ~(n6191 ^ n4935);
assign n13950 = ~(n10017 | n20349);
assign n2683 = n24435 | n21179;
assign n1598 = n21251 & n10830;
assign n10065 = ~(n9259 ^ n6456);
assign n4529 = ~(n27023 ^ n10818);
assign n25860 = n21845 | n8247;
assign n2896 = ~n16911;
assign n11000 = ~n20925;
assign n5724 = n25139 | n16696;
assign n16477 = ~n14723;
assign n2707 = n9509 | n6566;
assign n643 = ~(n8300 ^ n12761);
assign n7402 = ~(n14334 ^ n23393);
assign n14314 = ~(n2391 ^ n19647);
assign n13768 = n23111 | n18536;
assign n13423 = n4522 | n1579;
assign n22517 = ~n20621;
assign n1313 = ~(n21828 ^ n18227);
assign n11090 = n8856 | n19768;
assign n989 = n25931 & n1510;
assign n1391 = ~(n13734 ^ n18548);
assign n25587 = n22622 | n16535;
assign n11168 = ~(n1639 ^ n23842);
assign n27168 = ~(n26935 ^ n307);
assign n26750 = n11257 | n24121;
assign n10114 = ~(n18422 ^ n26816);
assign n16505 = n8711 | n17318;
assign n8241 = ~n13578;
assign n1353 = ~(n20138 ^ n10372);
assign n13859 = n2279 | n21232;
assign n1841 = ~(n11738 | n24024);
assign n25837 = n18227 & n21828;
assign n6139 = ~n16519;
assign n25399 = n12051 | n13813;
assign n14895 = ~(n26056 | n27151);
assign n20109 = ~n21916;
assign n26018 = ~(n12048 ^ n8210);
assign n14932 = n14618 & n10370;
assign n12358 = ~(n10001 ^ n21222);
assign n25057 = ~(n10400 ^ n15814);
assign n13091 = n1921 & n20309;
assign n5353 = ~(n403 | n509);
assign n695 = n25579 | n13592;
assign n22629 = n20257 & n26517;
assign n3877 = ~n17902;
assign n12171 = ~n4356;
assign n8552 = ~(n19270 | n19702);
assign n14431 = ~n26443;
assign n1123 = n23028 & n6539;
assign n14695 = ~n4409;
assign n22088 = n14530 & n19837;
assign n23993 = n5811 | n13437;
assign n13179 = ~(n13625 ^ n10989);
assign n496 = ~(n12439 ^ n15999);
assign n18676 = ~n2899;
assign n22202 = n22435 & n21479;
assign n16464 = ~n15636;
assign n3548 = n14283 & n12782;
assign n21361 = n26299 | n22535;
assign n98 = n2422 | n1562;
assign n17425 = ~(n16117 | n8891);
assign n25657 = n22209 | n9896;
assign n23264 = ~(n26978 ^ n1961);
assign n26213 = n23660 | n3671;
assign n16954 = ~(n1397 ^ n7783);
assign n22657 = n1275 | n7289;
assign n23436 = ~n6369;
assign n908 = n3388 & n18009;
assign n7726 = ~(n2247 | n19715);
assign n17228 = ~(n22247 ^ n19502);
assign n17990 = n26904 | n17266;
assign n8743 = ~(n19531 | n1999);
assign n18758 = ~(n5000 ^ n18282);
assign n25244 = ~(n20116 ^ n8245);
assign n20777 = ~n19399;
assign n23690 = ~(n23813 ^ n21968);
assign n25932 = n16077 | n21210;
assign n18608 = ~(n899 ^ n3564);
assign n7426 = ~(n1021 ^ n21604);
assign n10402 = n14078 | n4583;
assign n22677 = n26730 & n6823;
assign n2845 = ~(n13206 ^ n7421);
assign n7814 = n16053 | n1807;
assign n16847 = ~(n14680 ^ n16439);
assign n25907 = n8588 & n23404;
assign n13811 = n2973 & n19397;
assign n12041 = ~(n5617 ^ n20734);
assign n4019 = ~(n14254 ^ n11502);
assign n21807 = n1009 | n4999;
assign n5562 = n5401 & n3578;
assign n18827 = n26578 & n3999;
assign n24018 = ~n16482;
assign n9945 = ~n3465;
assign n13959 = ~(n11356 ^ n12587);
assign n1508 = n15429 & n23723;
assign n19448 = n4298 | n16290;
assign n26479 = ~(n20231 ^ n20201);
assign n10773 = ~n11455;
assign n26418 = n22089 | n20139;
assign n5483 = ~n16026;
assign n13716 = n14617 | n9786;
assign n4961 = ~(n2331 ^ n22879);
assign n15629 = ~(n18290 | n9455);
assign n2282 = ~(n25291 ^ n20558);
assign n3300 = ~(n2939 ^ n16960);
assign n4206 = n13910 | n20461;
assign n16915 = ~(n25126 ^ n21226);
assign n10100 = ~(n8694 | n20039);
assign n19563 = n11760 & n3816;
assign n19020 = ~(n18345 ^ n25168);
assign n18738 = n13596 & n10649;
assign n15557 = n1063 & n15394;
assign n14140 = ~n14692;
assign n22916 = n11635 & n13321;
assign n10234 = ~(n25144 ^ n11121);
assign n13431 = n21377 | n13299;
assign n6225 = n5037 | n17955;
assign n21322 = ~n18563;
assign n24675 = n10180 & n2865;
assign n9098 = ~n26972;
assign n3983 = ~(n14824 ^ n21315);
assign n21155 = ~(n14067 ^ n7468);
assign n13384 = ~(n20240 ^ n2845);
assign n355 = n18477 | n2060;
assign n23082 = n9733 | n13216;
assign n24416 = ~(n9223 | n4055);
assign n17246 = n14950 | n260;
assign n20615 = ~n17188;
assign n23023 = n9934 | n20290;
assign n18495 = ~n11537;
assign n26950 = n20062 | n6562;
assign n15107 = n3179 | n12658;
assign n13220 = ~(n3103 ^ n22471);
assign n27026 = n11390 | n7970;
assign n2741 = n22674 & n6378;
assign n21573 = ~(n21352 ^ n19057);
assign n14533 = ~(n18539 ^ n16818);
assign n10776 = n17534 & n19273;
assign n26851 = ~(n9676 ^ n26771);
assign n8258 = ~(n6403 ^ n4722);
assign n1765 = n5607;
assign n7835 = ~(n23005 | n11531);
assign n9020 = ~(n14718 | n8820);
assign n16924 = ~(n15591 ^ n10725);
assign n26064 = ~n16247;
assign n16309 = ~n2436;
assign n12075 = ~(n12333 ^ n18863);
assign n26186 = ~n7652;
assign n2393 = n15667 | n1983;
assign n3941 = n21502 | n5674;
assign n15530 = ~(n22491 | n22600);
assign n5526 = n21802 & n25294;
assign n11021 = n11566 | n10973;
assign n7954 = n19770 | n12022;
assign n4446 = ~(n8407 ^ n13491);
assign n9904 = n11903 & n14872;
assign n8446 = n25616 | n23246;
assign n20770 = ~(n5070 ^ n8734);
assign n26441 = n2012 & n6960;
assign n11493 = ~(n6115 ^ n2352);
assign n19623 = ~(n17376 ^ n7295);
assign n2183 = n21410 | n5862;
assign n20539 = ~(n5579 ^ n26054);
assign n7014 = n19173 | n8483;
assign n9319 = n24094 & n7922;
assign n18058 = ~n15053;
assign n25313 = n22176 | n19298;
assign n13159 = ~n2680;
assign n8085 = ~(n27002 ^ n18502);
assign n10656 = n10556 | n13846;
assign n18934 = ~(n23349 ^ n16759);
assign n14254 = ~n21073;
assign n20066 = n8945 | n16582;
assign n17646 = n22718 & n22957;
assign n17767 = n22719 & n24589;
assign n19257 = n14295 & n2720;
assign n25601 = n13026 | n13369;
assign n703 = ~(n8657 ^ n10593);
assign n737 = ~(n13339 ^ n4623);
assign n18559 = ~n26541;
assign n26212 = ~n22350;
assign n13459 = ~n20036;
assign n4311 = n12960 | n1344;
assign n19571 = ~(n5374 ^ n18649);
assign n17237 = ~(n23874 ^ n23923);
assign n13669 = ~(n24402 ^ n1230);
assign n11086 = ~n21768;
assign n7828 = ~(n12495 ^ n11479);
assign n5625 = ~(n16976 ^ n2880);
assign n25138 = n4887 & n5045;
assign n457 = ~(n23132 ^ n19204);
assign n3611 = ~(n21998 ^ n3945);
assign n17001 = n355 & n27077;
assign n9371 = ~(n16687 ^ n15213);
assign n7022 = n21811 & n2571;
assign n25085 = ~(n14254 | n6964);
assign n4866 = n99 & n1399;
assign n23810 = n26593 & n17374;
assign n20252 = ~(n26705 ^ n22061);
assign n18132 = n18774 | n22784;
assign n24611 = ~(n12454 | n5714);
assign n6967 = ~(n5492 ^ n19947);
assign n26259 = n23843 | n19486;
assign n213 = n2709 | n1093;
assign n25048 = n9248 & n14755;
assign n8164 = ~(n15704 ^ n21308);
assign n15850 = ~(n23533 ^ n9636);
assign n10882 = ~n21324;
assign n306 = ~n11201;
assign n14532 = ~n24042;
assign n24293 = n21987 & n8882;
assign n5480 = ~(n17906 | n24628);
assign n6123 = n15354 & n9721;
assign n3756 = n13172 | n23892;
assign n14817 = n23269 | n15848;
assign n17340 = n10376 & n3615;
assign n24935 = ~(n22528 ^ n20421);
assign n8635 = ~(n7508 ^ n12438);
assign n17590 = ~n4095;
assign n6486 = ~n6555;
assign n6669 = ~(n2910 ^ n19681);
assign n19419 = n2506 & n4465;
assign n641 = n21213 | n15392;
assign n22019 = n15891 | n9319;
assign n11069 = ~n20385;
assign n3994 = n16712 & n3706;
assign n21954 = n8675 | n18559;
assign n22572 = n14415 | n26717;
assign n17617 = ~n25018;
assign n21730 = n5338 | n16752;
assign n5614 = ~(n19312 ^ n24933);
assign n9324 = ~(n26170 ^ n19884);
assign n14034 = n19978 | n21111;
assign n5382 = n22055 | n9184;
assign n1385 = ~(n21949 ^ n24872);
assign n12777 = n8636 | n24591;
assign n6911 = ~(n10042 ^ n2686);
assign n13027 = ~n22321;
assign n22712 = n14060 & n16621;
assign n4281 = n23448 | n7325;
assign n6230 = n2080 & n13919;
assign n18131 = n10720 | n7285;
assign n25719 = ~(n20813 ^ n10423);
assign n25128 = ~(n5090 ^ n21674);
assign n18340 = ~(n21929 | n485);
assign n50 = ~(n16122 ^ n9022);
assign n10556 = n22585 & n23226;
assign n13135 = ~(n14630 ^ n7270);
assign n8693 = n5418 | n23847;
assign n1083 = n20090 & n8811;
assign n3614 = ~(n3205 ^ n24708);
assign n15618 = ~n25688;
assign n21505 = ~(n8959 ^ n3441);
assign n16280 = ~(n11504 ^ n752);
assign n18041 = n18690 | n7685;
assign n23168 = ~n11579;
assign n19915 = n9513 & n23417;
assign n10420 = ~(n4177 ^ n6545);
assign n4560 = ~(n12616 ^ n22879);
assign n3305 = ~(n2113 | n14345);
assign n22994 = ~(n25240 | n6510);
assign n22056 = n9554 | n9509;
assign n13845 = ~(n24600 | n3641);
assign n27164 = ~(n23475 ^ n13419);
assign n23015 = ~(n19940 | n10407);
assign n23158 = n23750 | n14963;
assign n8896 = ~(n23216 ^ n1324);
assign n1164 = ~(n7360 | n16482);
assign n8681 = ~(n14680 ^ n25240);
assign n25440 = n14040 & n8477;
assign n3732 = n6511 | n13738;
assign n10783 = ~(n15892 ^ n8448);
assign n16761 = n23750 | n7678;
assign n7651 = n52 | n23656;
assign n9741 = n21434 & n14301;
assign n23508 = n26474 & n24534;
assign n9042 = ~(n26633 ^ n20048);
assign n4349 = ~(n8713 ^ n21300);
assign n12883 = ~(n17600 ^ n6859);
assign n13834 = ~(n3414 ^ n20923);
assign n4984 = ~(n4446 ^ n24551);
assign n11797 = ~(n5055 ^ n14767);
assign n25479 = n5282 & n13720;
assign n10225 = ~(n2062 | n23191);
assign n25229 = n2015 & n309;
assign n24668 = n14897 | n6014;
assign n10205 = ~(n11302 | n2146);
assign n2654 = n23648 | n3646;
assign n9414 = n12943 & n797;
assign n6293 = ~n23882;
assign n19700 = n25769 & n15776;
assign n186 = ~(n14965 ^ n25465);
assign n25684 = ~(n13224 ^ n15041);
assign n11398 = ~(n15287 ^ n15140);
assign n6496 = n3403 | n3271;
assign n357 = ~(n23896 ^ n15909);
assign n8524 = n10439 & n12139;
assign n26250 = ~(n12331 ^ n23300);
assign n17858 = ~n8724;
assign n22063 = n20730 | n14453;
assign n19304 = ~(n602 | n19971);
assign n14380 = ~(n1489 ^ n19517);
assign n10502 = n6830 | n19773;
assign n25301 = n16009 | n12910;
assign n22521 = n11457 & n10266;
assign n2923 = ~(n14793 ^ n25375);
assign n2691 = n10752 & n21326;
assign n23661 = n1317 & n5202;
assign n26306 = ~(n13241 ^ n13998);
assign n9994 = n13576 | n25165;
assign n36 = n19472 | n8997;
assign n2197 = ~(n15283 ^ n8020);
assign n7516 = ~(n4924 ^ n25230);
assign n1177 = n17088 ^ n18472;
assign n14983 = ~(n21620 ^ n9404);
assign n8485 = ~(n4289 ^ n8178);
assign n23021 = n25674 | n16029;
assign n13436 = ~(n13606 ^ n7091);
assign n26348 = ~(n11356 ^ n2999);
assign n4891 = ~(n6906 ^ n26709);
assign n13779 = n13704 | n5240;
assign n34 = ~(n5796 ^ n25856);
assign n22143 = n9080 | n3609;
assign n26861 = n17531 | n8592;
assign n17957 = ~(n19978 | n24239);
assign n19395 = n19742 | n4867;
assign n6856 = n15529 | n11985;
assign n22663 = n2726 | n23179;
assign n8907 = n10946 | n18881;
assign n23777 = n18750 | n11609;
assign n20837 = ~(n22736 | n17390);
assign n5596 = n22919 | n19074;
assign n12997 = n4130 | n21740;
assign n24953 = ~(n9557 ^ n21832);
assign n18778 = n344 & n26205;
assign n7268 = ~(n1567 ^ n6412);
assign n15376 = ~(n13784 ^ n17959);
assign n4533 = ~(n840 | n7604);
assign n5175 = n3521 | n8323;
assign n2299 = ~(n7827 | n9505);
assign n3772 = n10218 ^ n22612;
assign n6969 = n17697 & n11599;
assign n18853 = ~(n3366 | n23456);
assign n14734 = ~(n7911 ^ n25983);
assign n21614 = n4902 | n928;
assign n16999 = n5611 | n9671;
assign n9854 = ~(n8785 ^ n14841);
assign n4353 = ~n15154;
assign n2103 = ~(n21209 | n25001);
assign n11846 = ~n4864;
assign n3893 = ~(n26046 ^ n21246);
assign n7034 = n1429 | n25555;
assign n8472 = ~n4917;
assign n21448 = ~(n19383 ^ n10422);
assign n6122 = ~n152;
assign n20054 = ~(n4588 ^ n27134);
assign n14693 = n21687 & n6458;
assign n7511 = ~n130;
assign n19242 = n20751 | n19845;
assign n8224 = ~n1138;
assign n18990 = ~(n24996 | n24488);
assign n5072 = ~(n15714 ^ n22364);
assign n926 = ~n12436;
assign n18751 = ~(n22356 ^ n4958);
assign n22287 = n3914 & n1717;
assign n4827 = n4974 | n26985;
assign n4459 = ~(n9156 ^ n9841);
assign n26353 = ~(n6698 ^ n1086);
assign n16624 = n8422 | n7100;
assign n25730 = ~(n21125 ^ n7377);
assign n25223 = ~(n7097 ^ n9469);
assign n24300 = n12923 | n23820;
assign n3372 = n13729 | n21674;
assign n19179 = n19362 & n15690;
assign n20738 = n17799 | n13917;
assign n187 = n24627 | n6374;
assign n21764 = ~n9124;
assign n19945 = n11980 | n9971;
assign n3088 = n21676 | n5135;
assign n23521 = n8835 | n2235;
assign n25419 = ~(n8892 ^ n2313);
assign n23407 = n9013 & n993;
assign n23602 = ~(n11718 ^ n13834);
assign n8537 = n8032 & n1343;
assign n3032 = n12437 | n17465;
assign n7911 = n16160 & n7113;
assign n15436 = n16818 | n13133;
assign n24198 = ~(n7566 ^ n19357);
assign n9617 = n3346 & n19311;
assign n1800 = n734 | n3321;
assign n904 = ~(n13482 ^ n10686);
assign n20944 = ~n19190;
assign n6907 = n5558 & n7481;
assign n1822 = ~(n14826 ^ n13549);
assign n15210 = ~(n8948 ^ n3470);
assign n24641 = n16842 | n23571;
assign n1790 = n9490 & n23693;
assign n13921 = n22892 & n5165;
assign n18611 = ~(n5517 ^ n21981);
assign n5290 = n5386 | n24326;
assign n9141 = ~(n14818 | n10158);
assign n16164 = n9098 | n6908;
assign n22178 = ~(n21867 | n7948);
assign n18294 = ~(n25764 | n17447);
assign n25840 = ~(n16344 ^ n26454);
assign n8361 = ~n19539;
assign n14689 = n18506 & n3994;
assign n25636 = ~(n21162 ^ n8614);
assign n26536 = ~n25748;
assign n20171 = ~(n363 ^ n21732);
assign n15356 = n4140 | n24882;
assign n3271 = ~(n12111 ^ n12668);
assign n24467 = n9628 | n21640;
assign n16149 = ~(n3909 ^ n19081);
assign n15344 = n18995 | n3614;
assign n6685 = ~n13300;
assign n2392 = n14992 | n22764;
assign n19795 = n9977 & n14956;
assign n14402 = ~(n6321 | n20349);
assign n16720 = ~(n22558 | n8155);
assign n10742 = n14978 & n26455;
assign n9954 = ~(n20127 ^ n13650);
assign n905 = n15723;
assign n17964 = n5316 | n7152;
assign n19043 = n23187 | n20833;
assign n23954 = ~(n7909 ^ n18636);
assign n25734 = n14374 | n8652;
assign n4196 = n9134 | n19412;
assign n12012 = ~(n27144 ^ n14692);
assign n22183 = ~(n17250 | n4409);
assign n3912 = n5039 | n8380;
assign n19176 = ~(n13415 ^ n6237);
assign n12756 = ~(n17128 ^ n21441);
assign n25305 = n22225 | n21620;
assign n3981 = n1913;
assign n22974 = ~(n20929 ^ n24620);
assign n25483 = n13865 | n4504;
assign n20790 = ~(n17360 ^ n14684);
assign n995 = n19898 | n17645;
assign n27186 = n20826 & n14532;
assign n18163 = ~(n17224 ^ n8526);
assign n13968 = ~(n13341 ^ n11251);
assign n12714 = ~n19803;
assign n23434 = ~(n719 ^ n25561);
assign n22834 = ~(n10571 | n9431);
assign n18136 = n25715 | n8343;
assign n24758 = ~(n10589 ^ n13698);
assign n12709 = ~n3223;
assign n780 = n10311 | n14713;
assign n21130 = n7730 & n15043;
assign n24037 = n11759 & n26836;
assign n19694 = ~(n23923 ^ n25119);
assign n2224 = n1901 & n12432;
assign n3314 = ~n26104;
assign n2124 = ~(n14078 ^ n18891);
assign n27132 = ~(n23731 ^ n5842);
assign n3903 = ~(n13132 ^ n17253);
assign n9703 = ~n3729;
assign n12029 = ~(n3447 ^ n10669);
assign n17966 = n8739 | n16693;
assign n26415 = n14972 & n5354;
assign n1080 = n26692 & n11015;
assign n10085 = ~(n13518 | n5743);
assign n13456 = ~(n9173 ^ n23148);
assign n21777 = ~n8107;
assign n10972 = n307 | n16046;
assign n20046 = n20965 | n8207;
assign n471 = n24285 | n6180;
assign n25270 = ~n14633;
assign n23737 = ~(n20104 | n15616);
assign n25000 = ~n27164;
assign n16108 = ~(n23216 ^ n15093);
assign n15011 = ~(n14368 ^ n16305);
assign n247 = n22196 | n20900;
assign n18935 = ~(n25494 ^ n6659);
assign n6018 = n15427 | n10168;
assign n15528 = n1013 & n25154;
assign n22432 = ~(n16476 | n15008);
assign n9571 = n23502 | n24567;
assign n18443 = n25857 & n14912;
assign n15232 = ~(n23476 ^ n19783);
assign n23148 = ~(n16559 ^ n6872);
assign n13198 = ~(n10708 ^ n20521);
assign n14909 = ~(n17069 | n16608);
assign n20114 = ~(n617 | n7798);
assign n22357 = n18853 | n3175;
assign n1677 = ~(n26064 | n10930);
assign n10735 = n13690 & n22927;
assign n24856 = n10112 & n21849;
assign n3766 = ~(n268 | n19265);
assign n14926 = ~n6765;
assign n12430 = ~(n2448 ^ n13296);
assign n1297 = n17346 & n13606;
assign n16341 = n26093 | n20138;
assign n10777 = ~(n22788 ^ n8427);
assign n1221 = n5271 & n11478;
assign n12812 = ~(n17686 ^ n4553);
assign n26579 = n26966 | n18063;
assign n21774 = ~n22552;
assign n6498 = n18870 & n12867;
assign n3610 = n12343 & n16357;
assign n8961 = n7014 & n23557;
assign n13568 = ~(n11382 ^ n16637);
assign n18865 = ~(n6167 ^ n13581);
assign n22325 = ~(n24362 ^ n17625);
assign n14857 = ~(n17600 ^ n16054);
assign n16061 = ~(n26553 | n23775);
assign n24419 = ~(n25877 ^ n26443);
assign n26767 = ~(n274 | n2618);
assign n16207 = ~(n14907 ^ n25238);
assign n8915 = n24019 | n24238;
assign n5114 = n16661 & n25859;
assign n14915 = n15249 | n19550;
assign n13025 = n10594 & n9355;
assign n23443 = ~n532;
assign n1444 = ~(n10529 ^ n22498);
assign n7867 = ~(n2849 ^ n20641);
assign n13688 = n22809 | n584;
assign n1910 = n18803 & n5327;
assign n3400 = ~(n12877 ^ n6094);
assign n25775 = ~(n11554 | n20734);
assign n1154 = ~(n21997 | n26962);
assign n1306 = n1804 | n15390;
assign n9366 = ~n24896;
assign n26857 = ~(n1445 ^ n18260);
assign n18666 = ~(n26452 | n3783);
assign n3666 = ~(n18934 | n9820);
assign n757 = ~(n10824 ^ n13761);
assign n18053 = n20530 | n4822;
assign n26841 = n21613 | n16807;
assign n25059 = n24638 | n26645;
assign n21976 = ~(n11333 ^ n11648);
assign n5563 = n16059 | n12737;
assign n3053 = ~n9972;
assign n19548 = n23590 | n20184;
assign n867 = ~n25365;
assign n13906 = ~(n26955 ^ n3478);
assign n3779 = ~n4404;
assign n26980 = ~(n252 | n20316);
assign n13663 = n11492 & n1347;
assign n19748 = n8108 & n24931;
assign n25016 = ~(n10514 ^ n4514);
assign n15668 = n10023 | n7216;
assign n22773 = ~n23268;
assign n1277 = ~(n16117 ^ n9832);
assign n6632 = ~n10022;
assign n23880 = n8227 & n11947;
assign n22026 = ~(n3382 ^ n18363);
assign n14634 = ~n11653;
assign n2265 = ~(n19222 ^ n1786);
assign n4652 = ~(n15912 ^ n19896);
assign n12947 = n6549 | n13108;
assign n19490 = n2404 | n9931;
assign n4412 = ~(n22095 | n713);
assign n23096 = ~n7505;
assign n27161 = n10118 & n2544;
assign n12445 = ~(n9137 ^ n5513);
assign n5099 = n18294 | n26383;
assign n12645 = n270 & n5198;
assign n1220 = n19074 | n6504;
assign n9266 = ~(n178 ^ n2042);
assign n10597 = n22091 & n18861;
assign n13687 = n18370 | n11289;
assign n17085 = n22529 & n179;
assign n26480 = n1437 | n17784;
assign n19165 = n1742 | n1798;
assign n14678 = n4511 & n19573;
assign n23234 = ~n11486;
assign n2561 = ~(n15044 ^ n6730);
assign n21062 = ~(n18923 ^ n22416);
assign n19487 = n16044 & n10772;
assign n24865 = n23211 | n14569;
assign n24078 = n20293 & n22006;
assign n21198 = ~(n3480 ^ n3136);
assign n2316 = ~(n26089 ^ n389);
assign n16893 = n4119 & n24746;
assign n16288 = n14879 | n16181;
assign n10602 = ~n16924;
assign n1721 = ~(n12542 ^ n25525);
assign n12863 = ~(n26312 | n23895);
assign n6246 = ~(n2865 ^ n21989);
assign n13310 = ~(n2705 ^ n18926);
assign n11790 = ~(n22110 | n25485);
assign n4806 = n2331 | n5506;
assign n12154 = n12343 | n16357;
assign n23704 = ~n11285;
assign n20851 = n27176 & n25633;
assign n7563 = n8680 & n7676;
assign n11823 = n14262 & n20884;
assign n24453 = ~(n13114 | n16283);
assign n10778 = n23479 | n1383;
assign n22310 = n3506 | n10658;
assign n1797 = ~(n6518 | n6410);
assign n18662 = ~n21287;
assign n26365 = n10164 | n21703;
assign n903 = n11156 & n595;
assign n13565 = ~(n5760 ^ n1754);
assign n5288 = ~(n13970 ^ n5805);
assign n7424 = ~(n11467 | n26015);
assign n16963 = ~(n3358 ^ n7108);
assign n10176 = n21546 & n24548;
assign n13521 = n17616 & n9966;
assign n25290 = n23163 | n10176;
assign n3068 = n16294 | n1380;
assign n16053 = ~(n3980 ^ n1716);
assign n8374 = n8673 & n26623;
assign n26727 = ~(n4789 ^ n14300);
assign n16130 = ~n25241;
assign n13209 = ~(n5861 ^ n10347);
assign n5756 = n7201 & n14403;
assign n23539 = ~n5905;
assign n2631 = n6422 | n24217;
assign n4344 = n23707 | n3730;
assign n5945 = n8322 | n19634;
assign n18284 = n4717 | n15813;
assign n9878 = n18060 | n19738;
assign n26043 = ~(n19951 | n20655);
assign n22791 = ~(n18926 | n6513);
assign n24259 = ~(n5313 ^ n24009);
assign n26602 = ~(n42 ^ n24648);
assign n3690 = ~n8507;
assign n24757 = n23521 & n21347;
assign n21280 = ~n24873;
assign n8512 = n5389 | n17313;
assign n5020 = ~(n2242 ^ n6225);
assign n22301 = n14251 | n10349;
assign n6450 = ~(n15659 ^ n18537);
assign n7892 = ~n22002;
assign n20177 = n3249 | n10936;
assign n22603 = n12429 & n15029;
assign n20901 = ~(n15468 ^ n4228);
assign n21459 = ~(n9098 ^ n25881);
assign n8855 = ~(n21392 ^ n18105);
assign n24996 = ~n3906;
assign n4555 = ~n22470;
assign n10459 = n14232 & n11264;
assign n6888 = ~(n5122 ^ n13821);
assign n24585 = ~(n13643 ^ n3038);
assign n11200 = n9986 | n3112;
assign n11537 = ~(n22429 ^ n6142);
assign n17275 = n9198 | n37;
assign n10554 = ~(n21110 ^ n3270);
assign n10601 = n25452 & n507;
assign n12944 = ~n2446;
assign n13862 = n8061 & n10972;
assign n24767 = ~(n24907 ^ n24485);
assign n26116 = ~(n20592 | n16833);
assign n12842 = ~(n926 ^ n21125);
assign n9092 = n26247 | n18135;
assign n19692 = n2172 & n17315;
assign n12809 = ~(n6003 ^ n21547);
assign n11294 = ~n12892;
assign n25819 = ~(n19630 | n16642);
assign n712 = n12919 & n3434;
assign n2759 = n7952 & n1365;
assign n23644 = ~n26851;
assign n16296 = ~(n25879 | n6295);
assign n20339 = ~(n5402 ^ n7361);
assign n13023 = ~n12209;
assign n25289 = ~(n25921 ^ n21753);
assign n9799 = n16775 & n22214;
assign n11189 = ~(n12950 | n949);
assign n17268 = n18994 | n2100;
assign n12275 = ~(n8097 ^ n17210);
assign n485 = ~(n12824 ^ n16342);
assign n1867 = n112 | n26264;
assign n24605 = n11011 & n16711;
assign n18463 = ~(n23849 ^ n2289);
assign n5798 = n5315 & n20387;
assign n21598 = ~(n16092 | n24536);
assign n15572 = ~n7191;
assign n529 = n3398 & n164;
assign n20505 = ~(n11042 ^ n24569);
assign n4940 = ~n8259;
assign n9766 = n13719 & n22342;
assign n7263 = n17872 | n9881;
assign n21844 = ~(n11881 | n10225);
assign n5635 = n23244 | n1801;
assign n20528 = n1200 | n15254;
assign n9838 = ~(n15568 ^ n5928);
assign n10965 = ~(n15784 ^ n25797);
assign n13480 = ~n21839;
assign n26937 = ~(n11734 ^ n22687);
assign n14747 = ~(n21780 | n816);
assign n15948 = n21292 | n654;
assign n9607 = n18714 | n24745;
assign n10367 = ~(n24244 ^ n11577);
assign n16419 = ~(n22233 ^ n13825);
assign n2968 = ~(n9700 ^ n9969);
assign n4483 = n9897 | n26711;
assign n1439 = n13400 & n18283;
assign n3339 = n23797 | n257;
assign n10942 = n21589 & n24075;
assign n15276 = ~n22805;
assign n8838 = ~n9368;
assign n10047 = ~(n19726 | n25583);
assign n5150 = n10200 & n22777;
assign n9477 = ~n24109;
assign n440 = ~(n23290 ^ n20002);
assign n8397 = n16939 | n968;
assign n19541 = ~n2113;
assign n17325 = ~(n19097 ^ n5333);
assign n26884 = ~(n24465 ^ n23647);
assign n3748 = ~(n14532 ^ n20826);
assign n23621 = n25318 | n21728;
assign n18768 = ~n5428;
assign n16 = ~(n851 ^ n17047);
assign n5280 = ~(n14033 | n22797);
assign n17517 = ~n15991;
assign n26427 = ~(n18649 ^ n3795);
assign n15075 = n16387 | n507;
assign n26715 = n3257 | n25243;
assign n18076 = n7344 | n26147;
assign n24447 = ~(n10614 ^ n21898);
assign n24688 = n4663 & n19390;
assign n24262 = n23440 & n25197;
assign n15951 = n22038 | n17548;
assign n5159 = n25946 & n18867;
assign n25157 = n24660 | n2787;
assign n19585 = ~(n14311 ^ n19895);
assign n25186 = n25508 & n10052;
assign n22769 = n26162 & n23556;
assign n14794 = ~n4959;
assign n9012 = ~(n25292 ^ n8765);
assign n14147 = ~(n19492 ^ n7145);
assign n8718 = ~(n21875 ^ n20610);
assign n18256 = ~n2518;
assign n1865 = ~(n2732 ^ n1432);
assign n6572 = n2003 | n6063;
assign n10988 = n3953 & n13996;
assign n26627 = n24537 | n11210;
assign n3222 = ~(n10534 ^ n9366);
assign n21111 = ~(n4945 ^ n8482);
assign n1331 = n11122 | n10849;
assign n18455 = ~(n24237 ^ n4017);
assign n20667 = ~n6356;
assign n8866 = n17558 | n1855;
assign n22245 = n14383 | n2107;
assign n5486 = n12543 | n5220;
assign n24102 = ~(n21672 ^ n19300);
assign n9943 = ~(n17447 ^ n25764);
assign n11884 = ~(n11056 | n18157);
assign n21063 = ~(n22626 | n26986);
assign n17442 = ~n3420;
assign n16698 = ~(n20700 | n932);
assign n13166 = ~(n26400 ^ n5453);
assign n20276 = n18483 | n16314;
assign n24292 = ~(n10925 ^ n22538);
assign n23297 = n15627 & n15896;
assign n9351 = ~(n9711 | n10980);
assign n25354 = n63 | n25240;
assign n13854 = n10282 & n4444;
assign n23845 = n1152 & n10917;
assign n6803 = n12160 & n10562;
assign n5759 = n9433 | n11858;
assign n16185 = ~(n17818 ^ n20144);
assign n24923 = ~n22704;
assign n21409 = ~(n1558 ^ n11566);
assign n6809 = ~n12070;
assign n4205 = ~(n5245 ^ n2326);
assign n19175 = n4721 & n13930;
assign n6759 = ~(n26834 | n5709);
assign n3767 = n7081 & n24213;
assign n10794 = ~(n21779 | n24392);
assign n17060 = n18629 & n19964;
assign n16668 = ~(n25324 | n14148);
assign n943 = n1896 | n4542;
assign n8204 = n6753 | n3220;
assign n10688 = n6778 | n21214;
assign n12683 = ~(n3591 ^ n3963);
assign n23623 = ~(n25389 | n13339);
assign n19496 = ~(n3497 ^ n3207);
assign n24352 = n16195 | n1853;
assign n7478 = ~(n26942 ^ n22634);
assign n17788 = n8634 & n893;
assign n25230 = ~(n7242 ^ n25277);
assign n17255 = ~(n17624 ^ n12632);
assign n9724 = n9880 | n1152;
assign n11613 = ~(n25724 ^ n24503);
assign n10962 = ~n20927;
assign n17189 = ~n4362;
assign n23470 = n15695 | n583;
assign n6932 = ~(n6154 | n21097);
assign n3522 = n9035 | n9494;
assign n1524 = ~(n6940 | n868);
assign n23460 = ~(n19993 ^ n10511);
assign n11849 = ~(n27203 ^ n1550);
assign n18678 = n14965 | n10389;
assign n15484 = n17175 & n3558;
assign n14554 = ~(n6161 | n21793);
assign n8413 = ~(n16600 | n11614);
assign n3593 = ~(n12149 ^ n7447);
assign n15776 = n26814 | n934;
assign n2918 = ~(n20275 ^ n26986);
assign n1826 = ~(n25558 | n21);
assign n21500 = n24733 | n2806;
assign n4660 = ~(n22096 ^ n20850);
assign n5297 = ~(n27142 | n2410);
assign n6681 = n21169 & n10717;
assign n979 = ~(n6841 | n13935);
assign n20905 = ~(n17287 | n21287);
assign n25777 = n10507 & n26205;
assign n3367 = n2812 | n17645;
assign n9970 = n14816 | n18318;
assign n6287 = ~(n19097 ^ n7949);
assign n20787 = ~(n16889 | n18105);
assign n26203 = n17358 | n7994;
assign n16368 = ~(n20542 ^ n25937);
assign n8351 = ~n12637;
assign n8396 = ~(n18925 | n25150);
assign n24217 = ~n16091;
assign n9908 = ~n17302;
assign n13764 = ~(n20204 ^ n14905);
assign n1772 = n24621 & n7196;
assign n22604 = n14044 & n91;
assign n8506 = n26428 | n1085;
assign n21246 = ~n23900;
assign n7654 = n21887 & n12061;
assign n11156 = n22865 | n12;
assign n1087 = n5331 | n24960;
assign n12049 = ~n13447;
assign n26267 = ~(n21416 | n4773);
assign n10319 = n12880 & n16229;
assign n17328 = ~(n12396 | n24937);
assign n1133 = n11624 | n14299;
assign n27004 = ~(n25493 ^ n7372);
assign n4936 = ~(n23697 ^ n19531);
assign n18635 = ~(n18380 ^ n22806);
assign n10680 = ~(n20811 ^ n19047);
assign n17125 = ~(n15365 | n1973);
assign n21725 = n6134 | n1707;
assign n5277 = n6385 & n23030;
assign n18011 = ~(n8398 ^ n710);
assign n5272 = n1406 | n19473;
assign n1175 = n5934 | n983;
assign n1953 = n7297 & n24102;
assign n7915 = ~n20957;
assign n24051 = ~(n10855 ^ n671);
assign n22700 = ~n2005;
assign n7119 = ~(n587 ^ n22452);
assign n16742 = n3393 & n1465;
assign n19008 = n17096 & n22950;
assign n17291 = ~(n5756 ^ n7467);
assign n9270 = ~(n20527 ^ n5880);
assign n7966 = ~n6127;
assign n13474 = ~n21759;
assign n23142 = ~(n7857 ^ n5060);
assign n8912 = n8630 | n18696;
assign n253 = ~(n24948 ^ n11322);
assign n25450 = ~(n10001 | n21263);
assign n21496 = ~(n16278 ^ n8259);
assign n21512 = ~(n16755 | n23493);
assign n4371 = ~n7191;
assign n25072 = n4748 | n21029;
assign n3399 = n23088 | n4668;
assign n24044 = ~n10763;
assign n20095 = n20205 | n4256;
assign n17321 = n1374 & n22728;
assign n2151 = ~n6686;
assign n22196 = ~(n13907 | n12493);
assign n3838 = n8552 | n17167;
assign n5853 = ~(n19360 ^ n19042);
assign n9233 = ~n19711;
assign n23309 = ~(n25877 ^ n22619);
assign n16649 = n14133 | n9570;
assign n8556 = n5605 | n23587;
assign n20631 = n15976 & n8093;
assign n26310 = n24359 | n19319;
assign n14376 = n5464 & n14065;
assign n13340 = ~(n11802 | n11502);
assign n20804 = ~(n2656 ^ n6851);
assign n18781 = ~n25906;
assign n16444 = ~(n1594 | n762);
assign n11484 = n17271 & n7159;
assign n25960 = n18012 | n10776;
assign n24431 = ~(n13020 ^ n19114);
assign n6813 = n11155 & n972;
assign n10895 = ~(n10625 ^ n11481);
assign n25599 = n26750 & n19538;
assign n13349 = ~n4319;
assign n7597 = ~n4872;
assign n25026 = n5097 & n3394;
assign n14605 = n21520 | n7536;
assign n17022 = ~n24315;
assign n25086 = ~(n21636 ^ n26107);
assign n6399 = n1977 & n5878;
assign n9668 = ~n25881;
assign n20798 = n11473 | n27;
assign n7653 = ~n18194;
assign n3458 = n14189 & n14795;
assign n3697 = ~(n8100 ^ n22211);
assign n13265 = n10627 & n18913;
assign n22025 = n18420 | n16532;
assign n9723 = ~n20557;
assign n7578 = ~n8657;
assign n26005 = n8579 | n27206;
assign n10174 = ~(n767 ^ n22793);
assign n6260 = n7066 | n9413;
assign n11935 = ~(n17409 ^ n10258);
assign n25729 = n7320 & n25560;
assign n15268 = ~(n3706 ^ n15539);
assign n25130 = ~(n8391 ^ n7917);
assign n4610 = n18325 & n14219;
assign n10561 = ~(n21689 ^ n16175);
assign n22552 = ~(n20999 ^ n24029);
assign n5206 = ~(n17060 ^ n26206);
assign n23956 = ~n25937;
assign n26634 = ~(n17222 ^ n2598);
assign n2073 = ~(n18821 ^ n9975);
assign n13623 = n13000 | n13997;
assign n16079 = n23800 & n1308;
assign n6642 = n11673 & n11948;
assign n3451 = ~(n8901 ^ n409);
assign n13240 = n24038 & n5894;
assign n15679 = ~(n1541 ^ n7524);
assign n6368 = n23529 | n10739;
assign n18575 = ~n9160;
assign n12561 = n2156 & n7402;
assign n370 = n20662 | n16533;
assign n23703 = n21420 | n21768;
assign n8648 = ~n12492;
assign n15233 = n5816 | n13981;
assign n20544 = ~n19042;
assign n15683 = ~(n6510 ^ n5031);
assign n20350 = n20474 | n19871;
assign n20363 = n26127 | n648;
assign n16271 = n14068 & n17335;
assign n22111 = n26197 | n19003;
assign n22276 = n20121 | n18235;
assign n10432 = ~(n16750 ^ n16981);
assign n13493 = ~(n8780 ^ n16479);
assign n20487 = n3297 | n13143;
assign n13036 = ~(n4388 ^ n23131);
assign n6519 = n4430 | n16666;
assign n26982 = ~(n15875 | n13352);
assign n7975 = ~(n26095 ^ n24461);
assign n2014 = n18777 & n8815;
assign n5399 = ~(n15686 ^ n5771);
assign n15225 = ~(n14487 ^ n4330);
assign n1925 = ~(n4755 ^ n25802);
assign n17881 = ~n3319;
assign n153 = n1437 & n12488;
assign n17697 = n7644 | n11235;
assign n45 = ~(n16476 | n19146);
assign n16851 = ~(n18537 ^ n4376);
assign n2764 = ~(n14686 ^ n2433);
assign n3438 = ~(n4967 | n26541);
assign n23584 = n23950 | n23002;
assign n20181 = ~n7083;
assign n25391 = n20338 | n13034;
assign n19489 = ~n3173;
assign n24716 = n2355 & n115;
assign n19661 = n1188 | n22427;
assign n15265 = ~n25073;
assign n7379 = n12490 & n19824;
assign n26228 = ~(n12991 ^ n24700);
assign n9355 = n14481 | n17145;
assign n11909 = n14936 & n15233;
assign n22544 = n4784 & n2603;
assign n15492 = n5869 & n19492;
assign n16678 = ~(n3138 | n2829);
assign n19552 = ~(n24420 ^ n12398);
assign n20331 = ~(n25289 ^ n5255);
assign n18482 = ~(n19416 ^ n14983);
assign n24421 = ~(n5045 ^ n7781);
assign n2061 = ~(n1710 ^ n23284);
assign n3302 = ~(n3266 | n3028);
assign n323 = ~(n26880 ^ n1693);
assign n17715 = ~(n5244 ^ n14852);
assign n3056 = ~(n18484 ^ n23855);
assign n15563 = n1329 | n1152;
assign n2096 = ~n14011;
assign n23564 = n22823 & n19213;
assign n24465 = ~(n26577 ^ n1074);
assign n14910 = n17728 & n18319;
assign n14272 = n12507 & n15739;
assign n14026 = n6753 | n3376;
assign n16736 = n26435 & n14903;
assign n4993 = n2429 | n15961;
assign n16124 = n4097 | n8527;
assign n12086 = ~(n5830 ^ n17288);
assign n20167 = n20993 | n22648;
assign n18643 = ~n19303;
assign n12143 = ~n19842;
assign n2457 = ~(n24327 ^ n4325);
assign n16840 = ~(n15443 ^ n15397);
assign n20517 = ~(n14871 ^ n23613);
assign n25526 = ~(n421 | n15272);
assign n20028 = n12735 | n11986;
assign n12749 = ~(n18915 ^ n6662);
assign n19688 = ~(n23645 | n22068);
assign n14039 = n23056 | n10371;
assign n4471 = n21517 & n8582;
assign n21084 = n23518 & n12830;
assign n10197 = n23213 | n4883;
assign n14100 = ~(n25268 | n20883);
assign n14236 = ~(n2886 ^ n1738);
assign n19252 = ~(n13263 ^ n21779);
assign n24092 = ~(n7500 ^ n19266);
assign n8841 = n11592 & n14003;
assign n7801 = n22170 | n4007;
assign n9931 = n12915 & n13012;
assign n20587 = n21100 | n17445;
assign n20083 = ~(n2473 | n20203);
assign n1404 = ~n22588;
assign n4864 = n279 & n9891;
assign n15623 = ~(n23849 | n2289);
assign n15664 = n12328 | n20663;
assign n25358 = ~(n15008 ^ n16476);
assign n3463 = ~(n11733 ^ n26789);
assign n20575 = ~(n2781 ^ n18102);
assign n1884 = ~(n18617 ^ n18452);
assign n689 = n10471 | n8600;
assign n13815 = n4040 | n16009;
assign n6049 = n15410 & n20969;
assign n6701 = ~n12900;
assign n786 = ~(n8419 | n17067);
assign n7752 = ~(n7150 ^ n2229);
assign n20372 = n6659 | n12991;
assign n3112 = ~n17412;
assign n26796 = ~(n5194 ^ n16743);
assign n7936 = n1882 | n12311;
assign n18677 = ~(n12112 | n9404);
assign n16293 = ~(n12426 | n11476);
assign n16355 = ~(n24620 | n7099);
assign n4911 = n14141 & n4827;
assign n20118 = ~(n9770 ^ n19143);
assign n1660 = ~(n27120 ^ n23065);
assign n14614 = ~n13303;
assign n16407 = ~(n20312 ^ n12352);
assign n10676 = n22830 | n7171;
assign n17870 = ~(n17135 ^ n16441);
assign n9401 = ~n7421;
assign n12574 = n20977 & n18076;
assign n25693 = ~(n96 ^ n8249);
assign n2271 = n20793 & n24528;
assign n12886 = ~(n9493 ^ n3918);
assign n14626 = n5253 | n20146;
assign n25304 = n21166 & n10811;
assign n4589 = n17711 | n8398;
assign n18960 = ~(n11542 | n18247);
assign n14617 = n7172 & n19806;
assign n7002 = ~(n16863 ^ n24816);
assign n2222 = n8739 & n23655;
assign n13468 = ~(n21464 ^ n14092);
assign n24186 = n2641 & n16036;
assign n13239 = ~(n7892 | n2718);
assign n22758 = n11116 | n7825;
assign n16015 = ~(n19472 | n24473);
assign n3062 = ~(n17111 ^ n6829);
assign n25678 = n7907 | n6455;
assign n5465 = ~n17299;
assign n17270 = n20216 | n3524;
assign n19145 = n23159 | n9161;
assign n9603 = ~n20595;
assign n13450 = ~(n11220 ^ n3425);
assign n7366 = ~(n2656 ^ n16929);
assign n1334 = ~n21398;
assign n6259 = n15060 & n10754;
assign n118 = n5298 | n2359;
assign n26655 = n1957 | n5197;
assign n20136 = n17945 | n5787;
assign n12592 = ~n1545;
assign n24132 = n8651 & n178;
assign n13461 = ~(n19061 | n9935);
assign n23342 = n1923 | n17129;
assign n13532 = n26988 | n21542;
assign n4401 = ~(n13678 ^ n1854);
assign n2767 = n21243 & n12331;
assign n7743 = ~n18274;
assign n8051 = n8361 | n1483;
assign n24145 = ~(n18267 ^ n17765);
assign n12460 = n25589 | n16831;
assign n17909 = ~n21674;
assign n18079 = ~n14809;
assign n14233 = n20733 | n7330;
assign n911 = ~(n839 ^ n6139);
assign n12140 = ~(n10683 | n23832);
assign n625 = n20370 & n3401;
assign n23711 = ~(n11184 | n19366);
assign n22264 = n24179 & n7998;
assign n550 = ~n9397;
assign n15906 = ~n24628;
assign n17025 = n2250 | n4324;
assign n27083 = n10552 | n2879;
assign n9176 = n9513 | n23417;
assign n18830 = ~(n8060 ^ n1695);
assign n4640 = ~(n10024 ^ n7347);
assign n14841 = ~(n6963 ^ n25974);
assign n10899 = ~(n6241 ^ n17462);
assign n21174 = ~(n8381 | n12889);
assign n24510 = ~n7765;
assign n2640 = ~(n19667 | n4272);
assign n22456 = ~(n20283 ^ n6939);
assign n18270 = n22855 | n26410;
assign n8033 = ~(n4930 ^ n21134);
assign n13746 = n13890 | n12336;
assign n7579 = ~(n7689 ^ n25115);
assign n1290 = n11321 | n3746;
assign n11628 = n14662 & n13187;
assign n5487 = n5842 | n13429;
assign n25754 = n11685 | n3890;
assign n24241 = n13378 | n13459;
assign n12471 = n25094 & n3049;
assign n10634 = ~n13905;
assign n2476 = n17351 & n21850;
assign n841 = n5431 | n13469;
assign n13831 = ~n23558;
assign n5899 = n14230 & n19922;
assign n973 = ~(n280 ^ n13875);
assign n1655 = ~n26011;
assign n19470 = n22166 | n23607;
assign n13232 = n18378 | n16504;
assign n23835 = ~(n19198 ^ n22684);
assign n10684 = ~n18322;
assign n2867 = n22164 & n19188;
assign n10655 = ~(n5266 | n11428);
assign n7238 = ~(n5001 ^ n7693);
assign n2897 = ~(n18360 ^ n11644);
assign n20170 = n23486 & n16663;
assign n21343 = n14337 | n4940;
assign n18913 = n20242 | n12724;
assign n11250 = n22656 | n3328;
assign n21388 = n21380 | n5211;
assign n13076 = n4376 | n19080;
assign n22982 = n5060 | n15380;
assign n10170 = n3709 | n8969;
assign n21359 = n22841 & n9935;
assign n16610 = n23910 | n21339;
assign n11107 = n20323 | n8564;
assign n1454 = ~(n48 | n8714);
assign n108 = ~(n17009 ^ n11376);
assign n22354 = n1826 | n22505;
assign n17227 = ~(n9125 ^ n10631);
assign n16141 = n21015 | n11452;
assign n16433 = ~(n16732 ^ n13056);
assign n4992 = n6379 | n10923;
assign n2998 = n1311 & n24270;
assign n10559 = n11425 | n19531;
assign n5714 = ~n2816;
assign n23902 = n16320 | n3304;
assign n16248 = n19850 | n24443;
assign n11942 = n13752 | n20304;
assign n7753 = ~(n6385 ^ n16223);
assign n22169 = n7725;
assign n4973 = n23075 | n18566;
assign n13801 = ~(n9476 ^ n21924);
assign n4369 = n16232 | n4509;
assign n22851 = ~n13677;
assign n5397 = n10403 | n21668;
assign n7825 = ~(n17520 ^ n5058);
assign n16348 = n18161 & n23205;
assign n11041 = n16211 | n7437;
assign n6780 = ~(n4780 | n21922);
assign n10208 = n13516 & n17761;
assign n13901 = ~(n7893 | n5400);
assign n9639 = n2160 | n27095;
assign n9730 = ~(n24705 ^ n21460);
assign n14365 = ~n8717;
assign n5257 = n23008 | n17640;
assign n26403 = n5655 & n26655;
assign n25763 = ~(n19868 | n19742);
assign n2482 = ~n16359;
assign n1139 = ~(n19328 | n16123);
assign n467 = n1847 | n18240;
assign n3291 = ~(n13696 ^ n7470);
assign n6004 = n11758 | n12457;
assign n17677 = ~n336;
assign n21231 = ~(n7775 ^ n6848);
assign n12512 = ~n14352;
assign n7195 = ~n1255;
assign n26432 = n1180 | n1206;
assign n18222 = n11870 | n184;
assign n14498 = ~n19475;
assign n510 = ~(n4326 ^ n3952);
assign n23017 = n1965 | n6220;
assign n7862 = n18403 & n18956;
assign n2135 = ~n20343;
assign n10902 = n12792 & n2064;
assign n6144 = n20913 | n5150;
assign n8238 = ~(n4769 | n11176);
assign n3629 = n12396 | n8297;
assign n1499 = ~(n15502 ^ n8553);
assign n17768 = ~(n9402 | n23209);
assign n13870 = n8678 & n3882;
assign n18261 = ~n25694;
assign n17576 = ~(n7057 ^ n12956);
assign n8158 = n19313 | n13354;
assign n10387 = ~(n25172 | n16545);
assign n18016 = ~n6475;
assign n5730 = n9187 | n4870;
assign n22283 = ~(n11616 ^ n18534);
assign n15010 = ~n6410;
assign n1459 = n21984 | n6255;
assign n14425 = n9588 | n14505;
assign n26771 = ~(n27089 ^ n12657);
assign n3521 = n26443 & n10017;
assign n16792 = ~n24543;
assign n26024 = ~(n14411 ^ n18243);
assign n22516 = n25556 | n7938;
assign n25055 = n15534 | n23885;
assign n6983 = ~(n22604 ^ n17589);
assign n15008 = ~n25805;
assign n13426 = ~(n25538 ^ n7305);
assign n24615 = ~n4590;
assign n12213 = n21766 | n9480;
assign n16352 = n24760 | n26721;
assign n14844 = n16894 & n25803;
assign n25498 = ~(n9365 ^ n23541);
assign n27118 = ~(n7854 ^ n6903);
assign n22036 = ~n7552;
assign n24144 = ~(n2815 ^ n10455);
assign n15680 = n3169 | n8622;
assign n17113 = n7109 | n19536;
assign n23386 = ~(n11045 | n19282);
assign n2009 = n2662 & n22969;
assign n3481 = n752 | n11504;
assign n2986 = ~(n23160 | n3570);
assign n3796 = ~(n3178 | n10614);
assign n2882 = n15551 & n25678;
assign n1547 = ~n13393;
assign n16199 = ~(n7430 ^ n11996);
assign n9241 = ~n25768;
assign n24643 = ~(n15047 ^ n8286);
assign n14741 = n10318 | n18752;
assign n9745 = n15096 | n10143;
assign n15180 = ~(n8755 ^ n26406);
assign n5354 = ~(n27137 ^ n26800);
assign n19899 = ~(n6934 ^ n14622);
assign n10415 = n17503 & n15833;
assign n23525 = ~n685;
assign n9744 = n5355 & n19962;
assign n3412 = n10083 | n18928;
assign n2450 = n9495 & n10073;
assign n20119 = n21424 & n1318;
assign n17122 = ~n25603;
assign n23078 = n10088 | n21185;
assign n11742 = n11394 | n5419;
assign n9514 = ~n7285;
assign n12205 = ~(n18027 ^ n19137);
assign n15721 = ~(n14958 ^ n17888);
assign n3848 = ~n2279;
assign n26371 = ~(n6666 ^ n10355);
assign n8741 = ~(n17323 | n5555);
assign n12242 = ~(n20000 | n20665);
assign n2263 = n24366 | n24695;
assign n11074 = n11630 | n18504;
assign n22511 = ~(n25035 ^ n10297);
assign n11462 = ~(n20537 ^ n21044);
assign n25817 = n13036 | n23307;
assign n24814 = n6649 & n17570;
assign n4816 = ~(n18895 ^ n26318);
assign n3923 = n15175 | n11098;
assign n1241 = n6653 | n15569;
assign n19367 = ~(n7687 ^ n23123);
assign n20477 = ~(n13193 ^ n5866);
assign n14386 = ~(n9385 ^ n25131);
assign n13937 = n14390 | n21684;
assign n15432 = n8068 & n1128;
assign n9126 = ~(n3625 ^ n13089);
assign n4515 = n17579 | n3320;
assign n4142 = n26915 | n8549;
assign n9105 = n613 | n8961;
assign n26336 = n4241 | n11160;
assign n12369 = n20998 | n2576;
assign n14502 = ~(n23144 | n8439);
assign n23222 = ~(n26495 ^ n23620);
assign n4062 = n744 & n18630;
assign n12166 = n5768 | n24988;
assign n7540 = n2974 & n16031;
assign n21675 = ~(n26797 ^ n24196);
assign n18546 = n20429 & n22909;
assign n2693 = ~(n3510 ^ n464);
assign n2333 = n13619 & n11886;
assign n13753 = ~(n24851 ^ n9251);
assign n2270 = n22566 | n19317;
assign n6363 = n26911 & n16566;
assign n2965 = ~(n5970 ^ n12570);
assign n12367 = ~(n2873 ^ n17813);
assign n16417 = ~(n18326 | n1230);
assign n21544 = ~(n15233 ^ n11920);
assign n8216 = n20599 | n2562;
assign n10211 = ~(n1293 | n25413);
assign n25002 = n20119 | n3168;
assign n11616 = n19704 | n6469;
assign n24342 = ~(n1556 ^ n15835);
assign n7265 = n24114 | n22067;
assign n22582 = n16624 & n9408;
assign n10370 = n27136 | n26270;
assign n26338 = n18818 | n24874;
assign n12190 = ~n7289;
assign n10333 = ~n5582;
assign n24200 = ~(n5038 ^ n20483);
assign n1577 = ~n13895;
assign n9563 = n9908 | n19843;
assign n85 = ~(n14465 | n15426);
assign n14304 = ~(n22626 ^ n8856);
assign n2798 = n9469 & n3237;
assign n9422 = ~(n25119 ^ n23529);
assign n4222 = n11501 & n22852;
assign n6566 = ~n26857;
assign n10734 = ~n2893;
assign n19802 = ~(n19331 ^ n23910);
assign n15666 = ~(n468 ^ n1255);
assign n14842 = n2514 | n26883;
assign n1592 = n21371 & n18106;
assign n17007 = n512 | n11571;
assign n16229 = ~n18446;
assign n14591 = n4823 & n10939;
assign n9369 = n22204 | n13589;
assign n10724 = n19970 | n3106;
assign n25014 = ~n1481;
assign n9562 = n8576 | n26243;
assign n12343 = ~n9140;
assign n4014 = ~(n14592 ^ n15278);
assign n22710 = ~(n2658 | n23172);
assign n9425 = n7184 & n20564;
assign n15203 = n14426 & n25159;
assign n9043 = ~(n23005 ^ n11531);
assign n17478 = ~(n23271 ^ n7670);
assign n27059 = n21386 | n23697;
assign n20000 = n6353 & n12391;
assign n2405 = n21156 & n24124;
assign n718 = ~(n8032 | n12161);
assign n14881 = ~n6679;
assign n14216 = ~(n15932 ^ n16163);
assign n26813 = ~(n20588 | n16131);
assign n26906 = n18954 | n23600;
assign n19662 = n26180 & n24700;
assign n6362 = ~(n7243 ^ n20963);
assign n4257 = ~(n2731 ^ n4376);
assign n2866 = n791 | n11322;
assign n5929 = ~(n23746 ^ n7269);
assign n24220 = n11583 | n1138;
assign n11226 = ~(n161 | n12780);
assign n5189 = ~(n7777 | n23751);
assign n9811 = n7807 | n13846;
assign n27094 = n8252 | n11850;
assign n17324 = n3059 & n17361;
assign n9370 = ~(n11600 ^ n16843);
assign n3715 = n7517 | n24318;
assign n697 = n15841 | n24808;
assign n13196 = n18380 & n25645;
assign n19653 = n6446 | n20060;
assign n15520 = n16935 & n16691;
assign n5444 = n12224 | n25829;
assign n3646 = n5554 & n21461;
assign n8223 = n7670 | n3253;
assign n14309 = ~(n21846 | n25370);
assign n1913 = ~(n24999 ^ n23594);
assign n21115 = ~(n5171 ^ n3550);
assign n13685 = ~(n26952 ^ n17504);
assign n17209 = ~(n22432 | n14808);
assign n19655 = n7969 & n9640;
assign n21953 = n22803 & n26873;
assign n6901 = n24226 | n3112;
assign n23653 = ~(n27164 ^ n7868);
assign n17214 = n17470 | n25998;
assign n26643 = n4041 | n3378;
assign n2925 = n408 & n19853;
assign n19347 = ~(n17198 | n2923);
assign n7222 = n4622 | n27089;
assign n19243 = n4542 | n2586;
assign n23928 = n6454 & n5476;
assign n1357 = ~(n3762 ^ n1862);
assign n3775 = n4897 | n26819;
assign n27034 = n16444 | n16284;
assign n27038 = n7841 & n4941;
assign n14611 = n436 | n13464;
assign n12584 = n13523 | n6917;
assign n26777 = n19531 & n21322;
assign n19348 = n9987 | n4094;
assign n15482 = ~n25210;
assign n19861 = n9053 | n8974;
assign n11088 = ~n9993;
assign n15589 = n22527 | n2268;
assign n1214 = ~(n3632 ^ n682);
assign n14622 = ~(n21997 ^ n19701);
assign n11430 = n2195 & n21197;
assign n2971 = ~(n12374 ^ n7695);
assign n17225 = ~(n6356 ^ n12956);
assign n19110 = n24131 & n1088;
assign n24532 = n20489 | n21693;
assign n2276 = n24762 | n21862;
assign n16114 = n14239 & n23672;
assign n8161 = n12543 | n23793;
assign n16620 = n4613 & n6561;
assign n13523 = ~n27015;
assign n19572 = ~(n11871 ^ n987);
assign n15400 = ~n14298;
assign n9946 = ~(n12993 ^ n23987);
assign n26262 = n23189 | n26535;
assign n24831 = n17678 | n12065;
assign n6975 = ~(n26595 ^ n22717);
assign n26223 = n1272 | n14247;
assign n2536 = ~(n23715 ^ n19584);
assign n14333 = n17778 & n17072;
assign n13204 = ~(n16352 ^ n9943);
assign n6039 = ~n1171;
assign n21889 = n1165 & n18342;
assign n1203 = ~(n13172 | n1881);
assign n25259 = ~(n14391 | n6293);
assign n4829 = n24995 & n3866;
assign n19203 = ~(n15636 ^ n24618);
assign n25648 = n3364 & n19199;
assign n12627 = ~(n10712 ^ n26512);
assign n7006 = ~(n2243 ^ n7658);
assign n23412 = ~n22878;
assign n16175 = ~(n24343 ^ n15767);
assign n12934 = n3857 | n3761;
assign n27143 = n20358 & n21379;
assign n24702 = n14864 | n6667;
assign n13273 = ~(n1828 ^ n14305);
assign n12452 = n3009 & n21729;
assign n2932 = n25507 | n14340;
assign n25830 = n15015 | n11216;
assign n220 = n3717 & n19031;
assign n26966 = n11454 & n19364;
assign n13237 = ~n25872;
assign n26319 = ~(n13152 | n15053);
assign n11020 = ~(n22061 | n26705);
assign n7584 = ~(n6265 | n1336);
assign n16039 = n26322 | n9962;
assign n5334 = n2511 | n21714;
assign n11947 = ~(n6301 ^ n6626);
assign n5478 = n8104 & n899;
assign n6649 = n3253 | n21021;
assign n8921 = n25586 | n23525;
assign n15151 = n12795 | n13315;
assign n6241 = ~n2128;
assign n26969 = ~(n26135 ^ n8119);
assign n13562 = ~(n11323 ^ n24504);
assign n10226 = n16669 | n13656;
assign n3604 = ~(n23254 | n27008);
assign n9343 = n12513 | n25568;
assign n16643 = n13460 | n5156;
assign n9966 = ~(n7353 ^ n20620);
assign n25689 = n6107 & n8725;
assign n17871 = ~n18075;
assign n24471 = ~(n16158 | n10204);
assign n27180 = n346 | n27138;
assign n9363 = ~n22201;
assign n25439 = ~(n14018 ^ n7735);
assign n6608 = n4520 | n1694;
assign n12320 = ~(n4061 | n9557);
assign n1276 = n21140 | n10241;
assign n25651 = n26810 & n12797;
assign n18042 = n5258 | n10415;
assign n26711 = ~n12456;
assign n16770 = ~(n20970 | n12961);
assign n2542 = n1458 | n19494;
assign n16192 = ~(n18371 | n21151);
assign n23518 = n20229 | n1936;
assign n2255 = n9436 & n3905;
assign n16657 = ~(n2035 ^ n26823);
assign n12232 = ~n23488;
assign n9687 = ~(n21321 ^ n1750);
assign n4577 = ~(n24355 | n11220);
assign n24201 = ~(n5031 ^ n11926);
assign n24007 = n4435 & n8533;
assign n22297 = n14226 | n23217;
assign n1573 = ~(n2276 ^ n9937);
assign n6810 = n3982 & n6439;
assign n6525 = ~(n10620 ^ n10255);
assign n4732 = n7866 & n13676;
assign n1120 = ~(n25065 ^ n6500);
assign n26644 = n7759 & n725;
assign n4136 = n15363 & n11704;
assign n21750 = ~(n16191 ^ n11296);
assign n4825 = n18652 | n11574;
assign n14197 = n12591 | n24254;
assign n26733 = ~(n22057 ^ n1523);
assign n5359 = n123 | n11130;
assign n17026 = ~n21998;
assign n3416 = ~(n19399 | n13848);
assign n19173 = ~(n528 | n17556);
assign n22211 = n2481 ^ n13650;
assign n11258 = ~n8165;
assign n20464 = n26822 & n5475;
assign n26672 = ~n10967;
assign n17772 = n12876 | n3287;
assign n12701 = ~(n4335 | n21544);
assign n24656 = ~(n17423 | n5101);
assign n6337 = n4684 | n16942;
assign n15982 = n4458 | n3415;
assign n1183 = ~(n25285 ^ n8293);
assign n6820 = n4844 & n16723;
assign n17404 = n16901 | n26171;
assign n11227 = n1458 | n21372;
assign n13969 = n4904 | n13829;
assign n8186 = ~n2978;
assign n14146 = n12149 | n19045;
assign n26475 = ~(n15190 | n182);
assign n1511 = n1155 | n11688;
assign n9128 = n26335 | n24099;
assign n1833 = ~(n19138 | n21114);
assign n10529 = n24851 | n2636;
assign n8508 = ~(n6599 ^ n19608);
assign n3502 = ~(n3254 ^ n14418);
assign n22889 = n7561 | n10797;
assign n614 = ~(n144 | n18290);
assign n8103 = ~(n14934 ^ n13881);
assign n20209 = ~n16520;
assign n7980 = ~(n9376 | n3045);
assign n17760 = n13638 | n22798;
assign n14142 = n6252 & n19329;
assign n6518 = ~n9961;
assign n19730 = ~(n18578 ^ n9090);
assign n8503 = n21432 | n26994;
assign n13344 = n5773 | n20464;
assign n24895 = n2339 | n908;
assign n11573 = n9206 | n24682;
assign n15990 = n26085 | n1245;
assign n6156 = n21125 & n926;
assign n2005 = ~(n13904 ^ n18463);
assign n20897 = ~n1339;
assign n5800 = ~(n6657 ^ n3513);
assign n25789 = n8603 & n18469;
assign n23501 = n6855 | n17217;
assign n9910 = ~n25120;
assign n26701 = n17316 | n1893;
assign n2958 = n4735 & n25811;
assign n26207 = n6094 | n12877;
assign n16399 = ~n24721;
assign n5885 = ~(n13297 | n11165);
assign n3598 = n2063 | n9621;
assign n9111 = ~(n23369 ^ n26572);
assign n18062 = n25913 | n10230;
assign n18991 = ~n5329;
assign n25394 = ~n2429;
assign n19558 = ~(n26673 | n19911);
assign n7147 = ~(n21442 ^ n8891);
assign n24194 = ~(n8469 ^ n5367);
assign n5872 = n10758 | n1717;
assign n6826 = ~(n22984 ^ n25173);
assign n22612 = n21672 & n19300;
assign n18459 = ~(n11970 ^ n1757);
assign n11794 = ~(n27104 ^ n19005);
assign n14382 = n13494 | n14031;
assign n13809 = ~(n5031 | n11926);
assign n6352 = n10795;
assign n8918 = n24823 | n20886;
assign n14464 = ~(n3357 ^ n20772);
assign n8473 = ~(n17308 ^ n8751);
assign n3674 = ~n23993;
assign n4193 = n16209 | n15836;
assign n19451 = n15761 | n11535;
assign n16636 = n25728 & n11629;
assign n10889 = n18504 | n17483;
assign n25372 = n24657 & n114;
assign n21503 = n8914 & n4666;
assign n26722 = ~(n4 ^ n23544);
assign n4499 = ~(n7196 ^ n1778);
assign n20643 = n1195 & n21412;
assign n13143 = n4274 & n20177;
assign n12497 = n10145 | n7846;
assign n16190 = n10995 & n1082;
assign n15991 = ~(n15372 ^ n17857);
assign n21651 = n18510 | n9888;
assign n7077 = ~(n12702 ^ n18105);
assign n12766 = ~(n8193 ^ n9914);
assign n6233 = ~(n23356 ^ n11129);
assign n19745 = n16720 | n23510;
assign n3218 = ~(n17789 ^ n10915);
assign n13417 = n25291 & n7061;
assign n23433 = ~(n22210 ^ n21149);
assign n2453 = ~n12875;
assign n3290 = ~(n22554 | n26318);
assign n5335 = n9040 & n26799;
assign n1758 = n26354 & n11873;
assign n1522 = ~(n16266 ^ n22458);
assign n13925 = ~n11335;
assign n25609 = n22920 & n11715;
assign n8989 = ~(n19890 | n6449);
assign n16909 = ~(n11486 ^ n18409);
assign n5356 = ~(n16633 | n22793);
assign n14418 = ~(n728 ^ n12029);
assign n1978 = n24358 & n20951;
assign n13452 = ~(n5512 ^ n16217);
assign n9072 = ~(n7755 ^ n21097);
assign n24376 = ~(n6255 ^ n6658);
assign n7741 = n2160 & n27095;
assign n4711 = ~(n16399 | n11603);
assign n16131 = n25207 & n1101;
assign n26094 = ~(n19634 | n19228);
assign n12332 = n3899 & n15263;
assign n21506 = ~n10472;
assign n265 = ~n501;
assign n12046 = ~(n1314 | n20967);
assign n24160 = ~(n7603 ^ n15111);
assign n19916 = ~(n18402 ^ n21816);
assign n3368 = n12640 | n18274;
assign n8317 = ~(n2739 ^ n4865);
assign n22129 = n10757 | n13811;
assign n4465 = n21598 | n10161;
assign n21292 = ~(n5559 | n7697);
assign n23882 = ~(n9355 ^ n3844);
assign n7658 = ~(n987 ^ n626);
assign n8814 = n17514 | n20960;
assign n16240 = n26625 | n14230;
assign n19295 = ~n1167;
assign n17164 = ~n23326;
assign n23295 = ~(n6631 ^ n12209);
assign n11109 = ~(n16401 ^ n7861);
assign n23016 = ~n24202;
assign n15488 = ~(n19978 ^ n4240);
assign n10359 = ~(n2813 ^ n23272);
assign n17477 = n18057 | n9362;
assign n23403 = n20638 | n5296;
assign n11443 = ~(n9215 | n15616);
assign n12172 = n4117 & n14188;
assign n19758 = ~n4368;
assign n26886 = n19541 & n14182;
assign n4292 = n4543 | n18860;
assign n21718 = ~(n1798 ^ n1742);
assign n13048 = ~(n394 ^ n18005);
assign n21594 = n1660 | n23634;
assign n10831 = ~n2651;
assign n16928 = ~n9700;
assign n18961 = ~(n14514 ^ n2279);
assign n7121 = n7876 | n11479;
assign n6953 = n24768 & n1019;
assign n25417 = n17365 | n6000;
assign n24484 = ~n12291;
assign n17525 = n604 | n13318;
assign n7213 = ~n13665;
assign n3428 = n3260 & n20512;
assign n23758 = ~(n15440 | n3147);
assign n7509 = n6206 | n11529;
assign n9971 = ~(n5754 ^ n27032);
assign n5380 = n3788 & n5920;
assign n18212 = n18451 & n27034;
assign n17821 = n6103 & n15211;
assign n10983 = ~(n10184 | n12366);
assign n15256 = n5519 & n20934;
assign n1159 = n17970 & n15250;
assign n627 = n7472 | n3288;
assign n10070 = n15202 & n17124;
assign n25555 = ~(n3032 ^ n11911);
assign n16661 = n22087 | n4824;
assign n16931 = ~(n10989 | n19017);
assign n26434 = n7893 | n20205;
assign n26783 = n13088 & n18987;
assign n16140 = ~(n25974 ^ n8399);
assign n18299 = n20684 | n16518;
assign n21444 = ~(n8190 ^ n19714);
assign n18941 = n25642 & n1133;
assign n240 = ~(n1205 | n8568);
assign n3519 = ~(n9851 | n10389);
assign n15227 = n24220 & n14191;
assign n8726 = n14766 | n8808;
assign n5766 = ~(n21749 | n919);
assign n14277 = ~(n10526 ^ n8665);
assign n17173 = ~n10405;
assign n2777 = ~(n2780 | n4665);
assign n24583 = n7818 | n18139;
assign n1763 = n18119 | n23827;
assign n16783 = n19175 | n12343;
assign n4960 = n15820 | n21824;
assign n5573 = n13920 | n5839;
assign n26587 = n24384 & n10528;
assign n1695 = ~(n4194 ^ n14643);
assign n22796 = n435 | n14494;
assign n15317 = ~(n14386 | n24051);
assign n9449 = n6877 & n17155;
assign n5153 = n2797 | n17742;
assign n7639 = ~n8876;
assign n2824 = n23772 | n23106;
assign n24896 = ~(n1038 ^ n15342);
assign n8998 = ~(n24202 | n9595);
assign n6301 = n6317 & n2670;
assign n13563 = ~(n5516 | n24085);
assign n16033 = n23211 | n24665;
assign n8812 = n8865 | n12946;
assign n14806 = n21924 | n9476;
assign n16728 = n3591 & n3963;
assign n11196 = ~(n3280 ^ n2038);
assign n11989 = ~n10051;
assign n15592 = n9880 | n13714;
assign n2468 = ~(n7107 ^ n26582);
assign n23409 = n17356 & n11716;
assign n8576 = ~(n8097 | n17210);
assign n13112 = ~(n2068 ^ n12219);
assign n24496 = n12210 & n17085;
assign n451 = n19557 | n9040;
assign n2720 = n11637 | n27058;
assign n5965 = n16751 | n27082;
assign n9321 = ~(n14996 ^ n7678);
assign n15940 = ~n9318;
assign n245 = ~(n8399 ^ n13708);
assign n60 = ~(n16364 ^ n7680);
assign n19401 = ~(n15708 ^ n16969);
assign n19868 = ~n1304;
assign n24899 = ~(n3694 | n14514);
assign n12731 = ~(n24112 ^ n15077);
assign n2200 = n26014 & n14144;
assign n984 = ~(n3321 ^ n14888);
assign n17640 = ~(n1075 ^ n24016);
assign n21643 = ~(n95 ^ n3851);
assign n25835 = ~n9362;
assign n8596 = ~(n25435 ^ n18);
assign n19890 = n9356 | n17373;
assign n13039 = ~(n11253 ^ n9208);
assign n11565 = ~(n20751 ^ n24593);
assign n16196 = ~(n23154 ^ n13788);
assign n16144 = n2088 & n6414;
assign n22104 = ~n10004;
assign n19716 = ~(n8067 | n3319);
assign n11228 = ~n12573;
assign n3184 = n4070 | n15479;
assign n10693 = n12991 | n24700;
assign n20480 = ~(n18759 ^ n16244);
assign n19940 = ~(n13101 ^ n19817);
assign n13034 = ~(n3944 ^ n941);
assign n25330 = ~n22138;
assign n910 = ~n3016;
assign n18612 = ~(n7769 | n25316);
assign n13103 = n25940 & n22325;
assign n121 = n4058 | n19534;
assign n8580 = ~(n15546 | n5629);
assign n4623 = ~(n20597 ^ n20055);
assign n6664 = ~(n5715 | n22918);
assign n13139 = ~(n20075 ^ n14386);
assign n9446 = n3348 & n202;
assign n9915 = ~(n1509 ^ n2517);
assign n23450 = ~(n6865 ^ n16378);
assign n21315 = ~(n18797 ^ n25799);
assign n20174 = n15864 | n1455;
assign n18819 = n20752 | n5458;
assign n4035 = n13775 & n8389;
assign n6964 = n4926 | n4517;
assign n6986 = n19650 | n21616;
assign n12310 = n16237 & n23003;
assign n5513 = ~(n13490 ^ n12446);
assign n19759 = n2038 & n2574;
assign n18297 = n6393 & n2028;
assign n18187 = ~(n15770 ^ n22881);
assign n24799 = n21634 & n16007;
assign n7015 = n11978 | n1194;
assign n9140 = n9681 | n16475;
assign n26962 = ~n7634;
assign n26211 = ~n7049;
assign n7252 = ~n5188;
assign n15998 = ~n2696;
assign n765 = ~(n9793 ^ n10250);
assign n16489 = n267 & n16317;
assign n23287 = ~(n24948 ^ n10514);
assign n13328 = ~(n7749 ^ n8681);
assign n13897 = ~n17035;
assign n24925 = ~n287;
assign n7872 = ~(n13633 ^ n19039);
assign n15099 = n25844 | n15552;
assign n15124 = n1330 & n14077;
assign n7545 = n22781 | n20394;
assign n12568 = n13481 | n11238;
assign n10272 = ~(n14510 ^ n16988);
assign n3042 = n6920 & n1286;
assign n6939 = ~(n15903 ^ n13468);
assign n2780 = ~n8309;
assign n19237 = n10171 & n10348;
assign n2755 = ~(n11207 ^ n22358);
assign n4713 = ~(n2420 ^ n22201);
assign n5248 = n9899 | n26952;
assign n4900 = n19894 & n22517;
assign n2006 = n9600 | n17870;
assign n25982 = ~n7707;
assign n5270 = n15554 & n66;
assign n11046 = n24044 | n22379;
assign n19244 = ~(n19654 ^ n21642);
assign n26524 = ~n22898;
assign n12038 = ~(n13089 | n3625);
assign n25493 = n13428 | n1368;
assign n17869 = ~n914;
assign n17633 = n2814 & n7651;
assign n5528 = n21051 & n16035;
assign n27003 = ~(n22874 | n9492);
assign n110 = ~(n333 ^ n15268);
assign n13944 = ~n10479;
assign n3322 = n17848 | n5863;
assign n24267 = ~(n20378 | n9493);
assign n8925 = ~n11254;
assign n15310 = n12894 | n25646;
assign n12611 = n25450 | n2128;
assign n8427 = ~(n16555 ^ n20040);
assign n14208 = n13159 & n15924;
assign n12492 = n1190 | n14721;
assign n8200 = n9496 | n22515;
assign n27019 = ~(n10110 ^ n22669);
assign n17130 = ~(n23507 ^ n16871);
assign n19139 = ~(n1163 | n2675);
assign n26527 = n17908 | n21550;
assign n18720 = ~(n26637 ^ n19866);
assign n24874 = n16372 & n10845;
assign n7035 = ~(n19789 | n21226);
assign n24655 = n13059 & n22913;
assign n21956 = ~(n23793 ^ n18);
assign n19705 = ~(n14444 | n1780);
assign n15654 = ~(n7428 ^ n19107);
assign n1426 = ~(n21079 ^ n369);
assign n25300 = n16770 | n12032;
assign n9113 = ~n27141;
assign n8894 = n6804 & n11768;
assign n8548 = n18666 | n26575;
assign n10023 = n23310;
assign n25122 = ~n7335;
assign n25844 = ~(n14736 | n22139);
assign n14797 = ~(n17122 ^ n23383);
assign n17765 = ~(n874 ^ n16949);
assign n19411 = n22320 & n6563;
assign n16579 = n9805 | n19055;
assign n20437 = ~n18416;
assign n21547 = n17152;
assign n1421 = ~n10039;
assign n3131 = ~(n6072 ^ n11706);
assign n23833 = ~(n8712 ^ n26620);
assign n2984 = n18074 & n26476;
assign n22269 = n23000 & n24908;
assign n3378 = ~n2965;
assign n23404 = n1250 | n8413;
assign n20626 = ~(n8672 ^ n26224);
assign n2869 = ~(n21948 ^ n20840);
assign n4282 = ~n21908;
assign n21060 = ~n14482;
assign n26651 = ~(n20700 ^ n932);
assign n14988 = ~(n18295 | n25974);
assign n10351 = n23141 & n3238;
assign n14555 = ~n25601;
assign n2963 = ~(n23895 ^ n5101);
assign n16606 = n19731 | n23993;
assign n1411 = n18379 & n21285;
assign n5880 = ~(n24624 ^ n23517);
assign n18457 = n15711 | n27124;
assign n22146 = n9373 | n7765;
assign n4153 = ~(n18640 ^ n3814);
assign n1551 = n9825 | n18612;
assign n14728 = ~(n9751 ^ n17353);
assign n24919 = ~(n26083 ^ n22734);
assign n17127 = n1937 | n1310;
assign n26844 = n7421 | n20044;
assign n17511 = ~n3509;
assign n17457 = n25156 | n2784;
assign n24943 = n6369 | n527;
assign n19136 = n4820 | n7745;
assign n15068 = n2976 | n10904;
assign n20593 = n17453 & n26783;
assign n21875 = n17464 & n4536;
assign n1635 = ~(n13422 | n685);
assign n12800 = ~(n24327 | n2768);
assign n17986 = n10175 & n22129;
assign n15697 = ~(n6750 | n63);
assign n276 = n3062 | n18047;
assign n22057 = n13756 | n7244;
assign n1001 = ~(n4625 ^ n20835);
assign n13386 = ~(n19515 | n10651);
assign n2995 = ~n13475;
assign n6834 = ~(n5488 ^ n7149);
assign n9255 = n13195 | n12217;
assign n20546 = ~(n20323 ^ n8564);
assign n23778 = ~(n23353 ^ n12702);
assign n6490 = n8325 & n13866;
assign n7896 = n25058 | n15487;
assign n26658 = ~n10053;
assign n2701 = n7681 | n2338;
assign n25922 = ~(n16795 | n17498);
assign n14861 = ~(n22281 | n18157);
assign n10720 = ~n1685;
assign n20354 = ~(n1478 ^ n12731);
assign n7637 = n26121 & n1409;
assign n18129 = n20228 & n8717;
assign n8765 = ~(n7430 ^ n18218);
assign n13833 = n23887 & n18989;
assign n25576 = ~(n23180 ^ n18690);
assign n18324 = n23097 | n7399;
assign n21648 = n9407 | n9109;
assign n24512 = ~(n2492 ^ n22175);
assign n14070 = ~(n9108 ^ n6877);
assign n21128 = ~(n21489 | n11062);
assign n15960 = ~(n18 ^ n22843);
assign n21985 = n9176 & n4907;
assign n6634 = ~(n9029 ^ n22711);
assign n4921 = n15785 & n16953;
assign n21369 = ~(n6187 | n25641);
assign n26056 = ~n14125;
assign n9985 = ~(n20151 | n19042);
assign n9834 = ~(n14472 | n26821);
assign n1039 = ~(n16396 | n8399);
assign n5857 = ~(n21101 ^ n16722);
assign n22887 = ~(n13941 | n6025);
assign n8874 = ~(n9003 ^ n6369);
assign n19190 = ~(n10919 ^ n8943);
assign n33 = n1557 | n5892;
assign n4348 = n23553 & n12643;
assign n24043 = ~n5733;
assign n5392 = ~(n3809 ^ n8719);
assign n4485 = n25242 & n8868;
assign n11411 = n23223 & n13785;
assign n831 = n20638 | n22986;
assign n3533 = n21201 & n26242;
assign n15764 = ~(n19990 ^ n18313);
assign n8400 = n25424 | n14432;
assign n21463 = n25510 | n4504;
assign n2823 = n16512 | n11340;
assign n25322 = ~(n16334 ^ n21784);
assign n24975 = ~(n17835 ^ n7026);
assign n14864 = ~(n20470 | n3366);
assign n6471 = ~(n17498 ^ n24989);
assign n8911 = ~(n27047 ^ n23698);
assign n16634 = n3959 & n25917;
assign n9500 = ~(n11802 ^ n15975);
assign n13182 = n17916 & n21624;
assign n18705 = ~(n19302 ^ n18875);
assign n26350 = ~n2954;
assign n17489 = n23998 & n17043;
assign n24429 = n11865 | n10876;
assign n9011 = ~(n246 ^ n17401);
assign n15968 = n18929 | n22036;
assign n27072 = ~(n25720 ^ n19834);
assign n4458 = n3199 & n3373;
assign n2881 = ~(n13958 ^ n15586);
assign n5069 = ~(n2470 | n10496);
assign n17012 = ~(n14886 ^ n17639);
assign n26439 = ~(n10128 ^ n16340);
assign n3234 = ~(n12508 ^ n22850);
assign n7735 = ~(n12379 ^ n8067);
assign n17239 = n19033 | n20724;
assign n10788 = ~n3968;
assign n21550 = n18879 & n25011;
assign n8057 = n23579 & n26223;
assign n19227 = n4956;
assign n9080 = ~(n16359 | n26149);
assign n5207 = n25248 & n13931;
assign n13086 = n13596 | n10649;
assign n7623 = ~(n26717 | n7963);
assign n14636 = ~(n1548 ^ n18661);
assign n1872 = n14684 | n21952;
assign n4018 = n9664 & n20122;
assign n22607 = ~(n13583 ^ n2963);
assign n14003 = ~(n24061 ^ n128);
assign n21345 = n26145 | n20360;
assign n10929 = ~(n13668 ^ n20923);
assign n22627 = ~(n26023 ^ n4692);
assign n23048 = ~(n14770 ^ n15234);
assign n3594 = ~(n3968 | n13980);
assign n27174 = n19862 | n16722;
assign n22719 = n3739 | n15892;
assign n14820 = n65 | n22464;
assign n10795 = n12779 & n18329;
assign n8070 = ~(n17221 ^ n6491);
assign n24434 = n19361 | n20060;
assign n15269 = ~n23784;
assign n1643 = n725 & n24804;
assign n21865 = ~(n19926 | n21295);
assign n12853 = n19869 | n20092;
assign n748 = n4913 | n13489;
assign n1851 = ~(n6486 ^ n15077);
assign n20447 = ~(n11589 ^ n4518);
assign n16052 = ~n21405;
assign n19793 = ~(n12657 ^ n23697);
assign n13164 = ~n4207;
assign n270 = n20249 | n9736;
assign n19224 = ~(n19754 ^ n20611);
assign n5192 = n17264 & n9128;
assign n10945 = n16474 & n15491;
assign n14098 = n14654 | n18519;
assign n1211 = n5055 | n1318;
assign n19620 = n23169 & n2823;
assign n23883 = ~(n2097 ^ n2869);
assign n24414 = n19144 & n5496;
assign n7530 = n25745 & n5291;
assign n340 = n19003 | n24475;
assign n4403 = ~(n12088 ^ n16029);
assign n5659 = n6796 & n1032;
assign n21672 = ~n18672;
assign n25702 = n19264 | n22088;
assign n6663 = n24098 | n23250;
assign n26017 = n16010 & n7984;
assign n2700 = ~(n3164 ^ n268);
assign n23098 = ~n7407;
assign n17756 = ~(n18191 ^ n21993);
assign n2081 = n13420 | n19337;
assign n16768 = ~(n16482 ^ n13074);
assign n3986 = ~(n26251 ^ n1630);
assign n21766 = n1742 & n25394;
assign n1624 = ~n7755;
assign n25096 = n17333 & n19247;
assign n19840 = n14963 & n19112;
assign n18576 = ~(n14935 ^ n9256);
assign n16771 = n1319 & n6864;
assign n21653 = n7215 | n23493;
assign n2670 = n10707 | n6535;
assign n25709 = n1812 | n15172;
assign n9077 = ~(n14652 ^ n9742);
assign n4077 = ~n6107;
assign n22222 = ~n1429;
assign n9600 = ~n10593;
assign n13588 = n10138 & n10105;
assign n888 = ~(n22824 | n23686);
assign n26694 = ~(n24868 ^ n13044);
assign n16523 = n18764 & n14175;
assign n3051 = n23094 & n24658;
assign n20861 = n6386 & n3501;
assign n13910 = ~(n18125 | n15131);
assign n25465 = ~(n19766 ^ n11557);
assign n27065 = ~n13476;
assign n23808 = ~(n8431 | n21547);
assign n2613 = ~(n26007 | n5621);
assign n10254 = n22071 & n26291;
assign n27166 = n8259 | n16551;
assign n20347 = n11645 & n17807;
assign n3255 = n2048 | n2607;
assign n25859 = n23030 | n4333;
assign n21737 = n25469 & n20631;
assign n316 = n11219 & n3088;
assign n11358 = n24012 | n12109;
assign n160 = n26408 | n1186;
assign n646 = ~(n14987 ^ n12959);
assign n18629 = n16474 | n18302;
assign n1280 = ~(n20667 | n26066);
assign n3374 = n3633 | n23389;
assign n24238 = n9255 & n7513;
assign n6469 = n5257 & n6876;
assign n10583 = n16159 | n22378;
assign n27194 = ~(n6114 ^ n1671);
assign n3163 = n17456 | n25653;
assign n20655 = ~n16907;
assign n9964 = ~n1451;
assign n13611 = ~(n21842 ^ n3828);
assign n13940 = ~(n15780 ^ n2387);
assign n25966 = ~(n25197 ^ n23498);
assign n25273 = n6554 & n25060;
assign n11526 = n15998 | n5142;
assign n9622 = ~(n21618 ^ n26337);
assign n8573 = ~(n24736 ^ n14603);
assign n25895 = n5245 | n11259;
assign n4398 = ~(n7249 | n10441);
assign n8236 = n3254 & n2738;
assign n12968 = ~n16264;
assign n1840 = ~(n18634 ^ n20470);
assign n13560 = ~(n1694 ^ n9909);
assign n4721 = ~n6105;
assign n24559 = ~n22314;
assign n24984 = n20325 | n5515;
assign n17236 = ~(n22263 ^ n9581);
assign n24005 = ~(n665 | n17599);
assign n3602 = n7973 ^ n8381;
assign n1007 = ~(n22349 ^ n13493);
assign n3857 = n16054 & n17600;
assign n14246 = n17598 | n17926;
assign n7157 = ~(n18255 ^ n23369);
assign n25594 = n21554 & n25158;
assign n26765 = ~(n11098 ^ n13912);
assign n3685 = ~(n12048 | n8210);
assign n17877 = ~(n9960 | n21482);
assign n6163 = n536 | n4848;
assign n4512 = n12006 & n21806;
assign n18510 = ~n11314;
assign n23710 = ~n8206;
assign n12397 = n3153 | n23459;
assign n266 = ~(n21591 ^ n13612);
assign n16919 = n20728 | n11483;
assign n6627 = n14514 | n3848;
assign n11436 = n26184 | n316;
assign n17293 = ~(n15265 | n12152);
assign n2356 = ~(n21014 ^ n8958);
assign n15858 = n109 & n6503;
assign n10039 = ~(n17979 ^ n22659);
assign n7839 = n10969 | n16470;
assign n2554 = n5586 | n19522;
assign n9258 = n524 | n25069;
assign n23391 = n25558 | n3414;
assign n18353 = ~(n24312 | n10847);
assign n14083 = n19043 & n1087;
assign n9581 = ~(n17953 ^ n12971);
assign n10074 = n340 & n700;
assign n14875 = ~n3019;
assign n12249 = ~n280;
assign n4895 = n13081 & n18729;
assign n21828 = ~(n13449 ^ n6381);
assign n21796 = ~n15126;
assign n25036 = ~n16173;
assign n13412 = ~(n7546 ^ n25846);
assign n15931 = ~(n15710 ^ n23309);
assign n23202 = ~(n20920 | n26851);
assign n6958 = n27104 | n15618;
assign n2592 = n3921 | n1894;
assign n850 = ~n12100;
assign n18747 = n13889 | n12123;
assign n3696 = n1438 & n11527;
assign n17701 = n17925 & n2270;
assign n3885 = n26683 & n16087;
assign n21454 = n7455 | n27200;
assign n18246 = n12277 | n10454;
assign n9793 = ~(n25683 ^ n15014);
assign n19538 = n26475 | n25364;
assign n4643 = n23126 & n10781;
assign n6850 = ~(n8006 ^ n15289);
assign n15281 = ~(n22492 ^ n9372);
assign n12860 = ~(n20876 ^ n24335);
assign n13448 = ~n21150;
assign n22174 = n20973 | n13539;
assign n5053 = ~(n16544 ^ n2160);
assign n17492 = n6026 | n8531;
assign n4678 = n11303 | n5948;
assign n22707 = n9378 | n10833;
assign n10365 = ~(n24897 | n24040);
assign n19549 = ~n25602;
assign n23510 = n13586 & n26950;
assign n188 = ~(n26522 ^ n1553);
assign n3963 = ~(n5644 ^ n827);
assign n1059 = ~(n25794 | n6944);
assign n3203 = ~n13195;
assign n16259 = n22727 | n17411;
assign n6804 = n7041 | n1924;
assign n4925 = ~(n21466 ^ n8598);
assign n7320 = ~n13914;
assign n25761 = n15888 | n1398;
assign n22212 = n2903 & n27041;
assign n21526 = n23337 | n16213;
assign n4655 = n3780 | n26311;
assign n21925 = n13443 | n10739;
assign n2847 = n8741 | n23919;
assign n6546 = n15274 | n16514;
assign n14004 = ~(n25789 ^ n2198);
assign n3346 = ~(n25275 ^ n18271);
assign n24244 = n15137 & n1305;
assign n21738 = n7956 & n4563;
assign n1632 = ~(n7561 ^ n8714);
assign n4592 = n11669 | n26523;
assign n22858 = ~(n4106 ^ n22398);
assign n20881 = ~(n2780 | n7910);
assign n2942 = ~(n8195 ^ n23757);
assign n15041 = ~n26109;
assign n22939 = ~(n15067 ^ n18075);
assign n16230 = ~(n27202 ^ n24482);
assign n7809 = ~(n1546 ^ n21532);
assign n18293 = n21213 & n4685;
assign n4573 = n21659 | n24914;
assign n15217 = ~n17250;
assign n3679 = ~(n11108 ^ n16794);
assign n20942 = n2863 & n21043;
assign n17309 = ~(n13286 ^ n14341);
assign n32 = ~n2127;
assign n13402 = n6764 | n2088;
assign n15732 = n9289 & n23152;
assign n24047 = ~(n22139 ^ n10343);
assign n19669 = n24671 | n10431;
assign n4758 = ~(n21839 ^ n22270);
assign n7662 = ~(n8492 | n8695);
assign n15285 = ~(n12049 ^ n9392);
assign n5473 = n14325 & n20063;
assign n13704 = ~(n9259 | n6456);
assign n12506 = n22230 | n20005;
assign n14161 = n23721 & n15849;
assign n23805 = ~n13277;
assign n19747 = ~(n27102 ^ n20250);
assign n17804 = ~(n17029 ^ n1416);
assign n25246 = ~n24161;
assign n27146 = ~(n16437 ^ n1129);
assign n7551 = ~(n9908 | n4576);
assign n22113 = ~(n2810 ^ n4929);
assign n23192 = ~(n18290 ^ n23529);
assign n8939 = n1178 | n1148;
assign n15046 = n13312 & n21706;
assign n962 = ~n1022;
assign n5858 = n2752 & n3678;
assign n10716 = ~(n349 | n12456);
assign n2664 = n6509 | n6080;
assign n1504 = n22901 & n16861;
assign n3996 = ~(n1205 | n13319);
assign n15899 = n22604 | n2093;
assign n5233 = n1186 & n12317;
assign n968 = ~(n10799 | n19326);
assign n2230 = ~n8381;
assign n12230 = ~(n18575 ^ n10430);
assign n19792 = ~(n13232 ^ n5507);
assign n24725 = n13339 | n13178;
assign n1843 = ~(n14265 | n15906);
assign n10537 = ~(n593 ^ n20036);
assign n8094 = ~n342;
assign n3385 = ~(n5095 | n24134);
assign n10727 = n25183 & n26531;
assign n459 = n17946 & n26697;
assign n26477 = ~n3196;
assign n26940 = ~(n16544 ^ n4319);
assign n7884 = ~(n14956 ^ n13622);
assign n11385 = n15265 | n9911;
assign n19560 = ~(n4921 ^ n15649);
assign n1817 = n12974 & n4332;
assign n8875 = n19162;
assign n19167 = n15522 | n21852;
assign n16018 = n18228 | n23651;
assign n11018 = ~(n25898 ^ n21674);
assign n8358 = ~(n17424 ^ n2370);
assign n12011 = ~(n16114 ^ n12195);
assign n11953 = ~(n4514 | n21698);
assign n14652 = ~n2020;
assign n11922 = n25178 | n9150;
assign n8919 = n2091 | n1940;
assign n25671 = n16386 & n5739;
assign n3246 = n5899 | n16567;
assign n16099 = ~(n24949 ^ n6199);
assign n14615 = ~n19683;
assign n23603 = ~(n8331 | n26216);
assign n6857 = ~n9851;
assign n17665 = n20249 | n26292;
assign n1749 = ~n9701;
assign n259 = ~(n20549 ^ n10551);
assign n24558 = ~(n6073 ^ n11344);
assign n18355 = ~n25617;
assign n9939 = n20290 | n21577;
assign n26610 = n22460 | n15788;
assign n23983 = ~n11351;
assign n21521 = ~(n26235 ^ n8146);
assign n19612 = n3440 | n6028;
assign n1448 = ~(n16482 ^ n5400);
assign n18427 = ~(n4858 ^ n23586);
assign n12481 = ~n9494;
assign n5603 = ~(n26558 ^ n23551);
assign n15094 = ~(n2075 ^ n11713);
assign n6361 = n16632 & n8460;
assign n2906 = ~n7162;
assign n25778 = ~(n16200 ^ n2743);
assign n15981 = ~(n12472 | n10397);
assign n16299 = ~(n4288 ^ n14902);
assign n6202 = n20014;
assign n20400 = ~(n8101 | n15109);
assign n12764 = ~(n6209 | n9507);
assign n3891 = ~(n10171 ^ n14499);
assign n6821 = n9988 | n21667;
assign n19811 = n23089 & n9830;
assign n24729 = n25316 & n8068;
assign n25920 = ~(n20957 | n25939);
assign n1896 = ~n18295;
assign n22189 = n8796 | n13833;
assign n21626 = ~(n16357 ^ n27187);
assign n15702 = n2985 | n13578;
assign n11260 = n7127 & n22013;
assign n5169 = ~(n2406 ^ n23251);
assign n4661 = ~(n21698 ^ n4514);
assign n13383 = ~(n8285 ^ n9323);
assign n6805 = ~n20384;
assign n21407 = n8575 & n5653;
assign n21240 = ~(n21028 ^ n4037);
assign n3815 = n6321 | n9802;
assign n12834 = n6227 & n14938;
assign n12745 = n15198 | n10848;
assign n4314 = n14858 | n12127;
assign n25390 = ~(n8589 | n3619);
assign n8115 = n323 | n5416;
assign n12391 = n9031 & n26430;
assign n25224 = n20085 & n13132;
assign n24361 = n25514 | n6254;
assign n7746 = ~(n13783 ^ n25119);
assign n2300 = ~n21529;
assign n3175 = n16790 & n26;
assign n7969 = n9425 | n22886;
assign n17657 = n25132 | n11546;
assign n9666 = n22982 & n1213;
assign n10145 = n20393 & n26832;
assign n7230 = ~(n6758 ^ n19585);
assign n6481 = ~(n3053 ^ n5436);
assign n23041 = n236 | n6540;
assign n13004 = ~(n23053 ^ n8612);
assign n12115 = n10514 & n24806;
assign n17815 = ~(n5052 ^ n21670);
assign n3684 = n15222 & n26579;
assign n13292 = ~n21733;
assign n13282 = ~n25442;
assign n2983 = n17895 & n4197;
assign n5275 = ~(n6789 ^ n26417);
assign n10796 = n21749 | n11676;
assign n20747 = ~(n24375 | n14625);
assign n19919 = ~(n24266 ^ n10493);
assign n24360 = n7909 & n16864;
assign n5764 = ~(n22895 ^ n17203);
assign n3843 = ~(n26051 ^ n18967);
assign n26972 = ~(n14166 ^ n25045);
assign n23768 = ~(n13237 | n12921);
assign n11640 = ~(n17174 ^ n26144);
assign n20601 = n20666 | n24251;
assign n21747 = n9211 & n24394;
assign n13617 = ~(n13899 ^ n21037);
assign n3072 = ~(n5175 ^ n15322);
assign n14961 = ~(n12960 | n6131);
assign n15917 = ~(n4222 ^ n25446);
assign n5135 = n18779 & n17905;
assign n14991 = ~n442;
assign n20328 = ~(n22660 ^ n26823);
assign n11472 = ~(n15177 ^ n13478);
assign n7094 = ~n18345;
assign n27184 = n26673 & n6820;
assign n17844 = n2141 | n5790;
assign n21625 = n25075 | n15564;
assign n24127 = ~(n19277 | n5213);
assign n17742 = n7736 & n18739;
assign n25232 = ~(n647 ^ n19941);
assign n12771 = ~(n11627 ^ n7593);
assign n16578 = n15832 | n19889;
assign n17641 = ~n2985;
assign n15901 = n5956;
assign n10722 = ~n1889;
assign n2969 = n9930 & n1062;
assign n20663 = n26537 & n25162;
assign n2844 = n10334 | n7557;
assign n13971 = n1461 | n5996;
assign n12987 = ~(n1983 ^ n622);
assign n11115 = ~(n4872 | n24009);
assign n6739 = n13039 | n6043;
assign n13304 = n4031 & n11697;
assign n6153 = n14492 | n1125;
assign n11571 = n21799 & n7620;
assign n21349 = ~(n23571 ^ n25104);
assign n5449 = ~n13069;
assign n12541 = ~(n14641 ^ n13499);
assign n7940 = ~(n23600 ^ n25887);
assign n8819 = ~n2698;
assign n23934 = n21663 | n11323;
assign n25833 = n12282 | n11003;
assign n16122 = n21814 & n19073;
assign n7056 = ~n14720;
assign n19833 = n16744 | n24383;
assign n24543 = n6712 & n15028;
assign n15898 = n26041 & n19135;
assign n15290 = n25663 | n9586;
assign n11421 = n5106 | n9666;
assign n18449 = n10947 | n23354;
assign n19394 = ~(n3044 ^ n23453);
assign n13253 = n14620 | n26914;
assign n19912 = ~(n15930 ^ n23207);
assign n11549 = n25466 | n16876;
assign n15294 = ~n24072;
assign n8493 = n18883 | n25146;
assign n7937 = ~(n2969 ^ n24742);
assign n7446 = n24521 | n35;
assign n2205 = n230 & n27109;
assign n22932 = n12909 & n12173;
assign n9338 = n13983 | n59;
assign n3790 = ~n11377;
assign n6893 = ~(n9507 ^ n10158);
assign n4429 = ~(n4825 ^ n22383);
assign n20625 = n17077 | n14620;
assign n3235 = ~(n22896 ^ n8848);
assign n18592 = ~(n1483 ^ n19539);
assign n4406 = n20654 | n5362;
assign n13323 = n7656 & n10104;
assign n14559 = ~(n19236 | n21930);
assign n7171 = n15638 & n11636;
assign n21543 = ~n9247;
assign n16212 = n11064 | n23524;
assign n977 = ~n17455;
assign n25470 = ~(n19009 ^ n4927);
assign n16471 = n16599 & n21202;
assign n10915 = ~(n15612 ^ n25884);
assign n18750 = ~(n23200 | n8391);
assign n14716 = ~(n6501 ^ n623);
assign n25616 = n12351 & n6503;
assign n8318 = n1502 & n22128;
assign n8344 = ~n2387;
assign n17381 = ~n5842;
assign n21034 = ~(n4951 | n26653);
assign n22485 = n18341 & n18262;
assign n16559 = ~n18826;
assign n7837 = n6907 | n23280;
assign n15016 = n8439 | n11106;
assign n1542 = n4011 & n26002;
assign n10031 = n16190 | n23696;
assign n21809 = ~(n2371 ^ n19255);
assign n9586 = ~n10577;
assign n12827 = ~(n2377 ^ n19633);
assign n19463 = n5986 | n23907;
assign n12117 = ~(n25877 | n5026);
assign n14682 = n5146 | n8957;
assign n7493 = n979 | n6968;
assign n8853 = ~n21858;
assign n11019 = n1284 & n8876;
assign n25070 = n21918 & n18974;
assign n14863 = n5826 | n23597;
assign n1569 = n16537 | n11783;
assign n26522 = ~(n24984 ^ n7275);
assign n4168 = ~(n2729 ^ n22298);
assign n12385 = ~(n22330 ^ n17913);
assign n7550 = n14790 | n5105;
assign n19388 = n22793 | n15016;
assign n19341 = n4841 & n2714;
assign n11081 = n14728 & n8570;
assign n7792 = ~(n7407 ^ n3030);
assign n26476 = n24963 | n10412;
assign n21316 = ~(n18409 ^ n5704);
assign n1781 = ~(n25049 | n23451);
assign n1095 = ~(n22892 | n5165);
assign n8370 = ~(n19762 | n9789);
assign n13777 = n18649 | n13968;
assign n14620 = ~(n4036 ^ n7330);
assign n15995 = n1558 & n17305;
assign n17997 = ~(n15236 ^ n23692);
assign n20612 = ~(n17047 | n851);
assign n23416 = n6924 & n18283;
assign n26308 = n23711 | n16785;
assign n20765 = n24457 | n19181;
assign n15206 = ~(n23061 ^ n21276);
assign n11417 = ~(n16712 | n10053);
assign n20949 = n1051 | n18365;
assign n27051 = ~(n18917 ^ n16368);
assign n18435 = n14338 & n18422;
assign n19512 = n10490 | n13324;
assign n10263 = ~(n10763 ^ n22379);
assign n3904 = ~(n6218 | n19652);
assign n23679 = n22879 | n12616;
assign n25979 = ~(n26264 ^ n21905);
assign n16380 = ~(n10501 | n5914);
assign n26058 = ~(n22935 ^ n4407);
assign n25827 = ~n10709;
assign n15510 = n16670 | n17247;
assign n21982 = ~n15652;
assign n24162 = ~(n20959 | n26947);
assign n13269 = ~n12385;
assign n19923 = ~(n9123 ^ n1632);
assign n19140 = n9490 | n4955;
assign n12925 = n18639 | n22399;
assign n13907 = ~n8319;
assign n20915 = ~(n18389 ^ n11401);
assign n15362 = ~(n3324 ^ n2272);
assign n2165 = ~n18638;
assign n11778 = n17061 | n25419;
assign n27006 = ~(n11486 ^ n13781);
assign n5079 = ~(n18934 | n11086);
assign n25529 = ~(n23677 | n19717);
assign n15588 = ~(n5773 ^ n20012);
assign n17884 = n17173 | n12236;
assign n22560 = n22313 | n761;
assign n18846 = ~n10785;
assign n4770 = ~(n24287 ^ n1225);
assign n195 = ~(n23878 ^ n1163);
assign n11332 = n24662 | n23046;
assign n15139 = ~(n5892 ^ n1231);
assign n10016 = n22971 | n20827;
assign n2291 = ~(n8602 ^ n3387);
assign n16956 = n8121 & n7723;
assign n1264 = ~(n1406 | n10372);
assign n19459 = ~(n23932 ^ n4939);
assign n4523 = ~(n25700 ^ n16803);
assign n24826 = ~(n13836 ^ n25652);
assign n22406 = ~(n15167 ^ n20036);
assign n21447 = n19026 & n20473;
assign n8471 = n2119 & n12982;
assign n11600 = ~(n10384 ^ n19575);
assign n8251 = ~(n25889 ^ n7885);
assign n22395 = ~(n21769 ^ n14779);
assign n2728 = ~(n26979 ^ n1152);
assign n1092 = ~(n21810 ^ n10235);
assign n18638 = n22720 & n1158;
assign n15720 = n13165 | n12689;
assign n16765 = ~(n12994 ^ n15594);
assign n13763 = n2045 | n9992;
assign n372 = n7204 | n19426;
assign n22822 = ~(n6309 ^ n15661);
assign n15873 = ~(n12956 ^ n1118);
assign n22085 = n3744 & n12248;
assign n6934 = n6228 & n16248;
assign n10687 = ~(n12070 | n3496);
assign n7074 = n5816 | n1329;
assign n21743 = ~n2813;
assign n13873 = ~n12702;
assign n20006 = ~n26463;
assign n22945 = ~(n13317 ^ n27104);
assign n17694 = n4028 | n21187;
assign n24933 = ~n19317;
assign n8209 = n12272 & n16709;
assign n6806 = n17710 | n3531;
assign n20490 = n2927 | n26677;
assign n26055 = ~(n20338 ^ n2756);
assign n6248 = ~(n9016 ^ n9120);
assign n12792 = n10037 | n678;
assign n3565 = ~(n17626 ^ n25241);
assign n4166 = ~(n11840 ^ n23059);
assign n15195 = n18773 | n1645;
assign n16540 = n771 & n23383;
assign n6711 = ~(n14997 ^ n8461);
assign n9857 = ~(n26882 | n19618);
assign n15125 = ~n26744;
assign n21162 = ~n513;
assign n5815 = n5127 & n21110;
assign n16042 = n2302 | n14535;
assign n11055 = ~(n5617 | n22414);
assign n13243 = ~(n20570 | n23962);
assign n9736 = ~n24684;
assign n10626 = ~(n17762 ^ n16247);
assign n17048 = n16658 | n20740;
assign n17536 = ~n14366;
assign n1710 = n19996 | n10421;
assign n2465 = n9068 | n24319;
assign n10755 = n25969 & n2447;
assign n15428 = ~(n17211 ^ n25509);
assign n12621 = ~(n10616 ^ n13060);
assign n25736 = n4878 | n2477;
assign n5148 = n22169 | n23783;
assign n7261 = ~(n1662 | n20946);
assign n11545 = n3455 | n14549;
assign n20387 = n17802 | n16487;
assign n21701 = ~n16249;
assign n17763 = n26633 & n2900;
assign n2888 = n2875 | n601;
assign n11383 = n4362 & n8514;
assign n8445 = n16048 & n7843;
assign n16133 = ~(n7071 | n14848);
assign n5984 = ~(n4484 ^ n2175);
assign n10981 = n13679 | n11811;
assign n25741 = n15138 | n26318;
assign n12837 = ~n3697;
assign n22733 = ~(n15905 | n23160);
assign n21937 = ~n27037;
assign n24213 = ~(n12233 ^ n2552);
assign n15715 = ~n11749;
assign n12428 = n8015 | n20255;
assign n26700 = n19382 & n26362;
assign n1275 = ~(n9076 | n704);
assign n26238 = n17396 & n19185;
assign n6978 = n25271 | n7566;
assign n27047 = n8764 & n5755;
assign n11585 = n631 & n12734;
assign n9658 = n21971 & n3640;
assign n26705 = ~(n9276 ^ n23199);
assign n21589 = n19488 | n2462;
assign n9735 = n18345 | n6179;
assign n19158 = ~(n16648 ^ n9602);
assign n14565 = n5611 & n20600;
assign n3936 = n18444 & n17028;
assign n5986 = ~(n17351 | n16468);
assign n14019 = n21543 | n3663;
assign n11923 = n20256 & n15567;
assign n5476 = n4020 | n4789;
assign n13566 = n5971 & n4742;
assign n1571 = ~n25736;
assign n4807 = ~(n15967 | n2783);
assign n4912 = n23225 | n3500;
assign n20756 = ~(n22442 ^ n3324);
assign n21854 = ~(n23974 ^ n24879);
assign n1226 = n13088 | n7674;
assign n24873 = ~(n5448 ^ n4026);
assign n3186 = ~(n10087 ^ n23534);
assign n13923 = ~(n11204 ^ n3806);
assign n22931 = n19616 | n8309;
assign n11925 = n9904 | n22921;
assign n11164 = n11369 & n17113;
assign n24550 = n17452 & n5683;
assign n14290 = n8216 & n10703;
assign n5307 = n21289 | n13418;
assign n21951 = ~n15023;
assign n16822 = ~n19184;
assign n4334 = ~(n1941 ^ n2659);
assign n16512 = ~(n1896 | n16396);
assign n26921 = ~(n24064 ^ n7764);
assign n15128 = ~(n20203 ^ n10705);
assign n17874 = n12321 & n21145;
assign n11506 = ~(n26987 ^ n23917);
assign n16107 = ~(n20423 ^ n13093);
assign n12489 = n13100 & n412;
assign n25239 = n13114 & n16641;
assign n2428 = ~(n14981 | n2718);
assign n9009 = n19298 | n22843;
assign n6624 = n26424 & n841;
assign n5864 = n21428 | n10550;
assign n17262 = n6396 | n22402;
assign n15669 = n371 | n25196;
assign n5033 = n7902 | n13926;
assign n19647 = n16762 & n1726;
assign n15019 = ~(n26485 ^ n14506);
assign n19072 = n3966 & n23077;
assign n5408 = ~(n5176 ^ n21771);
assign n378 = n16122 | n23050;
assign n2107 = n8536 & n13236;
assign n10498 = n26480 & n1546;
assign n9688 = n2060 | n6371;
assign n15516 = ~(n14790 ^ n604);
assign n13356 = ~(n17233 ^ n686);
assign n25898 = ~n5791;
assign n2191 = ~(n7409 ^ n21755);
assign n7368 = n20297 | n13603;
assign n7926 = n11144 | n23166;
assign n3847 = n22208 | n10902;
assign n3744 = ~n1696;
assign n25914 = ~n25240;
assign n8494 = n26582 | n7107;
assign n10020 = ~(n7785 ^ n1558);
assign n2452 = n3759 | n22682;
assign n5346 = n8611 & n10729;
assign n9852 = n14965 & n10389;
assign n20272 = n4033 | n8170;
assign n18687 = ~(n20585 ^ n21144);
assign n6680 = n155 & n22140;
assign n20703 = ~(n7678 ^ n11579);
assign n8486 = n26094 | n19735;
assign n26345 = n15901 | n21751;
assign n21597 = n6545 | n12271;
assign n22221 = n26207 & n6757;
assign n1131 = n8498 | n3656;
assign n15020 = n15880 | n10434;
assign n14014 = n6115 & n7385;
assign n3171 = n17287 & n16852;
assign n17038 = ~(n23307 ^ n13495);
assign n25742 = ~(n6356 | n1449);
assign n15534 = ~(n11940 ^ n9860);
assign n2605 = n5498 | n16886;
assign n22984 = n13513 | n5537;
assign n22574 = ~(n3468 ^ n15289);
assign n14390 = n17993 & n23145;
assign n25329 = n24245 | n3138;
assign n24763 = n16509 | n14945;
assign n22012 = ~n2489;
assign n6606 = ~(n6773 ^ n583);
assign n3777 = n23283 | n529;
assign n8830 = n12384 & n4667;
assign n20086 = n11131 | n21022;
assign n1995 = n21443 & n27014;
assign n18454 = ~(n8363 ^ n1222);
assign n15396 = n9961 | n15010;
assign n19796 = n2959 & n25493;
assign n11253 = n9951 & n19093;
assign n4570 = ~n8898;
assign n9280 = n26194 | n12299;
assign n3703 = n6304 | n14290;
assign n8617 = n18849 | n11066;
assign n4704 = n11993 & n8541;
assign n24383 = ~n21537;
assign n391 = ~(n6104 ^ n3945);
assign n3668 = ~(n19580 ^ n26829);
assign n3589 = ~(n189 | n5685);
assign n11412 = ~(n21232 ^ n2279);
assign n18947 = ~n16221;
assign n5343 = ~(n9114 ^ n27104);
assign n4112 = ~(n5048 ^ n25843);
assign n17188 = n4514 | n4122;
assign n3390 = ~(n22873 ^ n18760);
assign n25458 = ~(n8910 | n25018);
assign n9820 = ~n26573;
assign n15730 = ~n4587;
assign n19074 = ~n3618;
assign n2543 = n19429 | n14610;
assign n15191 = ~n5777;
assign n12953 = n25515 | n6949;
assign n9411 = n26255 & n14210;
assign n1093 = n10197 & n8800;
assign n15373 = ~(n3072 | n20145);
assign n842 = ~(n4923 | n14042);
assign n3466 = n20131 | n224;
assign n1952 = ~n1915;
assign n10080 = ~(n9598 ^ n7759);
assign n3284 = ~n8087;
assign n7641 = n15707 | n12174;
assign n5592 = n6616 & n17009;
assign n12958 = n6138 | n16965;
assign n23908 = n20768 | n25609;
assign n18073 = ~(n63 | n22359);
assign n8083 = ~n19210;
assign n19320 = n25534 & n5100;
assign n23402 = n19588 | n5211;
assign n20728 = ~(n10781 ^ n26512);
assign n27153 = ~(n8308 ^ n12522);
assign n14756 = n24300 & n21408;
assign n6517 = ~(n17212 ^ n16627);
assign n20649 = n20091 & n27050;
assign n19889 = n9292 & n14039;
assign n21073 = n6824 | n7624;
assign n10241 = ~(n25562 ^ n12216);
assign n25056 = n26878 | n6213;
assign n7244 = n3715 & n291;
assign n4746 = ~(n11382 ^ n20250);
assign n15760 = ~n11578;
assign n21327 = ~(n20826 | n18068);
assign n918 = n3276 & n13177;
assign n18336 = n20773 & n4750;
assign n23215 = ~(n4719 ^ n5822);
assign n8107 = n15364 | n10054;
assign n17248 = ~(n3306 | n21567);
assign n7677 = ~n18187;
assign n25617 = ~(n10678 ^ n25166);
assign n19863 = ~(n4317 ^ n22332);
assign n5434 = ~(n17902 | n20249);
assign n4210 = n20904 & n11573;
assign n2131 = ~(n1994 | n16559);
assign n25607 = ~(n4787 ^ n17405);
assign n7732 = n24827 | n297;
assign n23994 = n9948 | n308;
assign n6779 = ~n3603;
assign n6464 = ~n4410;
assign n9570 = ~n2783;
assign n10353 = ~n15305;
assign n19974 = ~(n20928 ^ n18315);
assign n1312 = n9038 & n13232;
assign n23649 = ~(n17902 ^ n337);
assign n17331 = n12341 & n13945;
assign n819 = ~(n14460 ^ n22026);
assign n14913 = ~(n19604 | n7359);
assign n412 = n11033 | n5699;
assign n10473 = n23016 | n25515;
assign n18343 = ~(n15270 ^ n11488);
assign n20402 = ~(n21901 ^ n5660);
assign n26137 = ~(n15271 ^ n12161);
assign n6679 = ~(n7978 ^ n10202);
assign n5052 = n20584 & n11795;
assign n15467 = n11143 | n8646;
assign n16648 = n1506 & n8039;
assign n8276 = ~(n8643 ^ n27168);
assign n15390 = n16385 & n25484;
assign n25325 = n22768 | n18915;
assign n13832 = ~(n13784 ^ n17302);
assign n10674 = n6332 & n12374;
assign n20690 = ~(n8526 ^ n17458);
assign n4506 = ~(n8647 ^ n18973);
assign n17424 = n22731 | n9087;
assign n14755 = n22925 | n13854;
assign n13046 = n8968 & n4126;
assign n4275 = ~(n3534 ^ n18756);
assign n23203 = ~(n19526 ^ n17863);
assign n11054 = ~(n788 ^ n16573);
assign n23706 = n3481 & n14054;
assign n12186 = ~(n12366 ^ n11736);
assign n8840 = ~(n25413 | n152);
assign n13534 = ~n24600;
assign n19736 = ~(n24190 ^ n20804);
assign n18757 = n25740 | n12045;
assign n7497 = ~(n10682 ^ n10234);
assign n19377 = ~(n5198 ^ n25501);
assign n12576 = ~n25345;
assign n23796 = ~(n18113 ^ n1467);
assign n22565 = n14685 | n13282;
assign n22409 = n25020 | n24385;
assign n12284 = n21462 | n19872;
assign n11838 = ~(n5405 ^ n23834);
assign n20291 = ~(n19665 ^ n10065);
assign n20983 = n16324 | n23688;
assign n17426 = n7068 & n2353;
assign n1225 = ~(n6471 ^ n10448);
assign n7780 = ~(n4968 ^ n500);
assign n1706 = ~(n11615 | n23779);
assign n21067 = ~(n13708 ^ n23775);
assign n17601 = ~n13367;
assign n3543 = ~(n7092 ^ n24486);
assign n18003 = ~(n20587 ^ n16457);
assign n15819 = n21605 | n21898;
assign n4646 = ~(n11833 ^ n4019);
assign n15445 = ~n4372;
assign n14207 = n1736 & n12243;
assign n21716 = n6204 & n23254;
assign n16096 = n16084 | n9557;
assign n2717 = n26382 & n1217;
assign n14580 = ~(n9892 ^ n23911);
assign n2498 = ~n18003;
assign n10808 = n23469 | n17666;
assign n26181 = n19710 & n7965;
assign n18289 = n22018 & n5979;
assign n14519 = ~n2547;
assign n16637 = ~n22537;
assign n26222 = ~(n15592 ^ n25009);
assign n19052 = n25004 | n1630;
assign n22747 = n25437 & n15098;
assign n22599 = ~(n2659 | n11926);
assign n17488 = n8851 & n4087;
assign n24792 = n1956 | n3877;
assign n17500 = ~(n24413 ^ n11054);
assign n23544 = ~(n6541 ^ n329);
assign n23030 = ~n8869;
assign n22810 = n7194 | n12180;
assign n14493 = ~(n26222 ^ n6944);
assign n20868 = ~(n1465 ^ n23304);
assign n17873 = ~(n11266 ^ n9926);
assign n26471 = ~n11910;
assign n2158 = n9870 & n4171;
assign n13221 = n14863 & n16578;
assign n5739 = ~(n11012 ^ n20118);
assign n1055 = ~(n15776 ^ n14009);
assign n20313 = n5475 | n3834;
assign n491 = n26116 | n1497;
assign n7309 = n10601 | n5845;
assign n12193 = n2257 | n21666;
assign n15944 = ~n1667;
assign n11933 = ~(n20434 ^ n3692);
assign n7365 = ~n1386;
assign n1509 = ~(n25565 ^ n21993);
assign n16239 = ~(n17048 ^ n22624);
assign n11556 = ~(n14397 ^ n16812);
assign n18598 = ~n4256;
assign n2773 = n4858 & n6895;
assign n17365 = ~(n1881 | n26857);
assign n4098 = n7991 & n4805;
assign n25516 = ~(n20548 ^ n4813);
assign n19540 = ~(n18076 ^ n19920);
assign n22930 = n24650 & n23729;
assign n26970 = ~(n22678 ^ n783);
assign n4530 = ~(n18295 | n23313);
assign n1538 = n22978 | n15228;
assign n14928 = n11477 | n22207;
assign n1100 = n11598 & n10042;
assign n23115 = n22105 | n5465;
assign n11740 = ~n647;
assign n11173 = n19883 & n21468;
assign n12855 = ~n20663;
assign n11127 = ~(n18648 ^ n23782);
assign n21291 = ~(n26130 ^ n16909);
assign n10403 = n18642 & n1899;
assign n411 = n19393 | n16982;
assign n15218 = ~n20950;
assign n13641 = ~(n22511 | n10251);
assign n20296 = n7343 | n11108;
assign n12825 = ~(n23476 | n12410);
assign n5498 = ~n12650;
assign n3402 = ~(n10250 | n13976);
assign n20038 = n16133 | n10675;
assign n1699 = n24 | n2876;
assign n12414 = n5942 & n7023;
assign n20442 = ~(n9462 ^ n17251);
assign n13574 = n11417 | n19700;
assign n26983 = n6186 | n2134;
assign n17761 = n12784 | n12887;
assign n10354 = ~(n16822 ^ n14661);
assign n9187 = ~n1350;
assign n21656 = n17473 & n24463;
assign n3335 = ~(n4859 | n2570);
assign n26278 = n6720 & n5396;
assign n10392 = n4239 ^ n11034;
assign n9281 = n4752 | n13114;
assign n14646 = ~(n25900 | n12697);
assign n6962 = ~n23253;
assign n8995 = n16186 | n2643;
assign n11773 = n24535 | n20052;
assign n19998 = n12760 | n20295;
assign n13229 = n10831 | n18500;
assign n19633 = ~n19309;
assign n13482 = n21057 | n13742;
assign n1560 = ~(n25637 ^ n19540);
assign n13995 = ~n5517;
assign n21575 = ~n13336;
assign n3943 = n19952 & n10178;
assign n10389 = ~n2599;
assign n14239 = n9494 | n21723;
assign n20993 = ~(n17549 | n20506);
assign n15144 = ~n23692;
assign n26252 = ~n11650;
assign n26386 = ~(n8391 ^ n23200);
assign n469 = n11303 | n10037;
assign n20148 = ~(n7769 ^ n26625);
assign n7713 = ~n25670;
assign n11015 = n19705 | n16021;
assign n12788 = ~n4160;
assign n5898 = ~(n14254 | n11502);
assign n14468 = ~(n17938 ^ n20966);
assign n18769 = n19165 & n41;
assign n21220 = n20643 | n12082;
assign n15971 = n5494 | n1487;
assign n15169 = n7007 & n8699;
assign n16986 = n24608 | n26016;
assign n9353 = n10597 | n10126;
assign n24940 = ~n5305;
assign n10495 = ~(n16349 | n604);
assign n7587 = ~(n22274 ^ n24129);
assign n15590 = ~(n25154 ^ n12323);
assign n15160 = ~(n12650 ^ n11220);
assign n204 = n6251 & n5092;
assign n6350 = n5205 | n6065;
assign n20555 = n7612 | n20883;
assign n18347 = ~(n20929 ^ n23068);
assign n350 = ~n22154;
assign n11080 = ~(n19823 ^ n2611);
assign n1021 = n26747 | n7923;
assign n5267 = n14826 & n20342;
assign n1442 = n26513 | n20902;
assign n15028 = n12125 | n7828;
assign n3692 = ~(n7809 ^ n25100);
assign n18080 = n23775 | n4601;
assign n10058 = n26140 | n843;
assign n25667 = ~(n8541 ^ n12826);
assign n19949 = ~n2659;
assign n6731 = ~n23602;
assign n23900 = ~(n4439 ^ n15281);
assign n22480 = ~(n15388 ^ n8046);
assign n1887 = ~(n27104 ^ n18295);
assign n6698 = ~n3937;
assign n8096 = n9514 | n17204;
assign n8403 = ~(n27107 ^ n7518);
assign n1516 = ~(n9017 ^ n25647);
assign n24770 = n6024 | n24334;
assign n5531 = ~(n4938 | n14130);
assign n14893 = n10805 & n247;
assign n16718 = n8101 & n3019;
assign n1402 = n15918 & n21021;
assign n20201 = ~(n16721 ^ n19941);
assign n9568 = n443 | n4797;
assign n18906 = ~(n2952 ^ n1639);
assign n24322 = ~(n15856 | n14357);
assign n14305 = ~(n182 ^ n15190);
assign n1044 = ~(n7965 ^ n6290);
assign n16730 = n1406 & n19473;
assign n9448 = ~(n16357 ^ n16880);
assign n9998 = n15365 & n1973;
assign n4107 = n4600 | n2264;
assign n800 = ~(n2995 ^ n18281);
assign n4840 = n12513 & n14106;
assign n9132 = n13985 | n12155;
assign n4308 = n18051 & n8124;
assign n2737 = n2895 | n16972;
assign n807 = ~(n11650 ^ n7750);
assign n21845 = ~(n2559 | n2117);
assign n12477 = ~n8649;
assign n23225 = ~(n2659 | n23704);
assign n20451 = n23413 | n14491;
assign n15197 = n16192 | n19795;
assign n17669 = n13876 & n9582;
assign n26229 = ~(n13585 ^ n9051);
assign n13686 = n22585 | n22527;
assign n8871 = ~(n17388 ^ n4242);
assign n3788 = n8571 | n11285;
assign n1268 = n26986 | n16832;
assign n26326 = ~n23851;
assign n21314 = n21380 | n16210;
assign n22594 = ~(n22895 | n17845);
assign n1970 = ~(n10057 ^ n8920);
assign n17898 = ~(n16267 ^ n9240);
assign n3038 = ~(n7082 ^ n21782);
assign n17588 = ~(n3734 | n14257);
assign n2262 = n17166 | n25989;
assign n22532 = n25135 & n20136;
assign n13741 = n24683 & n25801;
assign n2075 = n26772 & n15718;
assign n21356 = n25320 | n18836;
assign n2529 = n22041 & n5099;
assign n21850 = ~(n25117 ^ n25629);
assign n9612 = ~(n20132 | n2810);
assign n20457 = n748 & n7070;
assign n17583 = ~(n17324 ^ n23875);
assign n7515 = ~(n10275 ^ n25240);
assign n10993 = ~n13463;
assign n6212 = ~(n22607 | n15512);
assign n3997 = n13099 | n17545;
assign n12933 = ~(n15109 | n5532);
assign n24714 = ~(n16432 ^ n1667);
assign n16305 = ~(n15007 ^ n12281);
assign n4180 = ~(n1449 ^ n6356);
assign n13082 = ~(n10940 ^ n2240);
assign n9826 = ~n17970;
assign n12566 = ~(n11872 ^ n2532);
assign n20494 = ~(n5077 ^ n13914);
assign n27181 = ~(n11982 ^ n7931);
assign n9213 = ~(n19393 ^ n16982);
assign n16781 = ~(n16722 | n21101);
assign n11274 = ~(n12398 ^ n25694);
assign n12456 = n311 & n12721;
assign n9345 = ~(n14276 ^ n18035);
assign n26837 = n22176 | n10666;
assign n24570 = n16879 | n24235;
assign n7675 = n24325 | n23913;
assign n5457 = n7261 | n26601;
assign n12999 = ~(n11908 ^ n24538);
assign n12287 = ~(n8687 | n966);
assign n8056 = ~(n22436 | n11146);
assign n5901 = n21152 & n25496;
assign n23193 = n7279 & n23378;
assign n19251 = n3536 | n3109;
assign n14483 = n3116 | n16696;
assign n8870 = n15134 | n5179;
assign n9540 = ~(n23528 | n9099);
assign n25401 = n6581 | n17781;
assign n7442 = n7311 | n19944;
assign n6300 = ~n19524;
assign n26454 = ~(n2057 ^ n19603);
assign n18288 = ~(n25662 ^ n1482);
assign n20885 = n21741 & n6926;
assign n17685 = ~n11892;
assign n24489 = n23030 | n6385;
assign n16398 = ~(n22726 ^ n16451);
assign n6689 = ~(n26178 | n21290);
assign n20217 = n9518 & n14509;
assign n6466 = ~n3038;
assign n16426 = ~(n24630 ^ n6775);
assign n5501 = ~(n20796 | n21460);
assign n13454 = n15875 & n13352;
assign n18468 = n23195 & n8666;
assign n21404 = ~(n22437 ^ n5788);
assign n22437 = n5323 & n22258;
assign n24653 = n20260 | n18205;
assign n14999 = ~(n18607 ^ n22159);
assign n19617 = ~(n1068 ^ n7608);
assign n20716 = ~n18398;
assign n7877 = n4801 | n11970;
assign n12530 = ~n23035;
assign n17449 = ~(n16319 | n6293);
assign n22503 = ~(n12889 ^ n24298);
assign n10456 = ~(n3750 | n24397);
assign n17574 = n883 | n5452;
assign n6421 = ~(n3069 | n15289);
assign n10437 = ~(n21515 ^ n25000);
assign n25733 = ~(n9969 | n14705);
assign n8377 = n2192 | n12897;
assign n15471 = n486 & n18042;
assign n10369 = ~n17256;
assign n2960 = ~n14981;
assign n4531 = ~n24578;
assign n3887 = n26908 & n21552;
assign n15165 = ~(n12260 ^ n20997);
assign n14495 = n20841 | n13528;
assign n2766 = ~(n24608 | n428);
assign n21686 = ~(n21004 | n18265);
assign n10476 = n17596 | n22469;
assign n9228 = ~(n11749 ^ n14954);
assign n7739 = n22091 | n18861;
assign n8166 = ~(n10727 ^ n20932);
assign n13636 = n11521 | n22735;
assign n24082 = n13605 | n16365;
assign n8234 = ~(n12430 ^ n17780);
assign n12300 = ~(n20384 ^ n6659);
assign n7285 = ~(n24930 ^ n15515);
assign n16646 = n20572 | n21877;
assign n24139 = ~(n21222 ^ n26752);
assign n16724 = ~(n20816 ^ n6772);
assign n22636 = ~n15600;
assign n2747 = ~(n7164 ^ n17193);
assign n8009 = n18261 & n6413;
assign n3745 = ~(n26553 | n15041);
assign n2065 = ~(n1433 ^ n26344);
assign n6754 = n3130 | n5983;
assign n21406 = ~n13297;
assign n19481 = n16477 | n11697;
assign n22079 = ~(n25865 ^ n4403);
assign n19799 = n26162 | n6814;
assign n11822 = ~(n16702 ^ n7793);
assign n6360 = n7180 & n3333;
assign n12426 = ~(n7200 ^ n19307);
assign n26577 = n8493 & n865;
assign n6451 = ~(n25629 | n3795);
assign n14457 = ~(n940 ^ n17694);
assign n14129 = ~(n25376 | n18617);
assign n21705 = ~(n23068 ^ n18907);
assign n3316 = ~(n5083 ^ n4640);
assign n7173 = n23850 & n9101;
assign n6940 = n1406 & n1978;
assign n6500 = ~(n8773 ^ n18599);
assign n6617 = ~(n7260 | n13368);
assign n16095 = n4216 & n24069;
assign n12295 = ~(n23967 ^ n17251);
assign n13355 = n9284 | n25683;
assign n14668 = ~(n350 ^ n18004);
assign n8145 = n7772 | n10671;
assign n22346 = ~(n7963 | n6590);
assign n11469 = ~(n8224 ^ n20151);
assign n24389 = n5427 & n19633;
assign n24452 = ~(n10666 ^ n8656);
assign n21382 = n15530 | n2739;
assign n23094 = ~n13240;
assign n24046 = n14861 | n24697;
assign n11441 = n19962 | n22426;
assign n9417 = n9944 | n23842;
assign n4894 = n15442 & n18450;
assign n23617 = ~(n10593 | n4792);
assign n10604 = n2628 | n14345;
assign n9923 = n6841 & n4036;
assign n13964 = n23923 | n16608;
assign n25701 = ~n1869;
assign n24232 = n6574 | n14351;
assign n18209 = n21140 & n10241;
assign n25626 = n1089 | n5094;
assign n16428 = ~(n3034 ^ n16207);
assign n16753 = ~(n20326 ^ n5916);
assign n26071 = n20829 | n18171;
assign n10436 = ~(n24305 | n5012);
assign n23686 = ~n1047;
assign n16389 = ~(n6692 | n21249);
assign n11369 = n3078 | n15698;
assign n25772 = n11957 | n3873;
assign n11447 = ~(n7330 ^ n8439);
assign n10075 = ~n23310;
assign n18309 = n2230 | n16722;
assign n5956 = ~(n19893 ^ n15171);
assign n7632 = ~(n18398 | n25807);
assign n24959 = ~n1550;
assign n22382 = ~n18726;
assign n9115 = n3111 & n19671;
assign n16174 = ~(n11089 ^ n972);
assign n19101 = n13966 & n17441;
assign n10774 = ~(n15389 ^ n24468);
assign n21488 = ~(n3136 ^ n26913);
assign n26876 = n7634;
assign n11145 = ~(n1612 | n728);
assign n8779 = ~n26888;
assign n22802 = ~(n18880 | n2978);
assign n2177 = ~(n20192 ^ n21649);
assign n22050 = ~(n21821 ^ n10257);
assign n6478 = n3817 | n8761;
assign n26816 = ~(n14880 ^ n8210);
assign n5584 = ~(n16439 ^ n10275);
assign n19783 = ~(n8721 ^ n1040);
assign n4419 = n14514 | n26187;
assign n13486 = ~(n8726 ^ n24911);
assign n5292 = n2597 & n10682;
assign n23106 = n13675 & n12010;
assign n1247 = n3404 & n11943;
assign n16009 = ~(n14313 ^ n25180);
assign n26613 = n19429 & n23519;
assign n9604 = n5154 | n4138;
assign n4082 = n17878 & n7920;
assign n8139 = ~(n18250 ^ n7235);
assign n20536 = ~n25464;
assign n9124 = ~(n14558 ^ n12479);
assign n5247 = ~(n20948 ^ n1658);
assign n18356 = n7715 & n19528;
assign n3789 = ~(n1831 ^ n3320);
assign n2528 = ~(n6082 ^ n3228);
assign n4050 = ~n763;
assign n7253 = ~(n16750 ^ n20819);
assign n5651 = ~(n2858 | n26486);
assign n15179 = ~(n67 ^ n11494);
assign n4169 = n14628 | n16846;
assign n15518 = n23356 & n17801;
assign n199 = n3035 & n24997;
assign n2930 = ~(n8220 | n7361);
assign n15671 = ~(n19614 ^ n21222);
assign n17468 = n11666 & n17750;
assign n6654 = n8565 & n16363;
assign n6223 = ~(n22065 ^ n17865);
assign n14848 = ~n26016;
assign n17508 = ~(n3719 ^ n25119);
assign n25945 = n18560 | n2958;
assign n7245 = ~(n19849 | n18421);
assign n13288 = n2632 & n7368;
assign n6593 = ~(n27037 ^ n23913);
assign n15385 = ~n11769;
assign n7226 = n1577 & n22885;
assign n2607 = ~n11333;
assign n740 = ~(n11220 | n3425);
assign n16925 = ~(n22964 ^ n21060);
assign n18186 = n3591 | n3963;
assign n20722 = ~(n24054 ^ n10723);
assign n17199 = n25329 & n12676;
assign n17186 = ~(n8857 ^ n19578);
assign n11169 = ~(n26912 ^ n12895);
assign n21748 = n6318 & n96;
assign n11675 = n23910 & n21339;
assign n8369 = n2318 | n19038;
assign n4951 = ~(n26000 | n14725);
assign n14296 = n7206 & n6530;
assign n1393 = n18829 | n27090;
assign n23918 = ~(n15113 ^ n21957);
assign n6687 = n13577 | n26691;
assign n4794 = ~(n6104 ^ n24048);
assign n23823 = ~(n1451 ^ n16217);
assign n18887 = ~(n5646 ^ n2367);
assign n18958 = ~(n8244 ^ n6513);
assign n7009 = n1365 | n12315;
assign n23129 = n2331 & n13748;
assign n490 = n24653 | n10746;
assign n9602 = ~(n16707 ^ n13037);
assign n23167 = n6614 & n21305;
assign n15375 = ~(n3919 | n26105);
assign n7972 = n10657 & n1440;
assign n11975 = ~n26069;
assign n16028 = ~n24070;
assign n20833 = n8348 | n12625;
assign n5792 = n22401 & n17594;
assign n24498 = n24729 | n1846;
assign n25276 = ~n5727;
assign n645 = ~(n15930 ^ n14089);
assign n20515 = ~(n24312 ^ n5032);
assign n9582 = n2617 | n13911;
assign n23677 = ~(n25007 ^ n14083);
assign n1912 = ~(n22562 | n17412);
assign n13118 = n7292 | n14510;
assign n12138 = ~n24112;
assign n18180 = n18431 | n11295;
assign n6815 = n7692 & n16793;
assign n15741 = n25744 | n15218;
assign n15143 = n16827 & n7262;
assign n18110 = n1192 | n5569;
assign n24766 = ~n15440;
assign n5816 = ~n6611;
assign n25283 = ~(n20384 | n8008);
assign n12865 = n3820 & n3684;
assign n19104 = ~(n6990 ^ n26449);
assign n19810 = n7424 | n4052;
assign n22682 = ~(n14302 | n12837);
assign n21217 = n21846 | n24161;
assign n16904 = ~(n3472 | n25085);
assign n26182 = n11691 | n11073;
assign n10128 = ~n8387;
assign n16147 = ~n12241;
assign n15474 = ~n22270;
assign n13409 = ~(n10106 ^ n26072);
assign n24276 = ~(n4490 | n5261);
assign n11739 = ~(n11011 ^ n20179);
assign n11315 = ~(n5060 | n2808);
assign n2765 = ~(n22318 ^ n21626);
assign n9798 = n9003 | n1735;
assign n12918 = ~(n8008 | n14516);
assign n20726 = ~(n2160 ^ n11220);
assign n6602 = ~(n9666 ^ n6747);
assign n12402 = ~n12648;
assign n15533 = n21517 | n8582;
assign n630 = n22174 & n22277;
assign n13451 = ~n11792;
assign n24678 = n21016 | n21668;
assign n21960 = ~(n855 ^ n12234);
assign n21995 = n15850 & n22206;
assign n1847 = n7242 & n16123;
assign n1066 = ~(n14678 ^ n10938);
assign n18143 = ~(n18222 ^ n26518);
assign n23877 = ~n7134;
assign n5298 = ~(n5226 | n26724);
assign n13701 = n20169 | n8718;
assign n17550 = n13036 & n23307;
assign n22558 = ~n10201;
assign n24193 = ~(n17542 | n15146);
assign n9158 = n1715 | n15490;
assign n9073 = ~(n20032 | n4844);
assign n1407 = n11559 | n22861;
assign n13168 = ~(n22555 ^ n16287);
assign n6305 = n10519 & n11310;
assign n4386 = n11745 | n18249;
assign n19308 = ~(n9701 ^ n6076);
assign n11407 = ~(n20986 ^ n25471);
assign n5796 = ~n1204;
assign n21214 = n10264 & n21039;
assign n11314 = ~(n14689 ^ n20179);
assign n18714 = ~(n1337 ^ n26073);
assign n9722 = n8447 | n26254;
assign n3534 = n4493 | n768;
assign n23798 = ~n8769;
assign n18441 = n19827 | n17297;
assign n24266 = ~(n20041 ^ n7257);
assign n20839 = ~(n11649 ^ n9872);
assign n22613 = ~n2698;
assign n19278 = n5511 | n12270;
assign n12543 = ~n20658;
assign n5838 = ~(n9180 | n1262);
assign n20309 = n12841 | n16361;
assign n23554 = ~(n12561 | n11305);
assign n21837 = n3346 | n19311;
assign n10917 = ~(n2088 ^ n26979);
assign n15309 = ~n15127;
assign n26663 = n11292 & n3146;
assign n5039 = ~n11408;
assign n14694 = ~(n26452 ^ n5098);
assign n24999 = n10536 & n17650;
assign n21815 = n9770 | n26100;
assign n21669 = n11043 | n1252;
assign n16463 = n4910 & n1638;
assign n9861 = n7967 | n19154;
assign n23447 = n25822 & n13047;
assign n6774 = ~(n16726 ^ n20068);
assign n4302 = n25651 | n5921;
assign n2771 = ~(n22207 ^ n26851);
assign n1034 = ~(n21249 ^ n6692);
assign n955 = n1426 & n10105;
assign n25913 = n24565 & n3729;
assign n8882 = n7617 | n23706;
assign n6599 = ~n2730;
assign n11929 = ~(n13250 ^ n10685);
assign n1037 = ~(n22370 | n6034);
assign n21043 = n1643 | n20460;
assign n12037 = n22532 | n2260;
assign n8295 = ~n9313;
assign n26328 = n10558 & n18832;
assign n11832 = ~(n20099 ^ n3541);
assign n14602 = n1146 & n8469;
assign n13421 = ~(n17660 ^ n19758);
assign n15582 = ~n11448;
assign n3419 = ~(n15572 | n2989);
assign n10262 = ~(n47 ^ n12230);
assign n8777 = n18345 & n6179;
assign n6614 = n6321 | n5026;
assign n1713 = n13863 | n20134;
assign n5919 = ~(n22422 | n18648);
assign n23608 = ~n14984;
assign n11319 = n19380 & n13134;
assign n11049 = n25004 | n10158;
assign n25268 = ~n26000;
assign n5316 = ~(n1765 | n21309);
assign n2599 = ~(n11636 ^ n23673);
assign n23415 = ~n2778;
assign n25582 = ~n1872;
assign n26682 = n26914 | n26962;
assign n22711 = ~(n2729 ^ n9210);
assign n8247 = n26567 & n9385;
assign n1413 = ~(n9745 ^ n14900);
assign n3085 = ~(n7088 | n3132);
assign n18333 = ~(n2310 ^ n16769);
assign n20782 = ~(n19313 | n5974);
assign n25100 = ~(n16505 ^ n10080);
assign n7264 = n13419 | n14937;
assign n6933 = n15201 & n22705;
assign n5312 = n6790 | n10000;
assign n25076 = ~(n10083 ^ n13654);
assign n13158 = ~(n19295 ^ n22631);
assign n2043 = ~(n10109 ^ n26742);
assign n1150 = n533 & n24858;
assign n18017 = n18548 | n12239;
assign n26001 = ~(n25674 ^ n5585);
assign n10793 = ~(n18806 ^ n14518);
assign n5833 = ~(n16121 ^ n7366);
assign n3409 = ~(n21871 | n1314);
assign n10516 = ~(n23200 ^ n19116);
assign n22248 = n8910 | n22392;
assign n21147 = n22329 | n26369;
assign n20713 = ~(n15774 ^ n13947);
assign n13011 = n10514 | n24806;
assign n5924 = n9054;
assign n7007 = n13621 | n10114;
assign n15204 = ~n11824;
assign n11053 = ~(n17430 ^ n24311);
assign n18004 = ~n21636;
assign n5454 = n1398 ^ n9507;
assign n25875 = n19514 & n2415;
assign n1759 = ~n2189;
assign n10238 = n14285 & n2934;
assign n12050 = ~(n4742 ^ n870);
assign n24941 = n26643 & n383;
assign n19002 = n7126 & n24120;
assign n18034 = ~(n21222 ^ n26565);
assign n3487 = n17198 | n23882;
assign n18948 = n21437 | n3242;
assign n8699 = n21790 | n18815;
assign n21436 = ~n5462;
assign n14822 = n25237 | n21710;
assign n10588 = n11638 | n18382;
assign n16786 = ~(n25749 ^ n2113);
assign n4999 = ~(n21394 ^ n894);
assign n18845 = n25752 | n8173;
assign n15266 = ~n10658;
assign n26279 = n15229 | n20029;
assign n11553 = n17757 | n1150;
assign n25806 = n17368 & n2539;
assign n8650 = ~n17326;
assign n15311 = ~(n11559 | n2328);
assign n15407 = ~(n23928 ^ n8692);
assign n21435 = ~(n144 | n10710);
assign n10932 = n23736 | n8702;
assign n15887 = ~(n11898 | n23166);
assign n25424 = ~(n15766 | n6105);
assign n8082 = ~(n26961 | n864);
assign n11232 = ~(n6387 | n455);
assign n16302 = n17211 | n4345;
assign n16552 = n26279 & n23902;
assign n10221 = n9802 | n10017;
assign n9350 = ~(n8319 ^ n12493);
assign n3002 = ~(n2622 ^ n19500);
assign n3049 = ~(n8128 ^ n23766);
assign n11665 = ~(n8513 | n10709);
assign n23382 = n16698 | n26881;
assign n6781 = n2517 | n9194;
assign n1029 = n13293 & n17388;
assign n23794 = n10193 | n4755;
assign n1250 = ~(n13989 | n20138);
assign n18798 = ~n618;
assign n18931 = ~n25538;
assign n13274 = n17784 & n725;
assign n4865 = ~(n25115 ^ n22491);
assign n13615 = n14886 & n17639;
assign n11850 = n21855 & n13395;
assign n21665 = ~(n17242 ^ n24926);
assign n15212 = n1365 | n4087;
assign n1977 = n14431 | n8906;
assign n9712 = ~(n5719 | n7195);
assign n417 = ~n25289;
assign n24735 = n26380 & n18974;
assign n20941 = ~(n2462 ^ n19488);
assign n12851 = ~(n24069 ^ n13684);
assign n8393 = n24524 | n4069;
assign n11821 = n15682 | n4080;
assign n22125 = ~n26399;
assign n3321 = n26563 & n10809;
assign n16522 = ~(n26211 ^ n21219);
assign n21558 = n602 | n16963;
assign n19015 = ~(n16547 ^ n4085);
assign n8710 = n4285 | n16119;
assign n12274 = n21370 & n16083;
assign n8990 = n11745 & n6825;
assign n5156 = ~(n25377 ^ n16482);
assign n97 = ~(n11802 ^ n11502);
assign n19161 = n21541 & n16177;
assign n10062 = n22286 | n199;
assign n8612 = ~n23745;
assign n9890 = n13918 & n21595;
assign n25082 = ~(n14588 | n942);
assign n657 = ~(n10758 ^ n13562);
assign n18422 = n17550 | n14022;
assign n19301 = ~(n24898 ^ n22861);
assign n14354 = ~(n23616 ^ n18444);
assign n23060 = ~(n15135 ^ n18204);
assign n11608 = ~n14756;
assign n3763 = n3796 | n4416;
assign n150 = ~(n18066 ^ n20111);
assign n10740 = ~(n12366 | n23071);
assign n14410 = ~n3132;
assign n9174 = n378 | n5779;
assign n5564 = ~(n22011 ^ n17042);
assign n22330 = n11761 & n23496;
assign n20550 = ~n9625;
assign n19300 = n8504 | n24400;
assign n4427 = n11583 | n3190;
assign n1417 = n16748 | n14959;
assign n24049 = ~(n12543 ^ n15508);
assign n26188 = ~(n9240 | n16267);
assign n22313 = ~(n8367 | n2113);
assign n15801 = ~(n21478 ^ n833);
assign n7754 = ~(n23486 ^ n11734);
assign n656 = ~n9906;
assign n10340 = ~(n21690 ^ n9409);
assign n8658 = n3945 & n21998;
assign n15778 = n11322 | n26098;
assign n26200 = n10117 | n19825;
assign n11966 = n2926 | n25520;
assign n18516 = n4957 & n14979;
assign n13867 = n10877 & n8560;
assign n14669 = ~(n6262 ^ n11258);
assign n17530 = ~(n8816 ^ n21679);
assign n6264 = n19393 & n16982;
assign n16734 = ~(n20043 ^ n11071);
assign n10525 = n5631 | n13381;
assign n12629 = n6743 ^ n7713;
assign n5034 = n7524 | n8799;
assign n1458 = ~n20077;
assign n21768 = ~(n11716 ^ n12775);
assign n3075 = ~(n19656 ^ n16456);
assign n21204 = n9921 | n2736;
assign n18419 = ~(n3744 | n12248);
assign n6848 = ~(n18052 ^ n16073);
assign n17887 = ~(n1340 | n1099);
assign n19606 = n9127 & n8390;
assign n26632 = n10274 | n14168;
assign n13728 = n9701 & n6076;
assign n18626 = ~(n18171 ^ n1738);
assign n9515 = n21406 | n10034;
assign n16191 = n22369 & n11358;
assign n1146 = n13775 | n8389;
assign n11796 = n9942 | n2210;
assign n17482 = n17543 | n10445;
assign n26190 = n635 | n22415;
assign n17423 = ~n23895;
assign n9439 = n22585 & n26837;
assign n3835 = ~(n2859 ^ n608);
assign n27131 = ~(n19196 | n6122);
assign n3350 = n7778 | n4083;
assign n22910 = ~(n14105 ^ n1001);
assign n12454 = ~n8363;
assign n7274 = n22554 | n21890;
assign n11185 = ~(n1998 ^ n13230);
assign n18989 = n12715 | n10303;
assign n845 = n10990 | n2834;
assign n6531 = n795 & n10857;
assign n2589 = n246 | n8763;
assign n12844 = ~(n21380 | n24170);
assign n4720 = ~(n8236 | n728);
assign n17136 = n8244 | n8431;
assign n3141 = ~(n11697 ^ n19711);
assign n22753 = ~(n16401 ^ n9259);
assign n16621 = n7949 | n15562;
assign n4355 = n25432 | n21447;
assign n10598 = ~(n15268 | n333);
assign n21928 = ~n7710;
assign n2231 = ~n20631;
assign n12909 = n4342 | n9401;
assign n17481 = ~(n15693 ^ n24701);
assign n15312 = n16164 & n14221;
assign n7723 = n12965 | n17571;
assign n24753 = n20486 | n22556;
assign n18620 = n11087 | n16437;
assign n15322 = ~(n5822 ^ n7963);
assign n17201 = ~(n5055 ^ n3827);
assign n10152 = ~n16576;
assign n3046 = ~(n167 | n1339);
assign n22419 = n21125 | n926;
assign n21685 = ~(n14893 ^ n15919);
assign n3529 = n21644 & n18555;
assign n19725 = ~(n2109 ^ n963);
assign n17995 = ~n13189;
assign n22051 = n14963 | n10620;
assign n13059 = n16762 | n22662;
assign n950 = ~n1608;
assign n9221 = n4983 & n24045;
assign n25071 = ~n7212;
assign n20921 = ~n3839;
assign n19497 = ~(n16364 ^ n18891);
assign n26559 = n1558 | n17305;
assign n902 = ~(n14465 | n25074);
assign n10672 = ~(n23277 ^ n11975);
assign n22360 = ~(n12554 | n22871);
assign n22849 = ~n10096;
assign n499 = n19760 | n19994;
assign n17949 = n24705 & n26444;
assign n19183 = n21052 | n21576;
assign n19186 = ~n11945;
assign n20093 = n8202 | n14209;
assign n4728 = n7238 & n14923;
assign n24648 = ~(n17556 ^ n6896);
assign n1815 = n13951 & n24355;
assign n1693 = ~(n18649 ^ n3984);
assign n7820 = ~(n25289 ^ n4195);
assign n14904 = ~(n16722 | n13708);
assign n26322 = ~(n13333 | n15681);
assign n1209 = n16166 & n10407;
assign n11221 = ~(n17433 ^ n15574);
assign n13248 = n21462 & n19872;
assign n22343 = n5867 | n11930;
assign n9245 = ~(n14581 ^ n19187);
assign n22045 = n6992 & n2824;
assign n9548 = n11294 | n20608;
assign n2574 = ~(n8452 ^ n3141);
assign n18279 = ~n14061;
assign n13242 = n23886 | n13245;
assign n23959 = ~(n23589 ^ n12891);
assign n22008 = n17144 & n15641;
assign n11013 = ~n11651;
assign n16762 = ~n5048;
assign n18689 = ~(n22110 ^ n11378);
assign n20741 = n19878 & n20888;
assign n10863 = ~(n11381 | n4294);
assign n15753 = ~(n1118 ^ n4665);
assign n12744 = ~(n5425 ^ n1081);
assign n8352 = ~(n7482 ^ n16382);
assign n26323 = ~(n26580 ^ n13485);
assign n18856 = n9901 | n13447;
assign n10707 = ~(n20826 | n626);
assign n26294 = n20023 & n12734;
assign n19086 = n18811 & n21330;
assign n8176 = ~n23892;
assign n12418 = ~n24863;
assign n7059 = ~n20029;
assign n13399 = n338 & n10806;
assign n13871 = n6819 | n11671;
assign n16679 = ~n13425;
assign n8121 = n10527 | n5387;
assign n11543 = n19256 & n16941;
assign n21706 = n22042 | n6808;
assign n5908 = ~(n4149 | n22454);
assign n15121 = ~(n1222 | n8292);
assign n7088 = ~n21957;
assign n1020 = ~(n23633 ^ n24284);
assign n13723 = n2069 & n25315;
assign n15692 = n20614 & n8141;
assign n12979 = n20064 | n14345;
assign n9291 = n22002;
assign n12998 = ~(n12198 ^ n10405);
assign n9977 = n13844 | n19394;
assign n17531 = n24004 & n21081;
assign n13381 = n18191 & n18188;
assign n5081 = ~(n25738 ^ n6861);
assign n9772 = n12455 | n974;
assign n17852 = ~(n23568 ^ n27120);
assign n6208 = n10786 & n22922;
assign n14013 = n8244 | n22820;
assign n23077 = n191 | n18072;
assign n2811 = ~(n25872 | n2994);
assign n15581 = ~n15918;
assign n252 = ~(n26728 ^ n25655);
assign n19121 = ~(n17911 ^ n6814);
assign n16916 = n4999 | n27017;
assign n12952 = ~(n9249 | n14732);
assign n17445 = ~(n21843 | n20659);
assign n792 = n5710 & n4439;
assign n21370 = ~n22516;
assign n22836 = ~n9656;
assign n9995 = n11045 | n11220;
assign n11731 = ~(n9392 | n12049);
assign n24717 = ~n24764;
assign n13308 = ~n2964;
assign n19895 = ~n6254;
assign n6523 = ~(n1670 ^ n25087);
assign n16394 = ~(n3359 ^ n14570);
assign n7506 = ~(n3460 ^ n19477);
assign n20712 = n17975 | n4202;
assign n4067 = ~(n19 ^ n13803);
assign n6603 = ~(n11124 ^ n11469);
assign n10647 = ~(n18388 ^ n19851);
assign n17817 = ~(n17909 | n24650);
assign n4432 = ~(n7559 ^ n12484);
assign n20704 = ~(n8684 ^ n6783);
assign n292 = ~(n26443 | n23807);
assign n16989 = ~(n12016 ^ n14921);
assign n836 = ~(n5611 | n24420);
assign n23014 = ~(n3145 ^ n6745);
assign n24707 = n23360 & n12785;
assign n19044 = ~(n14980 ^ n9822);
assign n2248 = ~n15681;
assign n7734 = ~(n19441 ^ n26796);
assign n10382 = n17826 | n24620;
assign n4687 = ~n18909;
assign n17070 = ~(n16572 ^ n22385);
assign n13443 = ~n9942;
assign n13277 = ~(n15978 ^ n11949);
assign n10064 = ~(n15616 ^ n20104);
assign n15052 = n20228 | n13856;
assign n6751 = ~(n21997 ^ n18483);
assign n17582 = n23540 | n11923;
assign n13531 = n1792 | n19521;
assign n2732 = ~(n2851 ^ n4835);
assign n22484 = ~(n12629 ^ n10232);
assign n10579 = n323 | n8403;
assign n1205 = ~n15743;
assign n6276 = ~(n6343 ^ n9842);
assign n0 = n8660 | n8328;
assign n11155 = ~(n1974 ^ n17576);
assign n3488 = n19963 & n3432;
assign n19750 = n6836 & n23517;
assign n23825 = ~(n23166 ^ n4306);
assign n18426 = ~n17094;
assign n12962 = ~n13912;
assign n18141 = n18882 | n8856;
assign n6587 = ~(n4733 ^ n2699);
assign n7349 = ~(n14681 ^ n188);
assign n19695 = ~(n1531 | n7302);
assign n20205 = ~n18483;
assign n11457 = ~n16223;
assign n215 = n16848 & n19628;
assign n10024 = ~(n6074 ^ n15556);
assign n23417 = ~n24801;
assign n16896 = ~(n4831 ^ n21266);
assign n8019 = ~(n101 ^ n8416);
assign n23736 = n22808 & n7824;
assign n23531 = n4445 | n12574;
assign n25254 = ~(n16318 ^ n26118);
assign n13067 = n6695 & n499;
assign n14055 = ~(n15271 ^ n26748);
assign n14067 = n9363 | n11088;
assign n12790 = ~(n729 ^ n25692);
assign n55 = ~(n22776 ^ n2499);
assign n5220 = ~n6307;
assign n16663 = ~n6774;
assign n18534 = ~(n26211 ^ n15583);
assign n12221 = n21634 | n2035;
assign n10461 = n8948 | n9242;
assign n6414 = ~(n1152 ^ n25023);
assign n26488 = ~n18951;
assign n967 = n19911 & n26658;
assign n4079 = n16593 | n25191;
assign n4690 = n23455 | n25285;
assign n13153 = n15560 | n7006;
assign n10860 = n16695 | n6365;
assign n8778 = ~(n8241 ^ n2985);
assign n27020 = n4469 & n7212;
assign n23348 = n5144 | n5862;
assign n22172 = ~(n26216 ^ n8331);
assign n23179 = n15829 & n7690;
assign n26151 = n11921 | n1324;
assign n13681 = n22918 & n20719;
assign n10923 = ~n16948;
assign n1086 = ~(n21715 | n25615);
assign n7279 = n26695 | n23890;
assign n16628 = ~n5558;
assign n1434 = n3414 & n21465;
assign n20015 = ~n20003;
assign n26013 = ~n947;
assign n4953 = ~(n22206 ^ n5030);
assign n2639 = n9431 | n7592;
assign n24749 = ~(n22985 ^ n20182);
assign n24243 = ~n23344;
assign n9142 = ~(n22022 ^ n13832);
assign n9743 = ~(n13286 ^ n7096);
assign n24149 = n14751 | n7927;
assign n10534 = ~(n9041 ^ n7117);
assign n4586 = ~(n26318 | n18895);
assign n25567 = n14099 | n13526;
assign n2196 = ~(n6169 | n26302);
assign n2301 = ~(n6351 ^ n7731);
assign n20623 = ~(n22759 ^ n5435);
assign n26156 = ~(n1475 ^ n18694);
assign n3044 = n17942 & n17059;
assign n21376 = n26715 & n12690;
assign n22197 = ~n17900;
assign n23591 = n17933 | n25003;
assign n12025 = n27174 & n9866;
assign n17638 = ~(n7874 ^ n15399);
assign n7725 = ~(n26811 ^ n3895);
assign n16405 = ~(n2252 | n16672);
assign n11374 = ~n19876;
assign n14509 = n20541 | n21754;
assign n22806 = ~(n12513 ^ n8395);
assign n12434 = n26170 | n8635;
assign n15252 = ~(n7689 ^ n3827);
assign n10853 = n20427 | n13281;
assign n27165 = ~(n8176 ^ n9554);
assign n6639 = n9798 & n17672;
assign n21255 = n19684 & n14877;
assign n7750 = ~n20901;
assign n3411 = ~n19393;
assign n909 = ~(n17250 ^ n4409);
assign n21221 = n21982 & n2606;
assign n14473 = n11400 & n20130;
assign n10799 = ~(n7640 | n3509);
assign n3019 = ~(n22280 ^ n18522);
assign n6736 = ~(n6297 ^ n7272);
assign n8420 = ~n6456;
assign n16402 = n14336 | n18149;
assign n11026 = ~(n17579 | n6632);
assign n10558 = n24417 | n4719;
assign n9664 = n24417 | n24907;
assign n26254 = n5967 & n21835;
assign n15837 = n8732 & n4651;
assign n20230 = n3362 & n21695;
assign n16898 = ~(n18974 ^ n21918);
assign n8141 = n16668 | n5982;
assign n26561 = n522 | n20432;
assign n16003 = ~(n1205 | n7494);
assign n10061 = n26634 & n7314;
assign n5946 = ~(n26549 ^ n4482);
assign n7352 = n20395 & n11604;
assign n25769 = n26658 | n15539;
assign n10615 = n24231 | n9305;
assign n24010 = n10555 | n23291;
assign n21380 = ~n18537;
assign n4743 = n23615 & n4521;
assign n19707 = ~(n6566 ^ n10875);
assign n6127 = ~(n12824 ^ n7545);
assign n7621 = ~n8324;
assign n22602 = ~(n26963 | n22828);
assign n19346 = n11901 | n24044;
assign n12895 = ~(n10649 ^ n6289);
assign n8954 = n10726 & n124;
assign n13524 = n2411 & n9062;
assign n24803 = n3494 & n6211;
assign n5219 = n14723 | n12086;
assign n9059 = n27160 | n13948;
assign n18323 = ~(n64 ^ n5851);
assign n9795 = n10744 | n23243;
assign n23984 = ~(n24494 ^ n24359);
assign n14776 = n10883 & n19778;
assign n17386 = n2357 & n6008;
assign n20261 = ~(n23428 | n25282);
assign n17273 = ~(n27074 | n12208);
assign n5016 = n11758 & n12457;
assign n11830 = ~(n3574 ^ n10246);
assign n5507 = ~(n7297 ^ n304);
assign n25454 = ~(n16667 ^ n3460);
assign n24917 = n23974 | n26085;
assign n4791 = n25405 ^ n21627;
assign n24115 = ~n11018;
assign n23971 = n4815 | n22655;
assign n21455 = ~n2055;
assign n4528 = n12844 | n2158;
assign n22981 = ~n21907;
assign n15307 = ~(n23079 ^ n16040);
assign n465 = n23612 | n3906;
assign n13116 = ~(n13200 ^ n6147);
assign n7096 = ~n17758;
assign n4702 = n22752 & n16857;
assign n12098 = ~(n4314 ^ n15001);
assign n26265 = ~(n20030 ^ n337);
assign n8549 = ~n8438;
assign n23668 = ~(n9058 | n5925);
assign n15155 = ~(n2902 | n19809);
assign n16404 = n1358 | n12339;
assign n20608 = ~n12289;
assign n15247 = n15104 | n11123;
assign n20779 = n17354 | n23265;
assign n679 = ~(n9090 ^ n19107);
assign n16876 = n25105 & n10925;
assign n25174 = n25682 | n15457;
assign n6591 = ~n8730;
assign n6048 = n12199 & n14712;
assign n8810 = ~(n4957 ^ n25797);
assign n6598 = n11808 | n5645;
assign n18453 = ~(n5342 | n26919);
assign n6405 = n11583 | n18416;
assign n12711 = n4381 | n26809;
assign n2398 = n15129 | n541;
assign n16777 = n20675 | n18778;
assign n105 = n7142 | n3860;
assign n12876 = ~(n14603 | n24736);
assign n6113 = n16633 | n22379;
assign n15536 = ~n21390;
assign n954 = ~(n1099 | n6381);
assign n2502 = n11273 & n23086;
assign n24665 = ~n11479;
assign n25392 = n11737 | n14274;
assign n23185 = n22198 | n14424;
assign n24222 = n14633 | n2886;
assign n13847 = n15125 | n23587;
assign n26909 = n2121 | n10625;
assign n11860 = ~(n767 ^ n8806);
assign n13255 = ~(n12088 ^ n26483);
assign n26158 = n11919 | n12875;
assign n16323 = n1096 | n19879;
assign n25674 = ~n1777;
assign n4346 = ~(n7437 ^ n13367);
assign n3819 = ~(n23353 | n14881);
assign n15323 = n26677 | n21745;
assign n1335 = ~(n8546 | n10855);
assign n14234 = n8606 | n16282;
assign n21591 = n18264 | n14373;
assign n24444 = ~(n7525 ^ n11900);
assign n6990 = n20739 & n3864;
assign n8558 = n16498 & n13342;
assign n13993 = ~(n12928 ^ n12650);
assign n22717 = ~(n15132 ^ n4614);
assign n24838 = ~(n15655 | n12415);
assign n2194 = n13879;
assign n23598 = n3945 | n3393;
assign n2330 = n4256 & n20205;
assign n18601 = ~(n21086 ^ n2861);
assign n7215 = ~n8405;
assign n21560 = n19832 & n3201;
assign n5916 = ~n5694;
assign n21295 = ~(n11119 ^ n22279);
assign n6511 = ~(n13897 | n19515);
assign n19962 = ~n21993;
assign n1025 = ~n18250;
assign n12220 = n8372 | n17979;
assign n25188 = ~(n18438 | n26672);
assign n3990 = ~n2937;
assign n10971 = ~(n17485 | n17555);
assign n10653 = ~(n1303 ^ n4425);
assign n17118 = ~(n2815 | n4492);
assign n24944 = n3413 | n17762;
assign n2424 = n11487 & n2082;
assign n21783 = n15696 | n13071;
assign n3055 = n1561 & n13130;
assign n690 = ~(n10208 ^ n2290);
assign n4313 = n15121 | n4724;
assign n24790 = n1454 | n9123;
assign n15769 = ~n4836;
assign n27185 = ~(n9025 ^ n11032);
assign n14821 = ~(n10135 | n24863);
assign n4358 = n14404 | n25479;
assign n5061 = n25318 | n3955;
assign n12411 = n936 & n2584;
assign n161 = ~(n2359 ^ n25213);
assign n20045 = ~n21649;
assign n3275 = n3440 & n6028;
assign n3812 = n3553 | n5116;
assign n24272 = ~n686;
assign n6180 = n24492 & n17619;
assign n11387 = ~(n25523 ^ n26318);
assign n21980 = ~(n17467 ^ n16376);
assign n20841 = ~n4417;
assign n15440 = ~(n18733 ^ n565);
assign n5022 = ~(n13109 ^ n7731);
assign n25484 = n27093 | n6056;
assign n9601 = n22962 | n10567;
assign n4199 = n13951 | n19388;
assign n19874 = ~n13533;
assign n13827 = ~(n6847 ^ n2051);
assign n10126 = n24651 & n27162;
assign n18540 = n13964 & n26576;
assign n15394 = n12442 | n12677;
assign n13347 = ~(n7365 ^ n8495);
assign n5580 = ~n14570;
assign n15158 = ~(n17109 ^ n9686);
assign n10202 = ~(n25318 ^ n2645);
assign n7050 = ~(n8402 ^ n8589);
assign n4105 = n1611 | n21763;
assign n23782 = ~(n4856 ^ n3653);
assign n13393 = n926 & n14498;
assign n8279 = n5623 & n13181;
assign n9894 = n16331 | n5443;
assign n11468 = n994 & n19503;
assign n5100 = n21431 | n5529;
assign n7313 = ~(n25672 ^ n14280);
assign n16814 = n7739 & n9353;
assign n15791 = n11212 & n26033;
assign n394 = ~n15169;
assign n21714 = n3621 & n13002;
assign n6069 = n1918 | n16653;
assign n10453 = n9004 | n21014;
assign n21619 = n5825 | n8788;
assign n6250 = ~(n16822 ^ n17415);
assign n16601 = ~(n10882 | n8719);
assign n3626 = n13195 | n16051;
assign n14046 = ~(n12797 ^ n26810);
assign n11865 = n18171 & n24529;
assign n13582 = n5151 & n3191;
assign n23615 = n2960 | n1413;
assign n17556 = n21804 | n22272;
assign n5218 = n14281 & n8043;
assign n8679 = ~(n19199 ^ n3166);
assign n546 = ~n20442;
assign n25897 = ~(n14323 | n14071);
assign n21403 = n6320 | n8956;
assign n10375 = ~n17174;
assign n861 = ~(n3968 ^ n13980);
assign n7073 = n19880 | n2405;
assign n10005 = n20552 | n7841;
assign n5593 = ~(n20688 ^ n13421);
assign n5018 = n15025 | n23080;
assign n366 = ~(n16800 | n14678);
assign n1731 = ~(n11411 ^ n25195);
assign n16609 = ~(n258 ^ n7524);
assign n18326 = ~(n18457 ^ n9750);
assign n22902 = ~(n21517 ^ n16972);
assign n25124 = n9030 & n1789;
assign n15451 = ~n1400;
assign n6311 = ~(n6757 ^ n3400);
assign n12103 = n20809 | n7560;
assign n19366 = ~(n10115 ^ n17342);
assign n21102 = n18476 | n27042;
assign n4320 = ~n25848;
assign n13040 = n7170 & n19186;
assign n5344 = n14013 & n19656;
assign n460 = n26691 | n9496;
assign n8055 = n21487 & n10749;
assign n4374 = ~(n24012 ^ n18993);
assign n6319 = ~n18400;
assign n24882 = n19007 & n25002;
assign n9777 = ~(n9797 | n4240);
assign n24413 = n16405 | n1729;
assign n19788 = n7737 | n14218;
assign n358 = n19054 & n13331;
assign n392 = n9141 | n12533;
assign n3491 = n16713 | n17497;
assign n1464 = ~n1629;
assign n9256 = ~(n11428 ^ n5266);
assign n16725 = ~n5197;
assign n22144 = ~(n25118 ^ n3222);
assign n2922 = ~(n10077 ^ n4651);
assign n15603 = ~n9418;
assign n13894 = ~n11830;
assign n6346 = ~(n23843 ^ n25505);
assign n18685 = ~(n10761 ^ n14384);
assign n7033 = n19336 & n17111;
assign n13472 = ~(n1017 ^ n1011);
assign n23290 = ~n10603;
assign n12496 = n16980 & n5390;
assign n16879 = ~(n10125 | n7619);
assign n20087 = ~(n10124 ^ n1893);
assign n13014 = ~(n4119 ^ n5255);
assign n8414 = ~n6988;
assign n26485 = n1591 | n17621;
assign n13054 = ~(n19031 ^ n21142);
assign n10229 = ~(n17091 ^ n20288);
assign n6256 = ~(n19837 ^ n19686);
assign n15986 = ~(n13391 ^ n5193);
assign n6442 = ~n23773;
assign n19230 = ~(n7740 ^ n20429);
assign n2704 = n15572 & n27143;
assign n21297 = ~(n24116 | n1163);
assign n20854 = n4327 & n27045;
assign n14831 = n25494 | n10713;
assign n5418 = n13420 & n19337;
assign n12080 = n15847 | n24017;
assign n23326 = n12125 | n21224;
assign n12514 = ~n1855;
assign n5491 = ~(n5376 | n6037);
assign n5181 = n18921 & n1028;
assign n15188 = n4623 | n373;
assign n14124 = ~(n19146 ^ n16476);
assign n22035 = n6663 & n24253;
assign n1914 = n2874 & n25960;
assign n15240 = ~(n3917 ^ n23503);
assign n17606 = n9764 | n20082;
assign n17027 = n16929 | n1708;
assign n6317 = n15560 | n246;
assign n20834 = n25481 & n16323;
assign n23130 = n8449 & n14817;
assign n9014 = n6764 | n9964;
assign n15939 = ~(n9680 | n25360);
assign n1767 = n14972 | n5354;
assign n15248 = n5243 & n24961;
assign n17759 = n5445 | n17497;
assign n6021 = ~(n2750 ^ n25393);
assign n8261 = ~n21740;
assign n7810 = ~(n16429 | n6607);
assign n17727 = ~n1697;
assign n24422 = n4938 & n10999;
assign n6386 = n13190 | n15769;
assign n3988 = n18798 | n4723;
assign n8515 = n14887 | n4610;
assign n8277 = ~n8889;
assign n23792 = ~n8473;
assign n17315 = n7095 | n22665;
assign n3007 = ~n20233;
assign n22046 = n5711 | n26378;
assign n12706 = n23647 | n24465;
assign n5441 = n5926 & n2419;
assign n18322 = ~(n5203 ^ n26048);
assign n19435 = ~(n9814 ^ n12145);
assign n16599 = n3791 | n3710;
assign n5067 = ~n16217;
assign n23081 = n19652 | n22610;
assign n20475 = n3731 | n6176;
assign n1575 = ~(n7402 ^ n24367);
assign n6489 = ~n16875;
assign n6076 = ~(n24336 ^ n8986);
assign n9377 = ~(n16765 ^ n11650);
assign n14256 = ~(n23844 ^ n6328);
assign n11981 = ~n10833;
assign n24297 = ~(n17463 ^ n7210);
assign n9123 = n9484 & n18641;
assign n24065 = ~(n19406 | n2121);
assign n2458 = n17586 | n11295;
assign n6985 = ~(n17315 ^ n18489);
assign n15079 = ~n14071;
assign n19096 = n3312 | n2786;
assign n13572 = n3491 & n20677;
assign n7489 = n23646 & n17624;
assign n11 = n1950 | n17809;
assign n23822 = ~(n1153 ^ n24242);
assign n17506 = n22709 & n24895;
assign n20641 = ~n48;
assign n24291 = n18091 & n2400;
assign n19637 = n24904 | n2676;
assign n11171 = ~(n16544 | n1835);
assign n25673 = n23486 | n16663;
assign n1185 = n22232 & n4316;
assign n2308 = n12699 & n8688;
assign n14284 = ~(n1646 | n16638);
assign n25170 = ~(n16311 ^ n3356);
assign n3876 = n14150 | n23554;
assign n7974 = ~n8052;
assign n539 = n8004 & n26485;
assign n19111 = ~(n4328 ^ n9391);
assign n5910 = n22461 & n9074;
assign n6633 = ~(n15884 ^ n5211);
assign n26785 = n3883 & n4991;
assign n24277 = ~(n11048 | n3714);
assign n8050 = ~n2366;
assign n580 = ~(n2988 ^ n14769);
assign n8593 = n23437 & n16100;
assign n16490 = ~(n7600 ^ n5627);
assign n13195 = ~(n4534 ^ n10654);
assign n922 = n20517 | n16744;
assign n14283 = n5673 | n16146;
assign n19971 = ~n17000;
assign n5235 = n11378 | n853;
assign n13605 = ~(n4149 | n25523);
assign n17380 = ~(n24557 ^ n26820);
assign n17178 = n12404 & n7855;
assign n26096 = ~(n18623 ^ n10298);
assign n18362 = ~(n22373 ^ n25170);
assign n26168 = ~(n3640 ^ n20027);
assign n14645 = ~(n24517 | n26327);
assign n5656 = n18528 | n22544;
assign n137 = ~(n18745 | n11976);
assign n24045 = n12557 | n16489;
assign n2748 = n3753 | n11438;
assign n7204 = n13367 & n13074;
assign n11445 = n25376 | n4040;
assign n10178 = n19610 & n9159;
assign n14906 = n1234 | n15994;
assign n11737 = ~(n4416 ^ n24447);
assign n7154 = n8056 | n6358;
assign n3619 = ~(n6645 | n17379);
assign n2879 = n16169 & n25865;
assign n5251 = n16613 & n17783;
assign n19525 = ~(n13912 | n10684);
assign n25245 = ~(n1112 ^ n13190);
assign n1834 = ~(n1315 ^ n25635);
assign n19978 = ~n9797;
assign n18712 = n3230 | n589;
assign n2250 = ~(n5072 | n1132);
assign n16547 = ~(n18016 ^ n647);
assign n7861 = ~(n26171 ^ n4247);
assign n8966 = ~(n7731 | n23509);
assign n24557 = n25528 | n18556;
assign n10818 = ~(n5205 ^ n6065);
assign n15497 = n23732 & n17875;
assign n19129 = n16822 | n5963;
assign n9150 = ~n38;
assign n6041 = n4350 | n17216;
assign n2094 = ~(n22517 ^ n19894);
assign n7762 = n4878 | n15654;
assign n1954 = ~(n20213 | n7092);
assign n26912 = ~n7001;
assign n2445 = ~n17261;
assign n22561 = ~(n14563 | n23508);
assign n7051 = ~(n655 | n5386);
assign n7525 = n943 & n23811;
assign n26709 = ~(n14872 ^ n12553);
assign n9689 = ~(n21391 ^ n81);
assign n1362 = ~(n17771 | n14762);
assign n13973 = ~(n16022 ^ n18575);
assign n13789 = ~n24319;
assign n10257 = ~(n15498 ^ n16562);
assign n23795 = n23218 | n22266;
assign n7025 = ~(n2377 | n19633);
assign n12293 = ~n6184;
assign n446 = ~n16544;
assign n25637 = ~n12605;
assign n26548 = ~(n24301 | n2289);
assign n10939 = n16480 | n17001;
assign n22705 = n24595 | n17614;
assign n9033 = n5152 & n2097;
assign n17717 = ~(n20811 | n19047);
assign n830 = n25872 | n19262;
assign n3659 = ~n23754;
assign n22273 = ~n19222;
assign n808 = ~n11424;
assign n18025 = n8534 | n24550;
assign n14111 = ~n19236;
assign n20531 = n8472 | n23318;
assign n15709 = ~n4811;
assign n5669 = n19410 | n14035;
assign n3010 = ~(n13866 ^ n3973);
assign n5309 = n19150 | n25074;
assign n17376 = n6260 & n18448;
assign n8531 = n11992 & n11821;
assign n16607 = ~(n13960 | n12990);
assign n1665 = n5205 & n6065;
assign n26390 = ~(n20593 | n4174);
assign n11770 = ~(n7385 | n20241);
assign n21936 = ~(n11936 | n2756);
assign n1787 = n11585 | n5023;
assign n24357 = n11774 & n7250;
assign n19636 = ~(n7465 ^ n22550);
assign n10861 = ~n21726;
assign n23227 = n19902 | n15125;
assign n6542 = ~(n6187 ^ n25641);
assign n12898 = ~n16176;
assign n17040 = n2945 & n24946;
assign n13733 = n1211 & n16050;
assign n20019 = n15609 & n15915;
assign n18022 = n3576 & n26712;
assign n14562 = n2442 & n9041;
assign n25363 = n11020 | n24225;
assign n26877 = n20455 & n25099;
assign n18325 = n4315 | n3945;
assign n16146 = ~(n6166 ^ n22581);
assign n21270 = n17607 & n16470;
assign n23904 = n4359 | n10465;
assign n25226 = n8494 & n20762;
assign n2046 = ~(n13643 ^ n11707);
assign n19900 = n1473 & n7336;
assign n14076 = ~n409;
assign n13055 = n1439 | n13699;
assign n11498 = n18907 & n13033;
assign n1502 = n11745 | n10057;
assign n23154 = n21320 & n23785;
assign n10603 = ~(n22248 ^ n23567);
assign n15937 = n7335 | n11578;
assign n3301 = ~(n24017 ^ n10210);
assign n24348 = ~(n11321 | n964);
assign n3125 = ~(n23381 ^ n24679);
assign n308 = n21096 & n22044;
assign n15950 = ~(n23592 | n14226);
assign n2111 = ~(n27029 ^ n27028);
assign n23172 = n17187 | n17985;
assign n23387 = n1951 | n27008;
assign n7483 = n5280 | n19774;
assign n16306 = n21611 & n14585;
assign n2411 = n6692 | n10897;
assign n13645 = n5820 & n24445;
assign n7491 = ~(n2244 ^ n3465);
assign n20827 = n5041 & n7202;
assign n25314 = ~(n9259 | n16401);
assign n22266 = ~(n23977 ^ n2760);
assign n9295 = n2454 | n4970;
assign n25263 = ~(n16637 | n2776);
assign n19221 = ~(n19782 ^ n3565);
assign n4651 = ~(n21758 ^ n11461);
assign n1616 = n9790 & n3060;
assign n6370 = n13544 | n13570;
assign n24851 = ~n7428;
assign n23492 = n14685 & n13282;
assign n9173 = n15340 | n3048;
assign n8042 = ~(n10362 ^ n12498);
assign n18916 = ~(n14465 | n7057);
assign n346 = ~(n1055 | n12592);
assign n5326 = n10184 | n6284;
assign n1917 = ~(n2025 ^ n5053);
assign n5136 = n20106 | n4472;
assign n3274 = ~(n11819 ^ n6583);
assign n12557 = ~(n16890 | n3318);
assign n11059 = n7692 | n16793;
assign n1690 = ~(n7394 ^ n5579);
assign n6578 = ~(n16127 | n18918);
assign n2459 = n3460 & n24774;
assign n20821 = ~(n5065 | n12018);
assign n4795 = n7101 | n6990;
assign n14568 = n9592 | n19860;
assign n23829 = ~(n1078 ^ n13170);
assign n11198 = ~n21778;
assign n24179 = n6859 | n17600;
assign n4475 = n9725 | n19526;
assign n7588 = ~(n18716 ^ n26025);
assign n16315 = n11075 | n5858;
assign n13522 = n12159 & n23078;
assign n21693 = ~(n6820 ^ n24278);
assign n24837 = ~(n3354 ^ n12078);
assign n19930 = ~(n17807 ^ n8065);
assign n11105 = ~(n21674 ^ n22597);
assign n9996 = ~(n10684 ^ n13912);
assign n9876 = n11526 & n15199;
assign n853 = n15937 & n3704;
assign n12170 = n10317 | n23928;
assign n793 = ~(n5145 | n3675);
assign n11714 = ~n23873;
assign n6897 = ~(n22325 ^ n25940);
assign n17681 = ~(n25781 ^ n9469);
assign n20963 = ~(n22610 ^ n19652);
assign n12448 = ~(n20079 | n11406);
assign n1016 = ~(n10015 ^ n16262);
assign n22967 = n11633 | n14178;
assign n26440 = n25199 | n13955;
assign n11214 = n16081 & n21135;
assign n21300 = ~(n15320 ^ n245);
assign n26165 = n22837 & n18033;
assign n24507 = ~n25681;
assign n906 = ~(n26066 ^ n6356);
assign n19698 = ~(n10763 ^ n12657);
assign n14981 = ~(n22067 ^ n10516);
assign n21143 = ~(n15459 ^ n10585);
assign n12638 = ~n21165;
assign n8453 = ~(n2980 ^ n20601);
assign n17475 = ~(n23705 | n1759);
assign n24026 = n8599 | n10954;
assign n17344 = ~(n16172 ^ n21233);
assign n26941 = n2725 | n6389;
assign n5845 = n14435 & n1666;
assign n21390 = ~(n21348 ^ n21586);
assign n27025 = ~n14354;
assign n12539 = n5148 & n15412;
assign n22188 = n10495 | n8942;
assign n19013 = n4681 & n22037;
assign n25490 = ~(n7401 ^ n15964);
assign n16714 = ~(n17444 ^ n27037);
assign n26295 = ~n15625;
assign n24377 = n17173 | n4468;
assign n18998 = ~(n24134 ^ n5095);
assign n9719 = n1657 | n21672;
assign n25428 = n24699 & n17406;
assign n9112 = ~(n25621 | n6930);
assign n5027 = n21519 & n25709;
assign n3388 = n15883 | n14381;
assign n9941 = n16178 | n3955;
assign n8428 = n14487 & n27022;
assign n7976 = ~(n2482 ^ n7448);
assign n20103 = ~(n25269 ^ n24368);
assign n21888 = n11056 & n10181;
assign n6339 = ~(n7663 ^ n12790);
assign n4491 = n16569 & n19189;
assign n10916 = n23304 & n17069;
assign n1997 = ~n4042;
assign n3071 = n9560 & n14608;
assign n24832 = ~n19762;
assign n2062 = n24557 & n15630;
assign n15612 = n12492 & n21594;
assign n6474 = ~(n5998 ^ n12384);
assign n23990 = ~(n7510 ^ n13438);
assign n16929 = ~(n3585 ^ n6207);
assign n23127 = n19452 | n3527;
assign n12782 = n14803 | n1115;
assign n2657 = ~(n10988 ^ n3669);
assign n24472 = ~(n10163 ^ n20458);
assign n19906 = n11668 | n7332;
assign n19188 = n10958 | n19580;
assign n976 = ~(n14388 | n21575);
assign n10582 = ~(n1421 ^ n15378);
assign n24324 = ~(n27075 | n16239);
assign n7838 = ~(n23456 ^ n8964);
assign n2908 = ~n14762;
assign n27111 = ~n12713;
assign n4470 = n10892 | n419;
assign n23269 = ~(n17847 | n11394);
assign n7624 = n16515 | n9824;
assign n5384 = ~(n3276 | n2547);
assign n15903 = ~(n26576 ^ n5636);
assign n18384 = n25797 & n15784;
assign n19420 = ~(n9455 ^ n18290);
assign n23680 = ~(n10577 ^ n3279);
assign n7546 = ~n27046;
assign n24061 = n4662 & n25091;
assign n159 = ~(n19683 ^ n24048);
assign n5726 = n13277 | n19869;
assign n7248 = n23943 | n18723;
assign n4726 = n3248 | n11568;
assign n9521 = ~(n19377 ^ n17780);
assign n7232 = ~(n10631 | n9125);
assign n9161 = n20348 & n9724;
assign n18252 = ~(n7991 ^ n3133);
assign n3498 = ~n8974;
assign n24849 = ~(n22755 | n310);
assign n9240 = ~(n22108 ^ n22626);
assign n22075 = n17282 & n169;
assign n18797 = ~n9827;
assign n18224 = n5355 & n17659;
assign n15807 = ~(n439 ^ n16304);
assign n16697 = ~n22006;
assign n4251 = n4270 | n4438;
assign n18176 = n24654 | n22340;
assign n11213 = ~(n20196 ^ n25872);
assign n17160 = ~(n26270 ^ n19495);
assign n8854 = n26086 | n7149;
assign n15719 = ~(n21043 ^ n25963);
assign n10903 = ~(n14109 ^ n12357);
assign n26066 = ~n4067;
assign n19567 = ~(n22375 | n24815);
assign n21523 = n5119 & n6070;
assign n13900 = n13534 | n15500;
assign n7357 = n3840 | n24908;
assign n16860 = ~(n25164 ^ n16490);
assign n6176 = n25284 & n17823;
assign n20675 = n19754 & n11308;
assign n1270 = n9770 | n25676;
assign n18834 = n614 | n19075;
assign n2530 = n17532 & n1334;
assign n17304 = n14007 | n23144;
assign n11241 = ~(n557 ^ n19390);
assign n3166 = ~(n19914 ^ n23895);
assign n10835 = n16812 & n24402;
assign n17866 = ~(n24638 ^ n19327);
assign n22254 = ~n3570;
assign n26973 = n12058 | n285;
assign n11326 = ~(n8730 ^ n6130);
assign n5566 = n4278 | n15074;
assign n449 = n7676 | n9380;
assign n16944 = ~(n19471 | n11491);
assign n17631 = n5400 | n3149;
assign n4917 = ~(n20381 ^ n17218);
assign n17939 = ~(n985 | n19218);
assign n23194 = n26746 | n2224;
assign n26076 = ~(n8295 ^ n13037);
assign n1920 = n14785 | n480;
assign n3317 = ~n27181;
assign n1855 = ~(n16725 ^ n11973);
assign n22542 = ~(n14510 ^ n21649);
assign n10052 = n3417 | n12986;
assign n26312 = ~n8614;
assign n5162 = ~(n8472 ^ n6150);
assign n17399 = n504 | n26135;
assign n6438 = n16743 & n24081;
assign n26618 = n26611 & n4235;
assign n892 = n24081 | n16743;
assign n10764 = n7203 & n3989;
assign n10123 = ~(n1009 | n1293);
assign n2880 = ~(n2328 ^ n18274);
assign n17799 = ~(n24417 | n11363);
assign n6306 = ~(n19106 | n24879);
assign n17454 = ~n1418;
assign n17953 = ~n11116;
assign n17434 = n7030 | n23752;
assign n25936 = ~n16476;
assign n7369 = ~(n22820 ^ n7693);
assign n11348 = ~(n2047 ^ n19485);
assign n17573 = n25134 & n10865;
assign n5439 = ~(n17970 ^ n14324);
assign n14177 = n15463 | n13820;
assign n20547 = n17992 | n25137;
assign n2076 = ~(n16924 ^ n10984);
assign n7385 = n25483 & n1062;
assign n8723 = n1912 | n1160;
assign n5066 = ~n820;
assign n2962 = n19084 | n28;
assign n7198 = ~n14680;
assign n11677 = n4628 & n21769;
assign n22745 = ~(n20192 | n12481);
assign n6441 = n16380 | n886;
assign n25393 = ~n2023;
assign n10248 = ~(n22585 | n20986);
assign n23580 = ~n22215;
assign n20878 = n14293 | n2914;
assign n2787 = ~n12993;
assign n511 = n14026 & n15853;
assign n124 = n609 | n18070;
assign n22865 = ~n13489;
assign n26818 = n25029 | n10089;
assign n7602 = n24031 | n25261;
assign n20699 = n22102 & n3560;
assign n5075 = ~(n13062 ^ n21230);
assign n24087 = n23202 | n10813;
assign n7037 = n1191 | n14513;
assign n16873 = ~n5751;
assign n7181 = ~(n20925 ^ n23791);
assign n1684 = ~(n3883 ^ n18225);
assign n7873 = ~(n8856 ^ n4319);
assign n24113 = n18669 | n13891;
assign n17427 = ~(n11428 ^ n1181);
assign n24835 = ~(n25294 ^ n22474);
assign n14974 = ~n21309;
assign n5009 = n17660 | n26520;
assign n19012 = n10116 | n20485;
assign n8795 = ~n19111;
assign n19413 = n2321 | n11950;
assign n9143 = ~(n8531 ^ n5731);
assign n24140 = n25939 | n26947;
assign n19253 = n10940 | n1362;
assign n21188 = n13460 & n5156;
assign n9328 = n8412 & n12200;
assign n14152 = ~n18478;
assign n3091 = ~(n17835 | n8166);
assign n26746 = ~(n15918 | n21735);
assign n14936 = ~n27188;
assign n25347 = ~(n15979 | n15008);
assign n7441 = n15391 & n20816;
assign n23937 = n13912 & n11098;
assign n13262 = ~(n18369 ^ n21319);
assign n7400 = n2822 & n13090;
assign n20637 = n7301 & n26115;
assign n15461 = ~(n7734 | n5163);
assign n24370 = ~(n4859 | n5140);
assign n16738 = ~n23752;
assign n21412 = ~n11838;
assign n11461 = ~(n15998 ^ n5142);
assign n6162 = ~(n12875 ^ n26318);
assign n699 = ~(n17647 | n20146);
assign n8275 = n16427 | n1807;
assign n25066 = ~n26142;
assign n2630 = ~(n5673 ^ n19337);
assign n23340 = n22839 & n21419;
assign n5883 = ~(n5793 | n2782);
assign n2992 = ~(n14152 ^ n25987);
assign n13291 = ~(n26336 ^ n3264);
assign n22668 = n12893 | n2463;
assign n4283 = n4593 & n7694;
assign n26917 = n13918 ^ n26462;
assign n18155 = n15696 | n18800;
assign n610 = ~(n13783 ^ n22332);
assign n8561 = n12149 | n1915;
assign n24551 = ~n4734;
assign n14223 = ~(n16547 ^ n12900);
assign n26195 = ~(n18558 ^ n6556);
assign n11564 = ~(n26802 ^ n22172);
assign n18307 = ~(n20512 ^ n25726);
assign n27058 = n15729 & n24831;
assign n19067 = n18078 | n12543;
assign n9229 = n14660 & n14929;
assign n11963 = ~n20411;
assign n9066 = n3672 | n14886;
assign n7401 = n10559 & n10182;
assign n2136 = n11065 & n23334;
assign n3479 = ~(n1018 ^ n25808);
assign n17034 = n10374 | n22389;
assign n12661 = n9121 & n25343;
assign n20279 = ~(n5433 ^ n8807);
assign n23947 = n9739 & n4262;
assign n3920 = n15224 | n8877;
assign n26060 = n7796 & n13878;
assign n21961 = n16929 & n1708;
assign n17935 = n20357 & n998;
assign n2147 = ~(n3212 ^ n16251);
assign n26712 = n25553 | n2882;
assign n17329 = n12218 | n26637;
assign n5032 = n18353 | n24206;
assign n9315 = n3636 | n24889;
assign n16977 = n13575 | n19305;
assign n9962 = n3108 & n13805;
assign n4766 = ~(n10186 ^ n1539);
assign n5005 = n6353 | n12391;
assign n25732 = n9297 | n2767;
assign n5467 = n6032 | n15596;
assign n20262 = n6605 & n20322;
assign n8190 = n26526 & n7135;
assign n10959 = n15034 | n19408;
assign n731 = n24938 & n21618;
assign n20669 = ~(n26986 ^ n3425);
assign n5684 = ~(n24902 | n8623);
assign n2120 = n11155 | n972;
assign n23003 = n13306 | n7525;
assign n12226 = ~(n12592 ^ n1055);
assign n11199 = n2058 | n10112;
assign n7866 = n2169 | n7393;
assign n17446 = ~(n19895 | n14311);
assign n6151 = n53 | n18197;
assign n26867 = ~(n13708 ^ n24618);
assign n1878 = n3335 | n8057;
assign n455 = ~n14463;
assign n13520 = n17393 & n18457;
assign n21530 = n18180 & n5861;
assign n13548 = ~(n6806 ^ n2065);
assign n11510 = ~(n13651 ^ n20727);
assign n18942 = n3083 | n1564;
assign n23274 = ~(n18995 | n19357);
assign n1700 = ~(n6434 ^ n25956);
assign n14664 = n23108 & n17604;
assign n19821 = n21499 & n25753;
assign n1975 = n2868 | n881;
assign n23311 = n24828 & n19368;
assign n5869 = n25436 | n8395;
assign n17277 = ~(n25401 ^ n391);
assign n18863 = ~(n26789 ^ n342);
assign n20160 = ~n23889;
assign n10715 = n7652 | n18826;
assign n24983 = n26363 | n22047;
assign n2505 = n10947 & n23354;
assign n20530 = ~(n26792 ^ n21584);
assign n7978 = n9918 & n15420;
assign n12168 = n10712 | n14467;
assign n18061 = ~(n14817 ^ n13560);
assign n14708 = ~(n2568 | n13625);
assign n3478 = ~(n7439 ^ n3984);
assign n4357 = n11233 & n1990;
assign n6334 = ~(n966 ^ n8687);
assign n21816 = ~(n19974 ^ n23435);
assign n18285 = n26550 | n4768;
assign n10966 = ~n15424;
assign n4639 = n10826 | n16381;
assign n18438 = ~(n12415 ^ n16984);
assign n23254 = ~n19432;
assign n7235 = ~(n18046 ^ n14969);
assign n22922 = n3305 | n6538;
assign n17100 = ~(n7305 | n25538);
assign n22134 = ~(n24196 | n22049);
assign n21670 = ~(n9832 ^ n6513);
assign n12781 = n15658 | n1312;
assign n11853 = n24822 & n2772;
assign n24491 = ~(n8194 ^ n24093);
assign n5960 = ~n10739;
assign n12723 = ~(n15135 ^ n25712);
assign n17947 = ~(n8540 ^ n2146);
assign n12053 = ~(n14528 | n6713);
assign n26719 = ~(n8393 ^ n11298);
assign n1839 = ~n26141;
assign n26455 = n12847 | n2255;
assign n1811 = ~(n24475 | n19568);
assign n18659 = ~(n1960 | n18749);
assign n5149 = n11435 & n25670;
assign n11292 = n3284 | n2041;
assign n17779 = ~n2586;
assign n21076 = n6312 & n27083;
assign n8299 = ~(n25312 ^ n9206);
assign n1477 = n4801 & n9723;
assign n16681 = ~(n3298 ^ n26443);
assign n13102 = ~(n10378 | n2312);
assign n12939 = ~(n10031 ^ n23578);
assign n11224 = ~(n17211 ^ n20054);
assign n22875 = n23158 & n10880;
assign n22568 = ~(n22613 ^ n22631);
assign n19220 = ~(n3115 ^ n4523);
assign n24418 = ~(n17444 ^ n19652);
assign n11238 = ~(n1136 | n11667);
assign n17211 = ~n25498;
assign n12102 = ~(n8344 ^ n16217);
assign n16156 = n4760 & n24711;
assign n17829 = ~(n3161 ^ n21134);
assign n11465 = n19 | n26913;
assign n16946 = n24987 & n15584;
assign n3809 = ~(n2158 ^ n13830);
assign n23786 = n21021 & n18355;
assign n7170 = ~n20446;
assign n2828 = ~(n6341 ^ n13783);
assign n18603 = n25008 | n6501;
assign n24405 = ~(n9519 | n22330);
assign n3616 = ~(n14033 ^ n22554);
assign n11906 = n26530 | n25465;
assign n16633 = ~n767;
assign n16801 = ~(n13186 ^ n11611);
assign n11996 = ~(n18579 ^ n2177);
assign n25266 = n24892 | n8859;
assign n15102 = n10602 | n10984;
assign n13379 = ~n16526;
assign n24430 = n9673 | n13799;
assign n15718 = n9115 | n15461;
assign n11843 = ~(n8172 ^ n9086);
assign n5317 = ~(n23373 | n16732);
assign n23085 = ~n10179;
assign n13372 = ~(n7311 ^ n25023);
assign n3083 = ~(n19589 | n8935);
assign n14095 = ~(n850 ^ n6585);
assign n4267 = n26502 & n23332;
assign n10881 = ~(n24969 | n26544);
assign n23152 = ~n5969;
assign n24529 = ~(n10179 ^ n13708);
assign n17422 = n10425 | n18337;
assign n25318 = ~n1835;
assign n16078 = n17547 & n15524;
assign n19830 = ~(n14684 | n17360);
assign n22147 = n15240 | n14111;
assign n21566 = ~(n4602 | n12402);
assign n15189 = ~n8256;
assign n8881 = ~(n6656 ^ n9787);
assign n15333 = ~(n12759 ^ n26192);
assign n20082 = n3269 & n26843;
assign n21148 = ~(n27104 | n9114);
assign n9746 = n19644 | n25552;
assign n20378 = ~n3918;
assign n9164 = ~(n13913 ^ n5357);
assign n10851 = ~(n3342 ^ n11866);
assign n2427 = n1553 | n13774;
assign n25137 = n22890 & n23041;
assign n2369 = ~(n22077 | n26351);
assign n7452 = ~n23513;
assign n2245 = n9958 | n16538;
assign n14494 = n26850 & n213;
assign n23713 = n7747 | n9331;
assign n2321 = n4304 & n23876;
assign n5847 = ~(n20077 ^ n6794);
assign n24924 = ~(n10096 | n24511);
assign n2590 = ~(n24493 | n19200);
assign n6548 = n26613 | n4771;
assign n22697 = ~(n1126 ^ n7420);
assign n2089 = ~n24586;
assign n26305 = n14195 | n19874;
assign n3934 = ~(n17580 ^ n9760);
assign n19668 = ~(n8943 | n10919);
assign n12942 = ~(n26589 ^ n4647);
assign n4435 = ~(n12678 ^ n2700);
assign n25408 = ~(n12002 | n16890);
assign n1529 = n25257 | n24132;
assign n4092 = ~(n3472 ^ n10477);
assign n16930 = n14189 | n14795;
assign n5371 = ~(n25322 | n23329);
assign n15235 = n2389 | n20233;
assign n14081 = ~(n7044 ^ n6302);
assign n8202 = ~(n15415 | n12875);
assign n3818 = n3606 | n24643;
assign n7417 = ~n1243;
assign n13154 = ~n9493;
assign n11961 = n319 | n23032;
assign n17193 = ~(n22626 ^ n26986);
assign n23647 = ~(n22525 ^ n6121);
assign n13735 = ~(n115 ^ n22859);
assign n9993 = ~(n23477 ^ n21398);
assign n10552 = n16029 & n12088;
assign n3394 = n25882 | n19078;
assign n18567 = n7444 | n17076;
assign n23678 = ~n13354;
assign n24369 = n6259 | n14838;
assign n17969 = ~(n4722 ^ n14323);
assign n16324 = ~(n25842 ^ n13736);
assign n15296 = n18794 | n16038;
assign n1805 = n25629 | n2291;
assign n10515 = n3327 | n13120;
assign n25083 = ~(n24149 ^ n15965);
assign n11781 = n12511 | n4590;
assign n11247 = n25319 & n11250;
assign n761 = n20701 & n4447;
assign n10669 = ~(n5411 ^ n6729);
assign n8909 = ~(n1610 | n1500);
assign n12031 = n17826 | n13033;
assign n869 = n16722 & n2230;
assign n6789 = ~n5424;
assign n1534 = n2995 & n15678;
assign n3523 = n19547 | n12781;
assign n5511 = ~(n6352 | n424);
assign n1461 = ~(n3228 | n6082);
assign n12305 = n11921 & n1324;
assign n10817 = ~(n2717 ^ n5259);
assign n14670 = n25941 & n13958;
assign n13790 = n16211 | n2289;
assign n6257 = ~(n15132 ^ n23514);
assign n15660 = n3253 & n21021;
assign n8431 = ~n24744;
assign n2608 = ~(n3723 ^ n16823);
assign n4815 = ~(n16572 | n22012);
assign n1294 = n812 | n15498;
assign n17005 = n9196 | n13731;
assign n16238 = n7331 | n4356;
assign n14779 = ~(n18765 ^ n22626);
assign n15638 = n9693 | n10767;
assign n13567 = ~(n15486 ^ n11149);
assign n10858 = ~(n25637 ^ n27100);
assign n5793 = n4616;
assign n15500 = ~n3641;
assign n10925 = n25933 | n1323;
assign n19065 = n17208 | n12182;
assign n22296 = n653 & n13883;
assign n15865 = n21662 | n7568;
assign n16342 = n6547 | n4611;
assign n10352 = ~(n26397 ^ n13179);
assign n17630 = ~(n19565 ^ n10867);
assign n13479 = n17990 & n7037;
assign n16493 = ~(n27177 ^ n12005);
assign n15071 = ~(n17584 | n19282);
assign n5949 = ~n25966;
assign n3194 = n23662 & n22512;
assign n8457 = ~n7274;
assign n23358 = n11766 & n9530;
assign n9302 = ~(n7963 ^ n12161);
assign n875 = n7423 | n156;
assign n20342 = ~n17458;
assign n353 = ~(n24714 | n22501);
assign n18922 = n1587 | n1685;
assign n16275 = ~(n9604 ^ n16174);
assign n3556 = ~(n11485 ^ n19147);
assign n20781 = n15133 | n4289;
assign n953 = n21794 & n10332;
assign n19187 = ~(n7177 ^ n21828);
assign n17063 = n8416 & n101;
assign n11031 = ~(n20138 | n25073);
assign n1934 = ~n13562;
assign n11836 = n6451 | n10988;
assign n24168 = n3805 & n24159;
assign n23969 = ~(n5111 ^ n4514);
assign n11422 = n17642 | n26256;
assign n8514 = ~n26080;
assign n15315 = n4859 & n9793;
assign n17609 = n14818 | n17532;
assign n26366 = n18183 | n18466;
assign n8559 = n19938 | n11623;
assign n524 = ~n7693;
assign n17086 = n22754 | n13569;
assign n9308 = ~(n5444 ^ n8756);
assign n21331 = n20312 | n19567;
assign n5604 = ~n14899;
assign n7323 = ~(n3379 ^ n1099);
assign n24190 = n17272 | n13929;
assign n17555 = ~(n127 ^ n273);
assign n19482 = ~(n26556 ^ n12495);
assign n10613 = n4101 & n16435;
assign n25721 = ~(n19469 | n20235);
assign n16830 = ~n27104;
assign n26275 = n25959 | n20392;
assign n24727 = ~n4277;
assign n19475 = n7436 | n4606;
assign n13115 = ~(n715 ^ n9591);
assign n18684 = n21016 | n7966;
assign n6125 = ~(n11841 ^ n19701);
assign n16882 = ~n8441;
assign n8322 = ~n5213;
assign n15841 = ~(n4426 | n25246);
assign n6926 = n14789 | n3790;
assign n14743 = n11854 | n19807;
assign n7128 = n3634 | n9263;
assign n14166 = n22730 | n8235;
assign n15056 = n14830 & n6468;
assign n21466 = n16985 & n8833;
assign n14317 = n14133 & n7293;
assign n4139 = ~(n25739 ^ n8419);
assign n12252 = ~(n7334 ^ n20961);
assign n5201 = n11898 & n25063;
assign n327 = ~(n23898 ^ n15182);
assign n24479 = ~n8437;
assign n11060 = ~n12020;
assign n19610 = ~n16818;
assign n17430 = ~(n21362 ^ n25812);
assign n16201 = ~(n20390 ^ n12842);
assign n9008 = n5461 | n20529;
assign n25164 = ~(n23563 ^ n24979);
assign n20661 = ~(n594 ^ n9199);
assign n20573 = n17831 | n15475;
assign n22524 = n442 | n6319;
assign n4190 = n7689 | n22600;
assign n24600 = ~(n9701 ^ n19431);
assign n22240 = ~(n14907 | n26522);
assign n23887 = n14818 | n26491;
assign n31 = ~(n24305 ^ n2580);
assign n10326 = ~(n7199 ^ n10386);
assign n11057 = n21643 | n101;
assign n25095 = n14886 | n17639;
assign n21296 = n2556 | n8893;
assign n6638 = ~(n22198 | n5337);
assign n24942 = ~(n16713 | n15808);
assign n20725 = ~(n14272 | n1929);
assign n14814 = ~(n9108 | n530);
assign n14179 = n17385 | n27073;
assign n14666 = ~(n3324 ^ n16544);
assign n23451 = ~n5795;
assign n6740 = n23274 | n23689;
assign n21741 = n658 | n25339;
assign n21000 = ~(n9373 ^ n7677);
assign n20586 = n420 | n12535;
assign n22785 = n19353 & n6784;
assign n6447 = n8150 | n1328;
assign n12604 = n6691 | n19222;
assign n8177 = n2967 | n7099;
assign n507 = ~n3673;
assign n14108 = n13999 | n14376;
assign n12688 = ~(n1654 | n4256);
assign n15893 = n22991 & n467;
assign n4381 = n14923 & n12050;
assign n5551 = n16096 & n6952;
assign n319 = n5091 & n9743;
assign n14438 = n6691 & n21753;
assign n17786 = n12287 | n20299;
assign n16178 = ~n8182;
assign n25632 = ~(n11144 ^ n25500);
assign n26126 = ~(n22031 ^ n20824);
assign n9395 = ~n21195;
assign n10953 = n7548 | n9339;
assign n23837 = ~n21778;
assign n8062 = n22845 | n1655;
assign n6388 = ~(n23160 ^ n3570);
assign n13810 = n8713 & n6071;
assign n11844 = ~(n15546 ^ n14702);
assign n22086 = n24748 & n16170;
assign n21075 = n6291 | n5693;
assign n3213 = n25435 | n19527;
assign n9919 = ~(n5716 ^ n10280);
assign n16484 = ~(n23268 ^ n15282);
assign n13508 = ~(n18891 | n14078);
assign n3890 = ~n19575;
assign n17723 = ~(n21317 ^ n19196);
assign n16401 = ~n21577;
assign n19536 = n3855 & n1193;
assign n12027 = n3907 | n16586;
assign n3680 = n21271 | n15772;
assign n25142 = ~n20455;
assign n13210 = n16789 | n10962;
assign n6193 = ~n26483;
assign n14827 = ~(n8919 ^ n5819);
assign n6096 = ~(n3967 | n27054);
assign n7228 = n10181 | n5796;
assign n6236 = n7566 | n2389;
assign n18527 = ~n17854;
assign n1590 = ~(n4109 ^ n12827);
assign n19050 = ~(n18046 | n1025);
assign n10847 = ~n5171;
assign n12243 = n12666 | n7218;
assign n23635 = n24158 | n24785;
assign n14927 = ~(n20359 ^ n25240);
assign n23759 = n13559 | n4250;
assign n4249 = n22100 & n23482;
assign n5470 = ~(n23631 ^ n3365);
assign n4767 = ~n25076;
assign n1085 = n9055 & n21990;
assign n3443 = ~n1309;
assign n21006 = n23821 & n17769;
assign n13208 = ~(n17212 ^ n26725);
assign n12555 = ~(n11209 ^ n23250);
assign n14507 = ~n14603;
assign n3090 = ~n7822;
assign n26235 = ~n5285;
assign n25963 = ~(n21021 ^ n18355);
assign n707 = ~(n2776 | n4853);
assign n10000 = ~(n19957 ^ n26954);
assign n16672 = ~n22105;
assign n27122 = ~n4913;
assign n24304 = ~(n9988 | n17824);
assign n24567 = n27119 & n10656;
assign n21855 = n840 | n21001;
assign n10289 = ~(n19682 ^ n9133);
assign n5423 = n20852 | n26283;
assign n17114 = ~(n24802 ^ n19108);
assign n978 = ~n21964;
assign n15910 = ~(n11527 ^ n24365);
assign n22232 = ~n14045;
assign n23375 = n1511 & n19690;
assign n8109 = ~(n5979 ^ n18455);
assign n15341 = n2576 | n21276;
assign n9078 = n11650 | n20901;
assign n13088 = ~n21915;
assign n25312 = ~(n599 ^ n22888);
assign n7138 = ~(n10454 ^ n21856);
assign n16996 = n1458 | n22433;
assign n2323 = ~(n7601 ^ n4656);
assign n6865 = ~n6613;
assign n1067 = ~(n1843 | n25667);
assign n22899 = ~(n16882 ^ n16683);
assign n5171 = n25819 & n1050;
assign n1132 = ~n5200;
assign n11045 = ~n2160;
assign n26029 = n23923 | n23874;
assign n23025 = n22519 | n10734;
assign n26759 = n8605 | n8668;
assign n9526 = ~(n19108 | n24802);
assign n13234 = ~n6109;
assign n10048 = ~n224;
assign n18239 = n5238 | n26193;
assign n21014 = ~(n9746 ^ n22391);
assign n10998 = ~n15016;
assign n9231 = ~(n5420 | n14554);
assign n17285 = ~(n6343 ^ n25798);
assign n24003 = n16812 | n1279;
assign n19055 = ~n14918;
assign n3940 = ~n13455;
assign n4379 = n21563 | n8365;
assign n10765 = n13550 & n12062;
assign n7360 = ~n1654;
assign n25294 = n15763 | n5662;
assign n10383 = ~(n26991 ^ n1354);
assign n1424 = ~(n7057 | n7823);
assign n3244 = ~(n20309 ^ n14194);
assign n20283 = n21536 | n16491;
assign n21843 = n19201 | n23211;
assign n5342 = ~n24451;
assign n12938 = ~(n5072 ^ n1132);
assign n17505 = ~n22020;
assign n13165 = n19770 & n11451;
assign n24888 = n15542 | n8221;
assign n15781 = n26781 & n20738;
assign n25624 = ~(n14182 ^ n2113);
assign n25679 = ~(n14984 ^ n17954);
assign n22706 = n6393 & n19082;
assign n22696 = n26104 | n10527;
assign n4959 = ~(n1190 ^ n20353);
assign n25129 = n8773 & n11657;
assign n24504 = ~(n6834 ^ n8399);
assign n9669 = n23095 & n21704;
assign n20391 = ~(n21311 ^ n6216);
assign n21167 = n20570 | n1934;
assign n3807 = ~(n8875 | n19215);
assign n6187 = n24849 | n26785;
assign n21377 = ~(n18710 | n21796);
assign n12634 = n1624 | n23829;
assign n12824 = ~(n18338 ^ n17549);
assign n11561 = n18257 | n19905;
assign n8878 = ~(n8614 | n24705);
assign n20037 = ~(n24550 | n25405);
assign n3757 = n14988 | n8201;
assign n15999 = ~(n18735 ^ n14393);
assign n3661 = ~(n11486 | n18409);
assign n20850 = ~(n5296 ^ n8672);
assign n4378 = n2314 | n1163;
assign n25279 = ~(n8152 | n19695);
assign n25423 = ~(n26264 ^ n19454);
assign n17899 = ~(n6168 | n12151);
assign n16665 = ~n18584;
assign n19068 = n18150 & n21440;
assign n18338 = n20202 | n24633;
assign n7214 = n1031 & n8443;
assign n387 = ~(n3201 ^ n9085);
assign n2047 = n11861 & n22641;
assign n6982 = ~(n978 | n26946);
assign n6457 = ~(n14453 ^ n16860);
assign n18093 = n20612 | n21264;
assign n4752 = ~n19033;
assign n20994 = n26717 | n26748;
assign n15930 = ~n7684;
assign n1396 = ~n4024;
assign n10877 = n16711 | n2059;
assign n17560 = ~(n2289 ^ n18345);
assign n12656 = n18090 | n12474;
assign n21108 = n21643 & n101;
assign n8903 = n8106 | n10904;
assign n10346 = ~(n18480 ^ n9499);
assign n11700 = n25246 | n24728;
assign n17798 = ~(n16443 ^ n23996);
assign n9776 = n605 | n8691;
assign n25501 = ~(n20249 ^ n24684);
assign n4263 = ~(n26720 ^ n11832);
assign n3181 = n2465 & n13101;
assign n6324 = n20140 | n4308;
assign n22213 = ~(n4209 ^ n21212);
assign n21273 = n6341 | n21246;
assign n10786 = n19541 | n23863;
assign n958 = ~(n8420 | n10406);
assign n16310 = ~(n23983 ^ n20040);
assign n19122 = n15579 & n293;
assign n10992 = ~(n2915 | n12014);
assign n6562 = n7469 & n12608;
assign n15270 = n11951 & n18713;
assign n26803 = ~(n6696 ^ n23423);
assign n23005 = ~n23102;
assign n23752 = ~(n11150 ^ n4063);
assign n1401 = ~n14830;
assign n20323 = ~n23102;
assign n6851 = ~(n5551 ^ n22078);
assign n22729 = ~n10018;
assign n9047 = ~(n21714 ^ n14868);
assign n6686 = ~(n23141 ^ n20792);
assign n8877 = n11388 & n17161;
assign n23431 = ~(n10106 | n17379);
assign n24566 = n2719 | n15229;
assign n19450 = ~(n8686 ^ n25585);
assign n16914 = n23563 | n2434;
assign n456 = ~n6523;
assign n19152 = ~(n19494 ^ n2387);
assign n12311 = ~n2167;
assign n230 = n5065 | n8487;
assign n27129 = n23023 & n23520;
assign n17932 = ~n19820;
assign n26449 = ~(n10885 ^ n19276);
assign n24523 = n19531 & n11425;
assign n20424 = ~(n2969 | n3066);
assign n4793 = n19331 | n11675;
assign n15955 = ~(n2899 ^ n6485);
assign n7604 = ~n1469;
assign n3609 = n10670 & n19232;
assign n12020 = n10914 | n17685;
assign n8341 = n23492 | n22307;
assign n14352 = ~(n24129 ^ n9380);
assign n4631 = ~(n7532 ^ n17664);
assign n20845 = n13057 & n12391;
assign n19319 = n26420 | n21694;
assign n19980 = n19077 & n23149;
assign n14953 = ~(n22962 | n1715);
assign n21892 = n11178 | n1079;
assign n607 = n10948 | n10243;
assign n13264 = n20986 | n12212;
assign n22415 = n15184 & n16605;
assign n25117 = n13389 & n17695;
assign n11873 = n11456 | n25118;
assign n8891 = n22079;
assign n14846 = n20716 | n6708;
assign n8316 = n21222 | n18820;
assign n15849 = n16047 | n14167;
assign n18134 = ~(n3324 | n2272);
assign n23533 = n9235 & n24667;
assign n17889 = ~(n19744 ^ n24955);
assign n14363 = ~(n4293 | n5739);
assign n10832 = ~n115;
assign n22272 = ~(n6775 ^ n3925);
assign n17485 = ~(n10842 ^ n18571);
assign n26243 = n6966 & n27128;
assign n9138 = ~(n692 | n26015);
assign n12832 = ~(n8539 ^ n15975);
assign n14448 = n26264 | n5661;
assign n16784 = n7726 | n3550;
assign n5873 = n10325 & n8544;
assign n6980 = n2330 | n9188;
assign n24091 = ~n26927;
assign n1860 = ~(n2921 ^ n362);
assign n6648 = ~n14649;
assign n15904 = n16867 & n9173;
assign n16874 = ~(n11747 ^ n23400);
assign n22592 = ~(n20179 ^ n26823);
assign n8260 = n21646 & n22098;
assign n14096 = ~(n20153 ^ n13308);
assign n9758 = n24950 & n13416;
assign n8768 = n7016 & n12584;
assign n24473 = ~(n13433 ^ n16915);
assign n22347 = n53 | n14487;
assign n9096 = ~n21016;
assign n9139 = n21341 | n23780;
assign n3820 = n23516 & n17258;
assign n23006 = ~(n25906 ^ n22832);
assign n5073 = ~(n23509 ^ n23755);
assign n3345 = ~(n14826 | n13549);
assign n3878 = ~(n25862 ^ n9996);
assign n6146 = n5238 | n7351;
assign n24545 = n24383 & n6403;
assign n14063 = ~(n5320 ^ n24330);
assign n18411 = n15358 | n6182;
assign n23097 = ~n24475;
assign n18000 = ~(n20040 | n9396);
assign n5413 = n14859 & n3039;
assign n1074 = ~(n10086 ^ n25330);
assign n11607 = ~(n5558 ^ n7791);
assign n9975 = ~(n5065 ^ n6204);
assign n13425 = ~(n4677 ^ n3918);
assign n25823 = n1705 & n9456;
assign n13260 = n18159 | n8887;
assign n14705 = ~n10407;
assign n4476 = ~(n21440 ^ n17833);
assign n22029 = n13367 & n20970;
assign n7836 = ~(n23784 | n4127);
assign n25640 = n10452 | n22723;
assign n25661 = n16711 | n21753;
assign n3103 = n3129 & n26365;
assign n25740 = ~(n20751 | n24593);
assign n1365 = ~n18962;
assign n15327 = ~(n12340 ^ n16659);
assign n14023 = n25742 | n7312;
assign n13860 = ~(n24161 ^ n4426);
assign n22616 = n19466 | n25594;
assign n7301 = n21918 | n18974;
assign n18095 = n14119 | n7963;
assign n7008 = ~(n9395 ^ n7144);
assign n5776 = ~(n3624 ^ n10905);
assign n6415 = n24073 & n12170;
assign n22734 = ~(n19033 ^ n7674);
assign n4761 = n5226 | n11223;
assign n24412 = ~(n19143 ^ n5891);
assign n12633 = n18117 & n6997;
assign n11322 = n24451;
assign n19268 = n21924 & n9476;
assign n10138 = ~(n26185 ^ n4573);
assign n4988 = n2795 & n12796;
assign n2115 = ~(n2576 | n1682);
assign n14396 = n927 & n17165;
assign n23054 = ~(n9631 | n22879);
assign n20554 = ~n9445;
assign n3393 = ~n22972;
assign n25665 = ~(n5669 ^ n4358);
assign n19430 = n2850 | n14482;
assign n24482 = ~(n5934 ^ n23636);
assign n15479 = n10636 & n16362;
assign n824 = ~(n23559 ^ n21455);
assign n10729 = n10738 | n6934;
assign n9407 = ~(n23586 | n17728);
assign n10926 = n17435 & n2905;
assign n16317 = n2637 | n4248;
assign n5503 = ~(n25967 ^ n24327);
assign n5640 = n17579 & n12452;
assign n14419 = ~(n9605 ^ n11806);
assign n20273 = ~n6414;
assign n12042 = n21956 & n16076;
assign n9000 = ~(n22859 | n12859);
assign n25931 = ~n24150;
assign n17345 = n10480 | n23840;
assign n7868 = ~n17614;
assign n26493 = n6422 | n13503;
assign n8461 = ~(n22631 ^ n21078);
assign n18753 = ~(n17978 ^ n6456);
assign n5303 = n5255 | n6446;
assign n3258 = ~n3793;
assign n22323 = ~(n13152 | n2688);
assign n1768 = ~(n15602 | n8507);
assign n6072 = n25420 & n14807;
assign n20889 = n17449 | n568;
assign n24326 = ~(n16111 ^ n20109);
assign n26424 = n16029 | n4322;
assign n8873 = ~n18589;
assign n21790 = ~(n17626 | n2246);
assign n19727 = ~(n17098 ^ n11096);
assign n89 = n5427 | n19633;
assign n4962 = n11740 | n11816;
assign n5504 = n23718 | n17221;
assign n1056 = n12575 | n19325;
assign n17031 = n13529 | n20594;
assign n17184 = ~n21510;
assign n26858 = n18123 | n1697;
assign n15422 = ~n17771;
assign n24341 = ~(n18787 | n5944);
assign n533 = n3721 | n26403;
assign n17903 = ~(n5682 ^ n10468);
assign n21918 = ~(n12559 ^ n6620);
assign n10050 = ~(n20045 | n19357);
assign n15087 = ~(n17363 ^ n4758);
assign n17603 = n16496 | n17647;
assign n25315 = n15136 | n13051;
assign n2179 = n16128 | n1002;
assign n15587 = n116 & n16069;
assign n6494 = n6259 & n14838;
assign n5202 = n27140 | n19028;
assign n13 = ~n26038;
assign n25940 = ~(n1487 ^ n22928);
assign n1340 = ~n20409;
assign n13927 = n16983 & n14411;
assign n5695 = ~(n9711 ^ n11317);
assign n8464 = n20342 | n26830;
assign n16562 = ~(n5985 ^ n22514);
assign n13101 = n19688 | n7024;
assign n9520 = n14306 | n14400;
assign n9913 = ~(n395 | n19215);
assign n9695 = ~(n20943 ^ n17526);
assign n20197 = ~(n3257 ^ n3677);
assign n9625 = n10651 | n23639;
assign n24939 = ~n26565;
assign n26863 = n7997 | n15851;
assign n12908 = ~(n7241 ^ n10592);
assign n18447 = n483 | n8827;
assign n14477 = ~n19138;
assign n14897 = ~(n14878 | n16213);
assign n4819 = ~(n12956 | n1118);
assign n18763 = ~(n22219 ^ n4781);
assign n464 = ~(n17734 ^ n16900);
assign n9312 = n15505 | n5264;
assign n7409 = n17179 & n6035;
assign n16160 = n15127 | n26680;
assign n4093 = ~n4105;
assign n2342 = ~n3468;
assign n22300 = ~(n11824 ^ n5709);
assign n21037 = ~n26523;
assign n18976 = n13023 & n9548;
assign n17822 = n21268 | n14899;
assign n23709 = ~(n18111 ^ n2944);
assign n4755 = n24893 & n174;
assign n9483 = ~(n25345 ^ n23463);
assign n16136 = ~(n15099 ^ n8825);
assign n12420 = ~(n11397 ^ n12043);
assign n2034 = n21767 | n23985;
assign n22749 = n11611 & n13186;
assign n12201 = ~(n26947 ^ n4467);
assign n5426 = ~(n8000 | n13035);
assign n8001 = ~(n2186 ^ n19148);
assign n7080 = ~(n25512 | n23132);
assign n17789 = ~n16430;
assign n702 = n16820 | n18944;
assign n22150 = ~(n187 ^ n10549);
assign n3145 = n24735 | n26339;
assign n13875 = ~n16214;
assign n18379 = n22198 | n24493;
assign n1326 = n331 & n684;
assign n7905 = n25913 ^ n5490;
assign n5595 = n6288 | n14333;
assign n142 = ~(n20911 ^ n11576);
assign n3276 = ~n3164;
assign n26010 = n8175 & n13423;
assign n4490 = ~n20169;
assign n7277 = ~(n10462 ^ n25630);
assign n14977 = ~(n14655 ^ n13258);
assign n3245 = ~(n4557 ^ n3573);
assign n8597 = ~n24093;
assign n14460 = n18293 | n11444;
assign n405 = ~n26553;
assign n10517 = n1964 & n21387;
assign n17284 = n26997 | n6185;
assign n18434 = ~(n20679 ^ n15624);
assign n13656 = n22645 & n12711;
assign n22434 = ~(n26445 | n3881);
assign n10941 = n8363 & n2812;
assign n5013 = ~(n2659 | n9957);
assign n17418 = ~n4670;
assign n25514 = n11414;
assign n25194 = ~n2073;
assign n4004 = ~n25905;
assign n13702 = n2702 & n22863;
assign n10329 = n5076 & n22438;
assign n15531 = n23335 & n12678;
assign n19952 = ~n3541;
assign n4330 = ~n27022;
assign n22610 = ~(n22629 ^ n23735);
assign n9387 = ~n20822;
assign n25846 = n24932;
assign n18596 = ~(n8612 ^ n3324);
assign n12819 = ~(n10343 | n8997);
assign n2588 = ~n2425;
assign n6295 = n17182 & n21625;
assign n10107 = n15077 | n23412;
assign n20541 = n4893 & n21451;
assign n5222 = ~n19069;
assign n12878 = ~n11733;
assign n14348 = n14205 & n19998;
assign n6188 = n11055 | n9162;
assign n23769 = ~n8845;
assign n26963 = ~n379;
assign n13593 = n13900 & n19744;
assign n18680 = ~(n3968 ^ n16900);
assign n23804 = ~n15506;
assign n16135 = ~(n5172 | n16948);
assign n14199 = n7386 & n13242;
assign n4674 = ~(n26346 ^ n12194);
assign n6154 = ~(n17709 ^ n23747);
assign n25248 = n5498 | n16294;
assign n6554 = ~(n24067 ^ n20221);
assign n8451 = ~n6168;
assign n20773 = n14899 | n18496;
assign n27105 = ~(n8363 ^ n2145);
assign n14616 = n10488 | n2649;
assign n20406 = ~(n21283 ^ n20859);
assign n7013 = n18649 & n13968;
assign n5718 = n15950 | n4399;
assign n11099 = n6307 | n13079;
assign n11159 = ~(n10358 ^ n8484);
assign n11845 = ~(n18715 ^ n9247);
assign n23651 = n21090 & n1241;
assign n11839 = n19733 | n21338;
assign n18701 = n18095 & n18697;
assign n13487 = ~(n24120 ^ n24446);
assign n24191 = ~(n4887 ^ n15861);
assign n3930 = n1967 | n17334;
assign n296 = ~(n2857 | n13282);
assign n21330 = n10704 | n11908;
assign n4585 = ~(n4800 ^ n25846);
assign n9594 = ~n9323;
assign n22940 = ~(n3479 ^ n22386);
assign n1109 = ~(n5302 ^ n19116);
assign n25925 = ~(n20444 ^ n19313);
assign n5571 = n11027 | n7904;
assign n13364 = n24324 | n9437;
assign n17215 = ~(n6043 ^ n13039);
assign n2509 = ~n22654;
assign n2900 = ~(n21372 ^ n13276);
assign n20520 = n3931 | n20076;
assign n5668 = ~n10554;
assign n16303 = n8394 & n10801;
assign n1723 = ~(n6239 ^ n20209);
assign n25261 = ~(n2956 ^ n8985);
assign n2353 = n19596 | n15191;
assign n595 = n20605 | n1756;
assign n1801 = n26793 | n26470;
assign n17749 = ~(n10991 ^ n6463);
assign n1198 = ~(n400 | n2322);
assign n5311 = n25402 | n21084;
assign n2796 = n22909 | n19524;
assign n6991 = ~(n19514 ^ n2731);
assign n21136 = n7071 | n22122;
assign n8690 = ~n2420;
assign n2861 = ~(n5140 ^ n10250);
assign n15418 = n4469 | n7212;
assign n11752 = ~(n10041 ^ n10514);
assign n1346 = ~n24638;
assign n22447 = n7319 & n17224;
assign n475 = ~(n8451 | n17047);
assign n14237 = n22825 & n22689;
assign n9478 = n3092 | n18645;
assign n3187 = ~(n24129 ^ n26167);
assign n7705 = ~(n18514 | n16507);
assign n12017 = n18456 & n23530;
assign n9075 = ~(n16058 ^ n4846);
assign n3951 = n828 & n25757;
assign n22530 = n13918 ^ n11672;
assign n12360 = ~n15800;
assign n26647 = ~(n25624 ^ n19327);
assign n7715 = n21263 | n7376;
assign n11203 = n1734 | n5218;
assign n8833 = n7419 | n1126;
assign n16148 = n26436 & n15459;
assign n7782 = n7111 | n15546;
assign n15239 = ~n27042;
assign n20414 = n6769 | n3852;
assign n21405 = ~(n10642 ^ n23142);
assign n6292 = n11000 | n18037;
assign n18350 = ~(n20995 ^ n12680);
assign n7133 = ~n19491;
assign n20141 = n9574 & n1980;
assign n5040 = ~(n11355 | n12596);
assign n5300 = ~(n2806 ^ n4688);
assign n19279 = n25923 | n24184;
assign n11264 = n23431 | n25449;
assign n682 = n7636;
assign n24775 = n8228 | n5570;
assign n3240 = n8758 & n7591;
assign n20791 = ~(n5101 ^ n6659);
assign n13070 = ~(n8398 ^ n17711);
assign n20639 = ~n5874;
assign n17628 = ~(n617 | n20982);
assign n4228 = ~(n20354 ^ n18097);
assign n12195 = ~(n4499 ^ n21671);
assign n17393 = n15241 | n15146;
assign n67 = n1968 & n20223;
assign n8584 = ~(n25302 ^ n3440);
assign n4162 = n3773 & n6294;
assign n21269 = ~n24897;
assign n16104 = ~(n22413 ^ n18265);
assign n25642 = n10804 | n20901;
assign n26657 = n9985 | n14142;
assign n25547 = ~(n13006 ^ n6933);
assign n96 = n15727 | n16685;
assign n26210 = n26565 | n9142;
assign n1980 = n15700 & n5828;
assign n9506 = n10802 & n1719;
assign n16153 = n22808 | n7824;
assign n17539 = ~n987;
assign n19706 = ~(n3254 | n2738);
assign n4576 = ~(n21640 ^ n3492);
assign n5557 = ~n21622;
assign n13710 = ~(n6512 ^ n1723);
assign n23150 = n5505 | n27018;
assign n11676 = ~n16707;
assign n19963 = n25038 | n1380;
assign n11042 = n2476 | n25414;
assign n17740 = n25914 | n9242;
assign n16373 = ~(n1641 ^ n5093);
assign n20780 = ~(n2230 | n7973);
assign n3861 = ~(n443 ^ n18903);
assign n14260 = ~(n18662 | n12657);
assign n3823 = ~(n9279 ^ n5769);
assign n6181 = n17610 & n11327;
assign n1751 = n19061 & n13436;
assign n21002 = n7659 & n15563;
assign n21050 = ~(n5382 ^ n16226);
assign n16627 = ~n11653;
assign n1928 = n21277 & n1908;
assign n21166 = n18569 | n14635;
assign n12340 = n13807 | n301;
assign n15698 = ~(n5136 ^ n23388);
assign n24887 = ~(n7786 ^ n14446);
assign n3814 = ~(n12381 ^ n10557);
assign n25562 = n14250 & n25714;
assign n12182 = n26260 & n4214;
assign n22280 = n17851 | n2691;
assign n18283 = ~(n19167 ^ n26228);
assign n22011 = n22929 & n21844;
assign n9471 = n25629 & n2291;
assign n1730 = ~n6373;
assign n3130 = ~(n19222 | n1786);
assign n18939 = n3551 | n17259;
assign n21275 = ~(n23013 ^ n21622);
assign n1704 = ~n26860;
assign n13438 = ~(n17251 ^ n26107);
assign n9100 = ~n5661;
assign n2059 = ~(n16810 ^ n11739);
assign n1171 = n4918 | n5235;
assign n15083 = n23913 & n24325;
assign n8667 = n16213 | n6468;
assign n17050 = n20813 & n8290;
assign n18881 = n12656 & n26869;
assign n24499 = ~(n11871 ^ n18809);
assign n27127 = ~(n17728 ^ n22652);
assign n16094 = ~n3232;
assign n2953 = n16122 | n6522;
assign n10649 = n15695 | n11088;
assign n11188 = n15265 & n9911;
assign n5047 = n22003 & n7414;
assign n14115 = n11346 | n8902;
assign n12879 = n24125 | n15719;
assign n21971 = n6456 | n8881;
assign n23766 = ~(n9453 ^ n3959);
assign n26093 = ~n10372;
assign n8957 = n4992 & n26736;
assign n12609 = ~(n4325 | n21941);
assign n25432 = ~(n25915 | n13745);
assign n21028 = n21518 & n16338;
assign n8613 = n627 & n10579;
assign n14471 = ~(n15197 ^ n911);
assign n2749 = n24615 & n6181;
assign n20516 = ~n13115;
assign n26412 = n5646 | n16079;
assign n14235 = n21423 | n19781;
assign n4013 = n25347 | n20627;
assign n22459 = n22597 & n16473;
assign n20334 = ~(n656 | n3143);
assign n10042 = n14821 | n7714;
assign n5106 = ~(n1215 | n10486);
assign n19601 = n18518 | n8733;
assign n1186 = ~(n12778 ^ n10577);
assign n12383 = ~(n9714 ^ n8112);
assign n2652 = n26120 | n4116;
assign n12797 = ~n3903;
assign n20943 = n4223 | n4364;
assign n12043 = ~(n17911 ^ n25331);
assign n4120 = ~(n21316 ^ n25073);
assign n11516 = ~n14387;
assign n16111 = ~n19652;
assign n21103 = n3011 | n220;
assign n17666 = n12604 & n20766;
assign n335 = ~(n24612 ^ n21471);
assign n2153 = n11901 | n2281;
assign n19960 = n12764 | n26846;
assign n8288 = ~(n8836 | n22853);
assign n1813 = n13796 | n24740;
assign n18481 = ~(n8745 ^ n16476);
assign n15911 = n18269 & n10784;
assign n592 = ~(n22663 ^ n10737);
assign n4229 = n26421 | n25359;
assign n3040 = ~(n25229 ^ n25079);
assign n15415 = ~n26318;
assign n2973 = n7198 | n25914;
assign n24076 = ~(n26085 ^ n23974);
assign n21228 = ~(n333 ^ n13625);
assign n1457 = ~(n23160 ^ n2421);
assign n15989 = ~(n23141 | n5579);
assign n8610 = n15261 | n14630;
assign n5727 = ~(n14029 ^ n19203);
assign n18646 = ~(n15404 | n10610);
assign n22960 = ~(n16785 ^ n9702);
assign n22364 = ~(n461 ^ n8678);
assign n12806 = ~(n8414 ^ n17679);
assign n15872 = ~(n18 ^ n26808);
assign n8664 = n11694 | n18040;
assign n9306 = n22877 | n6582;
assign n15943 = ~(n6935 | n13249);
assign n4782 = ~(n15365 ^ n26545);
assign n13200 = n7459 & n19253;
assign n19135 = n17448 | n25167;
assign n17984 = ~(n8363 ^ n11481);
assign n9674 = n6091 & n11813;
assign n24355 = ~n12507;
assign n21367 = ~(n21099 ^ n17704);
assign n18023 = n4697 | n9311;
assign n20027 = ~(n10406 ^ n6456);
assign n13320 = n12543 | n25435;
assign n23962 = ~n1717;
assign n4117 = n24609 | n8044;
assign n7590 = ~(n11039 | n12679);
assign n23489 = ~n22198;
assign n16580 = n7198 | n8571;
assign n8760 = ~(n23686 ^ n7523);
assign n26422 = n8092 & n25278;
assign n16184 = n19599 & n24055;
assign n23996 = ~n13166;
assign n20417 = ~(n19145 ^ n14050);
assign n24804 = ~n25100;
assign n11702 = ~(n10637 | n4226);
assign n12007 = n25953 | n4429;
assign n10569 = n20732 | n23236;
assign n1764 = ~(n3078 ^ n26161);
assign n6136 = ~(n3623 | n22517);
assign n24762 = n9172 & n10571;
assign n15656 = n19692 | n4840;
assign n25757 = n12459 | n19324;
assign n15336 = ~(n4304 ^ n23876);
assign n2171 = ~n9509;
assign n21959 = n12004 | n12289;
assign n3185 = ~(n17276 | n3780);
assign n27068 = ~n12153;
assign n10391 = n25336 | n20433;
assign n21290 = n8351 & n11066;
assign n13099 = n1587 & n14008;
assign n18135 = n8627 & n9543;
assign n10956 = n5617 & n22414;
assign n15403 = n2684 & n3680;
assign n25965 = n10771 | n7033;
assign n4200 = n8678 | n16500;
assign n1686 = ~n3825;
assign n23374 = ~(n13529 ^ n7056);
assign n24268 = ~(n8570 ^ n14728);
assign n13778 = n20156 & n26440;
assign n4006 = n8839 & n22758;
assign n5894 = n22802 | n27087;
assign n8180 = ~(n456 | n15400);
assign n8619 = ~(n17630 ^ n18263);
assign n21268 = ~n7026;
assign n6296 = ~(n17122 ^ n14389);
assign n25480 = n14254 & n6964;
assign n1963 = n9004 & n21014;
assign n19953 = n9804 & n8663;
assign n19429 = ~n10477;
assign n7354 = ~(n19331 ^ n24187);
assign n16913 = ~n2517;
assign n11934 = n20871 | n9612;
assign n20009 = ~n14437;
assign n1943 = ~(n14713 ^ n10311);
assign n11901 = ~n6814;
assign n14852 = ~n24340;
assign n15748 = ~(n13044 | n8845);
assign n16058 = ~(n16231 ^ n17754);
assign n1191 = ~(n2570 | n7569);
assign n7702 = ~(n932 ^ n10739);
assign n19772 = ~(n27111 ^ n25265);
assign n6083 = n10491 & n22103;
assign n7389 = ~(n18558 | n6556);
assign n10511 = ~(n20442 ^ n16988);
assign n6629 = n18413 | n15591;
assign n23846 = n13239 | n22356;
assign n7799 = n212 & n17150;
assign n12946 = n8012 & n20870;
assign n23368 = n9756 | n24820;
assign n7956 = n13023 | n6631;
assign n6173 = ~n12113;
assign n5455 = ~(n339 | n11266);
assign n19452 = n25370 & n11603;
assign n3839 = n5763 | n23548;
assign n12856 = n2268 | n22417;
assign n12151 = ~n7555;
assign n5837 = n9537 & n4832;
assign n2239 = ~(n3506 | n9934);
assign n7500 = n3385 | n11990;
assign n18911 = n14572 | n25185;
assign n1531 = ~(n21739 | n24805);
assign n8936 = ~(n1807 ^ n16053);
assign n8114 = n1905 | n4618;
assign n6036 = n5516 | n20125;
assign n18078 = ~n9090;
assign n1469 = ~(n16711 ^ n14378);
assign n11621 = n11791 | n16255;
assign n20718 = ~(n7057 ^ n14570);
assign n1889 = n26855 & n23908;
assign n23220 = ~(n23044 ^ n1681);
assign n13672 = n26797 | n18234;
assign n9922 = ~(n6477 ^ n1118);
assign n16409 = n21700 | n1024;
assign n16604 = n18841 | n20183;
assign n1708 = ~(n17490 ^ n7053);
assign n7724 = n18058 | n12341;
assign n10591 = ~(n26216 ^ n16339);
assign n26836 = n5651 | n17683;
assign n26518 = ~(n19489 ^ n12405);
assign n19805 = ~n2723;
assign n23155 = n203 | n8035;
assign n10394 = ~n23224;
assign n26927 = ~(n18022 ^ n16746);
assign n26380 = ~(n11683 ^ n19015);
assign n7296 = ~(n13590 | n23923);
assign n556 = n5384 | n16899;
assign n20312 = n8664 & n22616;
assign n20253 = ~(n9507 ^ n18409);
assign n14657 = ~(n19985 ^ n6104);
assign n7803 = n14690 & n25399;
assign n1541 = ~(n21074 ^ n1470);
assign n12804 = n11107 & n17657;
assign n326 = n23860 | n18179;
assign n10701 = ~(n21660 ^ n23964);
assign n27054 = ~n1819;
assign n5394 = ~(n17610 | n4858);
assign n23143 = n5229 | n18889;
assign n5456 = n16057 | n12101;
assign n19443 = n14856 | n9107;
assign n18973 = ~n23454;
assign n20638 = ~n20213;
assign n24824 = ~n21508;
assign n23313 = ~n1238;
assign n21344 = ~(n14354 ^ n22335);
assign n8339 = ~(n12710 ^ n17149);
assign n9621 = n6087 & n13364;
assign n4237 = n468 | n1255;
assign n4481 = ~(n12477 ^ n26408);
assign n983 = ~(n8037 | n23636);
assign n6910 = n1705 & n5354;
assign n25905 = ~(n8344 ^ n21654);
assign n9267 = n932 | n2666;
assign n3971 = ~(n11941 ^ n8299);
assign n15370 = n7013 | n7803;
assign n5107 = n9677 & n12370;
assign n26241 = ~n11356;
assign n1004 = ~(n16524 ^ n13668);
assign n13339 = ~n23978;
assign n18040 = ~(n12255 ^ n14181);
assign n9118 = ~(n25914 | n10275);
assign n20640 = n162 | n20509;
assign n734 = n22912 & n7484;
assign n2056 = ~n24048;
assign n7822 = ~(n1451 ^ n26979);
assign n19115 = ~(n329 ^ n1163);
assign n16138 = n26297 & n18948;
assign n13612 = ~(n4801 ^ n11970);
assign n19742 = ~n3429;
assign n8908 = ~(n24487 | n17184);
assign n13948 = n5119 & n10639;
assign n5951 = n1329 | n1898;
assign n11375 = ~(n6913 ^ n9500);
assign n21133 = n10441 & n6727;
assign n15811 = n16156 | n18997;
assign n3170 = n15546 | n14702;
assign n2774 = ~(n14632 | n1507);
assign n109 = ~(n9336 ^ n17969);
assign n5038 = n20881 | n20492;
assign n3472 = ~(n11022 ^ n1955);
assign n26607 = n16743 & n20020;
assign n2877 = n4913 & n13489;
assign n26215 = ~n4867;
assign n1075 = n15647 | n13660;
assign n2614 = ~(n22173 ^ n12593);
assign n13858 = ~(n21974 ^ n22284);
assign n22980 = n13783 | n6341;
assign n26978 = n173 | n9380;
assign n15923 = ~(n5751 | n8730);
assign n5582 = ~(n26176 ^ n423);
assign n5652 = ~n19459;
assign n7916 = n15309 | n1934;
assign n17826 = ~n1163;
assign n11124 = n23532 & n16716;
assign n2769 = ~(n615 | n6944);
assign n22047 = ~(n19512 ^ n23984);
assign n14764 = ~n25652;
assign n21473 = n19831 & n15750;
assign n4454 = ~(n19926 ^ n21295);
assign n12573 = n27117 & n8725;
assign n6150 = ~n13841;
assign n16499 = ~(n13108 ^ n15258);
assign n17406 = n24189 | n13217;
assign n13984 = ~(n17606 ^ n24936);
assign n878 = n15138 | n22492;
assign n2022 = n18409 & n25004;
assign n3849 = ~(n25924 ^ n18962);
assign n16172 = n15357 & n14470;
assign n22489 = ~(n9795 ^ n2112);
assign n14569 = ~n25435;
assign n6273 = ~n9093;
assign n1048 = n1066 & n9502;
assign n15836 = n10056 & n20830;
assign n8066 = ~(n18145 | n26191);
assign n15608 = ~(n9398 | n24599);
assign n22350 = n8313 & n13371;
assign n2015 = n25888 | n24615;
assign n22894 = n19712 | n21080;
assign n14289 = n23411;
assign n22735 = n24958 & n10673;
assign n2055 = ~(n12901 ^ n27105);
assign n19193 = ~(n24143 ^ n12420);
assign n17198 = ~n16319;
assign n12608 = n18236 | n14069;
assign n21712 = n20422 | n12335;
assign n15097 = n19944 | n18962;
assign n14654 = ~n24196;
assign n16716 = n20496 | n15478;
assign n7278 = ~(n25302 ^ n19358);
assign n11588 = n6124 | n26236;
assign n2884 = ~(n13979 ^ n6385);
assign n7492 = ~(n17088 ^ n17832);
assign n2119 = n25324 | n12593;
assign n6636 = ~(n1630 ^ n9507);
assign n18801 = n18659 | n3929;
assign n26523 = ~(n21379 ^ n19731);
assign n15727 = ~(n2896 | n7773);
assign n18716 = n19022 & n875;
assign n8144 = ~(n5747 ^ n9963);
assign n16358 = n402 | n14380;
assign n18590 = n14862 & n16442;
assign n13385 = n10184 | n18006;
assign n24958 = n11580 | n1469;
assign n6411 = n23745 & n23053;
assign n13257 = ~(n24940 ^ n7719);
assign n1490 = n26789 & n11733;
assign n8568 = ~n2809;
assign n5274 = ~(n25114 ^ n16125);
assign n22478 = ~n26584;
assign n6734 = ~(n26960 ^ n1394);
assign n22312 = n13343 | n21286;
assign n25961 = n8555 & n19021;
assign n16615 = ~(n22433 ^ n10158);
assign n20672 = n10661 | n7076;
assign n17295 = ~n16807;
assign n687 = ~(n12068 ^ n4558);
assign n12 = ~n20575;
assign n20629 = ~(n23418 ^ n17207);
assign n9032 = ~(n22698 ^ n25147);
assign n21218 = n11630 & n18504;
assign n163 = n15122 | n16850;
assign n23385 = n13446 | n5676;
assign n25054 = ~(n9530 ^ n7596);
assign n8917 = n4100 | n26326;
assign n19001 = ~(n22554 ^ n26318);
assign n4537 = ~(n7699 ^ n4370);
assign n23475 = ~(n8102 ^ n20791);
assign n23671 = ~(n16203 ^ n12406);
assign n10570 = n21479 | n22435;
assign n7234 = n22347 | n24925;
assign n21087 = n15952 | n24986;
assign n2729 = ~n19751;
assign n133 = ~(n7769 ^ n25316);
assign n4173 = ~(n10980 ^ n5695);
assign n8657 = ~(n8457 ^ n23913);
assign n6942 = n4418 | n21018;
assign n2838 = n7048 | n13908;
assign n13104 = ~(n1836 ^ n5803);
assign n4909 = ~(n24939 ^ n24880);
assign n24562 = ~(n8067 | n11243);
assign n11596 = ~n8026;
assign n21703 = ~(n17090 | n27120);
assign n10781 = n3890 & n10384;
assign n19768 = n14130 | n1097;
assign n14855 = n20760 & n16151;
assign n18564 = n6444 | n4404;
assign n25865 = n23809 | n17209;
assign n17914 = n18381 | n22073;
assign n25622 = ~(n1875 ^ n21258);
assign n25486 = ~n11997;
assign n16001 = n8883 & n9624;
assign n25917 = ~(n17548 ^ n1620);
assign n25664 = n21517 | n16972;
assign n14409 = n14195 & n19874;
assign n22768 = n3984 & n22153;
assign n9220 = ~(n16804 ^ n22872);
assign n22256 = ~(n18925 | n15185);
assign n25288 = ~(n24557 ^ n15630);
assign n6228 = n13590 | n23529;
assign n19882 = ~(n17620 ^ n5330);
assign n14276 = ~n92;
assign n27074 = ~n4459;
assign n18585 = ~(n8830 ^ n11407);
assign n24764 = n647 | n6475;
assign n2221 = n18969 & n12206;
assign n11070 = ~(n24528 ^ n17487);
assign n7461 = n13367 | n20970;
assign n23350 = n24613 | n5269;
assign n15108 = ~(n20847 ^ n9415);
assign n5977 = ~(n24796 | n15536);
assign n267 = n1682 | n6427;
assign n18342 = n222 & n13396;
assign n5090 = ~(n427 ^ n22198);
assign n6558 = ~(n7993 ^ n23232);
assign n15704 = n5829 | n12344;
assign n18360 = ~n24756;
assign n14435 = n21678 | n684;
assign n1747 = n22232 | n19271;
assign n17714 = n19858 | n1984;
assign n11347 = ~(n10613 ^ n15721);
assign n16211 = ~n17077;
assign n949 = ~(n5209 ^ n21358);
assign n21088 = n21340 & n24266;
assign n15442 = ~n5207;
assign n21271 = n12562 & n12351;
assign n13994 = n18324 & n24308;
assign n25077 = n12840 & n26040;
assign n4280 = ~n4916;
assign n15889 = ~(n3550 ^ n2652);
assign n9660 = n24832 | n21050;
assign n7679 = ~(n23143 ^ n15783);
assign n26136 = ~(n21509 ^ n26090);
assign n20127 = ~n10141;
assign n17066 = ~n15282;
assign n26560 = n22537 | n15902;
assign n12624 = n26450 | n13088;
assign n23210 = n2868 | n13455;
assign n19383 = ~(n26244 ^ n17051);
assign n26141 = ~(n1569 ^ n4560);
assign n21952 = n6631 | n24732;
assign n19100 = n13748 | n22704;
assign n25150 = ~n23783;
assign n8938 = n24489 & n7848;
assign n26525 = n3813 | n8303;
assign n23393 = ~(n12878 ^ n22290);
assign n14801 = ~(n23944 ^ n2931);
assign n16121 = n4881 & n24888;
assign n16195 = n24646 & n4288;
assign n20896 = ~n8485;
assign n6214 = n18038 & n19627;
assign n7466 = ~(n7179 ^ n3229);
assign n1452 = n17747 & n21364;
assign n8388 = n20570 | n18474;
assign n4705 = n12416 & n11069;
assign n3991 = n23048 | n5795;
assign n26600 = ~(n7523 ^ n14440);
assign n15059 = n1587 & n13303;
assign n11309 = ~n21025;
assign n17450 = n9368 | n2297;
assign n23033 = n3815 & n12794;
assign n12651 = ~(n22335 | n14354);
assign n5028 = ~(n7188 ^ n21237);
assign n18398 = ~(n13201 ^ n1353);
assign n24271 = ~(n25913 ^ n15568);
assign n12628 = n16371 & n12523;
assign n4519 = ~(n10086 ^ n6175);
assign n12970 = n20708 | n1608;
assign n5749 = ~(n23506 ^ n19789);
assign n17780 = ~(n14427 ^ n78);
assign n21235 = ~(n4879 ^ n6460);
assign n4931 = n11157 & n8341;
assign n9930 = ~n21002;
assign n2557 = ~n16683;
assign n3294 = n144 | n21764;
assign n8016 = ~n19457;
assign n5063 = ~n5739;
assign n13586 = n10201 | n22379;
assign n23111 = ~(n23048 | n2872);
assign n5771 = ~(n3744 ^ n13990);
assign n18572 = ~(n8445 ^ n8488);
assign n15965 = ~(n1171 ^ n3407);
assign n5260 = ~(n14485 ^ n9483);
assign n23894 = ~(n8663 ^ n3708);
assign n17419 = n23436 & n21172;
assign n5942 = ~(n20766 ^ n21919);
assign n18235 = n1166 & n4187;
assign n2100 = ~n13216;
assign n5193 = ~(n26774 | n22177);
assign n17958 = ~(n20053 ^ n24984);
assign n5819 = ~(n12709 ^ n3776);
assign n24540 = ~(n7470 | n13696);
assign n12318 = n1182 | n11652;
assign n1830 = n4598 & n6771;
assign n26532 = n4999 & n27017;
assign n2198 = ~(n15850 ^ n4714);
assign n18640 = n20399 | n12695;
assign n8770 = ~(n17188 ^ n20225);
assign n21306 = ~n494;
assign n7572 = ~(n20228 ^ n27154);
assign n13920 = ~(n12464 | n20179);
assign n24146 = ~(n11453 ^ n21786);
assign n3868 = ~(n7334 | n5925);
assign n20830 = n9020 | n24957;
assign n537 = ~n5605;
assign n15171 = ~(n16696 ^ n8638);
assign n13975 = ~n15087;
assign n6190 = n5313 | n17156;
assign n3786 = ~(n9331 ^ n13794);
assign n423 = ~(n2090 ^ n11926);
assign n18273 = n6432 | n1045;
assign n1038 = n4035 | n14602;
assign n17885 = ~(n19230 ^ n11580);
assign n27175 = ~(n19778 ^ n6423);
assign n21430 = ~(n4732 ^ n5286);
assign n10815 = ~(n13349 | n13494);
assign n3875 = ~(n15271 ^ n26882);
assign n17154 = ~(n17835 ^ n8166);
assign n22740 = ~(n8088 | n8624);
assign n11998 = ~(n23209 ^ n4485);
assign n4692 = n15277;
assign n21414 = n5244 | n24340;
assign n17891 = ~(n725 ^ n17784);
assign n318 = n21438 | n2291;
assign n20600 = n832 & n19046;
assign n20988 = ~(n3984 | n7439);
assign n20065 = ~n23109;
assign n2831 = n23039 | n12734;
assign n25870 = ~(n11192 | n19805);
assign n1664 = n16728 | n21884;
assign n13306 = ~(n12956 | n11824);
assign n25217 = n26599 | n4343;
assign n20254 = n18603 & n13260;
assign n20263 = ~(n5668 ^ n1163);
assign n1998 = n17484 | n25141;
assign n17943 = n25282 & n25729;
assign n3585 = n9065 | n3667;
assign n9844 = n5624 | n14469;
assign n2388 = ~(n20310 ^ n551);
assign n17370 = ~(n16824 | n26295);
assign n19128 = ~n15250;
assign n176 = ~(n2886 | n1738);
assign n10455 = ~n13556;
assign n15733 = n8841 | n14780;
assign n132 = ~(n12762 ^ n3349);
assign n24187 = ~(n19765 ^ n19081);
assign n3770 = ~(n14497 ^ n23593);
assign n14754 = ~n17856;
assign n7190 = ~(n19491 ^ n6918);
assign n23961 = n13404 & n14169;
assign n8691 = n18122 & n6272;
assign n7081 = ~(n12855 ^ n13383);
assign n17420 = n23570 & n9265;
assign n16967 = ~n16739;
assign n25774 = n17273 | n26392;
assign n17624 = n17537 | n19280;
assign n3462 = n20313 & n11641;
assign n7103 = n19134 | n14385;
assign n9987 = ~(n18729 | n13081);
assign n20153 = ~(n11051 ^ n342);
assign n5554 = n6353 | n8434;
assign n12618 = n8068 | n4466;
assign n19210 = ~(n21339 ^ n19802);
assign n16862 = ~(n8732 ^ n9285);
assign n26226 = ~(n24750 ^ n7872);
assign n8004 = n2261 | n23653;
assign n15685 = n7902 & n13926;
assign n8418 = ~(n17310 ^ n23974);
assign n7909 = n14014 | n5189;
assign n25503 = ~(n8540 ^ n2399);
assign n6795 = n7893 | n26876;
assign n14598 = ~n17928;
assign n13021 = ~(n11044 ^ n4325);
assign n3660 = n4132 | n23849;
assign n23123 = ~(n14306 ^ n10389);
assign n16861 = n10788 | n21451;
assign n2161 = ~(n23700 ^ n26765);
assign n9627 = ~(n6385 | n18171);
assign n20382 = ~(n13246 ^ n15039);
assign n7220 = n11885 | n5361;
assign n6186 = n2146 & n20216;
assign n24830 = n21773 & n3375;
assign n18300 = ~n12546;
assign n17349 = n10903 | n20271;
assign n25436 = n9995 & n21677;
assign n7984 = n24516 | n2448;
assign n11619 = ~(n6502 ^ n19494);
assign n11691 = n22554 & n2628;
assign n21213 = ~n3382;
assign n3254 = n4684 | n7183;
assign n8947 = ~(n3134 ^ n16285);
assign n7771 = n18529 & n3858;
assign n26139 = n23244 & n1801;
assign n21554 = n25291 | n7061;
assign n23458 = n10598 | n26360;
assign n13782 = n18100 | n14155;
assign n12419 = ~(n19345 ^ n25574);
assign n19582 = n6568 | n7055;
assign n7805 = ~(n9349 ^ n15547);
assign n12333 = n24234 & n15460;
assign n12859 = ~n22960;
assign n19090 = ~n10903;
assign n1605 = ~n14384;
assign n680 = n16711 | n11011;
assign n24997 = n18172 | n26278;
assign n1450 = ~(n12057 ^ n24638);
assign n17388 = ~(n20636 ^ n5214);
assign n15569 = n14332 & n7916;
assign n4137 = n4242 | n17388;
assign n14599 = ~(n22470 ^ n11455);
assign n2808 = ~n8918;
assign n4796 = ~(n21997 | n18483);
assign n14892 = n141 | n7245;
assign n3134 = ~n20291;
assign n11949 = ~(n13976 ^ n23895);
assign n14065 = n3766 | n6074;
assign n17389 = n25821 & n15510;
assign n21551 = n88 | n14447;
assign n15700 = n9574 | n13623;
assign n21142 = ~(n2782 ^ n1387);
assign n20277 = n2371 & n14713;
assign n19469 = ~n6502;
assign n21958 = n13290 | n10730;
assign n10638 = ~(n3260 ^ n21832);
assign n14262 = n2407 | n7538;
assign n8825 = ~(n10785 ^ n19042);
assign n26899 = ~(n16803 | n25700);
assign n16481 = ~(n25488 ^ n17215);
assign n3347 = ~n20055;
assign n14274 = ~(n2748 ^ n13808);
assign n2538 = n13686 & n20034;
assign n534 = n26732 & n19434;
assign n9253 = n1718 & n20735;
assign n9480 = n7766 & n5992;
assign n4505 = ~(n5196 | n1878);
assign n13327 = ~(n19184 | n14580);
assign n2580 = n20638 & n10512;
assign n14469 = ~n6553;
assign n9618 = n24649 | n4426;
assign n10560 = n9979 | n25948;
assign n22444 = ~(n21840 ^ n1555);
assign n10103 = n21607 | n12726;
assign n1705 = ~(n16404 ^ n7323);
assign n10662 = n20214 | n23241;
assign n27061 = n25324 | n5951;
assign n18759 = ~n22380;
assign n17845 = ~(n25046 ^ n23473);
assign n24215 = n22436 & n100;
assign n17850 = n1975 & n26527;
assign n1757 = ~(n3894 ^ n14993);
assign n8848 = ~(n20059 ^ n216);
assign n15152 = ~(n19175 ^ n16880);
assign n5057 = ~(n17578 ^ n8653);
assign n14225 = ~(n17613 ^ n10593);
assign n20297 = ~(n19144 | n20210);
assign n281 = n2146 | n22455;
assign n7137 = ~n22092;
assign n25857 = n6230 | n25235;
assign n8476 = n27091 | n19317;
assign n2029 = n22506 | n6047;
assign n21265 = n14323 | n12351;
assign n7879 = ~n14192;
assign n6299 = ~(n12354 ^ n12121);
assign n13250 = n12134 | n21092;
assign n11948 = n5950 | n17893;
assign n19994 = n21454 & n4838;
assign n12985 = ~(n17242 ^ n336);
assign n11683 = n11522 | n9327;
assign n27189 = ~n23120;
assign n12697 = ~n4045;
assign n22375 = ~(n9703 ^ n25871);
assign n3095 = n17542 | n24402;
assign n13268 = ~(n25738 | n11314);
assign n11329 = n13986 & n23093;
assign n8385 = ~n1047;
assign n19296 = ~(n26486 ^ n2816);
assign n3892 = n3124 | n21832;
assign n16592 = n15923 | n9817;
assign n26456 = n23786 | n20942;
assign n9949 = n18000 | n4732;
assign n6723 = n13844 | n7516;
assign n26848 = ~(n3140 | n14103);
assign n3957 = ~(n7939 | n2925);
assign n17222 = n5262 | n22712;
assign n19189 = n3879 | n15978;
assign n14887 = ~(n22194 | n19116);
assign n17612 = ~(n5050 ^ n1558);
assign n3569 = n25491 & n26389;
assign n18170 = n5360 | n21340;
assign n12104 = ~(n11248 ^ n26318);
assign n25495 = n12150 & n11699;
assign n24100 = ~(n12098 ^ n21522);
assign n18944 = n19910 & n18822;
assign n12187 = n22324 & n18532;
assign n15430 = n26582 & n7107;
assign n21922 = n21127 | n20244;
assign n5943 = ~(n2701 ^ n9005);
assign n23092 = ~n9747;
assign n13042 = ~n24095;
assign n22880 = ~n23331;
assign n26611 = n13479 | n20343;
assign n27 = ~n17308;
assign n5691 = n12712 | n3003;
assign n8229 = ~(n14514 ^ n3694);
assign n11239 = ~(n21021 ^ n3253);
assign n14110 = ~(n26268 ^ n26285);
assign n3047 = n23099 | n24444;
assign n24163 = n21038 | n24645;
assign n26172 = n3136 & n11542;
assign n2109 = n15071 | n19748;
assign n13936 = ~(n26202 ^ n10712);
assign n22792 = ~(n27060 | n25543);
assign n5862 = ~(n19839 ^ n19979);
assign n5299 = ~n24922;
assign n6213 = n16892 & n14686;
assign n3599 = ~(n16544 | n4319);
assign n18971 = ~n801;
assign n4073 = ~(n10024 | n7347);
assign n8535 = ~(n1333 ^ n15927);
assign n1212 = ~(n17090 | n22173);
assign n18133 = ~(n914 ^ n26167);
assign n7293 = n18100 & n14569;
assign n15081 = ~(n13425 ^ n23580);
assign n25148 = n17027 & n23206;
assign n9924 = ~n16339;
assign n2988 = n23010 | n11139;
assign n23031 = n24078 | n21130;
assign n12160 = ~n16521;
assign n5416 = ~(n19841 ^ n25140);
assign n24659 = ~(n22588 | n13112);
assign n12631 = ~(n25038 | n22442);
assign n5621 = ~n15355;
assign n10906 = ~(n24042 ^ n17635);
assign n14133 = ~n15967;
assign n8800 = n22834 | n903;
assign n22393 = ~(n20409 ^ n18227);
assign n21124 = n3909 | n24200;
assign n17494 = ~(n11321 | n6703);
assign n12324 = ~(n24882 ^ n17312);
assign n5011 = ~(n18342 ^ n23045);
assign n13881 = ~(n25106 ^ n20921);
assign n6576 = ~(n25116 ^ n9346);
assign n951 = ~(n8964 | n1293);
assign n15347 = n7102 | n280;
assign n1540 = ~n23831;
assign n10374 = n26483 & n12088;
assign n2451 = n4462 | n26286;
assign n15064 = ~(n24058 ^ n21287);
assign n14858 = ~(n8155 | n767);
assign n12032 = n6376 & n18939;
assign n11343 = n13822 | n15077;
assign n16468 = ~n25261;
assign n6167 = n22713 | n7738;
assign n11471 = ~(n23018 ^ n11615);
assign n18793 = ~(n26818 ^ n14164);
assign n20369 = n8722 & n10791;
assign n10587 = ~(n18171 | n24529);
assign n2317 = n1254 & n9056;
assign n9902 = n20208 | n6732;
assign n13570 = n25272 & n9785;
assign n13057 = ~n3014;
assign n18997 = n5953 & n13211;
assign n19037 = ~n932;
assign n15238 = n18148 & n12906;
assign n11711 = ~n11473;
assign n4843 = n26552 | n3337;
assign n5998 = ~n25946;
assign n15805 = ~n1227;
assign n21557 = n12576 | n23463;
assign n12755 = n23489 | n22766;
assign n7371 = n19554 & n4281;
assign n7388 = ~(n12398 ^ n23586);
assign n22731 = ~(n26241 | n12587);
assign n15036 = ~(n11989 ^ n14087);
assign n6987 = n24862 | n14488;
assign n14908 = n25875 | n4852;
assign n4872 = ~(n14315 ^ n18626);
assign n162 = ~(n25430 ^ n8116);
assign n27081 = n6 | n21040;
assign n21522 = ~(n24087 ^ n20364);
assign n20985 = n18569 & n14635;
assign n1610 = n3090 & n16792;
assign n9912 = n10050 | n17669;
assign n16656 = ~(n8817 ^ n12440);
assign n26526 = n26495 | n26853;
assign n483 = ~n1881;
assign n8005 = n1444 | n3898;
assign n18821 = n545 | n519;
assign n11120 = ~(n19786 ^ n22448);
assign n1361 = n14714 | n3583;
assign n26850 = n18400 | n6270;
assign n26417 = n26303;
assign n17133 = n17632 | n16702;
assign n5345 = n15474 | n21839;
assign n18724 = ~(n11614 ^ n9454);
assign n16214 = ~(n16661 ^ n23410);
assign n23546 = ~(n4385 ^ n25814);
assign n17823 = n1443 | n7673;
assign n125 = ~n16619;
assign n9911 = n733 | n25067;
assign n8380 = ~(n8691 ^ n22546);
assign n24821 = ~n18337;
assign n16969 = ~(n18869 ^ n10741);
assign n10845 = n18986 | n2523;
assign n20035 = n5696 | n7871;
assign n17495 = ~n9269;
assign n8781 = ~(n23369 | n26572);
assign n22883 = n9840 | n20939;
assign n1078 = n17974 | n13025;
assign n7711 = ~(n25074 ^ n6556);
assign n25378 = n11678 & n6428;
assign n3337 = ~(n11767 ^ n18553);
assign n5536 = n24341 | n6848;
assign n15033 = ~(n24883 ^ n21696);
assign n22605 = n9671 | n12964;
assign n25861 = ~(n22515 ^ n12341);
assign n1750 = ~(n20408 ^ n23543);
assign n14399 = ~(n11736 ^ n22470);
assign n5500 = ~(n23697 ^ n9967);
assign n12565 = ~n3631;
assign n10521 = n24917 & n26983;
assign n22257 = n22800 & n8075;
assign n16391 = n10252 | n6102;
assign n6812 = n19298 | n21038;
assign n21484 = n3720 & n17262;
assign n12396 = ~n15546;
assign n14986 = ~(n4278 ^ n18687);
assign n13481 = n9365 | n1334;
assign n2709 = ~(n6319 | n19836);
assign n19903 = ~(n21972 | n9942);
assign n1950 = n21649 & n20192;
assign n4516 = n10576 | n11664;
assign n6480 = ~(n4685 ^ n21777);
assign n12413 = ~(n26722 ^ n18687);
assign n3058 = ~(n5201 | n9932);
assign n22814 = ~(n4719 | n12453);
assign n6396 = n582 & n3163;
assign n519 = n19288 & n12213;
assign n12036 = ~(n15008 ^ n15979);
assign n24208 = ~n24154;
assign n6138 = ~(n22032 ^ n17866);
assign n20968 = n6193 & n10070;
assign n10659 = ~n10712;
assign n12002 = ~n20250;
assign n26194 = ~(n9880 ^ n13714);
assign n1254 = n2818 | n21390;
assign n14738 = ~(n24907 ^ n5822);
assign n19263 = ~(n3277 ^ n13628);
assign n23089 = ~(n2727 ^ n12214);
assign n22042 = ~(n25475 | n13463);
assign n24476 = ~(n16526 ^ n4310);
assign n21949 = n17688 | n17389;
assign n23938 = n3047 & n10724;
assign n10891 = n15298 | n14855;
assign n9694 = ~(n26797 ^ n15077);
assign n8516 = n21101 | n13301;
assign n13941 = ~(n26379 ^ n19363);
assign n10438 = ~(n3299 | n17141);
assign n1266 = ~(n24868 ^ n13747);
assign n25196 = n12599 & n23777;
assign n11784 = ~n21286;
assign n11043 = ~n25629;
assign n16789 = n25570 | n21747;
assign n20286 = n23668 | n11769;
assign n10347 = ~(n22862 ^ n17663);
assign n14763 = ~(n10997 ^ n26619);
assign n14287 = n694 & n6217;
assign n5581 = ~(n22034 ^ n7476);
assign n22971 = ~(n5793 | n23710);
assign n21600 = n1720 | n26212;
assign n23224 = n7010 | n1547;
assign n22770 = ~(n15636 | n24618);
assign n16325 = ~n21240;
assign n2051 = ~(n23712 ^ n16753);
assign n5200 = ~(n19190 ^ n223);
assign n9879 = ~(n20146 ^ n5253);
assign n19126 = n3396 | n9397;
assign n4045 = ~(n11850 ^ n21189);
assign n27063 = n14633 & n2886;
assign n5657 = ~n13781;
assign n6443 = ~(n10451 ^ n13677);
assign n16966 = n2455 & n16564;
assign n13788 = ~(n2436 ^ n20391);
assign n6682 = ~n3253;
assign n21483 = ~(n14241 | n7418);
assign n23180 = ~(n10978 ^ n25126);
assign n6762 = n21632 & n19423;
assign n22448 = ~(n11714 ^ n10861);
assign n21929 = ~n21016;
assign n22250 = n22017 & n22671;
assign n3020 = ~(n24430 ^ n19908);
assign n9547 = ~(n15291 ^ n13401);
assign n3318 = ~n6427;
assign n22295 = ~n13241;
assign n8002 = ~n1483;
assign n6065 = ~(n18783 ^ n25908);
assign n26067 = ~(n23253 | n26641);
assign n16630 = ~(n11984 ^ n25815);
assign n25466 = n20411 & n17212;
assign n7993 = n26626 & n3073;
assign n14310 = ~(n13305 ^ n5377);
assign n9596 = n22065 | n9234;
assign n8566 = ~(n17826 | n329);
assign n13322 = n26294 | n15587;
assign n21408 = n9828 | n11979;
assign n25005 = n20142 | n17506;
assign n568 = n25912 & n18104;
assign n6302 = ~(n8378 ^ n10633);
assign n14074 = ~(n21739 ^ n704);
assign n9260 = n24054 & n14032;
assign n4177 = ~n12271;
assign n4814 = n739 | n4385;
assign n3363 = ~n16029;
assign n3707 = ~n12733;
assign n3348 = n20425 | n15498;
assign n18301 = ~(n26638 ^ n18933);
assign n21941 = ~n13161;
assign n7306 = ~(n2858 | n13907);
assign n20622 = n18662 | n9967;
assign n19048 = ~n20833;
assign n16583 = ~(n16833 ^ n18963);
assign n10154 = n9782 | n17520;
assign n18478 = ~(n13853 ^ n12274);
assign n6207 = ~(n7099 ^ n23068);
assign n20482 = ~n17541;
assign n14366 = ~(n10524 ^ n58);
assign n7474 = ~(n7170 ^ n11945);
assign n5846 = ~(n21929 | n6127);
assign n19521 = ~(n22735 ^ n21244);
assign n8513 = n16233 & n25566;
assign n11282 = n26996 & n6657;
assign n14052 = ~n9069;
assign n19579 = ~(n8614 | n12702);
assign n17597 = ~n24213;
assign n6570 = n13547 | n15601;
assign n3889 = n24945 & n1516;
assign n20423 = n19298 | n5816;
assign n7629 = n8878 | n19122;
assign n12668 = n4630 & n1073;
assign n21939 = n22281 | n26332;
assign n13258 = n20645 | n22577;
assign n24353 = ~(n5206 ^ n3990);
assign n8199 = n2217 & n15038;
assign n6024 = ~(n7893 | n18569);
assign n1397 = n5872 & n7945;
assign n17558 = n15156 & n21048;
assign n3651 = ~(n11890 ^ n27127);
assign n27005 = ~(n22173 ^ n583);
assign n9936 = n24315 | n8268;
assign n21776 = n22664 | n13524;
assign n6728 = ~(n5509 | n21363);
assign n22861 = n21900;
assign n14862 = n8568 | n13140;
assign n11879 = n2745 & n4637;
assign n26109 = ~(n14133 ^ n7293);
assign n12877 = ~(n10170 ^ n19217);
assign n25863 = ~(n3909 | n19081);
assign n25491 = n5119 | n6070;
assign n12835 = ~(n22379 ^ n15077);
assign n15456 = ~n21430;
assign n1827 = n25673 & n7512;
assign n15822 = ~(n12351 ^ n12562);
assign n22078 = ~(n25643 ^ n329);
assign n11883 = n17384 | n21077;
assign n17464 = n13577 | n19229;
assign n7541 = n2056 | n6104;
assign n19299 = n27006 | n7197;
assign n5505 = ~n15732;
assign n8125 = n17826 | n26660;
assign n19199 = n4286 | n14562;
assign n21604 = ~(n6729 ^ n11192);
assign n20570 = n11491 ^ n13826;
assign n20460 = n12326 & n8446;
assign n9051 = ~(n24102 ^ n860);
assign n2686 = ~(n18262 ^ n18341);
assign n12622 = ~(n5992 ^ n2456);
assign n10187 = ~(n9402 ^ n2439);
assign n22039 = n19898 | n17455;
assign n21755 = ~(n506 ^ n5386);
assign n13029 = n25559 & n15714;
assign n8661 = ~(n3287 ^ n8573);
assign n90 = ~(n6442 ^ n25265);
assign n2283 = ~(n13649 ^ n5842);
assign n18317 = ~(n7532 ^ n8745);
assign n11141 = n16054 | n17600;
assign n26292 = ~n21352;
assign n3590 = ~(n25064 ^ n26427);
assign n20462 = n7387;
assign n9430 = ~(n19787 ^ n10643);
assign n26030 = ~n13853;
assign n1023 = ~(n18495 ^ n2252);
assign n5372 = n24192 & n929;
assign n15535 = ~(n2385 ^ n7130);
assign n7445 = n9172 | n13665;
assign n9988 = ~n25336;
assign n5452 = n5966 & n13394;
assign n3639 = ~n6474;
assign n19094 = ~n24374;
assign n8809 = ~(n21376 ^ n4649);
assign n5435 = ~(n17255 ^ n17597);
assign n462 = n11501 & n25509;
assign n26373 = n11631 & n7398;
assign n11590 = n24828 | n19368;
assign n19307 = ~(n2409 ^ n7057);
assign n20992 = n1933 | n21200;
assign n2627 = n9438 | n22192;
assign n4926 = n8539 & n14610;
assign n24119 = ~(n8502 ^ n15488);
assign n11363 = ~n7963;
assign n9386 = n18995 | n7693;
assign n14120 = ~(n1403 ^ n5284);
assign n10327 = ~(n22184 ^ n11426);
assign n15670 = n26565 | n10787;
assign n11690 = ~(n5006 | n21117);
assign n11022 = ~(n23209 ^ n1319);
assign n16098 = ~(n23547 ^ n25569);
assign n11614 = n9251 & n8344;
assign n5407 = ~n21735;
assign n13852 = n320 | n4906;
assign n1384 = n1142 & n10294;
assign n12516 = ~(n24466 ^ n13595);
assign n11231 = n11828 | n14032;
assign n14810 = ~(n8352 ^ n12859);
assign n16100 = n4012 | n14264;
assign n25654 = ~(n5143 | n9337);
assign n24511 = ~(n18615 ^ n25872);
assign n7361 = n26866;
assign n15703 = ~(n19967 | n8245);
assign n24710 = n4022 | n1009;
assign n23357 = n8310 | n10309;
assign n18460 = n18077 | n11782;
assign n17861 = n6851 | n2656;
assign n19592 = ~n18793;
assign n502 = ~(n8481 ^ n11998);
assign n21132 = ~(n13490 ^ n10739);
assign n8411 = ~n11525;
assign n2825 = n7832 | n9527;
assign n1106 = ~n3447;
assign n16515 = n9259 & n12423;
assign n10295 = ~(n25657 ^ n11091);
assign n19826 = n8520 | n4375;
assign n8449 = n5793 | n20361;
assign n4055 = n19092 & n23734;
assign n6460 = ~(n7335 ^ n4319);
assign n7082 = n15913 | n2037;
assign n17720 = n25101 ^ n27075;
assign n13465 = n11748 & n7009;
assign n1343 = n18269 & n12354;
assign n25569 = n13049 | n5463;
assign n23854 = ~n20898;
assign n16447 = ~(n22110 ^ n25485);
assign n18937 = n8163 | n7173;
assign n1235 = n13912 | n11098;
assign n2964 = ~(n24429 ^ n8314);
assign n26301 = n7303 & n22946;
assign n4383 = ~(n4160 | n12770);
assign n20995 = n23351 | n24833;
assign n6697 = ~(n5689 | n11864);
assign n11303 = ~n8964;
assign n21415 = n17347 | n13939;
assign n14760 = ~n19404;
assign n24968 = n6882 | n719;
assign n23384 = n20420 & n23761;
assign n7850 = n16722 | n16165;
assign n25221 = ~(n3583 ^ n20328);
assign n1526 = ~(n8425 | n16184);
assign n24535 = ~(n20687 | n8415);
assign n4448 = ~(n17795 ^ n15051);
assign n8313 = ~(n9036 ^ n18878);
assign n3907 = ~(n7593 | n5101);
assign n26057 = n16085 | n14160;
assign n11782 = n753 & n20026;
assign n21720 = n4347 | n22916;
assign n6919 = ~(n12650 | n14765);
assign n12355 = ~(n18749 ^ n11980);
assign n21241 = n7348 | n4435;
assign n24647 = ~(n19062 | n14105);
assign n22853 = n2798 | n2319;
assign n5990 = ~n7338;
assign n19709 = ~(n20895 ^ n13373);
assign n15637 = n26841 & n7011;
assign n7372 = ~(n16672 ^ n302);
assign n4024 = ~(n26695 ^ n3742);
assign n24033 = n15503 | n8128;
assign n17052 = ~(n15442 | n17382);
assign n22192 = n18374 & n22966;
assign n26749 = ~(n14265 | n15445);
assign n1418 = ~(n7953 ^ n20908);
assign n19728 = ~(n6718 ^ n1611);
assign n19192 = ~n25261;
assign n22099 = ~(n12880 ^ n18446);
assign n26499 = ~n12973;
assign n19954 = n6726 | n18202;
assign n5782 = ~(n18009 ^ n13466);
assign n10413 = ~(n23878 | n5139);
assign n14415 = ~n15271;
assign n10449 = n10825 & n9304;
assign n17734 = ~n26641;
assign n22890 = n19875 | n9737;
assign n8832 = n24369 & n25894;
assign n19517 = ~(n7082 ^ n20593);
assign n17770 = ~n10232;
assign n14638 = n5159 | n11377;
assign n25497 = n20805 & n16289;
assign n27100 = ~(n12854 ^ n26867);
assign n1282 = n13719 | n22342;
assign n24442 = n9294 | n17568;
assign n21010 = n17098 | n12622;
assign n21860 = ~(n23952 ^ n4631);
assign n14596 = ~(n27203 | n24959);
assign n16395 = n353 | n22119;
assign n15871 = n25122 | n13349;
assign n22204 = ~(n5112 | n20954);
assign n1819 = ~(n22305 ^ n17102);
assign n104 = ~n17380;
assign n2186 = n16620 | n15599;
assign n14170 = ~(n7824 ^ n16654);
assign n22718 = n14718 | n20920;
assign n12586 = ~n21293;
assign n12969 = n1018 | n22306;
assign n26379 = n23560 | n21069;
assign n341 = n407 | n9717;
assign n19849 = ~n19163;
assign n15676 = ~(n24018 | n5400);
assign n24105 = ~(n11571 ^ n4725);
assign n19927 = ~(n7184 | n20564);
assign n2569 = n11628 | n2166;
assign n12752 = n15925 | n1123;
assign n619 = ~(n4348 ^ n13157);
assign n19298 = ~n583;
assign n6615 = n11581 | n14994;
assign n7123 = n23602 | n820;
assign n25814 = n26402 | n11879;
assign n10960 = n7185 & n5698;
assign n26991 = n5067 | n8344;
assign n21069 = n8081 & n21619;
assign n26616 = n14873 | n3644;
assign n12599 = n12258 | n1626;
assign n5952 = ~(n23566 | n9457);
assign n23931 = n612 & n17329;
assign n8864 = n6953 | n7282;
assign n20742 = n26180 | n24700;
assign n11153 = n22977 | n20923;
assign n22338 = n13892 & n16974;
assign n10318 = n5226 & n21205;
assign n9814 = ~n4675;
assign n9210 = ~(n12491 ^ n8154);
assign n21570 = ~(n20468 ^ n13453);
assign n16953 = n25463 | n20526;
assign n24505 = n15378 | n10039;
assign n11707 = n13349 & n24422;
assign n23471 = ~(n9629 ^ n1431);
assign n26034 = n3094 | n6284;
assign n24137 = n14647 & n23381;
assign n6721 = ~(n22644 | n10642);
assign n20032 = ~n19005;
assign n26681 = ~(n20580 ^ n19727);
assign n17385 = ~(n23863 | n25381);
assign n5263 = ~(n13130 ^ n24491);
assign n1857 = ~(n15404 ^ n18599);
assign n25375 = ~(n5443 ^ n1320);
assign n10708 = n8096 & n14748;
assign n14135 = ~(n17881 ^ n8067);
assign n9289 = ~(n14569 ^ n24732);
assign n15357 = n5122 | n12395;
assign n8460 = n12524 | n1287;
assign n4574 = ~n26180;
assign n6796 = n212 | n2783;
assign n8128 = n8967 & n26533;
assign n2083 = ~(n20970 ^ n12961);
assign n10220 = ~n17671;
assign n15308 = n25447 & n770;
assign n20244 = ~(n4588 ^ n22201);
assign n25285 = n16772 & n14286;
assign n4596 = ~(n23832 ^ n19238);
assign n14441 = ~(n7421 | n13206);
assign n9848 = n24357 | n3699;
assign n9546 = ~(n8614 | n21698);
assign n8609 = ~n24499;
assign n24420 = ~n25696;
assign n16932 = ~(n11802 | n7627);
assign n25724 = ~n26866;
assign n11679 = ~(n14774 | n26300);
assign n236 = n7973 & n15179;
assign n6192 = ~(n20036 | n22515);
assign n21425 = ~(n6865 ^ n6703);
assign n684 = ~n24616;
assign n26718 = ~(n22828 ^ n379);
assign n16429 = ~(n25772 | n21596);
assign n23341 = ~(n10270 ^ n13801);
assign n24776 = n3579 & n5667;
assign n17608 = n328 | n19387;
assign n9592 = ~(n1831 | n10250);
assign n5844 = ~(n16846 ^ n24101);
assign n4546 = n708 | n2781;
assign n14181 = ~(n3707 ^ n12802);
assign n19428 = n21272 | n8769;
assign n12980 = ~(n8725 ^ n15065);
assign n11815 = n13868 & n6441;
assign n25167 = n11612 & n27085;
assign n23891 = n12521 & n3787;
assign n18169 = n12091 | n25076;
assign n20776 = n2849 & n20641;
assign n3004 = n11001 & n22611;
assign n24998 = ~(n23933 ^ n17269);
assign n18046 = ~(n15097 ^ n6893);
assign n946 = ~(n13633 ^ n13171);
assign n12480 = n22515 & n10467;
assign n8562 = ~(n26695 | n22588);
assign n8528 = ~n6333;
assign n25950 = n26633 | n2900;
assign n8348 = ~(n13172 | n16252);
assign n25412 = ~(n5099 ^ n14216);
assign n4557 = n22396 | n17980;
assign n13596 = ~(n24032 ^ n22843);
assign n26051 = n19214 | n13705;
assign n24850 = ~n26882;
assign n12984 = n24890 & n18303;
assign n6131 = ~n18487;
assign n5938 = ~n6229;
assign n5755 = n5666 | n5232;
assign n22921 = n7381 & n16198;
assign n11689 = n6534 & n7009;
assign n11867 = n6854 & n26702;
assign n19663 = ~(n14060 ^ n6287);
assign n5285 = ~(n1544 ^ n7052);
assign n6023 = ~(n21226 | n586);
assign n22779 = ~(n6472 ^ n12938);
assign n21883 = ~(n3356 | n16311);
assign n1403 = ~n25470;
assign n6690 = n22001 & n3886;
assign n20484 = ~(n4665 ^ n8309);
assign n21337 = ~n8250;
assign n19174 = ~(n1607 ^ n3234);
assign n24470 = ~(n23572 | n18474);
assign n6868 = n25610 | n10984;
assign n3673 = ~(n26861 ^ n22160);
assign n7585 = ~(n627 ^ n4166);
assign n21773 = n21134 | n4930;
assign n22427 = ~(n8918 ^ n19365);
assign n1762 = n3346 & n8044;
assign n20654 = n7524 & n14133;
assign n2242 = ~n6498;
assign n22438 = n26391 | n2009;
assign n17896 = n16427 | n17888;
assign n24973 = ~(n18539 ^ n3366);
assign n23832 = ~n18201;
assign n1835 = ~(n19745 ^ n15160);
assign n26272 = n22197 | n21164;
assign n6830 = n5471 & n2864;
assign n832 = ~n19789;
assign n23042 = n26670 | n2206;
assign n1017 = n6177 | n22833;
assign n10758 = ~n20570;
assign n5276 = ~(n11011 | n20179);
assign n1301 = ~(n4873 ^ n23272);
assign n3701 = n2777 | n11517;
assign n23474 = ~(n342 | n26789);
assign n9806 = ~(n20735 ^ n3463);
assign n16682 = ~(n13342 ^ n25660);
assign n5121 = n25903 | n9659;
assign n787 = ~(n2383 | n15236);
assign n22622 = ~(n18452 | n6397);
assign n1725 = ~(n4844 | n13708);
assign n21582 = n13026 | n13906;
assign n4074 = n24236 & n19289;
assign n303 = ~(n832 ^ n19046);
assign n21427 = n23708 & n6013;
assign n7663 = n22223 | n731;
assign n8914 = n14991 | n24638;
assign n1383 = ~(n7389 | n7531);
assign n17266 = ~n7569;
assign n4571 = n7458 & n4763;
assign n16472 = ~(n11560 | n7080);
assign n8984 = n8166 | n7554;
assign n22130 = ~(n14103 ^ n19402);
assign n2180 = n13976 & n25419;
assign n10607 = n1224 | n10727;
assign n20686 = n26107 | n21636;
assign n23642 = ~n19240;
assign n814 = n889 | n13874;
assign n26314 = ~(n19457 | n1753);
assign n19545 = ~n18507;
assign n4634 = ~(n3480 ^ n19911);
assign n12330 = ~(n7173 ^ n13511);
assign n8555 = n17690 | n17235;
assign n24840 = ~(n14667 ^ n804);
assign n8979 = ~n21779;
assign n7467 = ~(n10406 ^ n8947);
assign n26665 = ~(n18737 ^ n2328);
assign n14809 = ~(n17579 ^ n12452);
assign n25242 = n3740 | n23683;
assign n1273 = ~(n25915 | n8024);
assign n25251 = n10930 ^ n10626;
assign n14228 = ~(n18690 | n1183);
assign n20207 = ~(n3498 ^ n3740);
assign n16082 = ~(n2291 ^ n21438);
assign n11459 = ~(n8064 ^ n1240);
assign n10160 = n21651 & n18460;
assign n2518 = ~(n11327 ^ n26752);
assign n6433 = ~(n13926 ^ n25864);
assign n58 = ~(n22660 ^ n11011);
assign n15404 = ~(n21109 ^ n5224);
assign n6957 = n8990 | n13108;
assign n4871 = ~(n19157 | n22793);
assign n623 = ~n25008;
assign n126 = ~n23801;
assign n18818 = ~(n16205 | n23068);
assign n5675 = ~n26303;
assign n8353 = n3386 & n22742;
assign n4648 = n15945 & n25824;
assign n24433 = ~(n21420 ^ n11086);
assign n21017 = ~(n26115 ^ n16898);
assign n20642 = ~(n9003 | n13453);
assign n22746 = n5766 | n12382;
assign n20211 = ~(n23273 | n10435);
assign n7710 = n5115 | n2548;
assign n4328 = n17921 & n4402;
assign n13999 = ~(n12587 | n10608);
assign n19091 = n12649 | n7865;
assign n16870 = ~(n9934 ^ n2272);
assign n19265 = ~n24156;
assign n3143 = ~(n24865 ^ n11040);
assign n24789 = n13238 & n17058;
assign n12423 = ~(n26039 ^ n9554);
assign n1574 = ~n8661;
assign n19025 = ~n13074;
assign n4511 = n5355 | n5000;
assign n8343 = ~n22253;
assign n4081 = ~(n9655 | n22700);
assign n3759 = n12042 & n11308;
assign n10549 = ~(n21737 ^ n24020);
assign n2719 = ~(n13357 ^ n11077);
assign n16877 = ~(n1095 | n1367);
assign n13868 = n9550 | n16203;
assign n1487 = n14329 & n26157;
assign n11452 = ~n20179;
assign n4683 = ~(n18754 | n19245);
assign n23700 = n26448 | n2200;
assign n25513 = ~(n5965 ^ n11241);
assign n20183 = n6743 | n5969;
assign n17013 = ~n24879;
assign n11245 = ~(n16749 ^ n20418);
assign n8201 = n23049 & n10621;
assign n4399 = n1661 & n15106;
assign n541 = n10862 & n26005;
assign n24871 = n22959 | n2529;
assign n12675 = ~n6894;
assign n24592 = ~(n27053 ^ n19501);
assign n12904 = n4208 | n20083;
assign n23101 = n21531 & n25098;
assign n6871 = ~(n9535 | n11846);
assign n15562 = ~n19097;
assign n9961 = ~(n21305 ^ n7544);
assign n16273 = ~(n11694 ^ n25810);
assign n10287 = ~(n9743 ^ n10296);
assign n23204 = n6190 & n21870;
assign n19311 = ~(n23906 ^ n8846);
assign n111 = ~n22738;
assign n8102 = n8501 | n25809;
assign n25527 = ~(n27199 | n6861);
assign n9899 = ~(n17458 | n20687);
assign n10919 = ~(n9582 ^ n299);
assign n7125 = n13682 & n22357;
assign n7178 = n7995 & n18917;
assign n20591 = n10189 & n23975;
assign n21453 = n157 | n16235;
assign n19519 = n859 | n24982;
assign n13703 = ~(n21567 ^ n3306);
assign n8632 = ~(n7524 ^ n19680);
assign n7205 = ~n4314;
assign n27066 = ~n6949;
assign n19024 = ~(n27037 | n13775);
assign n6665 = n22786 & n2921;
assign n11847 = ~(n21733 | n1753);
assign n9801 = n19157 | n6555;
assign n13639 = n13126 | n25103;
assign n19684 = n17115 | n2418;
assign n19957 = n22252 | n15256;
assign n13301 = ~n2586;
assign n20485 = ~(n21624 ^ n20944);
assign n2820 = ~n15124;
assign n3353 = n17292 | n5078;
assign n11118 = ~n21284;
assign n19022 = n12048 | n11688;
assign n18571 = ~(n12875 ^ n22492);
assign n2128 = n15419 & n12087;
assign n12244 = n11579 | n3962;
assign n8116 = n12933 | n4987;
assign n6404 = n25068 | n10620;
assign n8897 = ~n1893;
assign n26370 = ~(n20150 | n26187);
assign n20907 = ~n4748;
assign n8382 = ~(n6083 ^ n9922);
assign n16987 = n3959 | n25917;
assign n10530 = n16839 | n19030;
assign n24408 = n20615 & n20225;
assign n22127 = n12116 | n10742;
assign n11932 = n25698 | n10674;
assign n20972 = ~n5324;
assign n2926 = ~n1092;
assign n23347 = ~(n4894 | n2566);
assign n8433 = n19469 | n25625;
assign n5645 = ~(n23110 | n7058);
assign n23753 = ~(n9586 | n3279);
assign n16449 = ~(n5080 ^ n11262);
assign n4453 = n8455 | n24835;
assign n16981 = n12259 | n7197;
assign n26011 = n1127 | n17528;
assign n2429 = ~(n4111 ^ n17723);
assign n8371 = ~(n2749 ^ n25464);
assign n23184 = ~(n17819 | n23970);
assign n10612 = ~(n4256 ^ n18483);
assign n26800 = ~(n7787 ^ n10333);
assign n17625 = ~(n167 ^ n3554);
assign n12836 = ~(n17993 ^ n7674);
assign n15596 = n3068 & n17521;
assign n23840 = n11642 & n16042;
assign n13398 = n10276 | n23654;
assign n20324 = ~(n17454 | n8389);
assign n22495 = n83 | n13663;
assign n17635 = n18024;
assign n1692 = n5263 | n9160;
assign n18083 = n19310 | n7499;
assign n931 = n920 | n11618;
assign n11062 = ~n8823;
assign n23910 = ~(n24296 ^ n6174);
assign n16455 = ~(n7727 ^ n24363);
assign n24560 = ~n12086;
assign n12348 = ~(n5587 | n111);
assign n13915 = ~(n5947 ^ n14440);
assign n12277 = n21856 & n24163;
assign n7152 = n25212 & n127;
assign n261 = n8538 | n20971;
assign n21763 = n25094 | n24586;
assign n23218 = ~n1183;
assign n4820 = n3320 & n17579;
assign n9378 = ~(n5573 ^ n2201);
assign n23397 = n9872 | n26726;
assign n1788 = n6309 | n14999;
assign n5447 = n12446 | n966;
assign n1898 = ~n26556;
assign n20165 = ~(n25886 | n8399);
assign n22062 = ~(n10372 | n12152);
assign n20569 = n6086 | n3197;
assign n6160 = ~(n4786 ^ n25222);
assign n9533 = n16825 | n17703;
assign n12370 = n2299 | n5792;
assign n11073 = n6878 & n22280;
assign n21262 = ~(n21460 ^ n18079);
assign n18776 = ~(n15000 | n16106);
assign n18032 = ~n3299;
assign n12810 = ~n20906;
assign n16917 = n4897 & n26819;
assign n4096 = n15702 & n26500;
assign n19349 = n22522 & n17876;
assign n14712 = n26615 | n4025;
assign n10169 = ~(n23137 ^ n11617);
assign n17298 = ~(n25276 ^ n12341);
assign n18840 = ~(n21537 ^ n18031);
assign n19866 = ~(n13190 ^ n9318);
assign n13171 = ~(n16007 ^ n12821);
assign n11208 = n20329 | n6397;
assign n9332 = ~n9886;
assign n11148 = ~(n7437 ^ n1662);
assign n8983 = ~(n6877 | n874);
assign n10984 = ~(n21274 ^ n19191);
assign n22137 = n3660 & n8040;
assign n2754 = n21261 | n18204;
assign n13861 = n15796 | n12446;
assign n19722 = ~n5176;
assign n2552 = ~(n5313 ^ n14274);
assign n4467 = ~(n14134 ^ n20253);
assign n17674 = ~n8820;
assign n2606 = ~n4939;
assign n11454 = n13517 | n9522;
assign n15977 = n25926 & n9646;
assign n17476 = ~(n5938 ^ n7212);
assign n11913 = ~(n23244 | n5128);
assign n12214 = ~(n9345 ^ n19941);
assign n24627 = ~(n22755 | n7503);
assign n10219 = ~(n21211 ^ n917);
assign n1410 = ~(n20249 ^ n17902);
assign n26751 = n7353 | n19730;
assign n8669 = ~(n26660 ^ n18907);
assign n21386 = ~n12657;
assign n3386 = n25872 | n19618;
assign n17586 = ~n16543;
assign n10527 = ~n7276;
assign n20917 = ~(n12679 ^ n11039);
assign n22901 = n8960 | n12187;
assign n24801 = ~(n22757 ^ n24870);
assign n19769 = n8049 & n7446;
assign n8079 = ~(n19860 ^ n2785);
assign n16186 = ~(n26417 | n10509);
assign n16561 = ~n18227;
assign n2638 = n16161 & n2093;
assign n23813 = n2196 | n1059;
assign n23465 = n2669 | n347;
assign n19710 = n2187 | n5832;
assign n6592 = ~(n13590 | n1792);
assign n8706 = ~(n13960 ^ n9493);
assign n16927 = n1036 | n10967;
assign n9889 = ~(n10666 ^ n9489);
assign n3272 = n7017 | n1889;
assign n13509 = n3310 & n18627;
assign n26870 = ~(n26278 ^ n5042);
assign n18487 = ~(n23824 ^ n9730);
assign n16933 = n20984 & n250;
assign n8191 = ~(n23034 | n24684);
assign n21579 = ~(n14187 ^ n7162);
assign n3471 = ~(n17683 ^ n5552);
assign n20522 = n10565 | n23806;
assign n1126 = n6310 & n20672;
assign n17775 = n19344 & n14497;
assign n14501 = ~(n21162 ^ n10018);
assign n22520 = n26210 & n20380;
assign n8640 = n9600 | n7578;
assign n11986 = ~(n19693 ^ n20197);
assign n2623 = ~(n1662 ^ n3710);
assign n8996 = n22764 & n26830;
assign n5544 = n7238 | n14923;
assign n3845 = ~(n5342 ^ n17559);
assign n7481 = ~n7028;
assign n26196 = ~(n18183 ^ n23071);
assign n5624 = ~n12446;
assign n17334 = ~(n20077 | n3952);
assign n3860 = n25909 & n9153;
assign n12563 = ~n21725;
assign n8245 = n24983 & n19278;
assign n1877 = n4315 | n23200;
assign n16964 = n12038 | n22070;
assign n22684 = ~(n11822 ^ n12811);
assign n11829 = ~(n20455 | n2884);
assign n14868 = ~(n10097 ^ n9564);
assign n19648 = ~(n26275 ^ n26937);
assign n11390 = ~(n10902 ^ n9952);
assign n25021 = ~n19701;
assign n9541 = n22762 | n24846;
assign n19500 = ~(n5211 ^ n12811);
assign n2209 = ~(n23817 ^ n15299);
assign n20621 = ~(n15733 ^ n18692);
assign n24128 = ~(n5976 ^ n2694);
assign n14933 = ~(n23755 | n23509);
assign n23929 = n8566 | n24619;
assign n8956 = n26839 & n9667;
assign n19542 = ~(n3780 ^ n17276);
assign n18231 = ~(n13696 ^ n25514);
assign n5598 = n882 & n26097;
assign n6925 = ~(n13030 ^ n71);
assign n791 = ~(n19122 ^ n23632);
assign n21181 = ~(n10893 | n9817);
assign n3846 = ~(n4196 ^ n11415);
assign n6053 = n4871 | n815;
assign n18972 = ~(n23931 ^ n19020);
assign n10358 = n6773 & n20089;
assign n18018 = ~(n11630 | n3783);
assign n880 = ~n1513;
assign n23128 = n12541 & n3412;
assign n22929 = n20883 | n5859;
assign n18634 = ~(n23340 ^ n7570);
assign n17926 = ~n9218;
assign n16253 = n23981 | n17709;
assign n17232 = ~(n12026 ^ n10672);
assign n15295 = ~(n10405 | n8241);
assign n8307 = n17087 | n16092;
assign n17777 = n6325 | n27161;
assign n24225 = n14227 & n15968;
assign n17087 = ~n3694;
assign n7574 = n7724 & n3322;
assign n24760 = ~(n216 | n20059);
assign n7367 = n25139 | n7974;
assign n2410 = n18017 | n15582;
assign n11064 = n15766 & n7465;
assign n23727 = ~(n21393 ^ n3935);
assign n3532 = n5444 & n18748;
assign n17507 = ~(n25846 | n7546);
assign n13691 = ~(n10611 ^ n2680);
assign n26007 = ~(n21338 ^ n27010);
assign n11205 = n7099 & n18888;
assign n21717 = ~(n3609 ^ n24148);
assign n8859 = ~n17294;
assign n3810 = ~(n2161 ^ n5924);
assign n10279 = ~(n2410 ^ n6230);
assign n4520 = ~(n26535 ^ n4198);
assign n11910 = ~(n21033 ^ n9441);
assign n5151 = n16529 | n20005;
assign n1414 = ~(n474 ^ n12104);
assign n16985 = n3981 | n1741;
assign n12185 = n19056 & n22854;
assign n22744 = ~(n23155 ^ n14456);
assign n25849 = n20652 | n2890;
assign n942 = ~(n15258 | n2420);
assign n23476 = n22123 | n18078;
assign n26437 = ~n264;
assign n13538 = n7693 | n15644;
assign n9731 = n23629 | n25648;
assign n2212 = ~(n23234 | n20138);
assign n15659 = n3002;
assign n788 = ~n14816;
assign n24464 = ~(n26857 ^ n1881);
assign n18675 = n6915 | n15996;
assign n26612 = n212 | n2146;
assign n25264 = ~(n17716 ^ n25475);
assign n12796 = n25440 | n20644;
assign n20113 = ~(n15271 | n26748);
assign n14722 = n24638 & n19327;
assign n23893 = n15086 | n13927;
assign n15095 = n523 & n9912;
assign n9206 = ~(n20551 ^ n8283);
assign n17538 = ~(n21527 ^ n26174);
assign n18366 = n20544 | n22652;
assign n24088 = n1767 & n3250;
assign n18765 = ~(n22769 ^ n21839);
assign n21882 = n9657 & n19275;
assign n4341 = n19110 & n26753;
assign n8733 = n7225 & n26352;
assign n12517 = n2131 | n11809;
assign n4091 = n27092 | n2052;
assign n5203 = ~n7377;
assign n7473 = n14790 | n26075;
assign n2078 = ~(n24165 ^ n15842);
assign n16715 = n12309 & n4013;
assign n26160 = ~(n14487 ^ n53);
assign n7110 = n25544 & n18184;
assign n11003 = n18842 & n26487;
assign n4021 = n3025 | n9137;
assign n10928 = ~(n9570 | n1667);
assign n14385 = ~n9748;
assign n14785 = ~(n23863 | n14702);
assign n16658 = n10405 & n12198;
assign n26266 = n21652 & n5225;
assign n321 = ~(n16846 | n24101);
assign n22794 = ~(n9416 | n17587);
assign n3524 = ~(n12316 ^ n20340);
assign n18823 = n4085 & n16547;
assign n23306 = n9493 & n15507;
assign n10754 = ~(n11534 | n8659);
assign n9110 = ~(n25935 ^ n15817);
assign n26515 = ~(n26973 ^ n24533);
assign n1498 = ~(n7078 ^ n17012);
assign n23173 = ~(n18880 | n26594);
assign n10814 = n13326 | n2293;
assign n5922 = n16029 & n4322;
assign n23294 = n21558 & n18783;
assign n16213 = ~n18429;
assign n24203 = ~(n2576 ^ n15532);
assign n21236 = n6446 & n20060;
assign n21479 = ~(n347 ^ n4346);
assign n21663 = ~(n8399 | n6834);
assign n9856 = ~n24392;
assign n3377 = ~(n26667 ^ n16183);
assign n4677 = n12535 & n4705;
assign n7031 = ~(n4326 ^ n14148);
assign n10378 = ~n1090;
assign n6007 = n9018 | n18047;
assign n4927 = ~(n5330 ^ n919);
assign n19314 = ~(n6719 ^ n11967);
assign n18995 = ~n7566;
assign n1351 = ~(n10160 ^ n8229);
assign n3289 = ~(n14844 ^ n16862);
assign n6770 = n27202 | n15085;
assign n4393 = ~(n27095 ^ n2160);
assign n17243 = ~(n9408 ^ n11431);
assign n22385 = ~(n22012 ^ n13387);
assign n17992 = n19875 & n9737;
assign n13214 = ~n9170;
assign n16461 = n26370 | n10782;
assign n24067 = n15780 & n24358;
assign n16487 = n8880 & n5975;
assign n14870 = ~n12470;
assign n18549 = ~(n18799 ^ n10763);
assign n25992 = n15186 | n26928;
assign n25780 = n15712 | n12571;
assign n17115 = ~(n21185 ^ n27165);
assign n15371 = ~(n17790 | n9651);
assign n25467 = ~(n20411 ^ n9512);
assign n13814 = ~(n24116 | n23408);
assign n14520 = n20137 | n1662;
assign n22336 = n17162 & n868;
assign n23359 = ~n2979;
assign n13289 = n10323 | n25785;
assign n14174 = ~(n16425 ^ n19356);
assign n22667 = ~(n13249 ^ n25156);
assign n2448 = n12590 & n16270;
assign n26090 = ~n25608;
assign n22903 = ~(n20439 ^ n17114);
assign n8716 = ~(n4830 ^ n19740);
assign n10811 = n9791 | n13462;
assign n19479 = n25535 & n16546;
assign n26354 = n10534 | n24896;
assign n17808 = ~(n22748 ^ n24128);
assign n3121 = ~(n18888 ^ n7099);
assign n7224 = ~(n10124 | n8897);
assign n5876 = ~(n2036 ^ n23630);
assign n1240 = ~(n27120 ^ n11192);
assign n16215 = ~(n19637 ^ n11297);
assign n19445 = ~(n5682 | n10468);
assign n6920 = n22454 | n10710;
assign n1142 = n10191 | n15792;
assign n26574 = n14040 & n24711;
assign n10849 = ~n18551;
assign n19939 = n20032 | n19144;
assign n19060 = ~(n21387 ^ n12487);
assign n12141 = ~(n18438 ^ n26672);
assign n1395 = n22843 | n4155;
assign n19752 = ~(n835 ^ n13668);
assign n18090 = ~n18649;
assign n27154 = ~(n14365 ^ n2804);
assign n13211 = n26153 | n11372;
assign n20537 = ~n4597;
assign n7787 = ~(n21453 ^ n4273);
assign n810 = n3107 & n26941;
assign n10097 = ~n19589;
assign n20656 = n12007 & n23377;
assign n16113 = n4498 & n19766;
assign n5010 = n14012 & n7774;
assign n15196 = ~(n22240 | n2375);
assign n25140 = ~(n910 ^ n12891);
assign n14698 = ~(n1307 | n25219);
assign n6216 = ~(n19886 ^ n14091);
assign n2312 = ~n12687;
assign n23622 = n17137 | n11689;
assign n22009 = ~n24458;
assign n21635 = n14538 & n23862;
assign n15667 = ~(n10751 | n27009);
assign n17642 = ~(n21915 | n24919);
assign n1488 = n22559 | n19995;
assign n6284 = ~n2320;
assign n8655 = n16594 | n17351;
assign n13598 = n15026 | n5063;
assign n10834 = ~(n10187 ^ n26331);
assign n24517 = ~(n22840 ^ n11765);
assign n11491 = n13380 & n2067;
assign n19353 = n6543 | n1720;
assign n1348 = ~(n5220 ^ n6948);
assign n9005 = ~(n4572 ^ n23581);
assign n22015 = ~n21784;
assign n12128 = ~n25623;
assign n16529 = ~n16536;
assign n6644 = n7463 & n16821;
assign n4143 = ~n17415;
assign n10072 = n11805 | n20426;
assign n13298 = n16401 & n7861;
assign n5194 = ~n3072;
assign n21230 = ~n14058;
assign n21057 = ~(n25692 | n729);
assign n2326 = ~(n25052 ^ n25895);
assign n10071 = ~(n10267 | n12592);
assign n13697 = n8963 | n24041;
assign n4171 = n13337 | n7200;
assign n16566 = n23419 | n22951;
assign n11359 = n20410 | n7365;
assign n10143 = n937 & n15733;
assign n21897 = ~(n23920 ^ n5231);
assign n4902 = ~(n16524 | n20923);
assign n21707 = ~(n586 ^ n15274);
assign n15154 = n19019 & n16408;
assign n15472 = n3682 | n5339;
assign n2511 = ~(n19589 | n9564);
assign n21975 = ~n3955;
assign n10610 = ~n18599;
assign n21667 = n4087 | n808;
assign n17524 = ~(n3167 ^ n6001);
assign n6240 = ~n13090;
assign n5210 = n24598 & n14006;
assign n15870 = n3877 | n23034;
assign n19677 = n1573 | n4652;
assign n6732 = n22499 & n3331;
assign n2713 = ~n21471;
assign n17696 = ~(n18409 ^ n3952);
assign n23732 = n18027 | n4866;
assign n9974 = ~n5910;
assign n9573 = n17741 | n10451;
assign n20340 = ~(n16345 ^ n4542);
assign n23977 = n24891 & n7878;
assign n14811 = ~(n15442 ^ n6015);
assign n15935 = ~n5587;
assign n19511 = ~(n19646 | n8277);
assign n20771 = ~n8085;
assign n24533 = ~(n15236 ^ n2383);
assign n12815 = ~n3976;
assign n20031 = n22056 & n20817;
assign n13114 = ~n17037;
assign n25655 = ~(n26986 ^ n2272);
assign n9742 = ~(n13783 ^ n9942);
assign n10206 = n20365 | n14127;
assign n26469 = ~(n13898 | n25004);
assign n18268 = n5360 & n21340;
assign n19016 = n22976 & n21958;
assign n22059 = n9793 & n22361;
assign n12647 = n2933 & n372;
assign n25284 = n13044 | n4038;
assign n20394 = n5489 & n16342;
assign n7353 = ~n6307;
assign n26009 = n20346 & n9315;
assign n6406 = n543 & n2244;
assign n12258 = ~n23200;
assign n4046 = n22271 | n19417;
assign n13620 = n21265 & n23266;
assign n19991 = n14718 | n6814;
assign n13592 = n14955 & n13098;
assign n17731 = ~(n12875 ^ n7751);
assign n22055 = ~(n1685 | n9514);
assign n5383 = ~(n11056 ^ n20478);
assign n20321 = n22962 & n10567;
assign n24652 = n13967 | n18972;
assign n19369 = n1215 | n23715;
assign n14064 = ~(n5506 ^ n2331);
assign n5180 = ~n22698;
assign n7104 = n23836 & n7562;
assign n19365 = ~(n390 ^ n5060);
assign n22653 = n7763 & n1627;
assign n16797 = ~(n20437 ^ n26565);
assign n21283 = n9880 & n20273;
assign n11741 = ~(n24243 ^ n26044);
assign n588 = n16089 & n9316;
assign n27093 = ~(n144 | n5960);
assign n20774 = ~(n11588 ^ n21098);
assign n4133 = ~(n4194 | n8795);
assign n16886 = ~(n14287 ^ n585);
assign n13559 = n13117 & n20084;
assign n25697 = ~n2989;
assign n1619 = n22687 & n11734;
assign n16895 = ~(n22197 ^ n5927);
assign n21862 = n9644 & n17894;
assign n5688 = ~(n22379 | n22207);
assign n14950 = ~(n12137 | n10258);
assign n23871 = ~(n25100 ^ n23765);
assign n19845 = ~(n23604 ^ n15328);
assign n203 = ~(n21759 | n5445);
assign n26397 = n22331 & n9203;
assign n24857 = ~(n6002 ^ n20107);
assign n26739 = n25558 | n13668;
assign n24354 = n15995 | n516;
assign n6080 = n19799 & n15112;
assign n19877 = ~(n2783 ^ n6785);
assign n4941 = ~n20707;
assign n15916 = n7952 | n1136;
assign n3640 = n1300 | n14567;
assign n18777 = n13171 | n13633;
assign n3507 = n10147 | n15169;
assign n20306 = n16086 | n7105;
assign n1687 = ~n679;
assign n24123 = n25112 | n18084;
assign n19703 = ~(n1202 | n4246);
assign n11760 = n23920 | n23344;
assign n23604 = n20676 | n19400;
assign n20493 = n10693 & n19167;
assign n23575 = ~(n20409 ^ n1099);
assign n7270 = ~(n19123 ^ n18208);
assign n8626 = ~(n19508 ^ n21234);
assign n11591 = ~(n2654 ^ n10979);
assign n2718 = ~n1413;
assign n18698 = ~(n16793 ^ n18428);
assign n21759 = ~(n806 ^ n4051);
assign n14597 = ~(n23655 ^ n23755);
assign n9293 = ~(n4467 ^ n9752);
assign n14534 = ~(n2966 ^ n19627);
assign n11888 = ~(n18861 ^ n22091);
assign n14319 = ~(n7105 ^ n3543);
assign n6776 = n21089 & n13224;
assign n26385 = n16316 & n9279;
assign n24754 = ~(n25733 | n19498);
assign n9346 = ~(n7824 ^ n22808);
assign n17652 = ~(n2447 ^ n9089);
assign n21249 = ~n14999;
assign n19276 = ~(n16627 ^ n6765);
assign n13194 = ~(n3239 ^ n6648);
assign n14650 = n21138 | n14230;
assign n2132 = ~(n2939 ^ n6366);
assign n217 = n5719 | n14130;
assign n2628 = ~n25381;
assign n2244 = ~(n1496 ^ n7502);
assign n7314 = ~(n18785 ^ n14096);
assign n3525 = ~(n2858 | n5521);
assign n16745 = n8381 | n20382;
assign n25220 = ~n24988;
assign n25585 = ~(n3675 ^ n5145);
assign n2658 = n10522 & n23024;
assign n26463 = ~(n163 ^ n13015);
assign n22870 = ~(n26761 ^ n22080);
assign n10001 = ~(n22774 ^ n1611);
assign n21585 = ~(n11558 ^ n2280);
assign n11861 = n1923 | n9200;
assign n25952 = ~(n25015 ^ n15131);
assign n512 = n10565 & n23806;
assign n24275 = n3482 & n25374;
assign n23799 = ~(n11858 ^ n17885);
assign n19767 = ~(n16878 ^ n19835);
assign n24966 = ~(n18976 | n15090);
assign n19965 = n23867 | n12296;
assign n19132 = ~(n6165 ^ n12201);
assign n6782 = n1437 & n17784;
assign n17743 = ~(n115 ^ n2355);
assign n25306 = n19355 | n8153;
assign n6755 = n5233 | n7214;
assign n894 = ~(n1742 ^ n4590);
assign n11997 = ~(n5196 ^ n4491);
assign n19233 = ~(n20024 ^ n6088);
assign n18799 = ~(n7869 ^ n14968);
assign n2412 = ~n8041;
assign n25683 = n13644 & n3712;
assign n18263 = ~(n1148 ^ n17810);
assign n9550 = ~(n19952 ^ n10178);
assign n424 = ~n22047;
assign n11333 = n6394 & n9273;
assign n21517 = ~(n5959 ^ n9835);
assign n20463 = n2281 | n1047;
assign n19089 = ~(n12495 ^ n15780);
assign n15213 = ~(n8989 | n12162);
assign n3376 = ~n9455;
assign n25103 = ~n10229;
assign n6168 = ~(n16403 ^ n13008);
assign n2651 = ~(n9283 ^ n6633);
assign n15060 = n7593 | n25317;
assign n26623 = n5013 | n5305;
assign n11488 = ~(n15294 ^ n5538);
assign n11178 = ~n17485;
assign n2955 = n3161 | n18201;
assign n6835 = ~(n11931 ^ n17229);
assign n15466 = n4692 | n15775;
assign n13954 = n120 | n4939;
assign n25976 = n8891 | n7406;
assign n7212 = ~(n13554 ^ n7004);
assign n22826 = n6081 & n15434;
assign n8659 = n17776 & n8512;
assign n3237 = n793 | n12736;
assign n25319 = n11030 | n6141;
assign n10757 = ~(n8363 | n1222);
assign n5644 = n12365 & n20306;
assign n12767 = ~(n13378 ^ n10444);
assign n5775 = n1705 | n9456;
assign n7912 = n7391 | n24134;
assign n3312 = ~(n12522 | n8308);
assign n7610 = ~(n14929 ^ n2132);
assign n14439 = n1404 | n14684;
assign n5425 = n20893 & n18128;
assign n5127 = n24620 | n21753;
assign n20186 = n12398 | n25696;
assign n8753 = ~(n21138 ^ n20385);
assign n10753 = n5313 & n17156;
assign n94 = ~(n24808 ^ n13860);
assign n24483 = ~(n24034 ^ n26885);
assign n17484 = ~(n26471 | n22382);
assign n25717 = n21566 | n14343;
assign n717 = n8368 | n7504;
assign n7547 = ~(n6861 ^ n5255);
assign n23903 = ~(n17700 ^ n1728);
assign n6020 = ~(n8853 ^ n23036);
assign n5177 = n20120 | n9313;
assign n6272 = n7639 | n11703;
assign n3883 = n22288 | n24023;
assign n14263 = n14051 | n290;
assign n846 = ~(n13494 | n3425);
assign n14952 = ~(n22634 ^ n17816);
assign n6175 = ~(n10888 ^ n14176);
assign n6393 = ~n22619;
assign n23674 = n9773 & n26163;
assign n13629 = ~(n3659 | n17635);
assign n26504 = ~(n11694 ^ n18040);
assign n5126 = ~(n7935 ^ n18608);
assign n3870 = ~(n2462 ^ n21150);
assign n23836 = n16439 | n10275;
assign n772 = ~(n2498 ^ n14185);
assign n4741 = n10191 & n15792;
assign n20042 = ~(n5938 | n960);
assign n2154 = n25047 & n1381;
assign n22488 = ~(n27037 ^ n13775);
assign n2510 = ~(n21326 ^ n12623);
assign n9252 = n25855 ^ n24714;
assign n8962 = ~(n11146 ^ n17095);
assign n9473 = n21091 & n13415;
assign n25087 = ~(n14790 ^ n342);
assign n9714 = ~(n17590 ^ n17549);
assign n4757 = n13300 | n17000;
assign n13352 = ~(n652 ^ n16181);
assign n17973 = ~(n24187 | n19331);
assign n6563 = n8966 | n12128;
assign n4436 = ~(n769 ^ n16280);
assign n13068 = n23932 | n9380;
assign n19798 = ~(n10630 ^ n18876);
assign n12791 = n1838 | n14127;
assign n16134 = n5292 | n25144;
assign n1035 = n20853 | n10238;
assign n9155 = n19138 | n13066;
assign n5119 = ~n26641;
assign n21895 = n18345 | n22700;
assign n11366 = ~n8233;
assign n23019 = n16157 & n16343;
assign n22869 = n22775 | n20895;
assign n7447 = ~n19045;
assign n11956 = n18430 | n10764;
assign n11916 = n9654 | n23057;
assign n5261 = ~n8718;
assign n12520 = n22003 | n23705;
assign n16883 = n20319 & n25046;
assign n20351 = ~(n20049 ^ n12610);
assign n23573 = ~n7260;
assign n22506 = n7523 & n23686;
assign n24646 = ~(n8486 ^ n22592);
assign n1231 = ~(n4602 ^ n21337);
assign n25332 = ~(n23152 ^ n1909);
assign n16808 = ~(n19757 ^ n8126);
assign n19425 = ~(n6360 ^ n15970);
assign n1595 = n11186 | n23878;
assign n8747 = n15932 | n8728;
assign n18864 = ~(n25845 ^ n18497);
assign n14306 = ~n9851;
assign n12700 = n3790 ^ n11192;
assign n5051 = n1251 & n23595;
assign n19084 = ~n22154;
assign n6413 = n10966 & n3420;
assign n24218 = n24411 & n6957;
assign n1043 = n10414 | n23193;
assign n24165 = ~(n11948 ^ n652);
assign n24172 = ~(n2033 | n13706);
assign n14450 = n472 | n26752;
assign n3220 = ~(n5873 ^ n19001);
assign n6288 = ~(n21593 | n20972);
assign n23699 = n9048 | n14951;
assign n11546 = n18292 & n2029;
assign n2318 = ~(n18004 | n350);
assign n2834 = n8640 & n13065;
assign n10541 = ~n17048;
assign n9168 = n18523 & n9774;
assign n19352 = ~(n15258 ^ n4588);
assign n7341 = ~n22215;
assign n19657 = n14507 | n23208;
assign n3970 = ~(n9222 | n19143);
assign n8565 = n12924 | n23597;
assign n2740 = n9832 | n21240;
assign n20843 = n24783 | n5199;
assign n4833 = ~(n8856 | n8305);
assign n10063 = n2517 & n9194;
assign n14346 = ~n18234;
assign n16127 = ~(n8363 | n2816);
assign n19972 = n23362 | n13196;
assign n25029 = n16473 & n2111;
assign n4691 = n2371 & n19255;
assign n249 = ~(n10341 | n9855);
assign n25398 = ~(n7546 ^ n6831);
assign n21058 = n17609 & n12568;
assign n15714 = n7090 | n16855;
assign n9402 = ~n24692;
assign n19913 = ~(n23591 ^ n19465);
assign n16340 = ~(n252 ^ n20316);
assign n24086 = ~(n2146 ^ n19144);
assign n25690 = ~(n19469 | n27188);
assign n23548 = n1644 & n21612;
assign n25310 = ~(n7973 ^ n15179);
assign n13145 = n23522 & n7500;
assign n13695 = ~(n13376 ^ n4643);
assign n14783 = ~n13472;
assign n1816 = ~(n17568 | n26986);
assign n650 = ~(n23256 ^ n23287);
assign n10836 = ~(n9793 ^ n22361);
assign n22460 = ~(n24031 | n21915);
assign n19269 = n6350 & n27023;
assign n12814 = ~(n17993 ^ n23145);
assign n8152 = n21739 & n24805;
assign n11669 = n26208;
assign n26853 = ~(n9242 ^ n17541);
assign n24632 = ~(n8331 ^ n5743);
assign n26726 = ~(n7815 ^ n18210);
assign n2064 = n10211 | n19565;
assign n18410 = n16755 | n2816;
assign n5736 = n8948 & n3470;
assign n14648 = ~(n2984 ^ n25867);
assign n17581 = ~n14487;
assign n20465 = n2796 & n18984;
assign n13806 = n19373 & n23381;
assign n19106 = ~n10611;
assign n18394 = ~(n15959 | n10075);
assign n6540 = n15431 & n21105;
assign n23169 = n23487 | n12956;
assign n25834 = n4671 & n7128;
assign n17913 = ~(n13152 ^ n2688);
assign n10278 = ~(n151 ^ n21405);
assign n13653 = ~(n6351 | n354);
assign n11402 = ~(n23160 | n8067);
assign n15274 = ~n24473;
assign n15684 = ~(n6658 | n6255);
assign n18782 = ~(n1382 ^ n2356);
assign n11962 = n19697 & n11890;
assign n11427 = n7189 | n11255;
assign n3742 = ~n21952;
assign n23188 = ~(n11207 ^ n20986);
assign n26757 = n7026 | n17835;
assign n986 = n16045 | n7321;
assign n14600 = ~(n194 ^ n24696);
assign n1799 = ~n21001;
assign n10675 = n21917 & n16986;
assign n12483 = ~(n14573 ^ n25381);
assign n5094 = ~n474;
assign n17528 = ~(n2263 | n13857);
assign n4247 = ~(n3740 ^ n21784);
assign n9455 = ~(n10868 ^ n22554);
assign n2077 = ~n14954;
assign n9283 = n14203 | n26554;
assign n24325 = ~n16376;
assign n11259 = ~n26893;
assign n23520 = n14525 | n6818;
assign n6182 = ~n23357;
assign n11978 = ~(n2657 | n13073);
assign n16773 = n16443 | n23829;
assign n8192 = ~(n4040 | n13775);
assign n12552 = ~(n4329 ^ n8019);
assign n691 = ~(n17936 ^ n11971);
assign n5130 = n1681 & n9196;
assign n10388 = ~(n9271 ^ n21893);
assign n14699 = ~n1844;
assign n11370 = n19094 & n19156;
assign n11446 = n17479 | n26054;
assign n21007 = ~n9185;
assign n7484 = ~(n16037 ^ n18291);
assign n19211 = ~(n22557 | n7447);
assign n22649 = n19716 | n10269;
assign n3206 = ~(n13480 | n22270);
assign n12679 = ~(n10415 ^ n11299);
assign n3672 = ~n933;
assign n19986 = ~(n25043 | n25612);
assign n10646 = n17230 | n658;
assign n6853 = ~(n7248 ^ n12099);
assign n14054 = n22990 | n769;
assign n1284 = n5328 | n20273;
assign n20548 = n24366 & n14395;
assign n26556 = ~(n6764 ^ n1451);
assign n17465 = n1930 & n5681;
assign n10421 = ~(n18412 | n1837);
assign n17187 = ~(n2935 | n3203);
assign n2010 = ~(n7761 ^ n22222);
assign n10548 = ~(n446 | n3324);
assign n11093 = n12066 | n7788;
assign n6161 = ~(n11198 | n4384);
assign n3662 = ~(n13562 ^ n15127);
assign n16220 = n11389 & n9369;
assign n6068 = n25607;
assign n5097 = n4061 | n18473;
assign n2202 = ~(n19926 | n1243);
assign n25349 = n20272 & n20439;
assign n19485 = ~(n1066 ^ n21565);
assign n25280 = n4650 | n19008;
assign n25409 = ~(n2436 | n15502);
assign n16250 = n16931 | n26397;
assign n12558 = ~(n20179 ^ n3460);
assign n5002 = n23387 & n701;
assign n2514 = ~n12811;
assign n18630 = ~(n22919 ^ n3618);
assign n15298 = ~(n15897 | n24217);
assign n18376 = n7035 | n8529;
assign n25641 = ~(n7400 ^ n2124);
assign n4321 = ~(n17088 | n17832);
assign n3746 = ~(n2162 ^ n3486);
assign n18986 = ~(n18473 | n19514);
assign n11904 = n13088 | n12720;
assign n16163 = ~n3075;
assign n4845 = n8068 & n4466;
assign n8148 = ~(n16112 ^ n1034);
assign n14729 = n2563 | n19381;
assign n18373 = ~(n20289 ^ n12293);
assign n10874 = ~(n6973 ^ n21049);
assign n14318 = ~n219;
assign n11685 = ~n25126;
assign n10946 = ~(n10514 | n4514);
assign n14232 = n7883 | n8402;
assign n4578 = n16971 | n15600;
assign n2821 = ~(n21492 | n7776);
assign n22924 = ~(n8002 | n19539);
assign n19177 = ~(n1174 ^ n1109);
assign n19934 = n17013 | n18674;
assign n514 = n5802 | n19368;
assign n14656 = ~(n22342 ^ n13719);
assign n21801 = n10406 | n8947;
assign n5802 = ~(n10419 ^ n765);
assign n5913 = n16244 | n16264;
assign n19309 = ~(n893 ^ n13439);
assign n8110 = n8648 | n13287;
assign n5540 = n24325 | n6381;
assign n16038 = ~(n7851 ^ n10045);
assign n15140 = ~(n4294 ^ n11381);
assign n9896 = n15003 & n8995;
assign n18220 = ~n9259;
assign n13010 = ~(n20826 ^ n626);
assign n19473 = n24358 | n1898;
assign n21439 = n1154 | n20854;
assign n21553 = n10719 | n19958;
assign n9505 = ~n9266;
assign n8356 = n17682 & n3546;
assign n17778 = n15062 | n15985;
assign n22142 = n20974 & n2932;
assign n19643 = n17304 & n19212;
assign n24231 = ~(n16084 | n21691);
assign n1945 = ~(n10201 ^ n22379);
assign n19641 = ~(n10187 ^ n17165);
assign n11475 = n13283 | n24296;
assign n26710 = n27020 | n1567;
assign n9536 = n26857 | n13739;
assign n24695 = ~n25023;
assign n10191 = ~n3832;
assign n16226 = ~(n14996 ^ n9226);
assign n13325 = n7769 | n21436;
assign n9475 = n22333 | n5072;
assign n10299 = n16269 & n6314;
assign n15924 = n15944 & n16432;
assign n22494 = ~(n13741 ^ n15728);
assign n3539 = n7027 | n24436;
assign n7521 = n1720 & n6543;
assign n24481 = ~(n11332 ^ n25423);
assign n12235 = ~(n17869 ^ n4183);
assign n6106 = n13400 | n18283;
assign n16677 = n15778 & n18588;
assign n7834 = ~(n5870 ^ n6752);
assign n19099 = n17475 | n23262;
assign n21319 = ~(n8888 ^ n12871);
assign n3369 = ~(n1753 ^ n21733);
assign n25324 = ~n4326;
assign n9576 = ~n4762;
assign n25997 = n19806 | n5737;
assign n285 = n9016 & n26842;
assign n5643 = ~(n18568 ^ n674);
assign n3631 = n26194 & n12299;
assign n23053 = ~(n3433 ^ n13993);
assign n896 = ~(n17780 | n19377);
assign n11277 = ~(n2371 ^ n14713);
assign n13749 = n27199 | n19843;
assign n21682 = ~(n24868 ^ n23268);
assign n5366 = ~n27169;
assign n23648 = n6353 & n8434;
assign n3069 = ~n8006;
assign n11524 = n14220 & n24678;
assign n11895 = n420 & n18219;
assign n2163 = ~n26425;
assign n24077 = ~(n1642 | n18409);
assign n13275 = n13353 | n18035;
assign n23047 = ~(n3688 ^ n11206);
assign n4265 = n13960 & n19785;
assign n22702 = ~n20238;
assign n18451 = n20314 & n13348;
assign n19696 = ~(n8695 ^ n8492);
assign n21994 = ~(n23321 | n6300);
assign n18985 = n6036 & n20892;
assign n9803 = ~(n21838 ^ n25489);
assign n16308 = ~(n12249 | n13875);
assign n19850 = ~(n144 | n25119);
assign n2643 = n16912 & n7315;
assign n11149 = ~(n10027 ^ n5822);
assign n7614 = n21343 & n9710;
assign n9019 = n15187 & n5995;
assign n21384 = ~(n16524 ^ n20923);
assign n20990 = n26822 | n5475;
assign n21480 = n4030 & n13636;
assign n15952 = ~(n20517 | n26239);
assign n21022 = ~(n2704 | n7732);
assign n14823 = ~(n13291 | n2443);
assign n6333 = n22660 | n1596;
assign n17886 = n26296 | n25372;
assign n2023 = ~(n6000 ^ n24464);
assign n15511 = ~(n22556 ^ n7069);
assign n20496 = ~(n7693 | n22820);
assign n19598 = n22558 | n6814;
assign n12107 = n22118 | n7058;
assign n21998 = ~(n17830 ^ n10739);
assign n15874 = ~(n8052 ^ n23369);
assign n12846 = n7893 | n1654;
assign n18579 = n18896 | n3101;
assign n2406 = n12031 & n14752;
assign n3695 = n15507 | n19785;
assign n11800 = ~(n26947 ^ n12612);
assign n6858 = n18361 | n12439;
assign n9892 = n5356 | n5639;
assign n4322 = ~(n21928 ^ n11223);
assign n1041 = n1090 | n12687;
assign n3961 = n4041 & n3378;
assign n9530 = n17185 | n12747;
assign n20472 = ~(n23034 | n21352);
assign n9553 = n2567 & n4525;
assign n17207 = ~(n15242 ^ n11669);
assign n6688 = n25558 | n13748;
assign n5406 = ~(n6337 | n3686);
assign n535 = ~(n22114 ^ n268);
assign n2403 = ~(n21846 | n9493);
assign n8551 = n6528 | n16194;
assign n6652 = ~(n26254 ^ n8826);
assign n2143 = n315 & n25804;
assign n25139 = ~n11615;
assign n26971 = ~(n8272 | n17888);
assign n1924 = ~(n19418 ^ n3901);
assign n24693 = n3260 | n21832;
assign n18486 = ~(n9294 ^ n26022);
assign n10567 = n26661 | n8596;
assign n23783 = ~(n4302 ^ n3872);
assign n2050 = ~(n10097 ^ n8935);
assign n22066 = n9563 & n9903;
assign n1068 = n4188 & n12922;
assign n2017 = ~n9872;
assign n23776 = n17097 & n24909;
assign n21562 = n22442 & n25038;
assign n14713 = ~(n18093 ^ n25427);
assign n23444 = n3069 | n5211;
assign n12139 = n15076 | n13620;
assign n23743 = ~(n26028 ^ n17867);
assign n44 = n22115 & n22163;
assign n12146 = ~(n10299 ^ n24353);
assign n21237 = ~(n14749 ^ n856);
assign n23466 = ~n21782;
assign n12207 = ~n2226;
assign n10505 = n17653;
assign n17369 = ~n4909;
assign n10609 = n20758 & n5308;
assign n24697 = n15341 & n226;
assign n182 = ~n6445;
assign n15830 = ~(n27167 | n14804);
assign n17390 = ~n25113;
assign n23055 = ~(n19588 | n8322);
assign n3410 = ~(n17316 | n14750);
assign n3178 = ~n21898;
assign n594 = n1806 | n22185;
assign n18910 = n20712 & n12896;
assign n16224 = n22184 & n5962;
assign n17534 = n20929 | n23068;
assign n18215 = ~(n12657 ^ n21287);
assign n14002 = ~n22871;
assign n2810 = n7839 & n23363;
assign n1989 = n12871 | n8888;
assign n3720 = n6501 | n14941;
assign n12131 = ~(n2683 ^ n19071);
assign n430 = n4369 & n4336;
assign n1823 = ~(n16701 ^ n25144);
assign n26078 = ~n12860;
assign n16537 = n2117 & n6711;
assign n19528 = n20717 | n482;
assign n91 = ~(n25556 ^ n5328);
assign n20588 = ~(n10077 | n9285);
assign n26544 = ~n16724;
assign n15712 = ~(n4042 | n10833);
assign n17135 = n17839 & n2294;
assign n1854 = ~(n25953 ^ n12868);
assign n23437 = n7143 | n10728;
assign n4189 = ~(n23704 ^ n20359);
assign n25357 = n16742 | n12285;
assign n8974 = ~(n10157 ^ n22753);
assign n6373 = ~(n15988 ^ n5343);
assign n8014 = n8087 | n15643;
assign n22553 = n3046 | n19655;
assign n16457 = ~(n10096 ^ n26553);
assign n6077 = n3384 | n6244;
assign n10636 = n17122 | n26177;
assign n10631 = ~(n22037 ^ n20669);
assign n13599 = n9533 & n23794;
assign n8146 = ~(n25374 ^ n6532);
assign n2418 = ~(n12185 ^ n1301);
assign n24864 = ~(n399 | n13949);
assign n24362 = n18217 | n12718;
assign n22577 = ~(n7676 | n12512);
assign n18465 = n20532 & n7416;
assign n26756 = n11278 | n2815;
assign n14581 = n6156 | n19859;
assign n19197 = n776 | n21430;
assign n17733 = ~(n350 ^ n1882);
assign n24773 = n10119 | n2526;
assign n18140 = n9679 | n22626;
assign n16763 = n25760 | n18330;
assign n26667 = ~(n20855 ^ n5827);
assign n23170 = ~(n3888 ^ n2993);
assign n25143 = n4713 | n14067;
assign n19999 = n25772 | n22047;
assign n559 = n12160 | n10562;
assign n13840 = n12482 & n19441;
assign n16304 = ~(n17382 ^ n5207);
assign n277 = ~n10001;
assign n5728 = ~n23372;
assign n7016 = n11896 | n9384;
assign n6863 = ~(n4304 ^ n1563);
assign n13440 = n14437 | n16663;
assign n21694 = ~n1185;
assign n18825 = n24051 | n15996;
assign n1897 = n5641 | n1430;
assign n12850 = ~(n16325 ^ n9832);
assign n25472 = n543 | n2244;
assign n22004 = ~(n8933 ^ n6865);
assign n20320 = n7380 | n3226;
assign n15113 = ~n14156;
assign n11437 = n8436 & n16076;
assign n16622 = n16294 | n17568;
assign n6917 = ~n22993;
assign n7555 = ~(n8902 ^ n5902);
assign n17183 = ~(n6440 ^ n23420);
assign n9162 = ~(n10956 | n1598);
assign n1339 = ~(n12935 ^ n22162);
assign n738 = n7320 | n6381;
assign n2789 = n18280 | n5937;
assign n23265 = n26852 & n13213;
assign n2002 = ~(n1339 ^ n14633);
assign n14126 = ~(n10750 ^ n2086);
assign n4363 = n20667 | n12956;
assign n3230 = n19127 & n18200;
assign n23073 = ~(n8084 | n18755);
assign n27137 = n14422 | n16113;
assign n19951 = ~(n12745 ^ n22542);
assign n1063 = n20544 | n23586;
assign n1711 = n19606 | n14578;
assign n746 = n10470 & n4062;
assign n23059 = ~n8403;
assign n17991 = n10248 | n10358;
assign n14417 = n24611 | n6578;
assign n16091 = ~(n10765 ^ n2337);
assign n12301 = ~n17968;
assign n15938 = n23144 & n10306;
assign n591 = n12320 | n194;
assign n1868 = ~(n24327 | n4325);
assign n12665 = ~(n27069 ^ n4937);
assign n15379 = ~(n5226 ^ n11223);
assign n14556 = n12160 | n16994;
assign n20682 = n15425 & n19870;
assign n3270 = ~(n24620 ^ n21753);
assign n15573 = ~(n9862 ^ n19308);
assign n17549 = n7856;
assign n16907 = ~(n9390 ^ n11730);
assign n1991 = ~(n11163 ^ n19642);
assign n2188 = n9118 | n13661;
assign n26419 = ~(n16009 ^ n12910);
assign n3921 = ~n152;
assign n20914 = n16084 | n18537;
assign n22888 = ~(n23517 ^ n10369);
assign n22952 = n5622 & n12077;
assign n25687 = ~(n11454 ^ n19364);
assign n8136 = n15144 | n25359;
assign n17919 = n13109 | n24898;
assign n25438 = n3655 & n17924;
assign n7793 = ~(n26107 ^ n4376);
assign n22105 = ~(n12684 ^ n21683);
assign n15072 = n26925 & n9394;
assign n873 = ~(n22647 ^ n6402);
assign n6595 = ~n24949;
assign n12639 = ~n2272;
assign n10576 = n4338 & n24430;
assign n5184 = ~(n4754 ^ n13648);
assign n4111 = n16999 & n7370;
assign n13684 = ~(n24320 ^ n8256);
assign n2934 = n8802 | n16191;
assign n10503 = n11742 & n19600;
assign n24726 = ~(n17371 ^ n15506);
assign n20565 = n23144 | n22125;
assign n22431 = n7675 & n26182;
assign n9938 = ~(n21183 ^ n23364);
assign n14792 = n1076 & n5678;
assign n17042 = n33 & n999;
assign n4028 = n7923 & n11458;
assign n14726 = n5714 | n12531;
assign n14266 = n11026 | n13441;
assign n25589 = ~(n14719 | n1421);
assign n24796 = ~(n14674 ^ n10733);
assign n12124 = n24480 | n16627;
assign n20810 = n26462 | n2208;
assign n17569 = ~(n19805 ^ n11192);
assign n21556 = ~n7099;
assign n4642 = ~n19161;
assign n9986 = ~(n12336 ^ n11752);
assign n21978 = ~(n16665 | n19803);
assign n15693 = ~n9850;
assign n19006 = ~(n18105 | n21392);
assign n6422 = ~(n19048 ^ n16955);
assign n317 = ~(n24912 ^ n8490);
assign n444 = n26264 | n12911;
assign n26676 = n13013 | n14591;
assign n10938 = ~(n13224 ^ n11273);
assign n22281 = ~n21276;
assign n13495 = ~n13036;
assign n12981 = n24328 & n13616;
assign n8219 = ~(n456 ^ n15400);
assign n23051 = n7462 | n6524;
assign n305 = ~(n18737 | n15268);
assign n15984 = ~(n22425 | n14984);
assign n11291 = ~(n8138 | n21656);
assign n18037 = ~(n19387 ^ n14229);
assign n6807 = ~(n26536 ^ n19607);
assign n11973 = ~(n5207 ^ n21284);
assign n3805 = n16878 | n17883;
assign n11893 = ~(n14308 ^ n25979);
assign n15175 = ~(n26791 ^ n2457);
assign n14347 = n2120 & n877;
assign n24877 = ~(n537 | n8456);
assign n6191 = n12237 | n6639;
assign n6000 = n16598 & n2373;
assign n17730 = ~(n21941 ^ n4325);
assign n15214 = n10918 | n12105;
assign n21482 = n25717 & n26608;
assign n22595 = ~(n25475 | n17716);
assign n11072 = n15442 & n17382;
assign n19666 = n8671 & n17181;
assign n25934 = ~(n13541 ^ n12832);
assign n22479 = n21420 | n26573;
assign n19794 = n3909 & n13591;
assign n18969 = n20056 | n13356;
assign n22238 = ~(n14440 | n21287);
assign n18641 = n9177 | n18233;
assign n18374 = n1105 | n21175;
assign n13330 = n5480 | n1067;
assign n19739 = n17280 & n8312;
assign n7396 = ~n10529;
assign n4351 = n7341 | n2954;
assign n10789 = n6924 | n18283;
assign n23355 = ~(n8107 ^ n19891);
assign n6323 = ~(n261 ^ n12538);
assign n286 = ~n15360;
assign n8032 = ~n26748;
assign n1398 = ~(n14148 ^ n1152);
assign n11721 = n5799 & n20067;
assign n9065 = ~(n2514 | n19514);
assign n25990 = n644 | n154;
assign n7871 = ~(n16852 ^ n9967);
assign n14454 = ~(n14777 ^ n3236);
assign n19374 = n8337 & n2493;
assign n1005 = ~(n23847 ^ n2630);
assign n25610 = ~n8088;
assign n12127 = n6113 & n18733;
assign n23469 = n6691 & n19222;
assign n22361 = ~(n19937 ^ n20162);
assign n19699 = n9502 | n1066;
assign n6343 = ~(n24805 ^ n11321);
assign n6082 = ~(n6762 ^ n2289);
assign n20614 = n16937 | n19005;
assign n17591 = n18812 & n22408;
assign n22034 = ~n16582;
assign n19638 = n11562 & n2635;
assign n20902 = n9246 & n12955;
assign n5398 = n22468 | n5679;
assign n14082 = n11269 & n17025;
assign n5161 = ~(n21772 ^ n626);
assign n26801 = ~(n2824 ^ n13827);
assign n16556 = n2269 | n21689;
assign n4508 = ~n10750;
assign n7887 = ~(n25345 ^ n25475);
assign n23526 = n18345 & n20964;
assign n768 = n19279 & n6041;
assign n14491 = n9154 & n3658;
assign n10930 = n9095 | n7913;
assign n2419 = n13992 | n11722;
assign n17394 = n2915 | n10625;
assign n42 = ~n10746;
assign n5974 = ~n20933;
assign n1349 = ~n27055;
assign n9057 = ~(n3582 ^ n21784);
assign n22666 = ~n4108;
assign n4801 = ~(n21027 ^ n13555);
assign n1006 = n2483 & n6079;
assign n8250 = ~(n23191 ^ n25288);
assign n13904 = n11490 & n6856;
assign n16329 = n14490 & n2803;
assign n1002 = n9380 & n7676;
assign n16453 = ~(n17171 | n182);
assign n16710 = n5684 | n8558;
assign n4579 = ~(n10593 | n8657);
assign n23217 = ~n15064;
assign n22157 = ~(n13862 ^ n4015);
assign n24631 = ~(n6731 | n5066);
assign n24596 = ~(n8302 ^ n14545);
assign n23930 = n25371 & n17565;
assign n7854 = n18871 & n21614;
assign n14558 = n6398 | n5251;
assign n8195 = ~(n22615 ^ n14015);
assign n3405 = ~(n25361 ^ n5187);
assign n6537 = n2391 | n19886;
assign n13302 = n2967 | n20179;
assign n6645 = n6299 & n14341;
assign n24387 = ~(n19081 | n21400);
assign n22817 = ~(n7917 | n8391);
assign n11217 = ~n12668;
assign n22058 = ~(n17938 ^ n21455);
assign n22620 = ~(n4842 ^ n24634);
assign n18719 = ~(n17692 ^ n4877);
assign n7340 = n12600 & n3210;
assign n20618 = ~(n2167 ^ n17733);
assign n13191 = ~n25185;
assign n20426 = n5447 & n26811;
assign n3201 = n7898 | n27103;
assign n8865 = n13708 & n13842;
assign n20751 = ~n14153;
assign n8527 = n22707 & n7852;
assign n6211 = n13887 | n7786;
assign n18211 = n17031 & n11868;
assign n24252 = ~(n12762 | n25533);
assign n5707 = ~(n376 ^ n7721);
assign n26511 = ~(n14003 ^ n10920);
assign n14220 = n23153 | n16523;
assign n21638 = n8082 | n24864;
assign n19988 = ~(n9478 ^ n10032);
assign n10857 = n8055 | n12527;
assign n14900 = ~(n19521 ^ n3719);
assign n12646 = n22811 & n15485;
assign n10179 = n7682 & n733;
assign n16016 = n17869 | n24664;
assign n14105 = n13608 & n3768;
assign n13073 = ~n22548;
assign n14586 = n6498 | n5319;
assign n11651 = n6307 & n477;
assign n21025 = n19905 | n21501;
assign n24038 = n776 | n8186;
assign n23334 = n17856 | n21280;
assign n18709 = n12554 | n18295;
assign n23056 = ~(n6178 | n18715);
assign n25505 = ~n7435;
assign n9202 = ~n26075;
assign n11286 = n25591 & n23759;
assign n25502 = ~n10267;
assign n7650 = ~(n18444 ^ n26224);
assign n13633 = ~n5139;
assign n3800 = ~(n14111 ^ n14114);
assign n10309 = n9939 & n6899;
assign n8099 = ~(n7143 | n3625);
assign n20362 = n5673 & n16146;
assign n2757 = n15350 & n22451;
assign n7586 = ~(n3480 | n19911);
assign n23394 = n21650 & n7411;
assign n11572 = n12858 & n1436;
assign n16492 = ~(n21674 ^ n9172);
assign n8985 = ~(n15182 ^ n21915);
assign n688 = ~n6204;
assign n3067 = ~(n5497 ^ n15226);
assign n9786 = n19771 & n3910;
assign n25032 = ~(n19605 ^ n16448);
assign n23578 = ~(n15511 ^ n19192);
assign n3286 = n14288 | n6900;
assign n4039 = ~(n15967 | n1396);
assign n18508 = ~(n20715 | n25065);
assign n22923 = n1709 | n24961;
assign n10320 = n10038 | n23409;
assign n21478 = n9049 | n18524;
assign n14715 = n25335 & n20041;
assign n20248 = ~(n5400 ^ n21997);
assign n7898 = ~(n8509 | n4315);
assign n19907 = ~n19924;
assign n20648 = n22961 | n8342;
assign n8122 = ~(n8495 | n1386);
assign n21201 = n9603 | n10728;
assign n19832 = n3228 | n22470;
assign n17828 = n26725 | n17212;
assign n7324 = ~n3834;
assign n9264 = ~(n17143 | n3007);
assign n17471 = ~(n25345 | n9967);
assign n5722 = ~(n16410 ^ n13652);
assign n448 = ~(n13112 ^ n7707);
assign n17596 = ~(n22724 | n10001);
assign n6752 = ~(n25700 ^ n7281);
assign n17945 = ~(n2723 | n15650);
assign n22993 = ~(n25598 ^ n22503);
assign n18802 = ~(n3382 ^ n1668);
assign n8175 = n7940 | n6309;
assign n14758 = n5613 & n25193;
assign n19202 = ~(n24329 ^ n12683);
assign n16667 = ~(n20968 ^ n24768);
assign n11609 = n13749 & n15741;
assign n19565 = n18366 & n25580;
assign n1992 = ~(n20429 ^ n26054);
assign n13338 = ~(n23730 ^ n24900);
assign n22403 = ~(n26162 | n8806);
assign n4723 = ~(n21633 ^ n24376);
assign n11744 = ~(n3474 ^ n12075);
assign n23310 = ~(n13315 ^ n5503);
assign n10901 = n12849 | n25755;
assign n13819 = n20035 & n12559;
assign n3238 = ~n20792;
assign n25600 = n26252 | n16765;
assign n6251 = ~n19270;
assign n10616 = n5566 & n26676;
assign n4620 = n21644 | n20562;
assign n670 = n5906 & n21851;
assign n13866 = n7980 | n3065;
assign n1180 = ~(n8101 | n17250);
assign n19976 = ~n12395;
assign n291 = n2222 | n8567;
assign n5931 = ~(n2498 | n14185);
assign n23298 = n4764 & n6043;
assign n24825 = ~n13110;
assign n9400 = n21267 | n16874;
assign n26588 = n7452 | n21;
assign n11289 = n7700 & n13758;
assign n26874 = ~(n19215 ^ n8875);
assign n10419 = n18397 & n7720;
assign n21742 = n12164 & n4817;
assign n10360 = ~(n27114 ^ n17727);
assign n11581 = ~(n26951 | n22477);
assign n25297 = n26632 & n17049;
assign n13607 = ~(n17803 ^ n10201);
assign n7987 = ~(n22764 | n1536);
assign n24903 = n23089 & n12877;
assign n27151 = ~n25971;
assign n11937 = n15110 & n16701;
assign n7129 = n17846 | n12488;
assign n21578 = n11045 | n25122;
assign n23406 = n22604 & n2093;
assign n10324 = ~n18444;
assign n2649 = n16835 & n18757;
assign n11878 = n26473 & n16478;
assign n1853 = n19966 & n17281;
assign n20017 = ~(n6505 ^ n6249);
assign n25973 = ~(n15506 | n3246);
assign n27095 = ~(n10922 ^ n16870);
assign n8497 = ~(n2588 ^ n1654);
assign n11519 = n11393 | n3480;
assign n11560 = ~(n6478 | n17590);
assign n7760 = n26731 | n17764;
assign n26311 = ~(n8551 ^ n17071);
assign n10130 = ~(n10885 ^ n26725);
assign n22608 = n26374 | n14028;
assign n17976 = ~(n17606 ^ n9590);
assign n14206 = ~(n26629 ^ n22266);
assign n23716 = n19566 | n10300;
assign n16202 = n26898 & n1149;
assign n8342 = n12833 & n21009;
assign n25397 = n343 | n22302;
assign n15647 = ~n16167;
assign n8893 = n14019 & n651;
assign n14976 = ~(n1584 ^ n17690);
assign n20453 = n16711 | n12464;
assign n21823 = ~(n2446 | n2439);
assign n2770 = n3480 | n7373;
assign n23212 = ~(n3618 ^ n8581);
assign n11419 = ~(n25109 ^ n24514);
assign n10539 = n1322 | n17194;
assign n7664 = ~(n25490 | n12868);
assign n2334 = n14790 & n5105;
assign n4041 = n3652 | n22210;
assign n9903 = n15452 | n22022;
assign n20222 = ~(n18651 | n5855);
assign n244 = n5347 & n14663;
assign n19291 = ~(n3506 ^ n2743);
assign n5187 = n19875 ^ n7057;
assign n13015 = ~(n27102 ^ n21078);
assign n20218 = ~(n20925 ^ n17311);
assign n2506 = n23097 | n11365;
assign n15886 = n1401 | n22478;
assign n420 = ~n5330;
assign n17857 = ~(n11835 ^ n20044);
assign n26075 = n10096 | n22345;
assign n7070 = n11004 | n18081;
assign n7594 = n967 | n23511;
assign n473 = n22605 & n21648;
assign n14965 = ~(n13942 ^ n10222);
assign n19629 = n4567 & n19723;
assign n15556 = ~(n19265 ^ n268);
assign n18843 = ~(n9181 ^ n6928);
assign n19059 = n13863 & n5133;
assign n15209 = ~(n10156 | n20551);
assign n536 = n9003 & n23436;
assign n21085 = ~n21459;
assign n3577 = ~n8070;
assign n8108 = n11544 | n26986;
assign n9294 = ~n13494;
assign n14769 = ~(n15636 ^ n16223);
assign n12676 = n16256 | n12079;
assign n20064 = ~n14702;
assign n14508 = ~(n9093 | n17599);
assign n24025 = ~n23504;
assign n11764 = ~n2429;
assign n23095 = ~n7751;
assign n13478 = ~(n14830 ^ n6468);
assign n19441 = n12067 | n6067;
assign n8625 = ~(n4613 | n6561);
assign n23214 = n14707 | n6049;
assign n799 = n18872 | n5254;
assign n1842 = n11653 | n14926;
assign n789 = ~(n3196 ^ n2046);
assign n22027 = ~(n10238 ^ n3300);
assign n11701 = ~(n12142 ^ n6787);
assign n17137 = ~(n1642 | n10158);
assign n9783 = ~(n25456 ^ n4408);
assign n18049 = n20305 & n2179;
assign n14529 = n11159 | n10186;
assign n19763 = ~(n23966 | n13925);
assign n25698 = n26892 & n11623;
assign n9466 = n4514 & n5111;
assign n25169 = n13033 | n18907;
assign n3329 = ~(n2342 | n23430);
assign n13497 = ~n2117;
assign n19591 = n1663 & n3777;
assign n18413 = ~(n7237 | n25120);
assign n5347 = n1994 | n19556;
assign n25125 = n5589 & n7934;
assign n8134 = n14936 & n20423;
assign n18826 = ~(n20763 ^ n12013);
assign n18217 = n10335 & n10141;
assign n19505 = n11059 & n23948;
assign n9704 = n19461 | n6440;
assign n19687 = n13870 | n13029;
assign n6524 = n1157 & n20765;
assign n21151 = ~n19394;
assign n10252 = ~(n20462 | n7086);
assign n26205 = ~(n10335 ^ n9954);
assign n1644 = n16252 | n23166;
assign n3530 = n6927 | n5344;
assign n10745 = ~(n8614 ^ n12702);
assign n13072 = ~(n15497 ^ n26509);
assign n114 = n9325 | n17633;
assign n8181 = n19236 | n4275;
assign n23739 = n8068 | n25316;
assign n2830 = n12447 | n23599;
assign n6189 = ~(n14938 ^ n22497);
assign n770 = n13809 | n4512;
assign n23870 = n8158 & n2475;
assign n12435 = ~(n7882 | n24727);
assign n4115 = ~(n1173 ^ n583);
assign n3902 = ~(n7910 ^ n8309);
assign n15304 = ~(n23068 ^ n20179);
assign n478 = n8853 | n17652;
assign n11902 = n6379 | n3040;
assign n1342 = n25743 | n17751;
assign n9678 = ~n25426;
assign n1111 = ~(n8912 ^ n9474);
assign n10838 = ~(n7305 ^ n1204);
assign n13802 = ~(n26807 | n9273);
assign n19007 = n21424 | n1318;
assign n22464 = n7549 & n15247;
assign n7728 = n12420 | n24143;
assign n12674 = ~(n6810 ^ n9375);
assign n10964 = n7276;
assign n3328 = n5033 & n3177;
assign n11300 = ~(n19836 ^ n27121);
assign n24264 = ~(n20542 | n25937);
assign n23216 = ~(n518 ^ n18619);
assign n12158 = ~(n4262 ^ n20786);
assign n5589 = n13154 | n4426;
assign n221 = n12871 | n20411;
assign n23457 = n11144 & n25500;
assign n17565 = n26166 | n2106;
assign n4441 = ~(n6793 ^ n18459);
assign n7487 = ~(n14486 | n18031);
assign n11483 = ~n18438;
assign n13446 = n24226 & n3112;
assign n7420 = ~(n676 ^ n3981);
assign n15161 = n24869 & n1392;
assign n6778 = ~(n22170 | n5098);
assign n856 = ~n6129;
assign n21531 = n26227 | n21284;
assign n13651 = ~n18927;
assign n4088 = ~(n11065 ^ n13869);
assign n3437 = n24453 | n23844;
assign n12371 = ~n11209;
assign n26787 = n22591 | n24756;
assign n11717 = ~(n21140 ^ n10241);
assign n25791 = n19941 & n9345;
assign n10165 = ~(n17825 ^ n20574);
assign n1194 = n5881 & n4206;
assign n3146 = n18892 | n25482;
assign n9691 = ~(n18742 ^ n20409);
assign n17274 = n9383 | n21283;
assign n13222 = ~(n25915 ^ n8024);
assign n26828 = ~(n11615 | n8052);
assign n20831 = n18103 | n5182;
assign n23656 = ~(n11829 | n12935);
assign n18956 = n6623 | n2837;
assign n1506 = n9040 | n26799;
assign n22422 = ~n4856;
assign n14583 = ~(n15967 ^ n2783);
assign n25962 = ~(n12956 | n26913);
assign n26153 = n2895 & n16972;
assign n8689 = ~n10183;
assign n7870 = ~(n19905 | n14733);
assign n13528 = ~n17452;
assign n14736 = ~n19472;
assign n19427 = ~n17739;
assign n6981 = n20338 | n20477;
assign n373 = n16438 & n2569;
assign n10133 = n13715 | n10634;
assign n12564 = n7114 & n9746;
assign n9720 = n26802 & n18110;
assign n25947 = ~(n17987 ^ n15683);
assign n21879 = ~(n23291 ^ n14201);
assign n13644 = n688 | n3795;
assign n1908 = n26482 | n26089;
assign n15255 = ~(n12573 ^ n5614);
assign n20900 = n6198 & n9544;
assign n20855 = n8191 | n12645;
assign n21909 = ~(n21205 ^ n5226);
assign n7562 = n20400 | n13520;
assign n21689 = n17459 & n5216;
assign n11113 = ~n17233;
assign n10493 = ~(n17134 ^ n21573);
assign n12681 = n7255 & n22598;
assign n1709 = ~(n8951 ^ n9775);
assign n26147 = n17513 & n26490;
assign n22723 = ~n13668;
assign n8233 = ~(n13164 ^ n12060);
assign n5803 = ~(n22442 ^ n22253);
assign n24686 = ~n11458;
assign n17033 = n1743 & n25598;
assign n6328 = ~(n16283 ^ n17037);
assign n19141 = ~(n18393 ^ n5336);
assign n11111 = ~n7234;
assign n24964 = ~(n14761 ^ n6218);
assign n7345 = ~(n24599 ^ n9398);
assign n24454 = n4500 | n855;
assign n25891 = ~(n2463 ^ n5677);
assign n13405 = ~n8305;
assign n18642 = n25038 | n16544;
assign n11987 = ~(n10749 ^ n21487);
assign n5520 = n7960 & n7015;
assign n14590 = n26366 & n17080;
assign n19410 = n6659 & n20384;
assign n20935 = ~(n13057 ^ n17032);
assign n8583 = n14440 | n3504;
assign n10260 = ~(n22755 ^ n7503);
assign n782 = ~(n26437 | n25415);
assign n14185 = ~n26058;
assign n8404 = n7880 | n3389;
assign n22586 = ~(n19701 ^ n13074);
assign n18096 = n4468 | n2780;
assign n17161 = n9073 | n17044;
assign n25714 = n26995 | n25344;
assign n17737 = ~(n3890 | n12465);
assign n10028 = ~(n23865 | n19200);
assign n19764 = n19050 | n19130;
assign n27158 = ~(n10196 ^ n2234);
assign n5890 = ~(n20323 | n7835);
assign n10136 = n5580 | n19911;
assign n6194 = n16866 & n18066;
assign n19032 = n7524 & n10314;
assign n1663 = n18639 | n16097;
assign n23537 = ~n17183;
assign n2310 = n15063 & n16253;
assign n24598 = n25138 | n19784;
assign n21711 = n10109 | n4007;
assign n23734 = n26640 | n18175;
assign n27076 = ~n7592;
assign n1449 = ~n21927;
assign n16940 = ~(n4041 ^ n3378);
assign n11112 = ~(n17453 | n10250);
assign n12508 = ~(n11923 ^ n17237);
assign n8518 = ~(n16968 ^ n23120);
assign n4350 = n6790 & n10000;
assign n25758 = ~(n16197 ^ n9381);
assign n24950 = n25724 | n2173;
assign n6130 = ~(n5751 ^ n25184);
assign n25680 = ~(n20409 | n18227);
assign n762 = ~n25575;
assign n22639 = ~(n2058 ^ n5954);
assign n9485 = ~(n9311 ^ n12829);
assign n12775 = ~(n2510 ^ n8324);
assign n16279 = ~(n6326 ^ n2211);
assign n21374 = n11577 & n24244;
assign n25236 = n9823 | n25842;
assign n26273 = ~(n19039 | n13633);
assign n8941 = n14439 & n11661;
assign n11812 = ~(n8382 ^ n10352);
assign n3167 = n1766 & n25280;
assign n17151 = ~(n13453 | n14733);
assign n23339 = n2126 | n20624;
assign n1324 = ~(n26650 ^ n23422);
assign n24674 = n14336 | n9349;
assign n26095 = ~n24517;
assign n6733 = ~(n11572 ^ n23259);
assign n4933 = ~(n2518 ^ n1637);
assign n21593 = ~n23722;
assign n26817 = ~(n3737 | n25367);
assign n21394 = n14450 & n22866;
assign n4679 = n20289 | n25192;
assign n12803 = n20571 & n5595;
assign n8314 = ~(n22780 ^ n5752);
assign n5993 = ~n26420;
assign n6536 = ~(n8166 ^ n26413);
assign n12000 = ~(n13226 ^ n9324);
assign n13924 = ~(n23369 | n18255);
assign n23860 = ~(n25929 | n10013);
assign n21266 = ~(n10096 ^ n16824);
assign n26951 = ~n19709;
assign n6749 = n19530 & n23992;
assign n21493 = n8204 & n27094;
assign n22387 = ~n4112;
assign n9459 = ~(n23972 ^ n22004);
assign n26061 = ~(n21257 | n25935);
assign n18878 = ~(n14440 ^ n21287);
assign n7946 = ~(n26456 ^ n14973);
assign n1666 = n8360 | n18396;
assign n23408 = ~n21753;
assign n25605 = ~(n333 ^ n22091);
assign n25383 = n5487 & n14682;
assign n1796 = ~(n19852 | n23035);
assign n21723 = ~(n23127 ^ n22908);
assign n2417 = n12124 & n22429;
assign n21474 = n19555 & n21655;
assign n667 = n20044 | n11835;
assign n18739 = n13248 | n15219;
assign n13069 = ~(n7531 ^ n26195);
assign n7429 = ~n5915;
assign n16687 = ~n19890;
assign n8475 = n9267 & n10808;
assign n5653 = n15866 | n16552;
assign n16910 = n21562 | n3865;
assign n11950 = n7847 & n20195;
assign n9109 = n4420 & n26975;
assign n17278 = n5352 & n24339;
assign n5935 = n21867 | n8557;
assign n26352 = n17205 | n3042;
assign n18097 = ~n7134;
assign n11067 = n11680 | n24378;
assign n18357 = ~n14106;
assign n23063 = ~n20138;
assign n1545 = ~(n25051 ^ n13642);
assign n9841 = ~(n11918 ^ n20250);
assign n1640 = ~(n7058 ^ n22625);
assign n5123 = ~(n26994 ^ n4257);
assign n9863 = ~(n23612 | n8167);
assign n3446 = n21380 | n3018;
assign n2426 = ~(n8964 ^ n23200);
assign n18480 = n14842 & n11475;
assign n16842 = ~(n22933 | n11185);
assign n4617 = n23627 | n12165;
assign n6245 = ~(n3109 ^ n25786);
assign n893 = n2495 | n18804;
assign n25084 = n6780 | n961;
assign n19616 = ~n4665;
assign n10439 = n17784 | n725;
assign n25414 = ~(n18385 | n22840);
assign n14793 = n21978 | n19953;
assign n7844 = n21937 | n9219;
assign n82 = ~(n9251 ^ n16968);
assign n11429 = n17824 | n5955;
assign n7832 = ~n5559;
assign n4089 = ~(n6259 ^ n14665);
assign n25047 = n12762 | n4263;
assign n22645 = n13447 | n2072;
assign n1694 = ~n4616;
assign n11706 = ~(n20967 ^ n1314);
assign n18525 = n24625 | n11497;
assign n5252 = ~(n10135 ^ n552);
assign n15399 = ~(n2060 ^ n6660);
assign n25807 = n13753 & n16792;
assign n17771 = ~(n5863 ^ n20838);
assign n13368 = ~n6637;
assign n11150 = n9882 & n23338;
assign n11071 = ~(n17547 ^ n13755);
assign n4075 = ~(n12184 ^ n17322);
assign n15722 = ~(n2035 | n26823);
assign n18614 = n11999 & n5759;
assign n2891 = ~n12391;
assign n24644 = n20866 & n13574;
assign n15513 = ~(n6175 | n17967);
assign n2617 = ~(n7743 | n2328);
assign n22680 = n25123 & n15283;
assign n14210 = n16400 & n17561;
assign n701 = n11236 | n15231;
assign n18245 = n2743 | n1584;
assign n25235 = ~n9312;
assign n14867 = n22524 & n2276;
assign n15545 = n5929 | n24536;
assign n12412 = ~(n13368 ^ n7260);
assign n26040 = n68 | n25677;
assign n16571 = n922 & n13030;
assign n7004 = ~(n16642 ^ n8386);
assign n22670 = ~n2764;
assign n11504 = ~(n3175 ^ n24973);
assign n19883 = n25674 | n9992;
assign n12399 = ~(n10372 ^ n20235);
assign n1661 = n14130 | n12861;
assign n7048 = ~(n26695 | n15944);
assign n14547 = ~(n7615 ^ n6586);
assign n24034 = n11443 | n17303;
assign n24987 = n3506 | n26414;
assign n8542 = n8895 & n13727;
assign n2744 = n13159 | n10611;
assign n661 = ~(n16353 ^ n3485);
assign n18272 = ~(n3687 ^ n24879);
assign n6371 = ~(n12716 ^ n18862);
assign n3867 = ~(n7442 | n12485);
assign n23538 = n11349 | n20160;
assign n17068 = ~(n13381 ^ n6746);
assign n27187 = ~(n3610 | n25546);
assign n24404 = ~(n25998 ^ n17470);
assign n635 = ~(n6682 | n23084);
assign n26742 = n21853 & n20468;
assign n25768 = n19861 & n13397;
assign n7465 = ~n24399;
assign n4534 = n988 & n24642;
assign n15080 = n11380 | n5411;
assign n20187 = ~(n5653 ^ n23959);
assign n969 = n5544 & n1296;
assign n24318 = ~(n7744 ^ n2266);
assign n10645 = ~(n21412 ^ n1195);
assign n18117 = n2156 | n26332;
assign n1026 = ~n22640;
assign n24974 = ~n22068;
assign n17653 = ~(n5188 ^ n18481);
assign n16563 = n5123 | n15482;
assign n5948 = ~n22554;
assign n1604 = ~(n25164 ^ n9270);
assign n20446 = ~(n14240 ^ n5865);
assign n22911 = n17122 | n23383;
assign n1698 = ~(n863 ^ n25370);
assign n2786 = n9491 & n8392;
assign n26025 = ~(n15512 ^ n15147);
assign n11418 = n21083 | n8052;
assign n20852 = ~(n6750 | n14680);
assign n7144 = ~(n7146 ^ n3549);
assign n6455 = n9481 & n16741;
assign n8319 = ~(n11551 ^ n15393);
assign n16655 = n7689 | n10807;
assign n22073 = n15455 & n20310;
assign n15278 = ~(n154 ^ n7722);
assign n12637 = n26556 | n10917;
assign n859 = n19911 & n5580;
assign n4407 = ~(n1066 ^ n25872);
assign n24885 = n21997 | n15773;
assign n26696 = ~(n56 ^ n16472);
assign n6672 = ~(n8838 | n1987);
assign n6710 = n442 | n7445;
assign n7656 = n426 | n19943;
assign n23869 = n21632 | n13190;
assign n8712 = n6417 & n21899;
assign n9440 = ~(n22200 ^ n17805);
assign n4976 = n15901 | n9418;
assign n24949 = n18762 & n12027;
assign n5058 = ~(n16083 ^ n12161);
assign n3505 = n9465 | n4074;
assign n17830 = n23408 & n25921;
assign n26562 = ~(n162 ^ n19568);
assign n13895 = ~(n13781 ^ n9251);
assign n7535 = ~n11876;
assign n21781 = ~(n19090 | n17166);
assign n23632 = ~(n6705 ^ n8614);
assign n11331 = n6218 | n9296;
assign n17079 = n15767 | n26733;
assign n2463 = n26569 & n23465;
assign n9421 = n15826 & n21585;
assign n15789 = n8847 | n3651;
assign n22721 = ~(n25974 ^ n2355);
assign n11280 = n13340 | n24186;
assign n20678 = ~(n529 ^ n2488);
assign n8564 = ~n21284;
assign n16980 = n25738 | n6861;
assign n18204 = ~(n3949 ^ n5961);
assign n6504 = ~n15936;
assign n19660 = ~(n16933 ^ n15672);
assign n6758 = n13903 | n14073;
assign n1528 = ~(n17573 ^ n11029);
assign n15593 = ~(n15087 ^ n23272);
assign n18658 = n13546 | n9831;
assign n23681 = ~n789;
assign n4367 = n16462 | n10135;
assign n10937 = n2628 & n8786;
assign n4312 = ~(n14830 | n26584);
assign n24307 = ~(n12020 ^ n5164);
assign n4774 = ~(n15185 ^ n22169);
assign n22813 = n5221 | n2157;
assign n18125 = ~(n1453 ^ n27179);
assign n6521 = ~n5101;
assign n19557 = ~(n19673 | n5678);
assign n11557 = ~(n10767 ^ n4031);
assign n13432 = n15238 | n4571;
assign n7609 = n24665 | n1687;
assign n5672 = n20206 | n10250;
assign n21200 = n6621 & n10062;
assign n2597 = ~n11121;
assign n25530 = ~(n16562 | n15170);
assign n26692 = n12422 | n19087;
assign n20933 = ~(n5153 ^ n12548);
assign n26100 = ~n19143;
assign n16475 = ~(n15012 | n7401);
assign n13604 = n8177 & n3585;
assign n17416 = n23709 | n16267;
assign n22424 = n483 | n6566;
assign n20802 = ~(n2608 ^ n13553);
assign n12852 = ~(n4459 ^ n19391);
assign n2793 = n24876 | n24037;
assign n13466 = ~(n26289 ^ n14273);
assign n4242 = ~(n11361 ^ n13208);
assign n1802 = ~(n1456 ^ n10405);
assign n16316 = n2355 | n16223;
assign n25856 = n12921 & n17197;
assign n6070 = ~n16900;
assign n6244 = ~(n21880 | n9007);
assign n725 = ~(n7535 ^ n9003);
assign n1845 = ~(n20538 ^ n17873);
assign n5518 = ~(n14777 | n21442);
assign n1832 = n27202 | n15949;
assign n25175 = n25050 | n23281;
assign n4213 = n20554 & n25806;
assign n16143 = n364 | n6083;
assign n11414 = ~(n22916 ^ n11213);
assign n9199 = ~(n10861 ^ n21857);
assign n19079 = n12800 | n26498;
assign n12273 = ~(n19429 ^ n14610);
assign n21683 = ~(n17397 ^ n18227);
assign n18950 = ~(n6960 ^ n10150);
assign n12432 = n566 | n374;
assign n9041 = n10983 | n23562;
assign n21567 = ~(n23536 ^ n14899);
assign n10652 = n20232 & n12970;
assign n8823 = ~(n11816 ^ n24954);
assign n12354 = ~n8920;
assign n25146 = n2606 | n17211;
assign n16719 = ~(n20920 ^ n17911);
assign n21740 = ~(n9769 ^ n15955);
assign n20744 = n24255 & n9604;
assign n310 = ~n8729;
assign n23183 = n26947 | n15639;
assign n11733 = ~(n26924 ^ n24861);
assign n19588 = ~n15884;
assign n9701 = n23665 & n13355;
assign n19143 = ~(n7594 ^ n6991);
assign n21767 = ~(n23512 | n9124);
assign n15135 = ~(n16700 ^ n9321);
assign n3108 = n6580 | n11350;
assign n4034 = n11665 | n20211;
assign n3045 = ~n4618;
assign n14222 = ~(n20812 ^ n24596);
assign n17238 = n14117 | n5824;
assign n24469 = ~(n9502 | n2168);
assign n837 = n8745 | n8479;
assign n25773 = ~(n16076 ^ n1728);
assign n7583 = ~(n11841 ^ n17077);
assign n4293 = ~(n7451 ^ n8874);
assign n241 = n24426 & n3574;
assign n10977 = n3627 & n9367;
assign n21416 = n25494 & n10713;
assign n2974 = n26324 | n6359;
assign n7000 = ~(n23141 | n1370);
assign n5064 = ~(n568 ^ n14865);
assign n11729 = n11035 & n25266;
assign n3977 = ~(n25475 | n23697);
assign n14641 = n26793 | n25067;
assign n23072 = n921 & n10590;
assign n21811 = n12713 | n180;
assign n16659 = ~(n21613 ^ n6242);
assign n26467 = ~n560;
assign n11629 = n6234 | n14384;
assign n9797 = ~(n24770 ^ n13445);
assign n13869 = ~(n14754 ^ n26344);
assign n4876 = ~(n15182 | n26797);
assign n6116 = n20159 | n10884;
assign n21450 = ~n9110;
assign n21569 = n10578 | n5901;
assign n15826 = ~n23146;
assign n20348 = n13561 | n14148;
assign n26677 = ~n4335;
assign n12197 = n17128 | n26912;
assign n24829 = ~(n3131 ^ n22442);
assign n3151 = ~(n10057 ^ n5026);
assign n19901 = n11452 | n26823;
assign n4150 = ~(n13394 ^ n5997);
assign n24417 = ~n5822;
assign n8860 = n16755 | n20326;
assign n2938 = ~(n26799 ^ n12059);
assign n23535 = n2331 | n4587;
assign n11495 = n20133 | n5255;
assign n638 = ~(n2224 ^ n20603);
assign n6064 = n13351 | n7622;
assign n25320 = ~(n6724 | n6127);
assign n10711 = ~n19107;
assign n8187 = n5446 | n22647;
assign n25644 = ~(n811 | n13609);
assign n17387 = n18855 | n8787;
assign n8523 = ~(n3173 ^ n25393);
assign n1679 = n22290 & n12878;
assign n3097 = ~(n24350 ^ n6062);
assign n4356 = ~(n26773 ^ n19301);
assign n23245 = ~(n16687 | n20906);
assign n5405 = n18955 & n11887;
assign n6976 = n4471 | n8168;
assign n1124 = n14895 | n24409;
assign n15833 = n11622 | n9276;
assign n16538 = n20194 & n12089;
assign n25333 = n7953 | n13894;
assign n12614 = ~(n21823 | n11702);
assign n9999 = n26380 | n18974;
assign n13957 = n6898 | n6448;
assign n22972 = ~(n17656 ^ n25267);
assign n26307 = ~n14366;
assign n844 = ~(n11302 | n24786);
assign n21490 = n11339 | n5870;
assign n24066 = n2137 | n11085;
assign n3537 = n25674 | n21832;
assign n26541 = ~(n1010 ^ n9238);
assign n2080 = ~n8708;
assign n10654 = n3756 & n4354;
assign n9006 = ~(n3909 ^ n268);
assign n1649 = n20530 | n11394;
assign n11857 = n11544 | n2160;
assign n9117 = n4435 | n8533;
assign n19721 = n7804 & n4716;
assign n23036 = ~n21879;
assign n1208 = n21148 | n15988;
assign n17643 = ~(n3837 ^ n1040);
assign n18119 = ~(n22198 | n575);
assign n16337 = ~(n11580 ^ n2035);
assign n20146 = ~n4851;
assign n3344 = ~(n1370 ^ n26054);
assign n23865 = ~n24106;
assign n9648 = ~(n10871 ^ n17637);
assign n22168 = n10097 | n11974;
assign n17754 = ~(n19534 ^ n13319);
assign n18610 = ~(n1497 ^ n433);
assign n18740 = n10802 | n15903;
assign n263 = ~(n20311 | n20741);
assign n22630 = n2504 & n25860;
assign n17537 = ~(n15715 | n14954);
assign n24586 = n21538 | n6725;
assign n14060 = n13017 | n21483;
assign n16441 = ~(n23913 ^ n3710);
assign n16381 = n4761 & n8683;
assign n10448 = ~(n4018 ^ n19747);
assign n18354 = n10963 | n12969;
assign n24666 = ~n6606;
assign n660 = n17580 | n11008;
assign n24525 = n5888 & n4653;
assign n20452 = n14806 & n10270;
assign n18893 = n24494 & n14080;
assign n5778 = n21972 | n17120;
assign n1982 = ~(n10571 ^ n9172);
assign n23441 = ~n11266;
assign n8890 = n6611 & n26895;
assign n24117 = ~(n17564 ^ n26196);
assign n7071 = ~n24608;
assign n4714 = ~(n7488 ^ n13310);
assign n17395 = ~(n27170 ^ n1136);
assign n12663 = ~(n25691 ^ n13783);
assign n2742 = ~(n21912 ^ n9291);
assign n4804 = ~(n15267 ^ n2010);
assign n2841 = ~(n21075 ^ n16828);
assign n7791 = ~(n23280 ^ n4162);
assign n5514 = ~(n7130 | n2044);
assign n10 = n20201 & n20231;
assign n17342 = ~(n15053 ^ n3828);
assign n20945 = ~n12445;
assign n26331 = n3972 | n14396;
assign n8622 = ~(n2231 ^ n14070);
assign n24623 = ~(n12713 | n24701);
assign n13595 = ~(n5938 ^ n5987);
assign n3474 = ~(n3560 ^ n8863);
assign n17690 = ~(n272 ^ n19291);
assign n330 = ~(n6340 ^ n23667);
assign n9823 = ~(n7377 | n5629);
assign n1445 = n20261 | n13632;
assign n12747 = n24531 & n13852;
assign n13354 = ~(n8704 ^ n3488);
assign n7176 = n25342 | n16662;
assign n10298 = ~(n18601 ^ n13533);
assign n10648 = n11393 | n13359;
assign n1780 = ~n19087;
assign n25735 = ~(n9700 ^ n25210);
assign n18607 = ~n22826;
assign n9532 = ~(n23722 ^ n20972);
assign n1249 = ~(n12075 ^ n4957);
assign n19711 = ~(n22930 ^ n19327);
assign n21052 = ~(n24825 | n21317);
assign n14184 = ~(n3876 ^ n3748);
assign n22324 = n20820 | n16058;
assign n21613 = ~n23411;
assign n20819 = n10194 | n9597;
assign n20999 = ~(n2080 ^ n1319);
assign n8582 = ~n19904;
assign n4575 = ~n9545;
assign n22855 = ~(n21957 | n14156);
assign n12368 = n490 & n26755;
assign n13106 = ~(n25126 | n19575);
assign n8091 = n5044 | n10635;
assign n9249 = ~(n25797 | n15784);
assign n14812 = n25762 | n15612;
assign n17303 = n11362 & n6326;
assign n22320 = n11559 | n16693;
assign n8755 = n19706 | n4720;
assign n7318 = n4973 & n16815;
assign n9219 = ~(n17923 ^ n1752);
assign n11824 = ~(n20007 ^ n11799);
assign n6605 = n13898 | n6502;
assign n22848 = n19598 & n4251;
assign n19947 = ~(n10833 ^ n4042);
assign n9344 = ~(n14413 ^ n9175);
assign n11478 = n18224 | n6640;
assign n22957 = n8749 | n12972;
assign n6573 = n12022 | n8889;
assign n4103 = ~(n11164 ^ n22251);
assign n6915 = ~(n14876 ^ n2472);
assign n6458 = ~(n22176 ^ n19922);
assign n6201 = ~(n19439 | n22747);
assign n22531 = ~(n1690 ^ n1000);
assign n4803 = n3018 & n21380;
assign n21462 = ~(n12638 ^ n7026);
assign n22546 = ~(n23313 ^ n2586);
assign n24296 = n13128 & n10662;
assign n10314 = ~n1541;
assign n1179 = ~(n17705 | n22421);
assign n2940 = n23234 | n7682;
assign n18147 = n7290 | n18758;
assign n7529 = ~n2646;
assign n16032 = n2710 & n1124;
assign n18251 = n19652 | n21916;
assign n15300 = ~(n13599 ^ n564);
assign n19787 = n200 | n25247;
assign n17955 = n14586 & n14729;
assign n15200 = ~(n25041 | n25643);
assign n3332 = ~(n16123 ^ n497);
assign n11859 = n678 | n3921;
assign n2211 = ~(n15616 ^ n9215);
assign n3209 = ~(n6703 ^ n11321);
assign n26624 = n13406 | n8471;
assign n8671 = n21293 | n2926;
assign n6929 = ~(n10966 | n19789);
assign n27182 = ~(n20840 | n21948);
assign n10691 = ~n20210;
assign n2872 = ~n20731;
assign n15131 = ~n4890;
assign n2327 = ~(n17321 ^ n1053);
assign n25699 = n6222 & n9744;
assign n18560 = ~(n642 | n21194);
assign n1400 = n9594 & n5915;
assign n21940 = ~(n725 ^ n24804);
assign n25403 = ~n22008;
assign n13276 = ~(n19520 ^ n20077);
assign n5138 = n17457 & n10828;
assign n8932 = ~(n6915 | n9748);
assign n12994 = n1263 | n9885;
assign n6884 = ~(n4479 ^ n11986);
assign n12184 = ~n16494;
assign n2989 = ~(n4199 ^ n23101);
assign n12199 = n18511 | n14361;
assign n2578 = ~(n6761 ^ n7122);
assign n23062 = n2027 | n26942;
assign n16846 = ~(n5100 ^ n14200);
assign n9352 = n19836 | n3835;
assign n13249 = ~n2784;
assign n7939 = ~(n4801 | n9723);
assign n18469 = n15260 | n26148;
assign n4466 = n23932 | n10666;
assign n9572 = ~n16201;
assign n22018 = n10873 | n25250;
assign n15831 = ~(n20657 ^ n3799);
assign n749 = n24330 | n5320;
assign n12387 = n26565 & n9142;
assign n7310 = ~(n23921 ^ n11302);
assign n14835 = ~(n6011 ^ n13137);
assign n20310 = n18085 | n5157;
assign n19724 = ~(n1405 ^ n3317);
assign n7327 = ~n18988;
assign n11696 = ~(n16396 ^ n8399);
assign n9271 = n27155 | n10803;
assign n10027 = ~(n1123 ^ n26137);
assign n659 = n24755 | n22295;
assign n15453 = ~(n26363 | n1553);
assign n21346 = n25324 | n1642;
assign n12648 = ~(n5075 ^ n9241);
assign n675 = n20921 | n25106;
assign n2666 = ~(n21704 ^ n7751);
assign n10573 = ~(n19978 ^ n24239);
assign n9645 = ~(n2705 ^ n19551);
assign n226 = n718 | n7158;
assign n18386 = ~(n8351 | n11066);
assign n25176 = ~(n3382 | n18363);
assign n5719 = ~n468;
assign n11129 = ~(n455 ^ n6387);
assign n16937 = ~n7149;
assign n23801 = ~(n11579 ^ n3962);
assign n1615 = n11393 | n12956;
assign n22215 = ~(n1645 ^ n3978);
assign n11945 = ~(n20177 ^ n14946);
assign n18320 = n19905 | n2547;
assign n8367 = ~n25749;
assign n25537 = n18996 & n23461;
assign n7526 = ~(n19633 ^ n5427);
assign n16497 = ~(n677 | n24243);
assign n25262 = n24852 & n20487;
assign n13314 = n19042 | n18846;
assign n23550 = ~(n17602 ^ n14843);
assign n25151 = n12371 | n10534;
assign n9490 = ~n17653;
assign n5750 = ~(n13616 ^ n20263);
assign n22504 = n16309 | n20391;
assign n17093 = n22741 | n3944;
assign n5065 = ~n6819;
assign n12265 = ~(n21197 ^ n6125);
assign n13155 = ~(n10312 ^ n10013);
assign n26487 = n14079 | n5758;
assign n8992 = n14292 | n9876;
assign n7060 = ~(n5390 ^ n5081);
assign n6278 = ~(n14254 ^ n14610);
assign n5996 = n4179 & n10959;
assign n26509 = ~(n5852 ^ n19971);
assign n17153 = n26139 | n2952;
assign n4266 = ~(n17724 ^ n22633);
assign n22787 = ~(n7422 ^ n20917);
assign n13075 = ~(n23097 ^ n19568);
assign n22103 = n17551 | n8785;
assign n13105 = n19673 | n12416;
assign n3778 = ~n3859;
assign n23452 = ~(n17223 | n4488);
assign n12504 = n9766 | n16918;
assign n12787 = n10201 | n19691;
assign n3840 = ~n7797;
assign n15927 = ~(n5143 ^ n19625);
assign n26931 = ~(n23331 ^ n20604);
assign n20745 = n17088 & n5241;
endmodule
