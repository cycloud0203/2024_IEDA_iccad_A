// Benchmark "top_810026173_843396535_809698999_829556405_809567927" written by ABC on Mon Jul 15 23:49:29 2024

module top_810026173_843396535_809698999_829556405_809567927 ( 
    n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583, n604,
    n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099, n1112,
    n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279, n1288,
    n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536, n1558,
    n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689, n1738,
    n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035, n2088,
    n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210, n2272,
    n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421, n2479,
    n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809, n2816,
    n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030, n3136,
    n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324, n3349,
    n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582, n3618,
    n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945, n3952,
    n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306, n4319,
    n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665, n4722,
    n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026, n5031,
    n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211, n5213,
    n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438, n5443,
    n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752, n5822,
    n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369, n6379,
    n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556, n6590,
    n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785, n6790,
    n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149, n7305,
    n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524, n7566,
    n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721, n7731,
    n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949, n7963,
    n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285, n8305,
    n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581, n8614,
    n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806, n8827,
    n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246, n9251,
    n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460, n9493,
    n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872, n9926,
    n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096, n10117,
    n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411, n10514,
    n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739, n10763,
    n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201, n11220,
    n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473, n11479,
    n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630, n11667,
    n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113, n12121,
    n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384, n12398,
    n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626, n12650,
    n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892, n12900,
    n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190, n13263,
    n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490, n13494,
    n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781, n13783,
    n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148, n14230,
    n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576, n14603,
    n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826, n14899,
    n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258, n15271,
    n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539, n15546,
    n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884, n15918,
    n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223, n16247,
    n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521, n16524,
    n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911, n16968,
    n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090, n17095,
    n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911, n17954,
    n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171, n18227,
    n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483, n18496,
    n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745, n18880,
    n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081, n19107,
    n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282, n19327,
    n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515, n19531,
    n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701, n19770,
    n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036, n20040,
    n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250, n20259,
    n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470, n20478,
    n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929, n20946,
    n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276, n21287,
    n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654, n21674,
    n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839, n21898,
    n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043, n22068,
    n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290, n22309,
    n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470, n22492,
    n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660, n22764,
    n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065, n23068,
    n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304, n23333,
    n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586, n23657,
    n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895, n23912,
    n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093, n24129,
    n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374, n24485,
    n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937, n25023,
    n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168, n25240,
    n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381, n25435,
    n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629, n25643,
    n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923, n25926,
    n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180, n26191,
    n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510, n26512,
    n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748, n26752,
    n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037, n27089,
    n27104, n27120, n27134, n27188,
    n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194  );
  input  n18, n21, n196, n268, n329, n337, n342, n376, n442, n468, n583,
    n604, n626, n647, n655, n752, n767, n919, n932, n987, n1040, n1099,
    n1112, n1118, n1136, n1152, n1163, n1204, n1222, n1255, n1269, n1279,
    n1288, n1293, n1314, n1320, n1432, n1437, n1451, n1483, n1525, n1536,
    n1558, n1611, n1630, n1639, n1654, n1662, n1667, n1681, n1682, n1689,
    n1738, n1742, n1752, n1777, n1831, n1881, n1949, n1999, n2013, n2035,
    n2088, n2102, n2113, n2117, n2145, n2146, n2160, n2175, n2184, n2210,
    n2272, n2289, n2328, n2331, n2355, n2387, n2409, n2416, n2420, n2421,
    n2479, n2547, n2570, n2646, n2659, n2680, n2731, n2743, n2783, n2809,
    n2816, n2858, n2886, n2944, n2978, n2979, n2985, n2999, n3018, n3030,
    n3136, n3161, n3164, n3228, n3253, n3260, n3279, n3306, n3320, n3324,
    n3349, n3366, n3425, n3460, n3468, n3480, n3506, n3541, n3570, n3582,
    n3618, n3710, n3740, n3785, n3795, n3828, n3909, n3918, n3925, n3945,
    n3952, n3959, n3962, n3984, n4085, n4100, n4119, n4256, n4272, n4306,
    n4319, n4325, n4326, n4376, n4409, n4426, n4514, n4588, n4590, n4665,
    n4722, n4812, n4858, n4913, n4939, n4957, n4964, n4967, n5025, n5026,
    n5031, n5060, n5077, n5098, n5101, n5115, n5128, n5131, n5140, n5211,
    n5213, n5226, n5255, n5302, n5330, n5337, n5376, n5386, n5400, n5438,
    n5443, n5451, n5517, n5521, n5532, n5579, n5605, n5696, n5704, n5752,
    n5822, n5834, n5842, n5882, n6104, n6105, n6204, n6218, n6356, n6369,
    n6379, n6381, n6385, n6397, n6427, n6456, n6485, n6502, n6513, n6556,
    n6590, n6596, n6611, n6631, n6659, n6691, n6729, n6773, n6775, n6785,
    n6790, n6794, n6814, n6861, n6971, n7026, n7057, n7099, n7139, n7149,
    n7305, n7330, n7335, n7339, n7377, n7421, n7428, n7437, n7460, n7524,
    n7566, n7569, n7593, n7657, n7670, n7674, n7678, n7692, n7693, n7721,
    n7731, n7751, n7759, n7769, n7773, n7788, n7841, n7876, n7917, n7949,
    n7963, n8006, n8052, n8067, n8194, n8244, n8255, n8256, n8259, n8285,
    n8305, n8309, n8324, n8363, n8381, n8399, n8405, n8439, n8526, n8581,
    n8614, n8638, n8656, n8678, n8687, n8694, n8721, n8745, n8782, n8806,
    n8827, n8856, n8869, n8920, n8943, n8964, n9003, n9090, n9172, n9246,
    n9251, n9259, n9318, n9323, n9372, n9380, n9396, n9399, n9445, n9460,
    n9493, n9507, n9512, n9554, n9557, n9598, n9646, n9655, n9832, n9872,
    n9926, n9934, n9942, n9967, n10017, n10018, n10053, n10057, n10096,
    n10117, n10125, n10158, n10201, n10250, n10275, n10372, n10405, n10411,
    n10514, n10577, n10593, n10611, n10614, n10650, n10710, n10712, n10739,
    n10763, n10792, n11011, n11044, n11056, n11121, n11184, n11192, n11201,
    n11220, n11223, n11266, n11273, n11302, n11356, n11424, n11455, n11473,
    n11479, n11481, n11486, n11503, n11566, n11579, n11580, n11615, n11630,
    n11667, n11736, n11749, n11775, n11841, n11898, n11926, n11980, n12113,
    n12121, n12152, n12153, n12161, n12209, n12315, n12341, n12380, n12384,
    n12398, n12446, n12495, n12507, n12546, n12562, n12587, n12593, n12626,
    n12650, n12657, n12702, n12811, n12821, n12861, n12871, n12875, n12892,
    n12900, n12917, n12956, n13026, n13044, n13074, n13110, n13137, n13190,
    n13263, n13319, n13333, n13367, n13419, n13424, n13453, n13460, n13490,
    n13494, n13549, n13668, n13677, n13708, n13714, n13719, n13775, n13781,
    n13783, n13851, n13912, n13914, n13951, n14071, n14090, n14130, n14148,
    n14230, n14275, n14323, n14345, n14440, n14510, n14570, n14575, n14576,
    n14603, n14633, n14680, n14684, n14692, n14702, n14704, n14790, n14826,
    n14899, n14954, n15053, n15077, n15146, n15167, n15182, n15241, n15258,
    n15271, n15289, n15332, n15378, n15424, n15490, n15506, n15508, n15539,
    n15546, n15602, n15636, n15652, n15743, n15761, n15766, n15780, n15884,
    n15918, n15936, n15967, n15979, n16029, n16158, n16167, n16217, n16223,
    n16247, n16376, n16396, n16439, n16476, n16482, n16502, n16507, n16521,
    n16524, n16544, n16608, n16722, n16743, n16812, n16818, n16824, n16911,
    n16968, n16971, n16988, n16994, n17035, n17037, n17069, n17077, n17090,
    n17095, n17250, n17251, n17302, n17351, n17458, n17664, n17784, n17911,
    n17954, n17959, n17968, n18035, n18105, n18145, n18151, n18157, n18171,
    n18227, n18274, n18290, n18295, n18345, n18409, n18444, n18452, n18483,
    n18496, n18537, n18558, n18578, n18584, n18649, n18690, n18737, n18745,
    n18880, n18901, n18907, n18926, n18962, n19005, n19033, n19042, n19081,
    n19107, n19116, n19144, n19163, n19196, n19228, n19234, n19270, n19282,
    n19327, n19357, n19361, n19454, n19472, n19477, n19494, n19514, n19515,
    n19531, n19539, n19575, n19584, n19608, n19618, n19652, n19680, n19701,
    n19770, n19789, n19803, n19905, n19911, n19922, n19941, n20013, n20036,
    n20040, n20077, n20138, n20151, n20169, n20179, n20213, n20235, n20250,
    n20259, n20349, n20359, n20385, n20409, n20411, n20429, n20455, n20470,
    n20478, n20489, n20604, n20658, n20700, n20794, n20826, n20923, n20929,
    n20946, n20986, n21078, n21095, n21134, n21138, n21222, n21226, n21276,
    n21287, n21317, n21398, n21471, n21489, n21538, n21599, n21649, n21654,
    n21674, n21687, n21735, n21749, n21753, n21779, n21784, n21832, n21839,
    n21898, n21905, n21915, n21934, n21957, n21981, n21993, n21997, n22043,
    n22068, n22072, n22173, n22198, n22201, n22253, n22270, n22274, n22290,
    n22309, n22332, n22335, n22358, n22359, n22379, n22433, n22442, n22470,
    n22492, n22554, n22588, n22591, n22597, n22619, n22626, n22631, n22660,
    n22764, n22793, n22843, n22871, n22879, n22918, n23035, n23039, n23065,
    n23068, n23120, n23146, n23160, n23166, n23200, n23250, n23272, n23304,
    n23333, n23369, n23430, n23463, n23493, n23513, n23529, n23541, n23586,
    n23657, n23697, n23717, n23755, n23775, n23831, n23842, n23849, n23895,
    n23912, n23913, n23923, n23974, n24004, n24032, n24048, n24085, n24093,
    n24129, n24150, n24170, n24196, n24278, n24319, n24323, n24327, n24374,
    n24485, n24618, n24620, n24638, n24732, n24768, n24786, n24879, n24937,
    n25023, n25068, n25073, n25074, n25094, n25119, n25120, n25126, n25168,
    n25240, n25296, n25316, n25331, n25336, n25345, n25365, n25370, n25381,
    n25435, n25464, n25471, n25475, n25494, n25523, n25565, n25586, n25629,
    n25643, n25694, n25738, n25749, n25751, n25797, n25872, n25877, n25923,
    n25926, n25972, n25974, n26036, n26053, n26054, n26107, n26167, n26180,
    n26191, n26224, n26264, n26318, n26408, n26443, n26452, n26483, n26510,
    n26512, n26553, n26565, n26572, n26625, n26660, n26725, n26744, n26748,
    n26752, n26797, n26808, n26823, n26882, n26913, n26979, n26986, n27037,
    n27089, n27104, n27120, n27134, n27188;
  output n7, n50, n55, n108, n142, n175, n235, n242, n243, n248, n266, n298,
    n317, n332, n357, n422, n431, n457, n463, n491, n496, n498, n521, n548,
    n554, n567, n588, n597, n637, n646, n696, n723, n735, n779, n809, n819,
    n829, n849, n858, n873, n879, n887, n904, n948, n957, n980, n982, n984,
    n1005, n1016, n1020, n1044, n1060, n1069, n1111, n1119, n1120, n1196,
    n1237, n1239, n1302, n1332, n1357, n1371, n1385, n1498, n1501, n1518,
    n1527, n1580, n1586, n1590, n1602, n1634, n1636, n1684, n1701, n1703,
    n1721, n1760, n1791, n1808, n1821, n1832, n1859, n1860, n1861, n1891,
    n1925, n1942, n1972, n1981, n2004, n2007, n2061, n2092, n2095, n2105,
    n2122, n2147, n2209, n2214, n2238, n2327, n2343, n2361, n2363, n2374,
    n2388, n2440, n2444, n2513, n2515, n2533, n2535, n2537, n2553, n2555,
    n2560, n2561, n2573, n2578, n2582, n2602, n2619, n2661, n2693, n2703,
    n2706, n2711, n2761, n2774, n2779, n2826, n2853, n2860, n2887, n2929,
    n2948, n2961, n2971, n3010, n3017, n3020, n3067, n3076, n3089, n3125,
    n3126, n3208, n3219, n3235, n3244, n3263, n3289, n3301, n3316, n3332,
    n3340, n3343, n3390, n3426, n3451, n3459, n3502, n3516, n3528, n3555,
    n3561, n3563, n3617, n3642, n3649, n3665, n3679, n3725, n3733, n3755,
    n3758, n3760, n3781, n3794, n3842, n3850, n3869, n3871, n3891, n3932,
    n3934, n3971, n3983, n4000, n4010, n4014, n4071, n4088, n4089, n4103,
    n4123, n4134, n4146, n4150, n4151, n4152, n4153, n4165, n4172, n4173,
    n4176, n4186, n4204, n4205, n4215, n4221, n4224, n4231, n4266, n4340,
    n4374, n4401, n4424, n4432, n4441, n4451, n4476, n4478, n4529, n4552,
    n4595, n4624, n4646, n4674, n4693, n4731, n4745, n4747, n4766, n4770,
    n4777, n4785, n4804, n4810, n4814, n4850, n4891, n4925, n4947, n4952,
    n4966, n4972, n5011, n5020, n5024, n5046, n5062, n5064, n5082, n5120,
    n5158, n5168, n5184, n5228, n5256, n5265, n5273, n5274, n5300, n5325,
    n5351, n5353, n5399, n5403, n5430, n5439, n5472, n5485, n5524, n5564,
    n5593, n5603, n5609, n5634, n5643, n5680, n5687, n5700, n5732, n5742,
    n5765, n5776, n5782, n5833, n5840, n5841, n5850, n5903, n5904, n5911,
    n5936, n5943, n5964, n5980, n6012, n6022, n6031, n6044, n6046, n6084,
    n6160, n6171, n6183, n6189, n6223, n6233, n6245, n6248, n6256, n6271,
    n6276, n6308, n6311, n6323, n6330, n6339, n6354, n6375, n6383, n6407,
    n6431, n6437, n6457, n6465, n6470, n6476, n6506, n6514, n6542, n6558,
    n6560, n6567, n6576, n6587, n6612, n6628, n6630, n6634, n6652, n6655,
    n6669, n6671, n6673, n6674, n6684, n6706, n6707, n6736, n6791, n6802,
    n6826, n6835, n6853, n6862, n6863, n6867, n6965, n6967, n6975, n6983,
    n6985, n6998, n7032, n7038, n7079, n7190, n7229, n7230, n7233, n7236,
    n7253, n7256, n7268, n7277, n7280, n7298, n7308, n7313, n7346, n7349,
    n7363, n7390, n7403, n7408, n7432, n7475, n7477, n7507, n7514, n7558,
    n7572, n7575, n7585, n7588, n7598, n7607, n7610, n7616, n7630, n7643,
    n7647, n7679, n7686, n7698, n7708, n7780, n7794, n7811, n7830, n7834,
    n7884, n7937, n7943, n7950, n7959, n7968, n7992, n7999, n8027, n8031,
    n8042, n8095, n8103, n8109, n8127, n8130, n8135, n8139, n8148, n8149,
    n8159, n8179, n8215, n8267, n8276, n8288, n8306, n8320, n8321, n8339,
    n8376, n8408, n8417, n8432, n8453, n8480, n8489, n8505, n8510, n8519,
    n8535, n8550, n8563, n8594, n8608, n8620, n8637, n8662, n8716, n8744,
    n8803, n8809, n8821, n8824, n8849, n8861, n8862, n8884, n8909, n8911,
    n8971, n8982, n8993, n9012, n9032, n9042, n9046, n9047, n9104, n9129,
    n9146, n9164, n9166, n9182, n9191, n9217, n9220, n9261, n9287, n9308,
    n9344, n9364, n9371, n9382, n9403, n9419, n9423, n9430, n9435, n9451,
    n9458, n9459, n9508, n9552, n9556, n9558, n9616, n9622, n9626, n9633,
    n9635, n9648, n9689, n9695, n9699, n9726, n9753, n9761, n9763, n9767,
    n9771, n9778, n9783, n9803, n9833, n9838, n9867, n9890, n9917, n9919,
    n9938, n9946, n9968, n10009, n10010, n10019, n10021, n10055, n10101,
    n10111, n10165, n10236, n10239, n10244, n10261, n10262, n10287, n10295,
    n10321, n10326, n10327, n10330, n10340, n10345, n10356, n10385, n10387,
    n10388, n10390, n10404, n10409, n10420, n10432, n10484, n10489, n10525,
    n10540, n10561, n10564, n10588, n10595, n10617, n10628, n10647, n10653,
    n10692, n10694, n10701, n10756, n10775, n10780, n10817, n10834, n10851,
    n10874, n10924, n10943, n10961, n11005, n11023, n11025, n11063, n11078,
    n11080, n11094, n11101, n11103, n11120, n11127, n11132, n11134, n11138,
    n11182, n11234, n11245, n11261, n11275, n11290, n11313, n11325, n11326,
    n11330, n11347, n11348, n11352, n11375, n11379, n11386, n11391, n11398,
    n11403, n11419, n11439, n11462, n11470, n11472, n11496, n11506, n11515,
    n11538, n11548, n11564, n11591, n11607, n11647, n11674, n11682, n11710,
    n11712, n11724, n11741, n11770, n11771, n11818, n11837, n11842, n11843,
    n11905, n11965, n12000, n12003, n12011, n12072, n12131, n12146, n12157,
    n12158, n12179, n12192, n12223, n12225, n12228, n12235, n12302, n12304,
    n12324, n12325, n12329, n12330, n12346, n12349, n12364, n12383, n12397,
    n12408, n12449, n12461, n12462, n12467, n12469, n12515, n12516, n12540,
    n12545, n12552, n12566, n12569, n12607, n12620, n12621, n12654, n12665,
    n12670, n12707, n12725, n12727, n12740, n12742, n12746, n12756, n12783,
    n12801, n12812, n12816, n12843, n12864, n12865, n12870, n12873, n12904,
    n12941, n12942, n12978, n12980, n12985, n12987, n12992, n13005, n13043,
    n13048, n13054, n13082, n13096, n13116, n13122, n13141, n13144, n13168,
    n13198, n13199, n13204, n13209, n13270, n13273, n13285, n13338, n13407,
    n13409, n13456, n13457, n13477, n13484, n13486, n13487, n13500, n13501,
    n13506, n13548, n13551, n13602, n13626, n13683, n13710, n13722, n13754,
    n13764, n13798, n13835, n13850, n13922, n13923, n14004, n14036, n14059,
    n14081, n14095, n14107, n14121, n14126, n14136, n14147, n14174, n14190,
    n14211, n14222, n14267, n14271, n14277, n14294, n14310, n14326, n14342,
    n14353, n14364, n14375, n14412, n14414, n14457, n14464, n14471, n14475,
    n14541, n14546, n14547, n14593, n14636, n14701, n14734, n14746, n14763,
    n14772, n14801, n14819, n14827, n14839, n14849, n14891, n14931, n14944,
    n14977, n14989, n15002, n15004, n15011, n15019, n15031, n15033, n15052,
    n15082, n15094, n15118, n15128, n15139, n15145, n15165, n15176, n15180,
    n15205, n15230, n15255, n15275, n15300, n15307, n15327, n15345, n15353,
    n15366, n15382, n15407, n15428, n15435, n15438, n15465, n15467, n15470,
    n15477, n15481, n15496, n15501, n15555, n15558, n15559, n15570, n15573,
    n15588, n15590, n15598, n15614, n15662, n15716, n15749, n15762, n15793,
    n15812, n15815, n15816, n15831, n15846, n15859, n15869, n15885, n15889,
    n15917, n15922, n15947, n15956, n15958, n15986, n16013, n16060, n16062,
    n16068, n16080, n16098, n16110, n16142, n16185, n16196, n16206, n16215,
    n16218, n16219, n16230, n16243, n16275, n16279, n16322, n16327, n16350,
    n16367, n16379, n16398, n16406, n16407, n16419, n16424, n16428, n16433,
    n16440, n16445, n16460, n16481, n16493, n16506, n16516, n16517, n16527,
    n16554, n16583, n16584, n16589, n16596, n16617, n16630, n16640, n16656,
    n16674, n16682, n16684, n16688, n16733, n16798, n16834, n16837, n16841,
    n16885, n16905, n16951, n16954, n16989, n17006, n17068, n17070, n17075,
    n17084, n17104, n17106, n17119, n17130, n17138, n17163, n17168, n17202,
    n17219, n17232, n17236, n17243, n17263, n17285, n17320, n17337, n17344,
    n17359, n17387, n17391, n17392, n17421, n17432, n17436, n17440, n17450,
    n17461, n17466, n17493, n17500, n17524, n17529, n17557, n17583, n17592,
    n17638, n17687, n17721, n17735, n17738, n17746, n17749, n17820, n17855,
    n17877, n17889, n17912, n17927, n17931, n17948, n17956, n17963, n17976,
    n17998, n18025, n18043, n18045, n18059, n18061, n18071, n18143, n18152,
    n18193, n18232, n18238, n18241, n18254, n18288, n18301, n18304, n18310,
    n18311, n18323, n18332, n18343, n18350, n18362, n18377, n18405, n18414,
    n18418, n18437, n18439, n18445, n18467, n18482, n18509, n18513, n18515,
    n18572, n18574, n18576, n18582, n18583, n18610, n18635, n18653, n18679,
    n18693, n18708, n18721, n18725, n18751, n18780, n18782, n18802, n18830,
    n18831, n18843, n18858, n18859, n18864, n18865, n18886, n18887, n18919,
    n18940, n18945, n18970, n18977, n18982, n18999, n19044, n19125, n19141,
    n19164, n19174, n19176, n19202, n19220, n19221, n19223, n19224, n19233,
    n19244, n19314, n19315, n19323, n19333, n19348, n19354, n19367, n19385,
    n19389, n19401, n19414, n19424, n19450, n19458, n19467, n19496, n19523,
    n19570, n19602, n19617, n19623, n19641, n19648, n19664, n19736, n19749,
    n19756, n19767, n19780, n19792, n19798, n19873, n19909, n19916, n19923,
    n19930, n19968, n19988, n20004, n20017, n20033, n20061, n20069, n20086,
    n20096, n20103, n20126, n20149, n20187, n20279, n20287, n20301, n20330,
    n20333, n20355, n20366, n20388, n20402, n20403, n20424, n20436, n20441,
    n20445, n20450, n20490, n20495, n20515, n20533, n20582, n20590, n20602,
    n20609, n20623, n20629, n20661, n20673, n20678, n20680, n20685, n20691,
    n20696, n20704, n20705, n20709, n20713, n20722, n20723, n20748, n20761,
    n20774, n20788, n20795, n20803, n20869, n20879, n20915, n20935, n20936,
    n21008, n21017, n21034, n21046, n21062, n21093, n21094, n21123, n21154,
    n21157, n21168, n21173, n21176, n21182, n21193, n21203, n21225, n21238,
    n21254, n21298, n21302, n21349, n21365, n21367, n21396, n21399, n21404,
    n21446, n21472, n21525, n21549, n21615, n21628, n21637, n21645, n21665,
    n21680, n21685, n21717, n21719, n21750, n21765, n21800, n21820, n21874,
    n21943, n21960, n21976, n21986, n22016, n22027, n22050, n22063, n22076,
    n22090, n22107, n22113, n22124, n22126, n22130, n22144, n22150, n22157,
    n22213, n22283, n22311, n22317, n22341, n22353, n22444, n22467, n22484,
    n22489, n22494, n22533, n22584, n22589, n22620, n22623, n22697, n22714,
    n22761, n22779, n22787, n22819, n22858, n22870, n22891, n22897, n22903,
    n22907, n22910, n22914, n22939, n22998, n23006, n23007, n23009, n23014,
    n23047, n23058, n23066, n23067, n23238, n23247, n23248, n23270, n23289,
    n23305, n23341, n23342, n23355, n23371, n23401, n23414, n23429, n23433,
    n23434, n23450, n23471, n23480, n23546, n23550, n23585, n23588, n23619,
    n23624, n23628, n23637, n23663, n23669, n23684, n23690, n23714, n23719,
    n23748, n23856, n23883, n23888, n23899, n23903, n23924, n23935, n23942,
    n23954, n23958, n23986, n24002, n24039, n24052, n24092, n24096, n24097,
    n24105, n24119, n24133, n24141, n24145, n24146, n24155, n24160, n24167,
    n24172, n24177, n24228, n24258, n24260, n24289, n24297, n24307, n24342,
    n24345, n24347, n24373, n24406, n24415, n24421, n24431, n24472, n24476,
    n24483, n24501, n24512, n24558, n24576, n24579, n24602, n24604, n24626,
    n24629, n24636, n24715, n24723, n24749, n24758, n24784, n24807, n24826,
    n24840, n24841, n24853, n24857, n24887, n24934, n24998, n25006, n25032,
    n25062, n25083, n25097, n25133, n25155, n25181, n25200, n25209, n25215,
    n25244, n25254, n25256, n25293, n25328, n25332, n25337, n25356, n25362,
    n25412, n25460, n25468, n25499, n25513, n25518, n25532, n25539, n25550,
    n25611, n25614, n25619, n25665, n25706, n25719, n25756, n25758, n25773,
    n25784, n25792, n25816, n25826, n25839, n25840, n25873, n25934, n25938,
    n25985, n25994, n26084, n26096, n26111, n26113, n26156, n26159, n26179,
    n26220, n26229, n26237, n26250, n26274, n26287, n26317, n26353, n26375,
    n26396, n26429, n26431, n26439, n26492, n26515, n26538, n26590, n26598,
    n26605, n26656, n26674, n26675, n26681, n26696, n26698, n26707, n26719,
    n26727, n26729, n26745, n26775, n26780, n26794, n26795, n26801, n26815,
    n26847, n26900, n26902, n26905, n26921, n26923, n26929, n26930, n26943,
    n26970, n27004, n27011, n27019, n27031, n27051, n27072, n27079, n27096,
    n27110, n27112, n27130, n27145, n27158, n27163, n27194;
  wire new_n2349, new_n2350, new_n2351, new_n2352, new_n2353, new_n2354,
    new_n2355_1, new_n2356, new_n2357, new_n2358, new_n2359, new_n2360,
    new_n2361_1, new_n2362, new_n2363_1, new_n2364, new_n2365, new_n2366,
    new_n2367, new_n2368, new_n2369, new_n2370, new_n2371, new_n2372,
    new_n2373, new_n2374_1, new_n2375, new_n2376, new_n2377, new_n2378,
    new_n2379, new_n2380, new_n2381, new_n2382, new_n2383, new_n2384,
    new_n2385, new_n2386, new_n2387_1, new_n2388_1, new_n2389, new_n2390,
    new_n2391, new_n2392, new_n2393, new_n2394, new_n2395, new_n2396,
    new_n2397, new_n2398, new_n2399, new_n2400, new_n2401, new_n2402,
    new_n2403, new_n2404, new_n2405, new_n2406, new_n2407, new_n2408,
    new_n2409_1, new_n2410, new_n2411, new_n2412, new_n2413, new_n2414,
    new_n2415, new_n2416_1, new_n2417, new_n2418, new_n2419, new_n2420_1,
    new_n2421_1, new_n2422, new_n2423, new_n2424, new_n2425, new_n2426,
    new_n2427, new_n2428, new_n2429, new_n2430, new_n2431, new_n2432,
    new_n2433, new_n2434, new_n2435, new_n2436, new_n2437, new_n2438,
    new_n2439, new_n2440_1, new_n2441, new_n2442, new_n2443, new_n2444_1,
    new_n2445, new_n2446, new_n2447, new_n2448, new_n2449, new_n2450,
    new_n2451, new_n2452, new_n2453, new_n2454, new_n2455, new_n2456,
    new_n2457, new_n2458, new_n2459, new_n2460, new_n2461, new_n2462,
    new_n2463, new_n2464, new_n2465, new_n2466, new_n2467, new_n2468,
    new_n2469, new_n2470, new_n2471, new_n2472, new_n2473, new_n2474,
    new_n2475, new_n2476, new_n2477, new_n2478, new_n2479_1, new_n2480,
    new_n2481, new_n2482, new_n2483, new_n2484, new_n2485, new_n2486,
    new_n2487, new_n2488, new_n2489, new_n2490, new_n2491, new_n2492,
    new_n2493, new_n2494, new_n2495, new_n2496, new_n2497, new_n2498,
    new_n2499, new_n2500, new_n2501, new_n2502, new_n2503, new_n2504,
    new_n2505, new_n2506, new_n2507, new_n2508, new_n2509, new_n2510,
    new_n2511, new_n2512, new_n2513_1, new_n2514, new_n2515_1, new_n2516,
    new_n2517, new_n2518, new_n2519, new_n2520, new_n2521, new_n2522,
    new_n2523, new_n2524, new_n2525, new_n2526, new_n2527, new_n2528,
    new_n2529, new_n2530, new_n2531, new_n2532, new_n2533_1, new_n2534,
    new_n2535_1, new_n2536, new_n2537_1, new_n2538, new_n2539, new_n2540,
    new_n2542, new_n2543, new_n2544, new_n2545, new_n2546, new_n2548,
    new_n2549, new_n2550, new_n2551, new_n2552, new_n2554, new_n2555_1,
    new_n2556, new_n2557, new_n2558, new_n2559, new_n2560_1, new_n2561_1,
    new_n2562, new_n2563, new_n2564, new_n2565, new_n2566, new_n2567,
    new_n2568, new_n2569, new_n2570_1, new_n2571, new_n2572, new_n2573_1,
    new_n2574, new_n2575, new_n2576, new_n2577, new_n2578_1, new_n2579,
    new_n2580, new_n2581, new_n2582_1, new_n2583, new_n2584, new_n2585,
    new_n2586, new_n2587, new_n2588, new_n2589, new_n2590, new_n2591,
    new_n2592, new_n2593, new_n2594, new_n2595, new_n2596, new_n2597,
    new_n2598, new_n2599, new_n2600, new_n2601, new_n2602_1, new_n2603,
    new_n2604, new_n2605, new_n2606, new_n2607, new_n2608, new_n2609,
    new_n2610, new_n2611, new_n2612, new_n2613, new_n2614, new_n2615,
    new_n2616, new_n2617, new_n2618, new_n2619_1, new_n2620, new_n2621,
    new_n2622, new_n2623, new_n2624, new_n2625, new_n2626, new_n2627,
    new_n2628, new_n2629, new_n2630, new_n2631, new_n2632, new_n2633,
    new_n2634, new_n2635, new_n2636, new_n2637, new_n2638, new_n2639,
    new_n2640, new_n2641, new_n2642, new_n2643, new_n2644, new_n2645,
    new_n2646_1, new_n2647, new_n2648, new_n2649, new_n2650, new_n2651,
    new_n2652, new_n2653, new_n2654, new_n2655, new_n2656, new_n2657,
    new_n2658, new_n2659_1, new_n2660, new_n2661_1, new_n2662, new_n2663,
    new_n2664, new_n2665, new_n2666, new_n2667, new_n2668, new_n2669,
    new_n2670, new_n2671, new_n2672, new_n2673, new_n2674, new_n2675,
    new_n2676, new_n2677, new_n2678, new_n2679, new_n2680_1, new_n2681,
    new_n2682, new_n2683, new_n2684, new_n2685, new_n2686, new_n2687,
    new_n2688, new_n2689, new_n2690, new_n2691, new_n2692, new_n2693_1,
    new_n2694, new_n2695, new_n2696, new_n2697, new_n2698, new_n2699,
    new_n2700, new_n2701, new_n2702, new_n2703_1, new_n2704, new_n2705,
    new_n2706_1, new_n2707, new_n2708, new_n2709, new_n2710, new_n2711_1,
    new_n2712, new_n2713, new_n2714, new_n2715, new_n2716, new_n2717,
    new_n2718, new_n2719, new_n2720, new_n2721, new_n2722, new_n2723,
    new_n2724, new_n2725, new_n2726, new_n2727, new_n2728, new_n2729,
    new_n2730, new_n2731_1, new_n2732, new_n2733, new_n2734, new_n2735,
    new_n2736, new_n2737, new_n2738, new_n2739, new_n2740, new_n2741,
    new_n2742, new_n2743_1, new_n2744, new_n2745, new_n2746, new_n2747,
    new_n2748, new_n2749, new_n2750, new_n2751, new_n2752, new_n2753,
    new_n2754, new_n2755, new_n2756, new_n2757, new_n2758, new_n2759,
    new_n2760, new_n2761_1, new_n2762, new_n2763, new_n2764, new_n2765,
    new_n2766, new_n2767, new_n2768, new_n2769, new_n2770, new_n2771,
    new_n2772, new_n2773, new_n2774_1, new_n2775, new_n2776, new_n2777,
    new_n2778, new_n2779_1, new_n2780, new_n2781, new_n2782, new_n2783_1,
    new_n2784, new_n2785, new_n2786, new_n2787, new_n2788, new_n2789,
    new_n2790, new_n2791, new_n2792, new_n2793, new_n2794, new_n2795,
    new_n2796, new_n2797, new_n2798, new_n2799, new_n2800, new_n2801,
    new_n2802, new_n2803, new_n2804, new_n2805, new_n2806, new_n2807,
    new_n2808, new_n2809_1, new_n2810, new_n2811, new_n2812, new_n2813,
    new_n2814, new_n2815, new_n2816_1, new_n2817, new_n2818, new_n2819,
    new_n2820, new_n2821, new_n2822, new_n2823, new_n2824, new_n2825,
    new_n2826_1, new_n2827, new_n2828, new_n2829, new_n2830, new_n2831,
    new_n2832, new_n2833, new_n2834, new_n2835, new_n2836, new_n2837,
    new_n2838, new_n2839, new_n2840, new_n2841, new_n2842, new_n2843,
    new_n2844, new_n2845, new_n2846, new_n2847, new_n2849, new_n2850,
    new_n2851, new_n2852, new_n2853_1, new_n2854, new_n2855, new_n2856,
    new_n2857, new_n2858_1, new_n2859, new_n2860_1, new_n2861, new_n2862,
    new_n2863, new_n2864, new_n2865, new_n2866, new_n2867, new_n2868,
    new_n2869, new_n2870, new_n2871, new_n2872, new_n2873, new_n2874,
    new_n2875, new_n2876, new_n2877, new_n2878, new_n2879, new_n2880,
    new_n2881, new_n2882, new_n2883, new_n2884, new_n2885, new_n2886_1,
    new_n2887_1, new_n2888, new_n2889, new_n2890, new_n2891, new_n2892,
    new_n2893, new_n2894, new_n2895, new_n2896, new_n2897, new_n2898,
    new_n2899, new_n2900, new_n2901, new_n2902, new_n2903, new_n2904,
    new_n2905, new_n2906, new_n2907, new_n2908, new_n2909, new_n2910,
    new_n2911, new_n2912, new_n2913, new_n2914, new_n2915, new_n2916,
    new_n2917, new_n2918, new_n2919, new_n2920, new_n2921, new_n2922,
    new_n2923, new_n2924, new_n2925, new_n2926, new_n2927, new_n2928,
    new_n2929_1, new_n2930, new_n2931, new_n2932, new_n2933, new_n2934,
    new_n2935, new_n2936, new_n2937, new_n2938, new_n2939, new_n2940,
    new_n2941, new_n2942, new_n2943, new_n2944_1, new_n2945, new_n2946,
    new_n2947, new_n2948_1, new_n2949, new_n2950, new_n2951, new_n2952,
    new_n2953, new_n2954, new_n2955, new_n2956, new_n2957, new_n2958,
    new_n2959, new_n2960, new_n2961_1, new_n2962, new_n2963, new_n2964,
    new_n2965, new_n2966, new_n2967, new_n2968, new_n2969, new_n2970,
    new_n2971_1, new_n2972, new_n2973, new_n2974, new_n2975, new_n2976,
    new_n2977, new_n2978_1, new_n2979_1, new_n2980, new_n2981, new_n2982,
    new_n2983, new_n2984, new_n2985_1, new_n2986, new_n2987, new_n2988,
    new_n2989, new_n2990, new_n2991, new_n2992, new_n2993, new_n2994,
    new_n2995, new_n2996, new_n2997, new_n2998, new_n2999_1, new_n3000,
    new_n3001, new_n3002, new_n3003, new_n3004, new_n3005, new_n3006,
    new_n3007, new_n3008, new_n3009, new_n3010_1, new_n3011, new_n3012,
    new_n3013, new_n3014, new_n3015, new_n3016, new_n3017_1, new_n3018_1,
    new_n3019, new_n3020_1, new_n3021, new_n3022, new_n3023, new_n3024,
    new_n3025, new_n3026, new_n3027, new_n3028, new_n3029, new_n3030_1,
    new_n3031, new_n3032, new_n3033, new_n3034, new_n3035, new_n3036,
    new_n3037, new_n3038, new_n3039, new_n3040, new_n3041, new_n3042,
    new_n3043, new_n3044, new_n3045, new_n3046, new_n3047, new_n3048,
    new_n3049, new_n3050, new_n3051, new_n3052, new_n3053, new_n3054,
    new_n3055, new_n3056, new_n3057, new_n3058, new_n3059, new_n3060,
    new_n3061, new_n3062, new_n3063, new_n3064, new_n3065, new_n3066,
    new_n3067_1, new_n3068, new_n3069, new_n3070, new_n3071, new_n3072,
    new_n3073, new_n3074, new_n3075, new_n3076_1, new_n3077, new_n3078,
    new_n3079, new_n3080, new_n3081, new_n3082, new_n3083, new_n3084,
    new_n3086, new_n3087, new_n3088, new_n3089_1, new_n3090, new_n3091,
    new_n3092, new_n3093, new_n3094, new_n3095, new_n3096, new_n3097,
    new_n3098, new_n3099, new_n3100, new_n3101, new_n3102, new_n3103,
    new_n3104, new_n3105, new_n3106, new_n3107, new_n3108, new_n3109,
    new_n3110, new_n3111, new_n3112, new_n3113, new_n3114, new_n3115,
    new_n3116, new_n3117, new_n3118, new_n3119, new_n3120, new_n3121,
    new_n3122, new_n3123, new_n3124, new_n3125_1, new_n3126_1, new_n3127,
    new_n3128, new_n3129, new_n3130, new_n3131, new_n3132, new_n3133,
    new_n3134, new_n3135, new_n3136_1, new_n3137, new_n3138, new_n3139,
    new_n3140, new_n3141, new_n3142, new_n3143, new_n3144, new_n3145,
    new_n3146, new_n3147, new_n3148, new_n3149, new_n3150, new_n3151,
    new_n3152, new_n3153, new_n3154, new_n3155, new_n3156, new_n3157,
    new_n3158, new_n3159, new_n3160, new_n3161_1, new_n3162, new_n3163,
    new_n3164_1, new_n3165, new_n3166, new_n3167, new_n3168, new_n3169,
    new_n3170, new_n3171, new_n3172, new_n3173, new_n3174, new_n3175,
    new_n3176, new_n3177, new_n3178, new_n3179, new_n3180, new_n3181,
    new_n3182, new_n3183, new_n3184, new_n3185, new_n3186, new_n3187,
    new_n3188, new_n3189, new_n3190, new_n3191, new_n3192, new_n3193,
    new_n3194, new_n3195, new_n3196, new_n3197, new_n3198, new_n3199,
    new_n3200, new_n3201, new_n3202, new_n3203, new_n3204, new_n3205,
    new_n3206, new_n3207, new_n3208_1, new_n3209, new_n3210, new_n3211,
    new_n3212, new_n3213, new_n3214, new_n3215, new_n3216, new_n3217,
    new_n3218, new_n3219_1, new_n3220, new_n3221, new_n3222, new_n3223,
    new_n3224, new_n3225, new_n3226, new_n3227, new_n3228_1, new_n3229,
    new_n3230, new_n3231, new_n3232, new_n3233, new_n3234, new_n3235_1,
    new_n3236, new_n3237, new_n3238, new_n3239, new_n3240, new_n3241,
    new_n3242, new_n3243, new_n3244_1, new_n3245, new_n3246, new_n3247,
    new_n3248, new_n3249, new_n3250, new_n3251, new_n3252, new_n3253_1,
    new_n3254, new_n3255, new_n3256, new_n3257, new_n3258, new_n3259,
    new_n3260_1, new_n3261, new_n3262, new_n3263_1, new_n3264, new_n3265,
    new_n3266, new_n3267, new_n3268, new_n3269, new_n3270, new_n3271,
    new_n3272, new_n3273, new_n3274, new_n3275, new_n3276, new_n3277,
    new_n3278, new_n3279_1, new_n3280, new_n3281, new_n3282, new_n3283,
    new_n3284, new_n3285, new_n3286, new_n3287, new_n3288, new_n3289_1,
    new_n3290, new_n3291, new_n3292, new_n3293, new_n3294, new_n3295,
    new_n3296, new_n3297, new_n3298, new_n3299, new_n3300, new_n3301_1,
    new_n3302, new_n3303, new_n3304, new_n3305, new_n3306_1, new_n3307,
    new_n3308, new_n3309, new_n3310, new_n3311, new_n3312, new_n3313,
    new_n3314, new_n3315, new_n3316_1, new_n3317, new_n3318, new_n3319,
    new_n3320_1, new_n3321, new_n3322, new_n3323, new_n3324_1, new_n3325,
    new_n3326, new_n3327, new_n3328, new_n3329, new_n3330, new_n3331,
    new_n3332_1, new_n3333, new_n3334, new_n3335, new_n3336, new_n3337,
    new_n3338, new_n3339, new_n3340_1, new_n3341, new_n3342, new_n3343_1,
    new_n3344, new_n3345, new_n3346, new_n3347, new_n3348, new_n3349_1,
    new_n3350, new_n3351, new_n3352, new_n3353, new_n3354, new_n3355,
    new_n3356, new_n3357, new_n3358, new_n3359, new_n3360, new_n3361,
    new_n3362, new_n3363, new_n3364, new_n3365, new_n3366_1, new_n3367,
    new_n3368, new_n3369, new_n3370, new_n3371, new_n3372, new_n3373,
    new_n3374, new_n3375, new_n3376, new_n3377, new_n3378, new_n3379,
    new_n3380, new_n3381, new_n3382, new_n3383, new_n3384, new_n3385,
    new_n3386, new_n3387, new_n3388, new_n3389, new_n3390_1, new_n3391,
    new_n3392, new_n3393, new_n3394, new_n3395, new_n3396, new_n3397,
    new_n3398, new_n3399, new_n3400, new_n3401, new_n3402, new_n3403,
    new_n3405, new_n3406, new_n3407, new_n3408, new_n3409, new_n3410,
    new_n3411, new_n3412, new_n3413, new_n3414, new_n3415, new_n3416,
    new_n3417, new_n3418, new_n3419, new_n3420, new_n3421, new_n3422,
    new_n3423, new_n3424, new_n3425_1, new_n3426_1, new_n3427, new_n3428,
    new_n3429, new_n3430, new_n3431, new_n3432, new_n3433, new_n3434,
    new_n3435, new_n3436, new_n3437, new_n3438, new_n3439, new_n3440,
    new_n3441, new_n3442, new_n3443, new_n3444, new_n3445, new_n3446,
    new_n3447, new_n3448, new_n3449, new_n3450, new_n3451_1, new_n3452,
    new_n3453, new_n3454, new_n3455, new_n3456, new_n3457, new_n3458,
    new_n3459_1, new_n3460_1, new_n3461, new_n3462, new_n3463, new_n3464,
    new_n3465, new_n3466, new_n3467, new_n3468_1, new_n3469, new_n3470,
    new_n3471, new_n3472, new_n3473, new_n3474, new_n3475, new_n3476,
    new_n3477, new_n3478, new_n3479, new_n3480_1, new_n3481, new_n3482,
    new_n3483, new_n3484, new_n3485, new_n3486, new_n3487, new_n3488,
    new_n3489, new_n3490, new_n3491, new_n3492, new_n3493, new_n3494,
    new_n3495, new_n3496, new_n3497, new_n3498, new_n3499, new_n3500,
    new_n3501, new_n3502_1, new_n3503, new_n3504, new_n3505, new_n3506_1,
    new_n3507, new_n3508, new_n3509, new_n3510, new_n3511, new_n3512,
    new_n3513, new_n3514, new_n3515, new_n3516_1, new_n3517, new_n3518,
    new_n3519, new_n3520, new_n3521, new_n3522, new_n3523, new_n3524,
    new_n3525, new_n3526, new_n3527, new_n3528_1, new_n3529, new_n3530,
    new_n3531, new_n3532, new_n3533, new_n3534, new_n3535, new_n3536,
    new_n3537, new_n3538, new_n3539, new_n3540, new_n3541_1, new_n3542,
    new_n3543, new_n3544, new_n3545, new_n3546, new_n3547, new_n3548,
    new_n3549, new_n3550, new_n3551, new_n3552, new_n3553, new_n3554,
    new_n3555_1, new_n3556, new_n3557, new_n3558, new_n3559, new_n3560,
    new_n3561_1, new_n3562, new_n3563_1, new_n3564, new_n3565, new_n3566,
    new_n3567, new_n3568, new_n3569, new_n3570_1, new_n3571, new_n3572,
    new_n3573, new_n3574, new_n3575, new_n3576, new_n3577, new_n3578,
    new_n3579, new_n3580, new_n3581, new_n3582_1, new_n3583, new_n3584,
    new_n3585, new_n3586, new_n3587, new_n3588, new_n3589, new_n3590,
    new_n3591, new_n3592, new_n3593, new_n3594, new_n3595, new_n3596,
    new_n3597, new_n3598, new_n3599, new_n3600, new_n3601, new_n3602,
    new_n3603, new_n3604, new_n3605, new_n3606, new_n3607, new_n3608,
    new_n3609, new_n3610, new_n3611, new_n3612, new_n3613, new_n3614,
    new_n3615, new_n3616, new_n3617_1, new_n3618_1, new_n3619, new_n3620,
    new_n3621, new_n3622, new_n3623, new_n3624, new_n3625, new_n3626,
    new_n3627, new_n3628, new_n3629, new_n3630, new_n3631, new_n3632,
    new_n3633, new_n3634, new_n3635, new_n3636, new_n3637, new_n3638,
    new_n3639, new_n3640, new_n3641, new_n3642_1, new_n3643, new_n3644,
    new_n3645, new_n3646, new_n3647, new_n3648, new_n3649_1, new_n3650,
    new_n3651, new_n3652, new_n3653, new_n3654, new_n3655, new_n3656,
    new_n3657, new_n3658, new_n3659, new_n3660, new_n3661, new_n3662,
    new_n3663, new_n3664, new_n3665_1, new_n3666, new_n3667, new_n3668,
    new_n3669, new_n3670, new_n3671, new_n3672, new_n3673, new_n3674,
    new_n3675, new_n3676, new_n3677, new_n3678, new_n3679_1, new_n3680,
    new_n3681, new_n3682, new_n3683, new_n3684, new_n3685, new_n3686,
    new_n3687, new_n3688, new_n3689, new_n3690, new_n3691, new_n3692,
    new_n3693, new_n3694, new_n3695, new_n3696, new_n3697, new_n3698,
    new_n3699, new_n3700, new_n3701, new_n3702, new_n3703, new_n3704,
    new_n3705, new_n3706, new_n3707, new_n3708, new_n3709, new_n3710_1,
    new_n3711, new_n3712, new_n3713, new_n3714, new_n3715, new_n3716,
    new_n3717, new_n3718, new_n3719, new_n3720, new_n3721, new_n3722,
    new_n3723, new_n3725_1, new_n3726, new_n3727, new_n3728, new_n3729,
    new_n3730, new_n3731, new_n3732, new_n3733_1, new_n3734, new_n3735,
    new_n3736, new_n3737, new_n3738, new_n3739, new_n3740_1, new_n3741,
    new_n3742, new_n3743, new_n3744, new_n3745, new_n3746, new_n3747,
    new_n3748, new_n3749, new_n3750, new_n3751, new_n3752, new_n3753,
    new_n3754, new_n3755_1, new_n3756, new_n3757, new_n3758_1, new_n3759,
    new_n3760_1, new_n3761, new_n3762, new_n3763, new_n3764, new_n3765,
    new_n3766, new_n3767, new_n3768, new_n3769, new_n3770, new_n3771,
    new_n3772, new_n3773, new_n3774, new_n3775, new_n3776, new_n3777,
    new_n3778, new_n3779, new_n3780, new_n3781_1, new_n3782, new_n3783,
    new_n3784, new_n3785_1, new_n3786, new_n3787, new_n3788, new_n3789,
    new_n3790, new_n3791, new_n3792, new_n3793, new_n3794_1, new_n3795_1,
    new_n3796, new_n3797, new_n3798, new_n3799, new_n3800, new_n3801,
    new_n3802, new_n3803, new_n3804, new_n3805, new_n3806, new_n3807,
    new_n3808, new_n3809, new_n3810, new_n3811, new_n3812, new_n3813,
    new_n3814, new_n3815, new_n3816, new_n3817, new_n3818, new_n3819,
    new_n3820, new_n3821, new_n3822, new_n3823, new_n3824, new_n3825,
    new_n3826, new_n3827, new_n3828_1, new_n3829, new_n3830, new_n3831,
    new_n3832, new_n3833, new_n3834, new_n3835, new_n3836, new_n3837,
    new_n3838, new_n3839, new_n3840, new_n3841, new_n3842_1, new_n3843,
    new_n3844, new_n3845, new_n3846, new_n3847, new_n3848, new_n3849,
    new_n3850_1, new_n3851, new_n3852, new_n3853, new_n3854, new_n3855,
    new_n3856, new_n3857, new_n3858, new_n3859, new_n3860, new_n3861,
    new_n3862, new_n3863, new_n3864, new_n3865, new_n3866, new_n3867,
    new_n3868, new_n3869_1, new_n3870, new_n3871_1, new_n3872, new_n3873,
    new_n3874, new_n3875, new_n3876, new_n3877, new_n3878, new_n3879,
    new_n3880, new_n3881, new_n3882, new_n3883, new_n3884, new_n3885,
    new_n3886, new_n3887, new_n3888, new_n3889, new_n3890, new_n3891_1,
    new_n3892, new_n3893, new_n3894, new_n3895, new_n3896, new_n3897,
    new_n3898, new_n3899, new_n3900, new_n3901, new_n3902, new_n3903,
    new_n3904, new_n3905, new_n3906, new_n3907, new_n3908, new_n3909_1,
    new_n3910, new_n3911, new_n3912, new_n3913, new_n3914, new_n3915,
    new_n3916, new_n3917, new_n3918_1, new_n3919, new_n3920, new_n3921,
    new_n3922, new_n3923, new_n3924, new_n3925_1, new_n3926, new_n3928,
    new_n3929, new_n3930, new_n3931, new_n3932_1, new_n3933, new_n3934_1,
    new_n3935, new_n3936, new_n3937, new_n3938, new_n3939, new_n3940,
    new_n3941, new_n3942, new_n3943, new_n3944, new_n3945_1, new_n3946,
    new_n3947, new_n3948, new_n3949, new_n3950, new_n3951, new_n3952_1,
    new_n3953, new_n3954, new_n3955, new_n3956, new_n3957, new_n3958,
    new_n3959_1, new_n3960, new_n3961, new_n3962_1, new_n3963, new_n3964,
    new_n3965, new_n3966, new_n3967, new_n3968, new_n3969, new_n3970,
    new_n3971_1, new_n3972, new_n3973, new_n3974, new_n3975, new_n3976,
    new_n3977, new_n3978, new_n3979, new_n3980, new_n3981, new_n3982,
    new_n3983_1, new_n3984_1, new_n3985, new_n3986, new_n3987, new_n3988,
    new_n3989, new_n3990, new_n3991, new_n3992, new_n3993, new_n3994,
    new_n3995, new_n3996, new_n3997, new_n3998, new_n3999, new_n4000_1,
    new_n4001, new_n4002, new_n4003, new_n4004, new_n4005, new_n4006,
    new_n4007, new_n4008, new_n4009, new_n4010_1, new_n4011, new_n4012,
    new_n4013, new_n4014_1, new_n4015, new_n4016, new_n4017, new_n4018,
    new_n4019, new_n4020, new_n4021, new_n4022, new_n4023, new_n4024,
    new_n4025, new_n4026, new_n4027, new_n4028, new_n4029, new_n4030,
    new_n4031, new_n4032, new_n4033, new_n4034, new_n4035, new_n4036,
    new_n4037, new_n4038, new_n4039, new_n4040, new_n4041, new_n4042,
    new_n4043, new_n4044, new_n4045, new_n4046, new_n4047, new_n4048,
    new_n4049, new_n4050, new_n4051, new_n4052, new_n4053, new_n4054,
    new_n4055, new_n4056, new_n4057, new_n4058, new_n4059, new_n4060,
    new_n4061, new_n4062, new_n4063, new_n4064, new_n4065, new_n4066,
    new_n4067, new_n4068, new_n4069, new_n4070, new_n4071_1, new_n4072,
    new_n4073, new_n4074, new_n4075, new_n4076, new_n4077, new_n4078,
    new_n4079, new_n4080, new_n4081, new_n4082, new_n4083, new_n4084,
    new_n4085_1, new_n4086, new_n4087, new_n4088_1, new_n4089_1, new_n4090,
    new_n4091, new_n4092, new_n4093, new_n4094, new_n4095, new_n4096,
    new_n4097, new_n4098, new_n4099, new_n4100_1, new_n4101, new_n4102,
    new_n4103_1, new_n4104, new_n4106, new_n4107, new_n4108, new_n4109,
    new_n4110, new_n4111, new_n4112, new_n4113, new_n4114, new_n4115,
    new_n4116, new_n4117, new_n4118, new_n4119_1, new_n4120, new_n4121,
    new_n4122, new_n4123_1, new_n4124, new_n4125, new_n4126, new_n4127,
    new_n4128, new_n4129, new_n4130, new_n4131, new_n4132, new_n4133,
    new_n4134_1, new_n4135, new_n4136, new_n4137, new_n4138, new_n4139,
    new_n4140, new_n4141, new_n4142, new_n4143, new_n4144, new_n4145,
    new_n4146_1, new_n4147, new_n4148, new_n4149, new_n4150_1, new_n4151_1,
    new_n4152_1, new_n4153_1, new_n4154, new_n4155, new_n4156, new_n4157,
    new_n4158, new_n4159, new_n4160, new_n4161, new_n4162, new_n4163,
    new_n4165_1, new_n4166, new_n4167, new_n4168, new_n4169, new_n4170,
    new_n4171, new_n4172_1, new_n4173_1, new_n4174, new_n4175, new_n4176_1,
    new_n4177, new_n4178, new_n4179, new_n4180, new_n4181, new_n4182,
    new_n4183, new_n4184, new_n4185, new_n4186_1, new_n4187, new_n4188,
    new_n4189, new_n4190, new_n4191, new_n4192, new_n4193, new_n4194,
    new_n4195, new_n4196, new_n4197, new_n4198, new_n4199, new_n4200,
    new_n4201, new_n4202, new_n4203, new_n4204_1, new_n4205_1, new_n4206,
    new_n4207, new_n4208, new_n4209, new_n4210, new_n4211, new_n4212,
    new_n4213, new_n4214, new_n4215_1, new_n4216, new_n4217, new_n4218,
    new_n4219, new_n4220, new_n4221_1, new_n4222, new_n4223, new_n4224_1,
    new_n4225, new_n4226, new_n4227, new_n4228, new_n4229, new_n4230,
    new_n4231_1, new_n4232, new_n4233, new_n4234, new_n4235, new_n4236,
    new_n4237, new_n4238, new_n4239, new_n4240, new_n4241, new_n4242,
    new_n4243, new_n4244, new_n4245, new_n4246, new_n4247, new_n4248,
    new_n4249, new_n4250, new_n4251, new_n4252, new_n4253, new_n4254,
    new_n4255, new_n4256_1, new_n4257, new_n4258, new_n4259, new_n4260,
    new_n4261, new_n4262, new_n4263, new_n4264, new_n4265, new_n4266_1,
    new_n4267, new_n4268, new_n4269, new_n4270, new_n4271, new_n4272_1,
    new_n4273, new_n4274, new_n4275, new_n4276, new_n4277, new_n4278,
    new_n4279, new_n4280, new_n4281, new_n4282, new_n4283, new_n4284,
    new_n4285, new_n4286, new_n4287, new_n4288, new_n4289, new_n4290,
    new_n4291, new_n4292, new_n4293, new_n4294, new_n4295, new_n4296,
    new_n4297, new_n4298, new_n4299, new_n4300, new_n4301, new_n4302,
    new_n4303, new_n4304, new_n4305, new_n4306_1, new_n4307, new_n4308,
    new_n4309, new_n4310, new_n4312, new_n4313, new_n4314, new_n4315,
    new_n4316, new_n4317, new_n4318, new_n4319_1, new_n4320, new_n4321,
    new_n4322, new_n4323, new_n4324, new_n4325_1, new_n4326_1, new_n4327,
    new_n4328, new_n4329, new_n4330, new_n4331, new_n4332, new_n4333,
    new_n4334, new_n4335, new_n4336, new_n4337, new_n4338, new_n4339,
    new_n4340_1, new_n4341, new_n4342, new_n4343, new_n4344, new_n4345,
    new_n4346, new_n4347, new_n4348, new_n4349, new_n4350, new_n4351,
    new_n4352, new_n4353, new_n4354, new_n4355, new_n4356, new_n4357,
    new_n4358, new_n4359, new_n4360, new_n4361, new_n4362, new_n4363,
    new_n4364, new_n4365, new_n4366, new_n4367, new_n4368, new_n4369,
    new_n4370, new_n4371, new_n4372, new_n4373, new_n4374_1, new_n4375,
    new_n4376_1, new_n4377, new_n4378, new_n4379, new_n4380, new_n4381,
    new_n4382, new_n4383, new_n4384, new_n4385, new_n4386, new_n4387,
    new_n4388, new_n4389, new_n4390, new_n4391, new_n4392, new_n4393,
    new_n4394, new_n4395, new_n4396, new_n4397, new_n4398, new_n4399,
    new_n4400, new_n4401_1, new_n4402, new_n4403, new_n4404, new_n4405,
    new_n4406, new_n4407, new_n4408, new_n4409_1, new_n4410, new_n4411,
    new_n4412, new_n4413, new_n4414, new_n4415, new_n4416, new_n4417,
    new_n4418, new_n4419, new_n4420, new_n4421, new_n4422, new_n4423,
    new_n4424_1, new_n4425, new_n4426_1, new_n4427, new_n4428, new_n4429,
    new_n4430, new_n4431, new_n4432_1, new_n4433, new_n4434, new_n4435,
    new_n4436, new_n4437, new_n4438, new_n4439, new_n4440, new_n4441_1,
    new_n4442, new_n4443, new_n4444, new_n4445, new_n4446, new_n4447,
    new_n4448, new_n4449, new_n4450, new_n4451_1, new_n4452, new_n4453,
    new_n4454, new_n4455, new_n4456, new_n4457, new_n4458, new_n4459,
    new_n4460, new_n4461, new_n4462, new_n4463, new_n4464, new_n4465,
    new_n4466, new_n4467, new_n4468, new_n4469, new_n4470, new_n4471,
    new_n4472, new_n4473, new_n4474, new_n4475, new_n4476_1, new_n4477,
    new_n4478_1, new_n4479, new_n4480, new_n4481, new_n4482, new_n4483,
    new_n4484, new_n4485, new_n4486, new_n4487, new_n4488, new_n4489,
    new_n4490, new_n4491, new_n4492, new_n4493, new_n4494, new_n4495,
    new_n4496, new_n4497, new_n4498, new_n4499, new_n4500, new_n4501,
    new_n4502, new_n4503, new_n4504, new_n4505, new_n4506, new_n4507,
    new_n4508, new_n4509, new_n4510, new_n4511, new_n4512, new_n4513,
    new_n4514_1, new_n4515, new_n4516, new_n4517, new_n4518, new_n4519,
    new_n4520, new_n4521, new_n4522, new_n4523, new_n4524, new_n4525,
    new_n4526, new_n4527, new_n4528, new_n4529_1, new_n4530, new_n4531,
    new_n4532, new_n4533, new_n4534, new_n4535, new_n4536, new_n4537,
    new_n4538, new_n4539, new_n4540, new_n4541, new_n4542, new_n4543,
    new_n4544, new_n4545, new_n4546, new_n4547, new_n4548, new_n4549,
    new_n4550, new_n4551, new_n4552_1, new_n4553, new_n4554, new_n4555,
    new_n4556, new_n4557, new_n4558, new_n4559, new_n4560, new_n4561,
    new_n4562, new_n4563, new_n4564, new_n4565, new_n4566, new_n4567,
    new_n4568, new_n4569, new_n4570, new_n4571, new_n4572, new_n4573,
    new_n4574, new_n4575, new_n4576, new_n4577, new_n4578, new_n4579,
    new_n4580, new_n4581, new_n4582, new_n4583, new_n4584, new_n4585,
    new_n4586, new_n4587, new_n4588_1, new_n4589, new_n4590_1, new_n4591,
    new_n4592, new_n4593, new_n4594, new_n4595_1, new_n4596, new_n4597,
    new_n4598, new_n4599, new_n4600, new_n4601, new_n4602, new_n4603,
    new_n4604, new_n4605, new_n4606, new_n4607, new_n4608, new_n4609,
    new_n4610, new_n4611, new_n4613, new_n4614, new_n4615, new_n4616,
    new_n4617, new_n4618, new_n4619, new_n4620, new_n4621, new_n4622,
    new_n4623, new_n4624_1, new_n4625, new_n4626, new_n4627, new_n4628,
    new_n4629, new_n4630, new_n4631, new_n4632, new_n4633, new_n4634,
    new_n4635, new_n4636, new_n4637, new_n4638, new_n4639, new_n4640,
    new_n4641, new_n4642, new_n4643, new_n4644, new_n4645, new_n4646_1,
    new_n4647, new_n4648, new_n4649, new_n4650, new_n4651, new_n4652,
    new_n4653, new_n4654, new_n4655, new_n4656, new_n4657, new_n4658,
    new_n4659, new_n4660, new_n4661, new_n4662, new_n4663, new_n4664,
    new_n4665_1, new_n4666, new_n4667, new_n4668, new_n4669, new_n4670,
    new_n4671, new_n4672, new_n4673, new_n4674_1, new_n4675, new_n4676,
    new_n4677, new_n4678, new_n4679, new_n4680, new_n4681, new_n4682,
    new_n4683, new_n4684, new_n4685, new_n4686, new_n4687, new_n4688,
    new_n4689, new_n4690, new_n4691, new_n4692, new_n4693_1, new_n4694,
    new_n4695, new_n4696, new_n4697, new_n4698, new_n4699, new_n4700,
    new_n4701, new_n4702, new_n4703, new_n4704, new_n4705, new_n4706,
    new_n4707, new_n4708, new_n4709, new_n4710, new_n4711, new_n4712,
    new_n4713, new_n4714, new_n4715, new_n4716, new_n4717, new_n4718,
    new_n4719, new_n4720, new_n4721, new_n4722_1, new_n4723, new_n4724,
    new_n4725, new_n4726, new_n4727, new_n4728, new_n4729, new_n4730,
    new_n4731_1, new_n4732, new_n4733, new_n4734, new_n4735, new_n4736,
    new_n4737, new_n4738, new_n4739, new_n4740, new_n4741, new_n4742,
    new_n4743, new_n4744, new_n4745_1, new_n4746, new_n4747_1, new_n4748,
    new_n4749, new_n4750, new_n4751, new_n4752, new_n4753, new_n4754,
    new_n4755, new_n4756, new_n4758, new_n4759, new_n4760, new_n4761,
    new_n4762, new_n4763, new_n4764, new_n4765, new_n4766_1, new_n4767,
    new_n4768, new_n4769, new_n4770_1, new_n4771, new_n4772, new_n4773,
    new_n4774, new_n4775, new_n4776, new_n4777_1, new_n4778, new_n4779,
    new_n4780, new_n4781, new_n4782, new_n4783, new_n4784, new_n4785_1,
    new_n4786, new_n4787, new_n4788, new_n4789, new_n4790, new_n4791,
    new_n4792, new_n4793, new_n4794, new_n4795, new_n4796, new_n4797,
    new_n4798, new_n4799, new_n4800, new_n4801, new_n4802, new_n4803,
    new_n4804_1, new_n4805, new_n4806, new_n4807, new_n4808, new_n4809,
    new_n4810_1, new_n4811, new_n4812_1, new_n4813, new_n4814_1, new_n4815,
    new_n4816, new_n4817, new_n4818, new_n4819, new_n4820, new_n4821,
    new_n4822, new_n4823, new_n4824, new_n4825, new_n4826, new_n4827,
    new_n4828, new_n4829, new_n4830, new_n4831, new_n4832, new_n4833,
    new_n4834, new_n4835, new_n4836, new_n4837, new_n4838, new_n4839,
    new_n4840, new_n4841, new_n4842, new_n4843, new_n4844, new_n4845,
    new_n4846, new_n4847, new_n4848, new_n4849, new_n4850_1, new_n4851,
    new_n4852, new_n4853, new_n4854, new_n4855, new_n4856, new_n4857,
    new_n4858_1, new_n4859, new_n4860, new_n4861, new_n4862, new_n4863,
    new_n4864, new_n4865, new_n4866, new_n4867, new_n4868, new_n4869,
    new_n4870, new_n4871, new_n4872, new_n4873, new_n4874, new_n4875,
    new_n4876, new_n4877, new_n4878, new_n4879, new_n4880, new_n4881,
    new_n4882, new_n4883, new_n4884, new_n4885, new_n4886, new_n4887,
    new_n4888, new_n4889, new_n4890, new_n4891_1, new_n4892, new_n4893,
    new_n4894, new_n4895, new_n4896, new_n4897, new_n4898, new_n4899,
    new_n4900, new_n4901, new_n4902, new_n4903, new_n4904, new_n4905,
    new_n4906, new_n4907, new_n4908, new_n4909, new_n4910, new_n4911,
    new_n4912, new_n4913_1, new_n4914, new_n4915, new_n4916, new_n4917,
    new_n4918, new_n4919, new_n4920, new_n4921, new_n4922, new_n4923,
    new_n4924, new_n4925_1, new_n4926, new_n4927, new_n4928, new_n4929,
    new_n4930, new_n4931, new_n4932, new_n4933, new_n4934, new_n4935,
    new_n4936, new_n4937, new_n4938, new_n4939_1, new_n4940, new_n4941,
    new_n4942, new_n4943, new_n4944, new_n4945, new_n4946, new_n4947_1,
    new_n4948, new_n4949, new_n4950, new_n4951, new_n4952_1, new_n4953,
    new_n4954, new_n4955, new_n4956, new_n4957_1, new_n4958, new_n4959,
    new_n4960, new_n4961, new_n4962, new_n4963, new_n4964_1, new_n4965,
    new_n4966_1, new_n4967_1, new_n4968, new_n4969, new_n4970, new_n4971,
    new_n4972_1, new_n4973, new_n4974, new_n4975, new_n4976, new_n4977,
    new_n4978, new_n4979, new_n4980, new_n4981, new_n4982, new_n4983,
    new_n4984, new_n4985, new_n4986, new_n4987, new_n4988, new_n4989,
    new_n4990, new_n4991, new_n4992, new_n4993, new_n4994, new_n4995,
    new_n4996, new_n4997, new_n4998, new_n4999, new_n5000, new_n5001,
    new_n5002, new_n5003, new_n5004, new_n5005, new_n5006, new_n5007,
    new_n5008, new_n5009, new_n5010, new_n5011_1, new_n5012, new_n5013,
    new_n5014, new_n5015, new_n5016, new_n5017, new_n5018, new_n5019,
    new_n5020_1, new_n5021, new_n5022, new_n5023, new_n5024_1, new_n5025_1,
    new_n5026_1, new_n5027, new_n5028, new_n5030, new_n5031_1, new_n5032,
    new_n5033, new_n5034, new_n5035, new_n5036, new_n5037, new_n5038,
    new_n5039, new_n5040, new_n5041, new_n5042, new_n5043, new_n5044,
    new_n5045, new_n5046_1, new_n5047, new_n5048, new_n5049, new_n5050,
    new_n5051, new_n5052, new_n5053, new_n5054, new_n5055, new_n5056,
    new_n5057, new_n5058, new_n5059, new_n5060_1, new_n5061, new_n5062_1,
    new_n5063, new_n5064_1, new_n5065, new_n5066, new_n5067, new_n5068,
    new_n5069, new_n5070, new_n5071, new_n5072, new_n5073, new_n5074,
    new_n5075, new_n5076, new_n5077_1, new_n5078, new_n5079, new_n5080,
    new_n5081, new_n5082_1, new_n5083, new_n5084, new_n5085, new_n5086,
    new_n5087, new_n5088, new_n5090, new_n5091, new_n5092, new_n5093,
    new_n5094, new_n5095, new_n5096, new_n5097, new_n5098_1, new_n5099,
    new_n5100, new_n5101_1, new_n5102, new_n5103, new_n5104, new_n5105,
    new_n5106, new_n5107, new_n5108, new_n5109, new_n5110, new_n5111,
    new_n5112, new_n5113, new_n5114, new_n5115_1, new_n5116, new_n5117,
    new_n5118, new_n5119, new_n5120_1, new_n5121, new_n5122, new_n5123,
    new_n5124, new_n5125, new_n5126, new_n5127, new_n5128_1, new_n5129,
    new_n5130, new_n5131_1, new_n5132, new_n5133, new_n5134, new_n5135,
    new_n5136, new_n5137, new_n5138, new_n5139, new_n5140_1, new_n5141,
    new_n5142, new_n5143, new_n5144, new_n5145, new_n5146, new_n5147,
    new_n5148, new_n5149, new_n5150, new_n5151, new_n5152, new_n5153,
    new_n5154, new_n5155, new_n5156, new_n5157, new_n5158_1, new_n5159,
    new_n5160, new_n5161, new_n5162, new_n5163, new_n5164, new_n5165,
    new_n5166, new_n5167, new_n5168_1, new_n5169, new_n5170, new_n5171,
    new_n5172, new_n5173, new_n5174, new_n5175, new_n5176, new_n5177,
    new_n5178, new_n5179, new_n5180, new_n5181, new_n5182, new_n5183,
    new_n5184_1, new_n5185, new_n5186, new_n5187, new_n5188, new_n5189,
    new_n5190, new_n5191, new_n5192, new_n5193, new_n5194, new_n5195,
    new_n5196, new_n5197, new_n5198, new_n5199, new_n5200, new_n5201,
    new_n5202, new_n5203, new_n5204, new_n5205, new_n5206, new_n5207,
    new_n5208, new_n5209, new_n5210, new_n5211_1, new_n5212, new_n5213_1,
    new_n5214, new_n5215, new_n5216, new_n5217, new_n5219, new_n5220,
    new_n5221, new_n5222, new_n5223, new_n5224, new_n5225, new_n5226_1,
    new_n5227, new_n5228_1, new_n5229, new_n5230, new_n5231, new_n5232,
    new_n5233, new_n5234, new_n5235, new_n5236, new_n5237, new_n5238,
    new_n5239, new_n5240, new_n5241, new_n5242, new_n5243, new_n5244,
    new_n5245, new_n5246, new_n5247, new_n5248, new_n5249, new_n5250,
    new_n5251, new_n5252, new_n5253, new_n5254, new_n5255_1, new_n5256_1,
    new_n5257, new_n5258, new_n5259, new_n5260, new_n5261, new_n5262,
    new_n5263, new_n5264, new_n5265_1, new_n5266, new_n5267, new_n5268,
    new_n5269, new_n5270, new_n5271, new_n5272, new_n5273_1, new_n5274_1,
    new_n5275, new_n5276, new_n5277, new_n5278, new_n5279, new_n5280,
    new_n5281, new_n5282, new_n5283, new_n5284, new_n5285, new_n5286,
    new_n5287, new_n5288, new_n5289, new_n5290, new_n5291, new_n5292,
    new_n5293, new_n5294, new_n5295, new_n5296, new_n5297, new_n5298,
    new_n5299, new_n5300_1, new_n5301, new_n5302_1, new_n5303, new_n5304,
    new_n5305, new_n5306, new_n5307, new_n5308, new_n5309, new_n5310,
    new_n5311, new_n5312, new_n5313, new_n5314, new_n5315, new_n5316,
    new_n5317, new_n5318, new_n5319, new_n5320, new_n5321, new_n5322,
    new_n5323, new_n5324, new_n5325_1, new_n5326, new_n5327, new_n5328,
    new_n5329, new_n5330_1, new_n5331, new_n5332, new_n5333, new_n5334,
    new_n5335, new_n5336, new_n5337_1, new_n5338, new_n5339, new_n5340,
    new_n5341, new_n5342, new_n5343, new_n5344, new_n5345, new_n5346,
    new_n5347, new_n5348, new_n5349, new_n5350, new_n5351_1, new_n5352,
    new_n5353_1, new_n5354, new_n5355, new_n5356, new_n5357, new_n5358,
    new_n5359, new_n5360, new_n5361, new_n5362, new_n5363, new_n5364,
    new_n5365, new_n5366, new_n5367, new_n5368, new_n5369, new_n5370,
    new_n5371, new_n5372, new_n5373, new_n5374, new_n5375, new_n5376_1,
    new_n5377, new_n5378, new_n5379, new_n5380, new_n5381, new_n5382,
    new_n5383, new_n5384, new_n5385, new_n5386_1, new_n5387, new_n5388,
    new_n5389, new_n5390, new_n5391, new_n5392, new_n5393, new_n5394,
    new_n5395, new_n5396, new_n5397, new_n5398, new_n5399_1, new_n5400_1,
    new_n5401, new_n5402, new_n5403_1, new_n5404, new_n5405, new_n5406,
    new_n5407, new_n5408, new_n5409, new_n5410, new_n5411, new_n5412,
    new_n5413, new_n5414, new_n5415, new_n5416, new_n5417, new_n5418,
    new_n5419, new_n5420, new_n5421, new_n5422, new_n5423, new_n5424,
    new_n5425, new_n5426, new_n5427, new_n5428, new_n5429, new_n5430_1,
    new_n5431, new_n5432, new_n5433, new_n5434, new_n5435, new_n5436,
    new_n5437, new_n5438_1, new_n5439_1, new_n5440, new_n5441, new_n5442,
    new_n5443_1, new_n5444, new_n5445, new_n5446, new_n5447, new_n5448,
    new_n5449, new_n5450, new_n5451_1, new_n5453, new_n5454, new_n5455,
    new_n5456, new_n5457, new_n5458, new_n5459, new_n5460, new_n5461,
    new_n5462, new_n5463, new_n5464, new_n5465, new_n5466, new_n5467,
    new_n5468, new_n5469, new_n5470, new_n5471, new_n5472_1, new_n5473,
    new_n5474, new_n5475, new_n5476, new_n5477, new_n5478, new_n5479,
    new_n5480, new_n5481, new_n5482, new_n5483, new_n5484, new_n5485_1,
    new_n5486, new_n5487, new_n5488, new_n5489, new_n5490, new_n5491,
    new_n5492, new_n5493, new_n5494, new_n5495, new_n5496, new_n5497,
    new_n5498, new_n5499, new_n5500, new_n5501, new_n5502, new_n5503,
    new_n5504, new_n5505, new_n5506, new_n5507, new_n5508, new_n5509,
    new_n5510, new_n5511, new_n5512, new_n5513, new_n5514, new_n5515,
    new_n5516, new_n5517_1, new_n5518, new_n5519, new_n5520, new_n5521_1,
    new_n5522, new_n5523, new_n5524_1, new_n5525, new_n5526, new_n5527,
    new_n5528, new_n5529, new_n5530, new_n5531, new_n5532_1, new_n5533,
    new_n5534, new_n5535, new_n5536, new_n5537, new_n5538, new_n5539,
    new_n5540, new_n5541, new_n5542, new_n5543, new_n5544, new_n5545,
    new_n5546, new_n5547, new_n5548, new_n5549, new_n5550, new_n5551,
    new_n5552, new_n5553, new_n5554, new_n5555, new_n5556, new_n5557,
    new_n5558, new_n5559, new_n5560, new_n5561, new_n5562, new_n5563,
    new_n5564_1, new_n5565, new_n5566, new_n5567, new_n5568, new_n5569,
    new_n5570, new_n5571, new_n5572, new_n5573, new_n5574, new_n5575,
    new_n5576, new_n5577, new_n5578, new_n5579_1, new_n5580, new_n5581,
    new_n5582, new_n5583, new_n5584, new_n5585, new_n5586, new_n5587,
    new_n5588, new_n5589, new_n5590, new_n5591, new_n5592, new_n5593_1,
    new_n5594, new_n5595, new_n5596, new_n5597, new_n5598, new_n5599,
    new_n5600, new_n5601, new_n5602, new_n5603_1, new_n5604, new_n5605_1,
    new_n5606, new_n5607, new_n5608, new_n5609_1, new_n5610, new_n5611,
    new_n5612, new_n5613, new_n5614, new_n5615, new_n5616, new_n5617,
    new_n5618, new_n5619, new_n5620, new_n5621, new_n5622, new_n5623,
    new_n5624, new_n5625, new_n5626, new_n5627, new_n5628, new_n5629,
    new_n5630, new_n5631, new_n5632, new_n5633, new_n5634_1, new_n5635,
    new_n5636, new_n5637, new_n5638, new_n5639, new_n5640, new_n5641,
    new_n5642, new_n5643_1, new_n5644, new_n5645, new_n5646, new_n5647,
    new_n5648, new_n5649, new_n5650, new_n5651, new_n5652, new_n5653,
    new_n5654, new_n5655, new_n5656, new_n5657, new_n5658, new_n5659,
    new_n5660, new_n5661, new_n5662, new_n5663, new_n5664, new_n5665,
    new_n5666, new_n5667, new_n5668, new_n5669, new_n5670, new_n5671,
    new_n5672, new_n5673, new_n5674, new_n5675, new_n5676, new_n5677,
    new_n5678, new_n5679, new_n5680_1, new_n5681, new_n5682, new_n5683,
    new_n5684, new_n5685, new_n5686, new_n5687_1, new_n5688, new_n5689,
    new_n5690, new_n5691, new_n5692, new_n5693, new_n5694, new_n5695,
    new_n5696_1, new_n5697, new_n5698, new_n5699, new_n5700_1, new_n5701,
    new_n5702, new_n5703, new_n5704_1, new_n5705, new_n5706, new_n5707,
    new_n5708, new_n5709, new_n5710, new_n5711, new_n5712, new_n5713,
    new_n5714, new_n5715, new_n5716, new_n5717, new_n5718, new_n5719,
    new_n5720, new_n5721, new_n5722, new_n5723, new_n5724, new_n5725,
    new_n5726, new_n5727, new_n5728, new_n5729, new_n5730, new_n5731,
    new_n5732_1, new_n5733, new_n5734, new_n5735, new_n5736, new_n5737,
    new_n5738, new_n5739, new_n5740, new_n5741, new_n5742_1, new_n5743,
    new_n5744, new_n5745, new_n5746, new_n5747, new_n5748, new_n5749,
    new_n5750, new_n5751, new_n5752_1, new_n5753, new_n5754, new_n5755,
    new_n5756, new_n5757, new_n5758, new_n5759, new_n5760, new_n5761,
    new_n5762, new_n5763, new_n5764, new_n5765_1, new_n5766, new_n5767,
    new_n5769, new_n5770, new_n5771, new_n5772, new_n5773, new_n5774,
    new_n5775, new_n5776_1, new_n5777, new_n5778, new_n5779, new_n5780,
    new_n5781, new_n5782_1, new_n5783, new_n5784, new_n5785, new_n5786,
    new_n5787, new_n5788, new_n5789, new_n5790, new_n5792, new_n5793,
    new_n5794, new_n5795, new_n5798, new_n5799, new_n5800, new_n5801,
    new_n5802, new_n5803, new_n5804, new_n5805, new_n5806, new_n5807,
    new_n5808, new_n5809, new_n5810, new_n5811, new_n5812, new_n5813,
    new_n5814, new_n5815, new_n5816, new_n5817, new_n5818, new_n5819,
    new_n5820, new_n5821, new_n5822_1, new_n5823, new_n5825, new_n5826,
    new_n5827, new_n5828, new_n5829, new_n5830, new_n5831, new_n5832,
    new_n5833_1, new_n5834_1, new_n5835, new_n5836, new_n5837, new_n5838,
    new_n5839, new_n5840_1, new_n5841_1, new_n5842_1, new_n5843, new_n5844,
    new_n5845, new_n5846, new_n5847, new_n5848, new_n5849, new_n5850_1,
    new_n5851, new_n5853, new_n5856, new_n5857, new_n5858, new_n5859,
    new_n5860, new_n5861, new_n5862, new_n5863, new_n5864, new_n5865,
    new_n5866, new_n5867, new_n5868, new_n5869, new_n5870, new_n5871,
    new_n5872, new_n5873, new_n5874, new_n5875, new_n5876, new_n5877,
    new_n5878, new_n5879, new_n5880, new_n5881, new_n5882_1, new_n5883,
    new_n5884, new_n5885, new_n5886, new_n5887, new_n5888, new_n5889,
    new_n5890, new_n5891, new_n5892, new_n5893, new_n5894, new_n5895,
    new_n5896, new_n5897, new_n5898, new_n5899, new_n5900, new_n5901,
    new_n5902, new_n5903_1, new_n5904_1, new_n5905, new_n5906, new_n5907,
    new_n5908, new_n5909, new_n5910, new_n5911_1, new_n5912, new_n5913,
    new_n5914, new_n5915, new_n5916, new_n5917, new_n5918, new_n5919,
    new_n5920, new_n5921, new_n5922, new_n5923, new_n5924, new_n5925,
    new_n5926, new_n5927, new_n5928, new_n5929, new_n5930, new_n5931,
    new_n5932, new_n5933, new_n5934, new_n5935, new_n5936_1, new_n5937,
    new_n5938, new_n5939, new_n5940, new_n5941, new_n5942, new_n5943_1,
    new_n5944, new_n5945, new_n5946, new_n5947, new_n5948, new_n5949,
    new_n5950, new_n5951, new_n5952, new_n5953, new_n5954, new_n5955,
    new_n5956, new_n5957, new_n5958, new_n5959, new_n5960, new_n5961,
    new_n5962, new_n5963, new_n5964_1, new_n5965, new_n5966, new_n5967,
    new_n5968, new_n5969, new_n5970, new_n5971, new_n5972, new_n5973,
    new_n5974, new_n5975, new_n5976, new_n5977, new_n5978, new_n5979,
    new_n5980_1, new_n5981, new_n5982, new_n5983, new_n5984, new_n5985,
    new_n5986, new_n5987, new_n5988, new_n5989, new_n5990, new_n5991,
    new_n5992, new_n5993, new_n5994, new_n5995, new_n5996, new_n5997,
    new_n5998, new_n5999, new_n6000, new_n6001, new_n6002, new_n6003,
    new_n6004, new_n6005, new_n6006, new_n6007, new_n6008, new_n6009,
    new_n6010, new_n6011, new_n6012_1, new_n6013, new_n6014, new_n6015,
    new_n6016, new_n6017, new_n6018, new_n6019, new_n6020, new_n6021,
    new_n6022_1, new_n6023, new_n6024, new_n6025, new_n6026, new_n6027,
    new_n6028, new_n6029, new_n6030, new_n6031_1, new_n6032, new_n6033,
    new_n6034, new_n6035, new_n6036, new_n6037, new_n6038, new_n6039,
    new_n6040, new_n6041, new_n6042, new_n6043, new_n6044_1, new_n6045,
    new_n6046_1, new_n6047, new_n6048, new_n6049, new_n6050, new_n6051,
    new_n6052, new_n6053, new_n6054, new_n6055, new_n6056, new_n6057,
    new_n6058, new_n6059, new_n6060, new_n6061, new_n6062, new_n6063,
    new_n6064, new_n6065, new_n6066, new_n6067, new_n6068, new_n6069,
    new_n6070, new_n6071, new_n6072, new_n6073, new_n6074, new_n6075,
    new_n6076, new_n6077, new_n6078, new_n6079, new_n6080, new_n6081,
    new_n6082, new_n6083, new_n6084_1, new_n6085, new_n6086, new_n6087,
    new_n6088, new_n6089, new_n6090, new_n6091, new_n6092, new_n6093,
    new_n6094, new_n6095, new_n6096, new_n6097, new_n6098, new_n6099,
    new_n6100, new_n6101, new_n6102, new_n6103, new_n6104_1, new_n6105_1,
    new_n6106, new_n6107, new_n6108, new_n6109, new_n6110, new_n6111,
    new_n6112, new_n6113, new_n6114, new_n6115, new_n6116, new_n6117,
    new_n6118, new_n6119, new_n6120, new_n6121, new_n6122, new_n6123,
    new_n6124, new_n6125, new_n6126, new_n6127, new_n6128, new_n6129,
    new_n6130, new_n6131, new_n6132, new_n6133, new_n6134, new_n6135,
    new_n6136, new_n6137, new_n6138, new_n6139, new_n6140, new_n6141,
    new_n6142, new_n6143, new_n6144, new_n6145, new_n6146, new_n6147,
    new_n6148, new_n6149, new_n6151, new_n6152, new_n6153, new_n6154,
    new_n6155, new_n6156, new_n6157, new_n6158, new_n6159, new_n6160_1,
    new_n6161, new_n6162, new_n6163, new_n6164, new_n6165, new_n6166,
    new_n6167, new_n6168, new_n6169, new_n6170, new_n6171_1, new_n6172,
    new_n6173, new_n6174, new_n6175, new_n6176, new_n6177, new_n6178,
    new_n6179, new_n6180, new_n6181, new_n6182, new_n6183_1, new_n6184,
    new_n6185, new_n6186, new_n6187, new_n6188, new_n6189_1, new_n6190,
    new_n6191, new_n6192, new_n6193, new_n6194, new_n6195, new_n6196,
    new_n6197, new_n6198, new_n6199, new_n6200, new_n6201, new_n6202,
    new_n6203, new_n6204_1, new_n6205, new_n6206, new_n6207, new_n6208,
    new_n6209, new_n6210, new_n6211, new_n6212, new_n6213, new_n6214,
    new_n6215, new_n6216, new_n6217, new_n6218_1, new_n6219, new_n6220,
    new_n6221, new_n6222, new_n6223_1, new_n6224, new_n6225, new_n6226,
    new_n6227, new_n6228, new_n6229, new_n6230, new_n6231, new_n6232,
    new_n6233_1, new_n6234, new_n6235, new_n6236, new_n6237, new_n6238,
    new_n6239, new_n6240, new_n6241, new_n6242, new_n6243, new_n6244,
    new_n6245_1, new_n6246, new_n6247, new_n6248_1, new_n6249, new_n6250,
    new_n6251, new_n6252, new_n6253, new_n6254, new_n6255, new_n6256_1,
    new_n6257, new_n6258, new_n6259, new_n6260, new_n6261, new_n6262,
    new_n6263, new_n6264, new_n6265, new_n6266, new_n6267, new_n6268,
    new_n6269, new_n6270, new_n6271_1, new_n6272, new_n6273, new_n6274,
    new_n6275, new_n6276_1, new_n6277, new_n6278, new_n6279, new_n6280,
    new_n6281, new_n6282, new_n6283, new_n6284, new_n6285, new_n6286,
    new_n6287, new_n6288, new_n6289, new_n6290, new_n6291, new_n6292,
    new_n6293, new_n6294, new_n6295, new_n6296, new_n6297, new_n6298,
    new_n6299, new_n6300, new_n6301, new_n6302, new_n6303, new_n6304,
    new_n6305, new_n6306, new_n6307, new_n6308_1, new_n6309, new_n6310,
    new_n6311_1, new_n6312, new_n6313, new_n6314, new_n6315, new_n6316,
    new_n6317, new_n6318, new_n6319, new_n6320, new_n6321, new_n6322,
    new_n6323_1, new_n6324, new_n6325, new_n6326, new_n6327, new_n6328,
    new_n6329, new_n6330_1, new_n6331, new_n6332, new_n6333, new_n6334,
    new_n6335, new_n6336, new_n6337, new_n6338, new_n6339_1, new_n6340,
    new_n6341, new_n6342, new_n6343, new_n6344, new_n6345, new_n6346,
    new_n6347, new_n6348, new_n6349, new_n6350, new_n6351, new_n6352,
    new_n6353, new_n6354_1, new_n6355, new_n6356_1, new_n6357, new_n6358,
    new_n6359, new_n6360, new_n6361, new_n6362, new_n6363, new_n6364,
    new_n6365, new_n6366, new_n6367, new_n6368, new_n6369_1, new_n6370,
    new_n6371, new_n6372, new_n6373, new_n6374, new_n6375_1, new_n6376,
    new_n6377, new_n6378, new_n6379_1, new_n6380, new_n6381_1, new_n6382,
    new_n6383_1, new_n6384, new_n6385_1, new_n6386, new_n6387, new_n6388,
    new_n6389, new_n6390, new_n6391, new_n6392, new_n6393, new_n6394,
    new_n6395, new_n6396, new_n6397_1, new_n6398, new_n6399, new_n6400,
    new_n6401, new_n6402, new_n6403, new_n6404, new_n6405, new_n6406,
    new_n6407_1, new_n6408, new_n6409, new_n6410, new_n6411, new_n6412,
    new_n6413, new_n6414, new_n6415, new_n6416, new_n6417, new_n6418,
    new_n6419, new_n6420, new_n6421, new_n6422, new_n6423, new_n6425,
    new_n6426, new_n6427_1, new_n6428, new_n6429, new_n6430, new_n6431_1,
    new_n6432, new_n6433, new_n6434, new_n6435, new_n6436, new_n6437_1,
    new_n6438, new_n6439, new_n6440, new_n6441, new_n6442, new_n6443,
    new_n6444, new_n6445, new_n6446, new_n6447, new_n6448, new_n6449,
    new_n6450, new_n6451, new_n6452, new_n6453, new_n6454, new_n6455,
    new_n6456_1, new_n6457_1, new_n6458, new_n6459, new_n6460, new_n6461,
    new_n6462, new_n6463, new_n6464, new_n6465_1, new_n6466, new_n6467,
    new_n6468, new_n6469, new_n6470_1, new_n6471, new_n6472, new_n6473,
    new_n6474, new_n6475, new_n6476_1, new_n6477, new_n6478, new_n6479,
    new_n6480, new_n6481, new_n6482, new_n6483, new_n6484, new_n6485_1,
    new_n6486, new_n6487, new_n6488, new_n6489, new_n6490, new_n6491,
    new_n6492, new_n6493, new_n6494, new_n6495, new_n6496, new_n6497,
    new_n6498, new_n6499, new_n6500, new_n6501, new_n6502_1, new_n6503,
    new_n6504, new_n6505, new_n6506_1, new_n6507, new_n6508, new_n6509,
    new_n6510, new_n6511, new_n6512, new_n6513_1, new_n6514_1, new_n6515,
    new_n6516, new_n6517, new_n6518, new_n6519, new_n6520, new_n6521,
    new_n6522, new_n6523, new_n6524, new_n6525, new_n6526, new_n6527,
    new_n6528, new_n6529, new_n6530, new_n6531, new_n6532, new_n6533,
    new_n6534, new_n6535, new_n6536, new_n6537, new_n6538, new_n6539,
    new_n6540, new_n6541, new_n6542_1, new_n6543, new_n6544, new_n6545,
    new_n6546, new_n6547, new_n6548, new_n6549, new_n6550, new_n6551,
    new_n6552, new_n6553, new_n6554, new_n6555, new_n6556_1, new_n6557,
    new_n6558_1, new_n6559, new_n6560_1, new_n6561, new_n6562, new_n6563,
    new_n6564, new_n6565, new_n6566, new_n6567_1, new_n6568, new_n6569,
    new_n6570, new_n6571, new_n6572, new_n6573, new_n6574, new_n6575,
    new_n6576_1, new_n6577, new_n6578, new_n6579, new_n6580, new_n6581,
    new_n6582, new_n6583, new_n6585, new_n6586, new_n6587_1, new_n6589,
    new_n6590_1, new_n6591, new_n6592, new_n6593, new_n6594, new_n6595,
    new_n6596_1, new_n6597, new_n6598, new_n6599, new_n6600, new_n6601,
    new_n6602, new_n6603, new_n6604, new_n6605, new_n6606, new_n6607,
    new_n6608, new_n6609, new_n6610, new_n6611_1, new_n6612_1, new_n6613,
    new_n6614, new_n6615, new_n6616, new_n6617, new_n6618, new_n6619,
    new_n6620, new_n6621, new_n6622, new_n6623, new_n6624, new_n6625,
    new_n6626, new_n6627, new_n6628_1, new_n6629, new_n6630_1, new_n6631_1,
    new_n6632, new_n6633, new_n6634_1, new_n6635, new_n6636, new_n6637,
    new_n6638, new_n6639, new_n6640, new_n6641, new_n6642, new_n6643,
    new_n6644, new_n6645, new_n6646, new_n6647, new_n6648, new_n6649,
    new_n6650, new_n6651, new_n6652_1, new_n6653, new_n6654, new_n6655_1,
    new_n6656, new_n6657, new_n6658, new_n6659_1, new_n6660, new_n6661,
    new_n6662, new_n6663, new_n6664, new_n6665, new_n6666, new_n6667,
    new_n6668, new_n6669_1, new_n6670, new_n6671_1, new_n6672, new_n6673_1,
    new_n6675, new_n6676, new_n6677, new_n6678, new_n6679, new_n6680,
    new_n6681, new_n6682, new_n6683, new_n6684_1, new_n6685, new_n6686,
    new_n6687, new_n6688, new_n6689, new_n6690, new_n6691_1, new_n6692,
    new_n6693, new_n6694, new_n6695, new_n6696, new_n6697, new_n6698,
    new_n6699, new_n6700, new_n6701, new_n6702, new_n6703, new_n6704,
    new_n6705, new_n6706_1, new_n6707_1, new_n6708, new_n6709, new_n6710,
    new_n6711, new_n6712, new_n6713, new_n6714, new_n6715, new_n6716,
    new_n6717, new_n6718, new_n6719, new_n6720, new_n6721, new_n6722,
    new_n6723, new_n6724, new_n6725, new_n6726, new_n6727, new_n6728,
    new_n6729_1, new_n6730, new_n6731, new_n6732, new_n6733, new_n6734,
    new_n6735, new_n6736_1, new_n6737, new_n6738, new_n6739, new_n6740,
    new_n6741, new_n6742, new_n6744, new_n6745, new_n6746, new_n6747,
    new_n6748, new_n6749, new_n6750, new_n6751, new_n6752, new_n6753,
    new_n6754, new_n6755, new_n6756, new_n6757, new_n6758, new_n6759,
    new_n6760, new_n6761, new_n6762, new_n6763, new_n6764, new_n6765,
    new_n6766, new_n6767, new_n6768, new_n6769, new_n6770, new_n6771,
    new_n6772, new_n6773_1, new_n6774, new_n6775_1, new_n6776, new_n6777,
    new_n6778, new_n6779, new_n6780, new_n6781, new_n6782, new_n6783,
    new_n6784, new_n6785_1, new_n6786, new_n6787, new_n6788, new_n6789,
    new_n6790_1, new_n6791_1, new_n6792, new_n6793, new_n6794_1, new_n6795,
    new_n6796, new_n6797, new_n6798, new_n6799, new_n6800, new_n6801,
    new_n6802_1, new_n6803, new_n6804, new_n6805, new_n6806, new_n6807,
    new_n6808, new_n6809, new_n6810, new_n6811, new_n6812, new_n6813,
    new_n6814_1, new_n6815, new_n6816, new_n6817, new_n6818, new_n6819,
    new_n6820, new_n6821, new_n6822, new_n6823, new_n6824, new_n6825,
    new_n6826_1, new_n6827, new_n6828, new_n6829, new_n6830, new_n6831,
    new_n6832, new_n6833, new_n6834, new_n6835_1, new_n6836, new_n6837,
    new_n6838, new_n6839, new_n6840, new_n6841, new_n6842, new_n6843,
    new_n6844, new_n6845, new_n6846, new_n6847, new_n6848, new_n6849,
    new_n6850, new_n6851, new_n6852, new_n6853_1, new_n6854, new_n6855,
    new_n6856, new_n6857, new_n6858, new_n6859, new_n6860, new_n6861_1,
    new_n6862_1, new_n6863_1, new_n6864, new_n6865, new_n6866, new_n6867_1,
    new_n6868, new_n6869, new_n6870, new_n6871, new_n6872, new_n6873,
    new_n6874, new_n6875, new_n6876, new_n6877, new_n6878, new_n6879,
    new_n6880, new_n6881, new_n6882, new_n6883, new_n6884, new_n6885,
    new_n6886, new_n6887, new_n6888, new_n6889, new_n6890, new_n6891,
    new_n6892, new_n6893, new_n6894, new_n6895, new_n6896, new_n6897,
    new_n6898, new_n6899, new_n6900, new_n6901, new_n6902, new_n6903,
    new_n6904, new_n6905, new_n6906, new_n6907, new_n6908, new_n6909,
    new_n6910, new_n6911, new_n6912, new_n6913, new_n6914, new_n6915,
    new_n6916, new_n6917, new_n6918, new_n6919, new_n6920, new_n6921,
    new_n6922, new_n6923, new_n6924, new_n6925, new_n6926, new_n6927,
    new_n6928, new_n6929, new_n6930, new_n6931, new_n6932, new_n6933,
    new_n6934, new_n6935, new_n6936, new_n6937, new_n6938, new_n6939,
    new_n6940, new_n6941, new_n6942, new_n6943, new_n6944, new_n6945,
    new_n6946, new_n6947, new_n6948, new_n6949, new_n6950, new_n6951,
    new_n6952, new_n6953, new_n6954, new_n6955, new_n6956, new_n6957,
    new_n6958, new_n6959, new_n6960, new_n6961, new_n6962, new_n6963,
    new_n6964, new_n6966, new_n6967_1, new_n6968, new_n6969, new_n6970,
    new_n6971_1, new_n6972, new_n6973, new_n6974, new_n6975_1, new_n6976,
    new_n6977, new_n6978, new_n6979, new_n6980, new_n6981, new_n6982,
    new_n6983_1, new_n6984, new_n6985_1, new_n6986, new_n6987, new_n6988,
    new_n6989, new_n6990, new_n6991, new_n6992, new_n6993, new_n6994,
    new_n6995, new_n6996, new_n6997, new_n6998_1, new_n6999, new_n7000,
    new_n7001, new_n7002, new_n7003, new_n7004, new_n7005, new_n7006,
    new_n7007, new_n7008, new_n7009, new_n7010, new_n7011, new_n7012,
    new_n7013, new_n7014, new_n7015, new_n7016, new_n7017, new_n7018,
    new_n7019, new_n7020, new_n7021, new_n7022, new_n7023, new_n7024,
    new_n7025, new_n7026_1, new_n7027, new_n7028, new_n7029, new_n7030,
    new_n7031, new_n7032_1, new_n7033, new_n7034, new_n7035, new_n7036,
    new_n7037, new_n7038_1, new_n7039, new_n7040, new_n7041, new_n7042,
    new_n7043, new_n7044, new_n7045, new_n7046, new_n7047, new_n7048,
    new_n7049, new_n7050, new_n7051, new_n7052, new_n7053, new_n7054,
    new_n7055, new_n7056, new_n7057_1, new_n7058, new_n7059, new_n7060,
    new_n7061, new_n7062, new_n7063, new_n7064, new_n7065, new_n7066,
    new_n7067, new_n7068, new_n7069, new_n7070, new_n7071, new_n7072,
    new_n7073, new_n7074, new_n7075, new_n7076, new_n7077, new_n7078,
    new_n7079_1, new_n7080, new_n7081, new_n7082, new_n7083, new_n7084,
    new_n7085, new_n7086, new_n7087, new_n7088, new_n7089, new_n7090,
    new_n7091, new_n7092, new_n7093, new_n7094, new_n7095, new_n7096,
    new_n7097, new_n7098, new_n7099_1, new_n7100, new_n7101, new_n7102,
    new_n7103, new_n7104, new_n7105, new_n7106, new_n7107, new_n7108,
    new_n7109, new_n7110, new_n7111, new_n7112, new_n7113, new_n7114,
    new_n7115, new_n7116, new_n7117, new_n7118, new_n7119, new_n7120,
    new_n7121, new_n7122, new_n7123, new_n7124, new_n7125, new_n7126,
    new_n7127, new_n7128, new_n7129, new_n7130, new_n7131, new_n7132,
    new_n7133, new_n7134, new_n7135, new_n7136, new_n7137, new_n7138,
    new_n7139_1, new_n7140, new_n7141, new_n7142, new_n7143, new_n7144,
    new_n7145, new_n7146, new_n7147, new_n7148, new_n7149_1, new_n7150,
    new_n7151, new_n7152, new_n7153, new_n7154, new_n7155, new_n7156,
    new_n7157, new_n7158, new_n7159, new_n7160, new_n7161, new_n7162,
    new_n7163, new_n7164, new_n7165, new_n7166, new_n7167, new_n7168,
    new_n7169, new_n7170, new_n7171, new_n7172, new_n7173, new_n7174,
    new_n7175, new_n7176, new_n7177, new_n7178, new_n7179, new_n7180,
    new_n7181, new_n7182, new_n7183, new_n7184, new_n7185, new_n7186,
    new_n7187, new_n7188, new_n7189, new_n7190_1, new_n7191, new_n7192,
    new_n7193, new_n7194, new_n7195, new_n7196, new_n7198, new_n7199,
    new_n7200, new_n7201, new_n7203, new_n7204, new_n7205, new_n7206,
    new_n7207, new_n7208, new_n7209, new_n7210, new_n7211, new_n7212,
    new_n7213, new_n7214, new_n7215, new_n7216, new_n7217, new_n7218,
    new_n7219, new_n7220, new_n7221, new_n7222, new_n7223, new_n7224,
    new_n7225, new_n7226, new_n7227, new_n7228, new_n7229_1, new_n7230_1,
    new_n7231, new_n7232, new_n7233_1, new_n7234, new_n7235, new_n7236_1,
    new_n7237, new_n7238, new_n7239, new_n7240, new_n7241, new_n7242,
    new_n7243, new_n7244, new_n7245, new_n7246, new_n7247, new_n7248,
    new_n7249, new_n7250, new_n7251, new_n7252, new_n7253_1, new_n7254,
    new_n7255, new_n7256_1, new_n7257, new_n7258, new_n7259, new_n7260,
    new_n7261, new_n7262, new_n7263, new_n7264, new_n7265, new_n7266,
    new_n7267, new_n7268_1, new_n7269, new_n7270, new_n7271, new_n7272,
    new_n7273, new_n7274, new_n7275, new_n7276, new_n7277_1, new_n7278,
    new_n7279, new_n7280_1, new_n7281, new_n7282, new_n7283, new_n7284,
    new_n7285, new_n7286, new_n7287, new_n7288, new_n7289, new_n7290,
    new_n7291, new_n7292, new_n7293, new_n7294, new_n7295, new_n7296,
    new_n7297, new_n7298_1, new_n7299, new_n7300, new_n7301, new_n7302,
    new_n7303, new_n7304, new_n7305_1, new_n7306, new_n7307, new_n7308_1,
    new_n7309, new_n7310, new_n7311, new_n7312, new_n7313_1, new_n7314,
    new_n7315, new_n7316, new_n7317, new_n7318, new_n7319, new_n7320,
    new_n7321, new_n7322, new_n7323, new_n7324, new_n7325, new_n7326,
    new_n7327, new_n7328, new_n7329, new_n7330_1, new_n7331, new_n7332,
    new_n7333, new_n7334, new_n7335_1, new_n7336, new_n7337, new_n7338,
    new_n7339_1, new_n7340, new_n7341, new_n7342, new_n7343, new_n7344,
    new_n7345, new_n7346_1, new_n7347, new_n7348, new_n7349_1, new_n7350,
    new_n7351, new_n7352, new_n7353, new_n7354, new_n7355, new_n7356,
    new_n7357, new_n7358, new_n7359, new_n7360, new_n7361, new_n7362,
    new_n7363_1, new_n7364, new_n7365, new_n7366, new_n7367, new_n7368,
    new_n7369, new_n7370, new_n7371, new_n7372, new_n7373, new_n7374,
    new_n7375, new_n7376, new_n7377_1, new_n7378, new_n7379, new_n7380,
    new_n7381, new_n7382, new_n7383, new_n7384, new_n7385, new_n7386,
    new_n7387, new_n7388, new_n7389, new_n7390_1, new_n7391, new_n7392,
    new_n7393, new_n7394, new_n7395, new_n7396, new_n7397, new_n7398,
    new_n7399, new_n7400, new_n7401, new_n7402, new_n7403_1, new_n7404,
    new_n7405, new_n7406, new_n7407, new_n7408_1, new_n7409, new_n7410,
    new_n7411, new_n7412, new_n7413, new_n7414, new_n7415, new_n7416,
    new_n7417, new_n7418, new_n7419, new_n7420, new_n7421_1, new_n7422,
    new_n7423, new_n7424, new_n7425, new_n7426, new_n7427, new_n7429,
    new_n7430, new_n7431, new_n7432_1, new_n7433, new_n7434, new_n7435,
    new_n7436, new_n7437_1, new_n7438, new_n7439, new_n7440, new_n7441,
    new_n7442, new_n7443, new_n7444, new_n7445, new_n7446, new_n7447,
    new_n7448, new_n7449, new_n7450, new_n7451, new_n7452, new_n7453,
    new_n7454, new_n7455, new_n7456, new_n7457, new_n7458, new_n7459,
    new_n7460_1, new_n7461, new_n7462, new_n7463, new_n7464, new_n7465,
    new_n7466, new_n7467, new_n7468, new_n7469, new_n7470, new_n7471,
    new_n7472, new_n7473, new_n7474, new_n7475_1, new_n7476, new_n7477_1,
    new_n7478, new_n7479, new_n7480, new_n7481, new_n7482, new_n7483,
    new_n7484, new_n7485, new_n7486, new_n7487, new_n7488, new_n7489,
    new_n7490, new_n7491, new_n7492, new_n7493, new_n7494, new_n7495,
    new_n7496, new_n7497, new_n7498, new_n7499, new_n7500, new_n7501,
    new_n7502, new_n7503, new_n7504, new_n7505, new_n7506, new_n7507_1,
    new_n7508, new_n7509, new_n7510, new_n7511, new_n7512, new_n7513,
    new_n7514_1, new_n7515, new_n7516, new_n7517, new_n7518, new_n7519,
    new_n7520, new_n7521, new_n7522, new_n7523, new_n7524_1, new_n7525,
    new_n7526, new_n7527, new_n7528, new_n7529, new_n7530, new_n7531,
    new_n7532, new_n7533, new_n7534, new_n7535, new_n7536, new_n7537,
    new_n7538, new_n7539, new_n7540, new_n7541, new_n7542, new_n7543,
    new_n7544, new_n7545, new_n7546, new_n7547, new_n7548, new_n7549,
    new_n7550, new_n7551, new_n7552, new_n7553, new_n7554, new_n7555,
    new_n7556, new_n7557, new_n7558_1, new_n7559, new_n7560, new_n7561,
    new_n7562, new_n7563, new_n7564, new_n7565, new_n7566_1, new_n7567,
    new_n7568, new_n7569_1, new_n7570, new_n7571, new_n7572_1, new_n7573,
    new_n7574, new_n7575_1, new_n7576, new_n7577, new_n7578, new_n7579,
    new_n7580, new_n7581, new_n7582, new_n7583, new_n7584, new_n7585_1,
    new_n7586, new_n7587, new_n7588_1, new_n7589, new_n7590, new_n7591,
    new_n7592, new_n7593_1, new_n7594, new_n7595, new_n7596, new_n7597,
    new_n7598_1, new_n7599, new_n7600, new_n7601, new_n7602, new_n7603,
    new_n7604, new_n7605, new_n7606, new_n7608, new_n7609, new_n7610_1,
    new_n7611, new_n7612, new_n7613, new_n7614, new_n7615, new_n7616_1,
    new_n7617, new_n7618, new_n7619, new_n7620, new_n7621, new_n7622,
    new_n7623, new_n7624, new_n7625, new_n7626, new_n7627, new_n7628,
    new_n7629, new_n7630_1, new_n7631, new_n7632, new_n7633, new_n7634,
    new_n7635, new_n7636, new_n7637, new_n7638, new_n7639, new_n7640,
    new_n7641, new_n7642, new_n7643_1, new_n7644, new_n7645, new_n7646,
    new_n7647_1, new_n7648, new_n7649, new_n7650, new_n7651, new_n7652,
    new_n7653, new_n7654, new_n7655, new_n7656, new_n7657_1, new_n7658,
    new_n7659, new_n7660, new_n7661, new_n7662, new_n7663, new_n7664,
    new_n7665, new_n7666, new_n7667, new_n7668, new_n7669, new_n7670_1,
    new_n7671, new_n7672, new_n7673, new_n7674_1, new_n7675, new_n7676,
    new_n7677, new_n7678_1, new_n7679_1, new_n7680, new_n7681, new_n7682,
    new_n7683, new_n7684, new_n7685, new_n7686_1, new_n7687, new_n7688,
    new_n7689, new_n7690, new_n7691, new_n7692_1, new_n7693_1, new_n7694,
    new_n7695, new_n7696, new_n7697, new_n7698_1, new_n7699, new_n7700,
    new_n7701, new_n7702, new_n7703, new_n7704, new_n7705, new_n7706,
    new_n7707, new_n7708_1, new_n7709, new_n7710, new_n7711, new_n7712,
    new_n7713, new_n7714, new_n7715, new_n7716, new_n7717, new_n7718,
    new_n7719, new_n7720, new_n7721_1, new_n7722, new_n7723, new_n7724,
    new_n7725, new_n7726, new_n7727, new_n7728, new_n7729, new_n7730,
    new_n7731_1, new_n7732, new_n7733, new_n7734, new_n7735, new_n7736,
    new_n7737, new_n7738, new_n7739, new_n7740, new_n7741, new_n7742,
    new_n7743, new_n7744, new_n7745, new_n7746, new_n7747, new_n7748,
    new_n7749, new_n7750, new_n7751_1, new_n7752, new_n7753, new_n7754,
    new_n7755, new_n7756, new_n7757, new_n7758, new_n7759_1, new_n7760,
    new_n7761, new_n7762, new_n7763, new_n7764, new_n7765, new_n7766,
    new_n7767, new_n7768, new_n7769_1, new_n7770, new_n7771, new_n7772,
    new_n7773_1, new_n7774, new_n7775, new_n7776, new_n7777, new_n7778,
    new_n7779, new_n7780_1, new_n7781, new_n7782, new_n7783, new_n7784,
    new_n7785, new_n7786, new_n7787, new_n7788_1, new_n7789, new_n7790,
    new_n7791, new_n7792, new_n7793, new_n7794_1, new_n7795, new_n7796,
    new_n7797, new_n7798, new_n7799, new_n7800, new_n7801, new_n7802,
    new_n7803, new_n7804, new_n7805, new_n7806, new_n7807, new_n7808,
    new_n7809, new_n7810, new_n7811_1, new_n7812, new_n7813, new_n7814,
    new_n7815, new_n7816, new_n7817, new_n7818, new_n7819, new_n7820,
    new_n7821, new_n7822, new_n7823, new_n7824, new_n7825, new_n7826,
    new_n7827, new_n7828, new_n7829, new_n7830_1, new_n7831, new_n7832,
    new_n7833, new_n7834_1, new_n7835, new_n7836, new_n7837, new_n7838,
    new_n7839, new_n7840, new_n7841_1, new_n7842, new_n7843, new_n7844,
    new_n7845, new_n7846, new_n7847, new_n7848, new_n7849, new_n7850,
    new_n7851, new_n7852, new_n7853, new_n7854, new_n7855, new_n7856,
    new_n7857, new_n7858, new_n7859, new_n7860, new_n7861, new_n7862,
    new_n7863, new_n7864, new_n7865, new_n7866, new_n7867, new_n7868,
    new_n7869, new_n7870, new_n7871, new_n7872, new_n7873, new_n7874,
    new_n7875, new_n7876_1, new_n7877, new_n7878, new_n7879, new_n7880,
    new_n7881, new_n7882, new_n7883, new_n7884_1, new_n7885, new_n7886,
    new_n7887, new_n7888, new_n7889, new_n7890, new_n7891, new_n7892,
    new_n7893, new_n7894, new_n7895, new_n7896, new_n7897, new_n7898,
    new_n7899, new_n7900, new_n7901, new_n7902, new_n7903, new_n7904,
    new_n7905, new_n7906, new_n7907, new_n7908, new_n7909, new_n7910,
    new_n7911, new_n7912, new_n7913, new_n7914, new_n7915, new_n7916,
    new_n7918, new_n7919, new_n7920, new_n7921, new_n7922, new_n7923,
    new_n7924, new_n7925, new_n7926, new_n7927, new_n7928, new_n7929,
    new_n7930, new_n7931, new_n7932, new_n7933, new_n7934, new_n7935,
    new_n7936, new_n7937_1, new_n7938, new_n7939, new_n7940, new_n7941,
    new_n7942, new_n7943_1, new_n7944, new_n7945, new_n7946, new_n7947,
    new_n7948, new_n7949_1, new_n7950_1, new_n7951, new_n7952, new_n7953,
    new_n7954, new_n7955, new_n7956, new_n7957, new_n7958, new_n7959_1,
    new_n7960, new_n7961, new_n7962, new_n7963_1, new_n7964, new_n7965,
    new_n7966, new_n7967, new_n7968_1, new_n7969, new_n7970, new_n7971,
    new_n7972, new_n7973, new_n7974, new_n7975, new_n7976, new_n7977,
    new_n7978, new_n7979, new_n7980, new_n7981, new_n7982, new_n7983,
    new_n7984, new_n7985, new_n7986, new_n7987, new_n7988, new_n7989,
    new_n7990, new_n7991, new_n7992_1, new_n7993, new_n7994, new_n7995,
    new_n7996, new_n7997, new_n7998, new_n7999_1, new_n8000, new_n8001,
    new_n8002, new_n8003, new_n8004, new_n8005, new_n8006_1, new_n8007,
    new_n8008, new_n8009, new_n8010, new_n8011, new_n8012, new_n8013,
    new_n8014, new_n8015, new_n8016, new_n8017, new_n8018, new_n8019,
    new_n8020, new_n8021, new_n8022, new_n8023, new_n8024, new_n8025,
    new_n8026, new_n8027_1, new_n8028, new_n8029, new_n8030, new_n8031_1,
    new_n8032, new_n8033, new_n8034, new_n8035, new_n8036, new_n8037,
    new_n8038, new_n8039, new_n8040, new_n8041, new_n8042_1, new_n8043,
    new_n8044, new_n8045, new_n8046, new_n8047, new_n8048, new_n8049,
    new_n8050, new_n8051, new_n8052_1, new_n8053, new_n8054, new_n8055,
    new_n8056, new_n8057, new_n8058, new_n8059, new_n8060, new_n8061,
    new_n8062, new_n8063, new_n8064, new_n8065, new_n8066, new_n8067_1,
    new_n8068, new_n8069, new_n8070, new_n8071, new_n8072, new_n8073,
    new_n8074, new_n8075, new_n8076, new_n8077, new_n8078, new_n8079,
    new_n8080, new_n8081, new_n8082, new_n8083, new_n8084, new_n8085,
    new_n8086, new_n8087, new_n8088, new_n8089, new_n8090, new_n8091,
    new_n8092, new_n8093, new_n8094, new_n8095_1, new_n8096, new_n8097,
    new_n8098, new_n8099, new_n8100, new_n8101, new_n8102, new_n8103_1,
    new_n8104, new_n8105, new_n8106, new_n8107, new_n8108, new_n8109_1,
    new_n8110, new_n8111, new_n8112, new_n8113, new_n8114, new_n8115,
    new_n8116, new_n8117, new_n8118, new_n8119, new_n8120, new_n8121,
    new_n8122, new_n8123, new_n8124, new_n8125, new_n8126, new_n8127_1,
    new_n8128, new_n8129, new_n8130_1, new_n8131, new_n8132, new_n8133,
    new_n8134, new_n8135_1, new_n8136, new_n8137, new_n8138, new_n8139_1,
    new_n8140, new_n8141, new_n8142, new_n8143, new_n8144, new_n8145,
    new_n8146, new_n8147, new_n8148_1, new_n8149_1, new_n8150, new_n8151,
    new_n8152, new_n8153, new_n8154, new_n8155, new_n8156, new_n8157,
    new_n8158, new_n8159_1, new_n8160, new_n8161, new_n8162, new_n8163,
    new_n8164, new_n8165, new_n8166, new_n8167, new_n8168, new_n8169,
    new_n8170, new_n8171, new_n8172, new_n8173, new_n8174, new_n8175,
    new_n8176, new_n8177, new_n8178, new_n8179_1, new_n8180, new_n8181,
    new_n8182, new_n8183, new_n8184, new_n8185, new_n8186, new_n8187,
    new_n8188, new_n8189, new_n8190, new_n8191, new_n8192, new_n8193,
    new_n8194_1, new_n8195, new_n8196, new_n8197, new_n8198, new_n8199,
    new_n8200, new_n8201, new_n8202, new_n8203, new_n8204, new_n8205,
    new_n8208, new_n8209, new_n8210, new_n8211, new_n8212, new_n8213,
    new_n8214, new_n8215_1, new_n8216, new_n8217, new_n8218, new_n8219,
    new_n8220, new_n8221, new_n8222, new_n8223, new_n8224, new_n8225,
    new_n8226, new_n8227, new_n8228, new_n8229, new_n8230, new_n8231,
    new_n8232, new_n8233, new_n8234, new_n8235, new_n8236, new_n8237,
    new_n8238, new_n8239, new_n8240, new_n8241, new_n8242, new_n8243,
    new_n8244_1, new_n8245, new_n8246, new_n8247, new_n8248, new_n8249,
    new_n8250, new_n8251, new_n8252, new_n8253, new_n8254, new_n8255_1,
    new_n8256_1, new_n8257, new_n8258, new_n8259_1, new_n8260, new_n8261,
    new_n8262, new_n8263, new_n8264, new_n8265, new_n8266, new_n8267_1,
    new_n8268, new_n8269, new_n8270, new_n8271, new_n8272, new_n8273,
    new_n8274, new_n8275, new_n8276_1, new_n8277, new_n8278, new_n8279,
    new_n8280, new_n8281, new_n8282, new_n8283, new_n8284, new_n8285_1,
    new_n8286, new_n8287, new_n8288_1, new_n8289, new_n8290, new_n8291,
    new_n8292, new_n8293, new_n8294, new_n8295, new_n8296, new_n8297,
    new_n8298, new_n8299, new_n8300, new_n8301, new_n8302, new_n8303,
    new_n8304, new_n8305_1, new_n8306_1, new_n8307, new_n8308, new_n8309_1,
    new_n8310, new_n8311, new_n8312, new_n8313, new_n8314, new_n8315,
    new_n8316, new_n8317, new_n8318, new_n8319, new_n8320_1, new_n8321_1,
    new_n8322, new_n8323, new_n8324_1, new_n8325, new_n8326, new_n8327,
    new_n8328, new_n8329, new_n8330, new_n8331, new_n8332, new_n8333,
    new_n8334, new_n8335, new_n8336, new_n8337, new_n8338, new_n8339_1,
    new_n8340, new_n8341, new_n8342, new_n8343, new_n8344, new_n8345,
    new_n8346, new_n8347, new_n8348, new_n8349, new_n8350, new_n8351,
    new_n8352, new_n8353, new_n8354, new_n8355, new_n8356, new_n8357,
    new_n8358, new_n8359, new_n8360, new_n8361, new_n8362, new_n8363_1,
    new_n8364, new_n8365, new_n8366, new_n8367, new_n8368, new_n8369,
    new_n8370, new_n8371, new_n8372, new_n8373, new_n8374, new_n8375,
    new_n8376_1, new_n8377, new_n8378, new_n8379, new_n8380, new_n8381_1,
    new_n8382, new_n8383, new_n8384, new_n8385, new_n8386, new_n8387,
    new_n8388, new_n8389, new_n8390, new_n8391, new_n8393, new_n8394,
    new_n8395, new_n8396, new_n8397, new_n8398, new_n8399_1, new_n8400,
    new_n8401, new_n8402, new_n8403, new_n8404, new_n8405_1, new_n8406,
    new_n8407, new_n8408_1, new_n8409, new_n8410, new_n8411, new_n8412,
    new_n8413, new_n8414, new_n8415, new_n8416, new_n8417_1, new_n8418,
    new_n8419, new_n8420, new_n8421, new_n8422, new_n8423, new_n8424,
    new_n8425, new_n8426, new_n8427, new_n8428, new_n8429, new_n8430,
    new_n8432_1, new_n8433, new_n8434, new_n8435, new_n8436, new_n8437,
    new_n8438, new_n8439_1, new_n8440, new_n8441, new_n8442, new_n8443,
    new_n8444, new_n8445, new_n8446, new_n8447, new_n8448, new_n8449,
    new_n8450, new_n8451, new_n8452, new_n8453_1, new_n8454, new_n8455,
    new_n8456, new_n8457, new_n8458, new_n8459, new_n8460, new_n8461,
    new_n8462, new_n8463, new_n8464, new_n8465, new_n8466, new_n8467,
    new_n8468, new_n8469, new_n8470, new_n8471, new_n8472, new_n8473,
    new_n8474, new_n8476, new_n8477, new_n8478, new_n8479, new_n8480_1,
    new_n8481, new_n8482, new_n8483, new_n8484, new_n8485, new_n8486,
    new_n8487, new_n8488, new_n8489_1, new_n8490, new_n8491, new_n8492,
    new_n8493, new_n8494, new_n8495, new_n8496, new_n8497, new_n8498,
    new_n8499, new_n8500, new_n8501, new_n8502, new_n8503, new_n8504,
    new_n8505_1, new_n8506, new_n8507, new_n8508, new_n8509, new_n8510_1,
    new_n8511, new_n8512, new_n8513, new_n8514, new_n8515, new_n8516,
    new_n8517, new_n8518, new_n8519_1, new_n8520, new_n8521, new_n8522,
    new_n8523, new_n8524, new_n8525, new_n8526_1, new_n8527, new_n8528,
    new_n8529, new_n8530, new_n8531, new_n8532, new_n8533, new_n8534,
    new_n8535_1, new_n8536, new_n8537, new_n8538, new_n8539, new_n8540,
    new_n8541, new_n8542, new_n8543, new_n8544, new_n8545, new_n8546,
    new_n8547, new_n8548, new_n8549, new_n8550_1, new_n8551, new_n8552,
    new_n8553, new_n8554, new_n8555, new_n8556, new_n8557, new_n8558,
    new_n8559, new_n8560, new_n8561, new_n8562, new_n8563_1, new_n8564,
    new_n8565, new_n8566, new_n8567, new_n8568, new_n8569, new_n8570,
    new_n8572, new_n8573, new_n8574, new_n8575, new_n8576, new_n8577,
    new_n8578, new_n8579, new_n8580, new_n8581_1, new_n8582, new_n8583,
    new_n8584, new_n8585, new_n8586, new_n8587, new_n8588, new_n8589,
    new_n8590, new_n8591, new_n8592, new_n8593, new_n8594_1, new_n8595,
    new_n8596, new_n8597, new_n8598, new_n8599, new_n8600, new_n8601,
    new_n8602, new_n8603, new_n8604, new_n8605, new_n8606, new_n8607,
    new_n8608_1, new_n8609, new_n8610, new_n8611, new_n8612, new_n8613,
    new_n8614_1, new_n8615, new_n8616, new_n8617, new_n8618, new_n8619,
    new_n8620_1, new_n8621, new_n8622, new_n8623, new_n8624, new_n8625,
    new_n8626, new_n8627, new_n8628, new_n8629, new_n8630, new_n8631,
    new_n8632, new_n8633, new_n8634, new_n8635, new_n8636, new_n8637_1,
    new_n8638_1, new_n8639, new_n8640, new_n8641, new_n8642, new_n8643,
    new_n8645, new_n8646, new_n8647, new_n8648, new_n8649, new_n8650,
    new_n8651, new_n8652, new_n8653, new_n8654, new_n8655, new_n8656_1,
    new_n8657, new_n8658, new_n8659, new_n8660, new_n8661, new_n8662_1,
    new_n8663, new_n8664, new_n8665, new_n8666, new_n8667, new_n8668,
    new_n8669, new_n8670, new_n8671, new_n8672, new_n8673, new_n8674,
    new_n8675, new_n8676, new_n8677, new_n8678_1, new_n8679, new_n8680,
    new_n8681, new_n8682, new_n8683, new_n8684, new_n8685, new_n8686,
    new_n8687_1, new_n8688, new_n8689, new_n8690, new_n8691, new_n8692,
    new_n8693, new_n8694_1, new_n8695, new_n8696, new_n8697, new_n8698,
    new_n8699, new_n8700, new_n8701, new_n8702, new_n8703, new_n8704,
    new_n8705, new_n8706, new_n8707, new_n8708, new_n8709, new_n8710,
    new_n8711, new_n8712, new_n8713, new_n8714, new_n8715, new_n8716_1,
    new_n8717, new_n8718, new_n8719, new_n8720, new_n8721_1, new_n8722,
    new_n8723, new_n8724, new_n8725, new_n8726, new_n8727, new_n8728,
    new_n8729, new_n8730, new_n8731, new_n8732, new_n8733, new_n8734,
    new_n8735, new_n8736, new_n8737, new_n8738, new_n8739, new_n8740,
    new_n8741, new_n8742, new_n8743, new_n8744_1, new_n8745_1, new_n8746,
    new_n8747, new_n8748, new_n8749, new_n8750, new_n8751, new_n8752,
    new_n8753, new_n8754, new_n8755, new_n8756, new_n8757, new_n8758,
    new_n8759, new_n8760, new_n8761, new_n8762, new_n8763, new_n8764,
    new_n8765, new_n8766, new_n8767, new_n8768, new_n8769, new_n8770,
    new_n8771, new_n8772, new_n8773, new_n8774, new_n8775, new_n8776,
    new_n8777, new_n8778, new_n8779, new_n8780, new_n8781, new_n8782_1,
    new_n8783, new_n8784, new_n8785, new_n8786, new_n8787, new_n8788,
    new_n8789, new_n8790, new_n8791, new_n8792, new_n8793, new_n8794,
    new_n8795, new_n8796, new_n8797, new_n8798, new_n8799, new_n8800,
    new_n8801, new_n8802, new_n8803_1, new_n8804, new_n8805, new_n8806_1,
    new_n8807, new_n8808, new_n8809_1, new_n8810, new_n8811, new_n8812,
    new_n8813, new_n8814, new_n8815, new_n8816, new_n8817, new_n8818,
    new_n8819, new_n8820, new_n8821_1, new_n8822, new_n8823, new_n8824_1,
    new_n8825, new_n8826, new_n8827_1, new_n8828, new_n8829, new_n8830,
    new_n8831, new_n8832, new_n8833, new_n8834, new_n8835, new_n8836,
    new_n8837, new_n8838, new_n8839, new_n8840, new_n8841, new_n8842,
    new_n8843, new_n8844, new_n8845, new_n8846, new_n8847, new_n8848,
    new_n8849_1, new_n8850, new_n8851, new_n8852, new_n8853, new_n8854,
    new_n8855, new_n8856_1, new_n8857, new_n8858, new_n8859, new_n8860,
    new_n8861_1, new_n8862_1, new_n8863, new_n8864, new_n8865, new_n8866,
    new_n8867, new_n8868, new_n8869_1, new_n8870, new_n8871, new_n8872,
    new_n8873, new_n8874, new_n8875, new_n8876, new_n8877, new_n8878,
    new_n8879, new_n8880, new_n8881, new_n8882, new_n8883, new_n8884_1,
    new_n8885, new_n8886, new_n8887, new_n8888, new_n8889, new_n8890,
    new_n8891, new_n8892, new_n8893, new_n8894, new_n8895, new_n8896,
    new_n8897, new_n8898, new_n8899, new_n8900, new_n8901, new_n8902,
    new_n8903, new_n8904, new_n8905, new_n8906, new_n8907, new_n8908,
    new_n8909_1, new_n8911_1, new_n8912, new_n8913, new_n8915, new_n8916,
    new_n8917, new_n8918, new_n8919, new_n8920_1, new_n8921, new_n8922,
    new_n8923, new_n8924, new_n8925, new_n8926, new_n8927, new_n8928,
    new_n8929, new_n8930, new_n8931, new_n8932, new_n8933, new_n8934,
    new_n8935, new_n8936, new_n8937, new_n8938, new_n8939, new_n8940,
    new_n8941, new_n8942, new_n8943_1, new_n8944, new_n8945, new_n8946,
    new_n8947, new_n8948, new_n8949, new_n8950, new_n8951, new_n8952,
    new_n8953, new_n8954, new_n8955, new_n8956, new_n8957, new_n8958,
    new_n8959, new_n8960, new_n8961, new_n8962, new_n8963, new_n8964_1,
    new_n8965, new_n8966, new_n8967, new_n8968, new_n8969, new_n8970,
    new_n8971_1, new_n8972, new_n8973, new_n8974, new_n8975, new_n8976,
    new_n8977, new_n8978, new_n8979, new_n8980, new_n8981, new_n8982_1,
    new_n8983, new_n8984, new_n8985, new_n8986, new_n8987, new_n8988,
    new_n8989, new_n8990, new_n8991, new_n8992, new_n8993_1, new_n8994,
    new_n8995, new_n8996, new_n8997, new_n8998, new_n8999, new_n9000,
    new_n9001, new_n9002, new_n9003_1, new_n9004, new_n9005, new_n9006,
    new_n9007, new_n9008, new_n9009, new_n9010, new_n9011, new_n9012_1,
    new_n9013, new_n9014, new_n9015, new_n9016, new_n9017, new_n9018,
    new_n9019, new_n9020, new_n9021, new_n9022, new_n9023, new_n9024,
    new_n9025, new_n9026, new_n9027, new_n9028, new_n9029, new_n9030,
    new_n9031, new_n9032_1, new_n9033, new_n9034, new_n9035, new_n9036,
    new_n9037, new_n9038, new_n9039, new_n9040, new_n9041, new_n9042_1,
    new_n9043, new_n9044, new_n9045, new_n9046_1, new_n9047_1, new_n9048,
    new_n9049, new_n9050, new_n9051, new_n9052, new_n9053, new_n9054,
    new_n9055, new_n9056, new_n9057, new_n9058, new_n9059, new_n9061,
    new_n9062, new_n9063, new_n9064, new_n9065, new_n9066, new_n9067,
    new_n9068, new_n9069, new_n9070, new_n9071, new_n9072, new_n9073,
    new_n9074, new_n9075, new_n9076, new_n9077, new_n9078, new_n9079,
    new_n9080, new_n9081, new_n9082, new_n9083, new_n9084, new_n9085,
    new_n9086, new_n9087, new_n9088, new_n9089, new_n9090_1, new_n9091,
    new_n9092, new_n9093, new_n9094, new_n9095, new_n9096, new_n9097,
    new_n9098, new_n9099, new_n9100, new_n9101, new_n9102, new_n9103,
    new_n9104_1, new_n9105, new_n9106, new_n9107, new_n9108, new_n9109,
    new_n9110, new_n9111, new_n9112, new_n9113, new_n9114, new_n9115,
    new_n9116, new_n9117, new_n9118, new_n9119, new_n9120, new_n9121,
    new_n9122, new_n9123, new_n9124, new_n9125, new_n9126, new_n9127,
    new_n9128, new_n9129_1, new_n9130, new_n9131, new_n9132, new_n9133,
    new_n9134, new_n9135, new_n9136, new_n9137, new_n9138, new_n9139,
    new_n9140, new_n9141, new_n9142, new_n9143, new_n9144, new_n9145,
    new_n9146_1, new_n9147, new_n9148, new_n9149, new_n9150, new_n9151,
    new_n9152, new_n9153, new_n9154, new_n9155, new_n9156, new_n9157,
    new_n9158, new_n9159, new_n9160, new_n9161, new_n9162, new_n9163,
    new_n9164_1, new_n9165, new_n9166_1, new_n9167, new_n9168, new_n9169,
    new_n9170, new_n9171, new_n9172_1, new_n9173, new_n9174, new_n9175,
    new_n9176, new_n9177, new_n9178, new_n9179, new_n9180, new_n9181,
    new_n9182_1, new_n9183, new_n9184, new_n9185, new_n9186, new_n9187,
    new_n9188, new_n9189, new_n9190, new_n9191_1, new_n9192, new_n9193,
    new_n9194, new_n9195, new_n9196, new_n9197, new_n9198, new_n9199,
    new_n9200, new_n9201, new_n9202, new_n9203, new_n9204, new_n9205,
    new_n9206, new_n9207, new_n9208, new_n9209, new_n9210, new_n9211,
    new_n9212, new_n9213, new_n9214, new_n9215, new_n9216, new_n9217_1,
    new_n9218, new_n9219, new_n9220_1, new_n9221, new_n9226, new_n9227,
    new_n9228, new_n9229, new_n9230, new_n9231, new_n9232, new_n9233,
    new_n9234, new_n9235, new_n9236, new_n9237, new_n9238, new_n9239,
    new_n9240, new_n9241, new_n9242, new_n9243, new_n9244, new_n9245,
    new_n9246_1, new_n9247, new_n9248, new_n9249, new_n9250, new_n9251_1,
    new_n9252, new_n9253, new_n9254, new_n9255, new_n9256, new_n9257,
    new_n9258, new_n9259_1, new_n9260, new_n9261_1, new_n9262, new_n9263,
    new_n9264, new_n9265, new_n9266, new_n9267, new_n9268, new_n9269,
    new_n9270, new_n9271, new_n9272, new_n9273, new_n9274, new_n9275,
    new_n9276, new_n9277, new_n9278, new_n9279, new_n9280, new_n9281,
    new_n9282, new_n9283, new_n9284, new_n9285, new_n9286, new_n9287_1,
    new_n9288, new_n9289, new_n9290, new_n9291, new_n9292, new_n9293,
    new_n9294, new_n9295, new_n9296, new_n9297, new_n9298, new_n9299,
    new_n9300, new_n9301, new_n9302, new_n9303, new_n9304, new_n9305,
    new_n9306, new_n9307, new_n9308_1, new_n9309, new_n9310, new_n9311,
    new_n9312, new_n9313, new_n9314, new_n9315, new_n9316, new_n9317,
    new_n9318_1, new_n9319, new_n9320, new_n9321, new_n9322, new_n9323_1,
    new_n9324, new_n9325, new_n9326, new_n9327, new_n9328, new_n9329,
    new_n9330, new_n9331, new_n9332, new_n9333, new_n9334, new_n9335,
    new_n9336, new_n9337, new_n9338, new_n9339, new_n9340, new_n9341,
    new_n9342, new_n9343, new_n9344_1, new_n9345, new_n9346, new_n9347,
    new_n9348, new_n9349, new_n9350, new_n9351, new_n9352, new_n9353,
    new_n9354, new_n9355, new_n9356, new_n9357, new_n9358, new_n9359,
    new_n9360, new_n9361, new_n9362, new_n9363, new_n9364_1, new_n9365,
    new_n9366, new_n9367, new_n9368, new_n9369, new_n9370, new_n9371_1,
    new_n9372_1, new_n9373, new_n9374, new_n9375, new_n9376, new_n9377,
    new_n9378, new_n9379, new_n9380_1, new_n9381, new_n9382_1, new_n9383,
    new_n9384, new_n9385, new_n9386, new_n9387, new_n9388, new_n9389,
    new_n9390, new_n9391, new_n9393, new_n9394, new_n9395, new_n9396_1,
    new_n9397, new_n9398, new_n9399_1, new_n9400, new_n9401, new_n9402,
    new_n9403_1, new_n9404, new_n9405, new_n9406, new_n9407, new_n9408,
    new_n9409, new_n9410, new_n9411, new_n9412, new_n9413, new_n9414,
    new_n9415, new_n9416, new_n9417, new_n9418, new_n9419_1, new_n9420,
    new_n9421, new_n9422, new_n9423_1, new_n9424, new_n9425, new_n9426,
    new_n9427, new_n9428, new_n9429, new_n9430_1, new_n9431, new_n9432,
    new_n9433, new_n9434, new_n9435_1, new_n9436, new_n9437, new_n9438,
    new_n9439, new_n9440, new_n9441, new_n9442, new_n9443, new_n9444,
    new_n9445_1, new_n9446, new_n9447, new_n9448, new_n9449, new_n9450,
    new_n9451_1, new_n9452, new_n9453, new_n9454, new_n9455, new_n9456,
    new_n9457, new_n9458_1, new_n9459_1, new_n9460_1, new_n9461, new_n9462,
    new_n9463, new_n9464, new_n9465, new_n9466, new_n9467, new_n9468,
    new_n9469, new_n9470, new_n9471, new_n9472, new_n9473, new_n9476,
    new_n9477, new_n9478, new_n9479, new_n9480, new_n9481, new_n9482,
    new_n9483, new_n9484, new_n9485, new_n9486, new_n9487, new_n9488,
    new_n9489, new_n9490, new_n9491, new_n9492, new_n9493_1, new_n9494,
    new_n9495, new_n9496, new_n9497, new_n9498, new_n9499, new_n9500,
    new_n9501, new_n9502, new_n9503, new_n9504, new_n9505, new_n9506,
    new_n9507_1, new_n9508_1, new_n9509, new_n9510, new_n9511, new_n9512_1,
    new_n9513, new_n9514, new_n9515, new_n9516, new_n9517, new_n9518,
    new_n9519, new_n9520, new_n9521, new_n9522, new_n9523, new_n9524,
    new_n9525, new_n9526, new_n9527, new_n9528, new_n9529, new_n9530,
    new_n9531, new_n9532, new_n9533, new_n9534, new_n9535, new_n9536,
    new_n9537, new_n9538, new_n9539, new_n9540, new_n9541, new_n9542,
    new_n9543, new_n9544, new_n9545, new_n9546, new_n9547, new_n9548,
    new_n9549, new_n9550, new_n9551, new_n9552_1, new_n9553, new_n9554_1,
    new_n9555, new_n9556_1, new_n9557_1, new_n9558_1, new_n9559, new_n9560,
    new_n9561, new_n9562, new_n9563, new_n9564, new_n9565, new_n9566,
    new_n9567, new_n9569, new_n9570, new_n9571, new_n9572, new_n9573,
    new_n9574, new_n9575, new_n9576, new_n9577, new_n9578, new_n9579,
    new_n9580, new_n9581, new_n9582, new_n9583, new_n9584, new_n9585,
    new_n9586, new_n9587, new_n9588, new_n9589, new_n9590, new_n9591,
    new_n9592, new_n9593, new_n9594, new_n9595, new_n9596, new_n9597,
    new_n9598_1, new_n9599, new_n9600, new_n9601, new_n9602, new_n9603,
    new_n9604, new_n9605, new_n9606, new_n9607, new_n9608, new_n9609,
    new_n9610, new_n9611, new_n9612, new_n9613, new_n9614, new_n9615,
    new_n9616_1, new_n9617, new_n9618, new_n9619, new_n9620, new_n9621,
    new_n9622_1, new_n9623, new_n9624, new_n9625, new_n9626_1, new_n9627,
    new_n9628, new_n9629, new_n9630, new_n9631, new_n9632, new_n9633_1,
    new_n9634, new_n9635_1, new_n9636, new_n9637, new_n9638, new_n9639,
    new_n9640, new_n9641, new_n9642, new_n9643, new_n9644, new_n9645,
    new_n9646_1, new_n9647, new_n9648_1, new_n9649, new_n9650, new_n9651,
    new_n9652, new_n9653, new_n9654, new_n9655_1, new_n9656, new_n9657,
    new_n9658, new_n9659, new_n9660, new_n9661, new_n9662, new_n9663,
    new_n9664, new_n9665, new_n9666, new_n9667, new_n9668, new_n9669,
    new_n9670, new_n9671, new_n9672, new_n9673, new_n9674, new_n9675,
    new_n9676, new_n9677, new_n9678, new_n9679, new_n9680, new_n9681,
    new_n9682, new_n9683, new_n9684, new_n9685, new_n9686, new_n9687,
    new_n9688, new_n9689_1, new_n9690, new_n9691, new_n9692, new_n9693,
    new_n9694, new_n9695_1, new_n9696, new_n9697, new_n9698, new_n9699_1,
    new_n9700, new_n9701, new_n9702, new_n9703, new_n9705, new_n9707,
    new_n9708, new_n9709, new_n9710, new_n9712, new_n9713, new_n9714,
    new_n9715, new_n9716, new_n9717, new_n9718, new_n9719, new_n9720,
    new_n9721, new_n9722, new_n9723, new_n9724, new_n9725, new_n9726_1,
    new_n9727, new_n9729, new_n9731, new_n9732, new_n9733, new_n9734,
    new_n9735, new_n9736, new_n9737, new_n9738, new_n9739, new_n9740,
    new_n9741, new_n9742, new_n9743, new_n9744, new_n9745, new_n9746,
    new_n9747, new_n9748, new_n9749, new_n9750, new_n9751, new_n9752,
    new_n9753_1, new_n9754, new_n9755, new_n9756, new_n9757, new_n9758,
    new_n9759, new_n9760, new_n9761_1, new_n9762, new_n9763_1, new_n9764,
    new_n9765, new_n9766, new_n9767_1, new_n9768, new_n9769, new_n9770,
    new_n9771_1, new_n9772, new_n9773, new_n9774, new_n9775, new_n9776,
    new_n9777, new_n9778_1, new_n9779, new_n9780, new_n9781, new_n9782,
    new_n9783_1, new_n9784, new_n9785, new_n9786, new_n9787, new_n9788,
    new_n9789, new_n9790, new_n9791, new_n9792, new_n9793, new_n9794,
    new_n9795, new_n9796, new_n9797, new_n9798, new_n9799, new_n9800,
    new_n9801, new_n9802, new_n9803_1, new_n9804, new_n9805, new_n9806,
    new_n9807, new_n9808, new_n9809, new_n9810, new_n9811, new_n9812,
    new_n9813, new_n9814, new_n9815, new_n9816, new_n9817, new_n9818,
    new_n9819, new_n9820, new_n9821, new_n9822, new_n9823, new_n9824,
    new_n9825, new_n9826, new_n9827, new_n9828, new_n9829, new_n9830,
    new_n9831, new_n9832_1, new_n9833_1, new_n9834, new_n9835, new_n9836,
    new_n9837, new_n9838_1, new_n9839, new_n9840, new_n9841, new_n9842,
    new_n9843, new_n9844, new_n9845, new_n9846, new_n9847, new_n9848,
    new_n9849, new_n9850, new_n9851, new_n9852, new_n9853, new_n9854,
    new_n9855, new_n9856, new_n9857, new_n9858, new_n9859, new_n9860,
    new_n9861, new_n9862, new_n9863, new_n9864, new_n9865, new_n9866,
    new_n9867_1, new_n9868, new_n9869, new_n9870, new_n9871, new_n9872_1,
    new_n9873, new_n9874, new_n9875, new_n9876, new_n9877, new_n9878,
    new_n9879, new_n9880, new_n9881, new_n9882, new_n9883, new_n9884,
    new_n9885, new_n9886, new_n9887, new_n9888, new_n9889, new_n9890_1,
    new_n9891, new_n9892, new_n9893, new_n9894, new_n9895, new_n9896,
    new_n9897, new_n9898, new_n9899, new_n9900, new_n9901, new_n9902,
    new_n9903, new_n9904, new_n9905, new_n9906, new_n9907, new_n9908,
    new_n9909, new_n9910, new_n9911, new_n9912, new_n9913, new_n9914,
    new_n9915, new_n9916, new_n9917_1, new_n9918, new_n9919_1, new_n9920,
    new_n9921, new_n9922, new_n9923, new_n9924, new_n9925, new_n9926_1,
    new_n9927, new_n9928, new_n9929, new_n9930, new_n9931, new_n9932,
    new_n9933, new_n9934_1, new_n9935, new_n9936, new_n9937, new_n9938_1,
    new_n9939, new_n9940, new_n9941, new_n9942_1, new_n9943, new_n9944,
    new_n9945, new_n9946_1, new_n9947, new_n9948, new_n9949, new_n9950,
    new_n9951, new_n9952, new_n9953, new_n9954, new_n9955, new_n9956,
    new_n9957, new_n9958, new_n9959, new_n9960, new_n9961, new_n9962,
    new_n9963, new_n9964, new_n9965, new_n9966, new_n9967_1, new_n9968_1,
    new_n9969, new_n9970, new_n9971, new_n9972, new_n9973, new_n9974,
    new_n9975, new_n9976, new_n9977, new_n9978, new_n9979, new_n9980,
    new_n9981, new_n9982, new_n9983, new_n9984, new_n9985, new_n9986,
    new_n9988, new_n9989, new_n9990, new_n9991, new_n9992, new_n9993,
    new_n9994, new_n9995, new_n9996, new_n9997, new_n9998, new_n9999,
    new_n10000, new_n10001, new_n10002, new_n10003, new_n10004, new_n10005,
    new_n10006, new_n10007, new_n10008, new_n10009_1, new_n10010_1,
    new_n10011, new_n10012, new_n10013, new_n10014, new_n10015, new_n10016,
    new_n10017_1, new_n10018_1, new_n10019_1, new_n10020, new_n10021_1,
    new_n10022, new_n10023, new_n10024, new_n10025, new_n10026, new_n10027,
    new_n10028, new_n10029, new_n10030, new_n10031, new_n10032, new_n10033,
    new_n10034, new_n10035, new_n10036, new_n10037, new_n10038, new_n10039,
    new_n10040, new_n10041, new_n10042, new_n10043, new_n10044, new_n10045,
    new_n10046, new_n10047, new_n10048, new_n10049, new_n10050, new_n10051,
    new_n10052, new_n10053_1, new_n10054, new_n10055_1, new_n10056,
    new_n10057_1, new_n10058, new_n10059, new_n10060, new_n10061,
    new_n10062, new_n10063, new_n10064, new_n10065, new_n10066, new_n10067,
    new_n10068, new_n10069, new_n10070, new_n10071, new_n10072, new_n10073,
    new_n10074, new_n10075, new_n10076, new_n10077, new_n10078, new_n10079,
    new_n10080, new_n10081, new_n10082, new_n10083, new_n10084, new_n10085,
    new_n10086, new_n10087, new_n10088, new_n10089, new_n10090, new_n10091,
    new_n10092, new_n10093, new_n10094, new_n10095, new_n10096_1,
    new_n10097, new_n10098, new_n10099, new_n10100, new_n10101_1,
    new_n10102, new_n10103, new_n10104, new_n10105, new_n10106, new_n10107,
    new_n10108, new_n10109, new_n10110, new_n10111_1, new_n10112,
    new_n10113, new_n10114, new_n10115, new_n10116, new_n10117_1,
    new_n10118, new_n10119, new_n10120, new_n10121, new_n10122, new_n10123,
    new_n10124, new_n10125_1, new_n10126, new_n10127, new_n10128,
    new_n10129, new_n10130, new_n10131, new_n10132, new_n10133, new_n10134,
    new_n10135, new_n10136, new_n10137, new_n10138, new_n10139, new_n10140,
    new_n10141, new_n10142, new_n10143, new_n10144, new_n10145, new_n10146,
    new_n10147, new_n10148, new_n10149, new_n10150, new_n10151, new_n10152,
    new_n10153, new_n10154, new_n10155, new_n10156, new_n10157,
    new_n10158_1, new_n10159, new_n10160, new_n10161, new_n10162,
    new_n10163, new_n10165_1, new_n10166, new_n10167, new_n10168,
    new_n10169, new_n10170, new_n10171, new_n10172, new_n10173, new_n10174,
    new_n10175, new_n10176, new_n10177, new_n10178, new_n10179, new_n10180,
    new_n10181, new_n10182, new_n10183, new_n10184, new_n10185, new_n10186,
    new_n10187, new_n10188, new_n10189, new_n10190, new_n10191, new_n10192,
    new_n10193, new_n10194, new_n10195, new_n10196, new_n10197, new_n10198,
    new_n10199, new_n10200, new_n10201_1, new_n10202, new_n10203,
    new_n10204, new_n10205, new_n10206, new_n10207, new_n10208, new_n10209,
    new_n10210, new_n10211, new_n10212, new_n10213, new_n10214, new_n10215,
    new_n10216, new_n10217, new_n10218, new_n10219, new_n10220, new_n10221,
    new_n10222, new_n10223, new_n10224, new_n10225, new_n10226, new_n10227,
    new_n10228, new_n10229, new_n10230, new_n10231, new_n10232, new_n10233,
    new_n10234, new_n10235, new_n10236_1, new_n10237, new_n10238,
    new_n10239_1, new_n10240, new_n10241, new_n10242, new_n10243,
    new_n10244_1, new_n10245, new_n10246, new_n10247, new_n10248,
    new_n10249, new_n10250_1, new_n10251, new_n10252, new_n10253,
    new_n10254, new_n10255, new_n10256, new_n10257, new_n10258, new_n10259,
    new_n10260, new_n10261_1, new_n10262_1, new_n10263, new_n10264,
    new_n10265, new_n10266, new_n10267, new_n10268, new_n10269, new_n10270,
    new_n10271, new_n10272, new_n10273, new_n10274, new_n10275_1,
    new_n10276, new_n10277, new_n10278, new_n10279, new_n10280, new_n10281,
    new_n10282, new_n10283, new_n10284, new_n10285, new_n10286,
    new_n10287_1, new_n10288, new_n10289, new_n10290, new_n10291,
    new_n10292, new_n10293, new_n10294, new_n10295_1, new_n10296,
    new_n10297, new_n10298, new_n10299, new_n10300, new_n10301, new_n10302,
    new_n10303, new_n10304, new_n10305, new_n10306, new_n10307, new_n10308,
    new_n10309, new_n10310, new_n10311, new_n10312, new_n10313, new_n10314,
    new_n10315, new_n10316, new_n10317, new_n10318, new_n10319, new_n10320,
    new_n10321_1, new_n10322, new_n10323, new_n10324, new_n10325,
    new_n10326_1, new_n10327_1, new_n10328, new_n10329, new_n10330_1,
    new_n10331, new_n10332, new_n10333, new_n10334, new_n10335, new_n10336,
    new_n10337, new_n10338, new_n10339, new_n10340_1, new_n10341,
    new_n10342, new_n10343, new_n10344, new_n10345_1, new_n10346,
    new_n10347, new_n10348, new_n10349, new_n10350, new_n10351, new_n10352,
    new_n10353, new_n10354, new_n10355, new_n10356_1, new_n10357,
    new_n10358, new_n10359, new_n10360, new_n10361, new_n10362, new_n10363,
    new_n10364, new_n10365, new_n10366, new_n10367, new_n10368, new_n10369,
    new_n10370, new_n10371, new_n10372_1, new_n10373, new_n10374,
    new_n10375, new_n10376, new_n10377, new_n10378, new_n10379, new_n10380,
    new_n10381, new_n10382, new_n10383, new_n10384, new_n10385_1,
    new_n10386, new_n10387_1, new_n10388_1, new_n10389, new_n10390_1,
    new_n10391, new_n10392, new_n10393, new_n10394, new_n10395, new_n10396,
    new_n10397, new_n10398, new_n10399, new_n10400, new_n10401, new_n10402,
    new_n10403, new_n10404_1, new_n10405_1, new_n10406, new_n10407,
    new_n10408, new_n10409_1, new_n10410, new_n10412, new_n10413,
    new_n10414, new_n10415, new_n10416, new_n10417, new_n10418, new_n10419,
    new_n10420_1, new_n10421, new_n10422, new_n10423, new_n10424,
    new_n10425, new_n10426, new_n10427, new_n10428, new_n10429, new_n10430,
    new_n10431, new_n10432_1, new_n10433, new_n10434, new_n10435,
    new_n10436, new_n10437, new_n10438, new_n10439, new_n10440, new_n10441,
    new_n10442, new_n10443, new_n10444, new_n10445, new_n10446, new_n10447,
    new_n10448, new_n10449, new_n10450, new_n10451, new_n10452, new_n10453,
    new_n10454, new_n10455, new_n10456, new_n10457, new_n10458, new_n10459,
    new_n10460, new_n10461, new_n10462, new_n10463, new_n10464, new_n10465,
    new_n10466, new_n10467, new_n10468, new_n10469, new_n10470, new_n10471,
    new_n10472, new_n10473, new_n10474, new_n10475, new_n10476, new_n10477,
    new_n10478, new_n10479, new_n10480, new_n10481, new_n10482, new_n10483,
    new_n10484_1, new_n10485, new_n10486, new_n10487, new_n10488,
    new_n10489_1, new_n10490, new_n10491, new_n10492, new_n10493,
    new_n10494, new_n10495, new_n10496, new_n10497, new_n10498, new_n10499,
    new_n10500, new_n10501, new_n10502, new_n10503, new_n10505, new_n10506,
    new_n10507, new_n10508, new_n10509, new_n10510, new_n10511, new_n10512,
    new_n10513, new_n10514_1, new_n10515, new_n10516, new_n10517,
    new_n10518, new_n10519, new_n10520, new_n10521, new_n10522, new_n10523,
    new_n10524, new_n10525_1, new_n10526, new_n10527, new_n10528,
    new_n10529, new_n10530, new_n10531, new_n10532, new_n10533, new_n10534,
    new_n10535, new_n10536, new_n10537, new_n10538, new_n10539,
    new_n10540_1, new_n10541, new_n10542, new_n10543, new_n10544,
    new_n10545, new_n10546, new_n10547, new_n10548, new_n10549, new_n10550,
    new_n10551, new_n10552, new_n10553, new_n10554, new_n10555, new_n10556,
    new_n10557, new_n10558, new_n10559, new_n10560, new_n10561_1,
    new_n10562, new_n10563, new_n10564_1, new_n10565, new_n10566,
    new_n10567, new_n10568, new_n10569, new_n10570, new_n10571, new_n10572,
    new_n10573, new_n10574, new_n10575, new_n10576, new_n10577_1,
    new_n10578, new_n10579, new_n10580, new_n10581, new_n10582, new_n10583,
    new_n10584, new_n10585, new_n10586, new_n10587, new_n10588_1,
    new_n10589, new_n10590, new_n10591, new_n10592, new_n10593_1,
    new_n10594, new_n10595_1, new_n10596, new_n10597, new_n10598,
    new_n10599, new_n10600, new_n10601, new_n10602, new_n10603, new_n10604,
    new_n10605, new_n10607, new_n10608, new_n10609, new_n10610,
    new_n10611_1, new_n10612, new_n10613, new_n10614_1, new_n10615,
    new_n10616, new_n10617_1, new_n10618, new_n10619, new_n10620,
    new_n10621, new_n10622, new_n10623, new_n10624, new_n10625, new_n10626,
    new_n10627, new_n10628_1, new_n10629, new_n10630, new_n10631,
    new_n10632, new_n10633, new_n10634, new_n10635, new_n10636, new_n10637,
    new_n10638, new_n10639, new_n10640, new_n10641, new_n10642, new_n10643,
    new_n10644, new_n10645, new_n10646, new_n10647_1, new_n10648,
    new_n10649, new_n10650_1, new_n10651, new_n10652, new_n10653_1,
    new_n10654, new_n10655, new_n10656, new_n10657, new_n10658, new_n10659,
    new_n10660, new_n10661, new_n10662, new_n10663, new_n10664, new_n10665,
    new_n10666, new_n10667, new_n10668, new_n10669, new_n10670, new_n10671,
    new_n10672, new_n10673, new_n10674, new_n10675, new_n10676, new_n10677,
    new_n10678, new_n10679, new_n10680, new_n10681, new_n10682, new_n10683,
    new_n10684, new_n10685, new_n10686, new_n10687, new_n10688, new_n10689,
    new_n10690, new_n10691, new_n10692_1, new_n10693, new_n10694_1,
    new_n10695, new_n10696, new_n10697, new_n10698, new_n10699, new_n10700,
    new_n10701_1, new_n10702, new_n10703, new_n10704, new_n10705,
    new_n10706, new_n10707, new_n10708, new_n10709, new_n10710_1,
    new_n10711, new_n10712_1, new_n10713, new_n10714, new_n10715,
    new_n10716, new_n10717, new_n10718, new_n10719, new_n10720, new_n10721,
    new_n10722, new_n10723, new_n10724, new_n10725, new_n10726, new_n10727,
    new_n10728, new_n10729, new_n10730, new_n10731, new_n10732, new_n10733,
    new_n10734, new_n10735, new_n10736, new_n10737, new_n10738,
    new_n10739_1, new_n10740, new_n10741, new_n10742, new_n10743,
    new_n10744, new_n10745, new_n10746, new_n10747, new_n10748, new_n10749,
    new_n10750, new_n10751, new_n10752, new_n10753, new_n10754, new_n10755,
    new_n10756_1, new_n10757, new_n10758, new_n10759, new_n10760,
    new_n10761, new_n10762, new_n10763_1, new_n10764, new_n10765,
    new_n10766, new_n10767, new_n10768, new_n10769, new_n10770, new_n10771,
    new_n10772, new_n10773, new_n10774, new_n10775_1, new_n10777,
    new_n10778, new_n10779, new_n10781, new_n10782, new_n10783, new_n10784,
    new_n10785, new_n10786, new_n10787, new_n10788, new_n10789, new_n10790,
    new_n10791, new_n10792_1, new_n10793, new_n10794, new_n10795,
    new_n10796, new_n10797, new_n10798, new_n10799, new_n10800, new_n10801,
    new_n10802, new_n10803, new_n10804, new_n10805, new_n10806, new_n10807,
    new_n10808, new_n10809, new_n10810, new_n10811, new_n10812, new_n10813,
    new_n10814, new_n10815, new_n10816, new_n10817_1, new_n10818,
    new_n10819, new_n10820, new_n10821, new_n10822, new_n10823, new_n10824,
    new_n10825, new_n10826, new_n10827, new_n10828, new_n10829, new_n10830,
    new_n10831, new_n10832, new_n10833, new_n10834_1, new_n10835,
    new_n10836, new_n10837, new_n10838, new_n10839, new_n10840, new_n10841,
    new_n10842, new_n10843, new_n10844, new_n10845, new_n10846, new_n10847,
    new_n10848, new_n10849, new_n10850, new_n10851_1, new_n10852,
    new_n10853, new_n10854, new_n10855, new_n10856, new_n10857, new_n10858,
    new_n10859, new_n10860, new_n10861, new_n10862, new_n10863, new_n10864,
    new_n10865, new_n10866, new_n10867, new_n10868, new_n10870, new_n10871,
    new_n10872, new_n10873, new_n10874_1, new_n10875, new_n10876,
    new_n10877, new_n10878, new_n10879, new_n10880, new_n10881, new_n10882,
    new_n10883, new_n10884, new_n10885, new_n10886, new_n10887, new_n10888,
    new_n10889, new_n10890, new_n10891, new_n10892, new_n10893, new_n10894,
    new_n10895, new_n10896, new_n10897, new_n10898, new_n10899, new_n10900,
    new_n10901, new_n10902, new_n10903, new_n10904, new_n10905, new_n10906,
    new_n10907, new_n10908, new_n10909, new_n10910, new_n10911, new_n10912,
    new_n10913, new_n10914, new_n10915, new_n10916, new_n10917, new_n10918,
    new_n10919, new_n10920, new_n10921, new_n10922, new_n10923,
    new_n10924_1, new_n10925, new_n10926, new_n10927, new_n10928,
    new_n10929, new_n10930, new_n10931, new_n10932, new_n10933, new_n10934,
    new_n10935, new_n10936, new_n10937, new_n10938, new_n10939, new_n10940,
    new_n10941, new_n10942, new_n10943_1, new_n10944, new_n10945,
    new_n10946, new_n10947, new_n10948, new_n10949, new_n10950, new_n10951,
    new_n10952, new_n10953, new_n10954, new_n10955, new_n10956, new_n10957,
    new_n10958, new_n10959, new_n10960, new_n10961_1, new_n10962,
    new_n10963, new_n10964, new_n10965, new_n10966, new_n10967, new_n10968,
    new_n10969, new_n10970, new_n10971, new_n10972, new_n10973, new_n10974,
    new_n10975, new_n10976, new_n10977, new_n10978, new_n10979, new_n10980,
    new_n10981, new_n10982, new_n10983, new_n10984, new_n10985, new_n10986,
    new_n10987, new_n10988, new_n10989, new_n10990, new_n10991, new_n10992,
    new_n10993, new_n10994, new_n10995, new_n10996, new_n10997, new_n10998,
    new_n10999, new_n11000, new_n11001, new_n11002, new_n11003, new_n11004,
    new_n11005_1, new_n11006, new_n11007, new_n11008, new_n11009,
    new_n11010, new_n11011_1, new_n11012, new_n11013, new_n11014,
    new_n11015, new_n11016, new_n11017, new_n11018, new_n11019, new_n11020,
    new_n11021, new_n11022, new_n11023_1, new_n11024, new_n11025_1,
    new_n11026, new_n11027, new_n11028, new_n11029, new_n11030, new_n11031,
    new_n11032, new_n11033, new_n11034, new_n11035, new_n11036, new_n11037,
    new_n11038, new_n11039, new_n11040, new_n11041, new_n11042, new_n11043,
    new_n11044_1, new_n11045, new_n11046, new_n11047, new_n11048,
    new_n11049, new_n11050, new_n11051, new_n11052, new_n11053, new_n11054,
    new_n11055, new_n11056_1, new_n11057, new_n11058, new_n11059,
    new_n11060, new_n11061, new_n11062, new_n11063_1, new_n11064,
    new_n11065, new_n11066, new_n11067, new_n11068, new_n11069, new_n11070,
    new_n11071, new_n11072, new_n11073, new_n11074, new_n11075, new_n11076,
    new_n11077, new_n11078_1, new_n11079, new_n11080_1, new_n11081,
    new_n11082, new_n11083, new_n11084, new_n11085, new_n11086, new_n11087,
    new_n11088, new_n11089, new_n11090, new_n11092, new_n11093,
    new_n11094_1, new_n11095, new_n11096, new_n11097, new_n11098,
    new_n11099, new_n11100, new_n11101_1, new_n11102, new_n11103_1,
    new_n11104, new_n11105, new_n11106, new_n11107, new_n11108, new_n11109,
    new_n11110, new_n11111, new_n11112, new_n11113, new_n11114, new_n11115,
    new_n11116, new_n11117, new_n11118, new_n11119, new_n11120_1,
    new_n11121_1, new_n11122, new_n11123, new_n11124, new_n11125,
    new_n11126, new_n11127_1, new_n11128, new_n11129, new_n11130,
    new_n11131, new_n11132_1, new_n11133, new_n11134_1, new_n11135,
    new_n11136, new_n11137, new_n11138_1, new_n11139, new_n11140,
    new_n11141, new_n11142, new_n11143, new_n11144, new_n11145, new_n11147,
    new_n11148, new_n11149, new_n11150, new_n11151, new_n11152, new_n11154,
    new_n11155, new_n11156, new_n11157, new_n11158, new_n11159, new_n11160,
    new_n11161, new_n11162, new_n11163, new_n11164, new_n11165, new_n11166,
    new_n11167, new_n11168, new_n11169, new_n11170, new_n11171, new_n11172,
    new_n11173, new_n11174, new_n11175, new_n11176, new_n11177, new_n11178,
    new_n11179, new_n11180, new_n11181, new_n11182_1, new_n11183,
    new_n11184_1, new_n11185, new_n11186, new_n11187, new_n11188,
    new_n11189, new_n11190, new_n11191, new_n11192_1, new_n11193,
    new_n11194, new_n11195, new_n11196, new_n11197, new_n11198, new_n11199,
    new_n11200, new_n11201_1, new_n11202, new_n11203, new_n11204,
    new_n11205, new_n11206, new_n11207, new_n11208, new_n11209, new_n11210,
    new_n11211, new_n11212, new_n11213, new_n11214, new_n11215, new_n11216,
    new_n11217, new_n11218, new_n11219, new_n11220_1, new_n11221,
    new_n11222, new_n11223_1, new_n11224, new_n11225, new_n11226,
    new_n11227, new_n11228, new_n11229, new_n11230, new_n11231, new_n11232,
    new_n11233, new_n11234_1, new_n11235, new_n11236, new_n11237,
    new_n11238, new_n11239, new_n11240, new_n11241, new_n11242, new_n11243,
    new_n11244, new_n11245_1, new_n11246, new_n11247, new_n11248,
    new_n11249, new_n11250, new_n11251, new_n11252, new_n11253, new_n11254,
    new_n11255, new_n11256, new_n11257, new_n11258, new_n11259, new_n11260,
    new_n11261_1, new_n11262, new_n11263, new_n11264, new_n11265,
    new_n11266_1, new_n11267, new_n11272, new_n11273_1, new_n11274,
    new_n11275_1, new_n11276, new_n11277, new_n11278, new_n11279,
    new_n11280, new_n11281, new_n11282, new_n11283, new_n11284, new_n11285,
    new_n11286, new_n11287, new_n11288, new_n11289, new_n11290_1,
    new_n11291, new_n11292, new_n11293, new_n11294, new_n11295, new_n11296,
    new_n11297, new_n11298, new_n11299, new_n11300, new_n11301,
    new_n11302_1, new_n11303, new_n11304, new_n11305, new_n11306,
    new_n11307, new_n11308, new_n11309, new_n11310, new_n11311, new_n11312,
    new_n11313_1, new_n11314, new_n11315, new_n11316, new_n11317,
    new_n11318, new_n11319, new_n11320, new_n11321, new_n11322, new_n11323,
    new_n11324, new_n11325_1, new_n11326_1, new_n11327, new_n11328,
    new_n11329, new_n11330_1, new_n11331, new_n11332, new_n11333,
    new_n11334, new_n11335, new_n11336, new_n11337, new_n11338, new_n11339,
    new_n11340, new_n11341, new_n11342, new_n11343, new_n11344, new_n11345,
    new_n11346, new_n11347_1, new_n11348_1, new_n11349, new_n11350,
    new_n11351, new_n11352_1, new_n11353, new_n11354, new_n11355,
    new_n11356_1, new_n11357, new_n11358, new_n11359, new_n11360,
    new_n11361, new_n11362, new_n11363, new_n11364, new_n11365, new_n11366,
    new_n11367, new_n11368, new_n11369, new_n11370, new_n11371, new_n11372,
    new_n11373, new_n11374, new_n11375_1, new_n11376, new_n11377,
    new_n11378, new_n11379_1, new_n11380, new_n11381, new_n11382,
    new_n11383, new_n11384, new_n11385, new_n11386_1, new_n11387,
    new_n11388, new_n11389, new_n11390, new_n11391_1, new_n11392,
    new_n11393, new_n11394, new_n11395, new_n11396, new_n11397,
    new_n11398_1, new_n11399, new_n11400, new_n11401, new_n11402,
    new_n11403_1, new_n11404, new_n11405, new_n11406, new_n11407,
    new_n11408, new_n11409, new_n11410, new_n11411, new_n11412, new_n11413,
    new_n11415, new_n11416, new_n11417, new_n11418, new_n11419_1,
    new_n11420, new_n11421, new_n11422, new_n11423, new_n11424_1,
    new_n11425, new_n11426, new_n11427, new_n11428, new_n11429, new_n11430,
    new_n11431, new_n11432, new_n11433, new_n11434, new_n11435, new_n11436,
    new_n11437, new_n11438, new_n11439_1, new_n11440, new_n11441,
    new_n11442, new_n11443, new_n11444, new_n11445, new_n11446, new_n11447,
    new_n11448, new_n11449, new_n11450, new_n11451, new_n11452, new_n11453,
    new_n11454, new_n11455_1, new_n11456, new_n11457, new_n11458,
    new_n11459, new_n11460, new_n11461, new_n11462_1, new_n11463,
    new_n11464, new_n11465, new_n11466, new_n11467, new_n11468, new_n11469,
    new_n11470_1, new_n11471, new_n11472_1, new_n11473_1, new_n11474,
    new_n11475, new_n11476, new_n11477, new_n11478, new_n11479_1,
    new_n11480, new_n11481_1, new_n11482, new_n11483, new_n11484,
    new_n11485, new_n11486_1, new_n11487, new_n11488, new_n11489,
    new_n11490, new_n11491, new_n11492, new_n11493, new_n11494, new_n11495,
    new_n11496_1, new_n11497, new_n11498, new_n11499, new_n11500,
    new_n11501, new_n11502, new_n11503_1, new_n11504, new_n11505,
    new_n11506_1, new_n11507, new_n11508, new_n11509, new_n11510,
    new_n11511, new_n11512, new_n11513, new_n11514, new_n11515_1,
    new_n11516, new_n11517, new_n11518, new_n11519, new_n11520, new_n11521,
    new_n11522, new_n11523, new_n11524, new_n11525, new_n11526, new_n11527,
    new_n11528, new_n11529, new_n11530, new_n11531, new_n11532, new_n11533,
    new_n11534, new_n11535, new_n11536, new_n11537, new_n11538_1,
    new_n11539, new_n11540, new_n11541, new_n11542, new_n11543, new_n11544,
    new_n11545, new_n11546, new_n11547, new_n11548_1, new_n11549,
    new_n11550, new_n11551, new_n11552, new_n11553, new_n11554, new_n11555,
    new_n11556, new_n11557, new_n11558, new_n11559, new_n11560, new_n11561,
    new_n11562, new_n11563, new_n11564_1, new_n11565, new_n11566_1,
    new_n11567, new_n11568, new_n11569, new_n11570, new_n11571, new_n11572,
    new_n11573, new_n11574, new_n11575, new_n11576, new_n11577, new_n11578,
    new_n11579_1, new_n11580_1, new_n11581, new_n11582, new_n11583,
    new_n11584, new_n11585, new_n11586, new_n11590, new_n11591_1,
    new_n11592, new_n11593, new_n11594, new_n11595, new_n11596, new_n11597,
    new_n11598, new_n11599, new_n11600, new_n11603, new_n11605, new_n11606,
    new_n11607_1, new_n11608, new_n11609, new_n11610, new_n11611,
    new_n11612, new_n11613, new_n11614, new_n11615_1, new_n11616,
    new_n11617, new_n11618, new_n11619, new_n11620, new_n11621, new_n11622,
    new_n11623, new_n11624, new_n11625, new_n11626, new_n11627, new_n11628,
    new_n11629, new_n11630_1, new_n11631, new_n11634, new_n11635,
    new_n11636, new_n11637, new_n11638, new_n11639, new_n11640, new_n11641,
    new_n11642, new_n11643, new_n11644, new_n11645, new_n11646,
    new_n11647_1, new_n11648, new_n11649, new_n11650, new_n11651,
    new_n11652, new_n11653, new_n11654, new_n11655, new_n11656, new_n11657,
    new_n11658, new_n11659, new_n11660, new_n11661, new_n11662, new_n11663,
    new_n11664, new_n11665, new_n11666, new_n11667_1, new_n11668,
    new_n11669, new_n11670, new_n11671, new_n11672, new_n11673,
    new_n11674_1, new_n11675, new_n11676, new_n11677, new_n11678,
    new_n11679, new_n11680, new_n11681, new_n11682_1, new_n11683,
    new_n11684, new_n11685, new_n11686, new_n11687, new_n11688, new_n11689,
    new_n11690, new_n11691, new_n11692, new_n11693, new_n11694, new_n11695,
    new_n11696, new_n11697, new_n11698, new_n11699, new_n11700, new_n11701,
    new_n11702, new_n11703, new_n11704, new_n11705, new_n11706, new_n11707,
    new_n11708, new_n11709, new_n11710_1, new_n11711, new_n11712_1,
    new_n11713, new_n11714, new_n11715, new_n11716, new_n11717, new_n11718,
    new_n11719, new_n11720, new_n11721, new_n11722, new_n11723,
    new_n11724_1, new_n11725, new_n11726, new_n11727, new_n11728,
    new_n11729, new_n11730, new_n11731, new_n11732, new_n11733, new_n11734,
    new_n11735, new_n11736_1, new_n11737, new_n11738, new_n11739,
    new_n11740, new_n11741_1, new_n11742, new_n11743, new_n11744,
    new_n11745, new_n11746, new_n11747, new_n11748, new_n11749_1,
    new_n11750, new_n11751, new_n11752, new_n11753, new_n11754, new_n11755,
    new_n11756, new_n11757, new_n11758, new_n11759, new_n11760, new_n11761,
    new_n11762, new_n11763, new_n11764, new_n11765, new_n11766, new_n11767,
    new_n11768, new_n11769, new_n11770_1, new_n11771_1, new_n11772,
    new_n11773, new_n11774, new_n11775_1, new_n11776, new_n11777,
    new_n11778, new_n11779, new_n11780, new_n11781, new_n11782, new_n11783,
    new_n11784, new_n11785, new_n11786, new_n11787, new_n11788, new_n11789,
    new_n11792, new_n11793, new_n11794, new_n11795, new_n11796, new_n11797,
    new_n11798, new_n11799, new_n11800, new_n11801, new_n11802, new_n11803,
    new_n11804, new_n11805, new_n11806, new_n11807, new_n11808, new_n11809,
    new_n11810, new_n11811, new_n11812, new_n11813, new_n11814, new_n11815,
    new_n11816, new_n11817, new_n11818_1, new_n11819, new_n11820,
    new_n11821, new_n11822, new_n11823, new_n11824, new_n11825, new_n11826,
    new_n11827, new_n11828, new_n11829, new_n11830, new_n11831, new_n11832,
    new_n11833, new_n11834, new_n11835, new_n11836, new_n11837_1,
    new_n11838, new_n11839, new_n11840, new_n11841_1, new_n11842_1,
    new_n11843_1, new_n11844, new_n11845, new_n11846, new_n11847,
    new_n11848, new_n11849, new_n11850, new_n11851, new_n11852, new_n11853,
    new_n11854, new_n11855, new_n11856, new_n11857, new_n11858, new_n11859,
    new_n11860, new_n11861, new_n11862, new_n11863, new_n11864, new_n11865,
    new_n11866, new_n11867, new_n11868, new_n11869, new_n11870, new_n11871,
    new_n11872, new_n11873, new_n11874, new_n11875, new_n11876, new_n11877,
    new_n11878, new_n11879, new_n11880, new_n11881, new_n11882, new_n11883,
    new_n11884, new_n11885, new_n11886, new_n11887, new_n11888, new_n11889,
    new_n11890, new_n11891, new_n11892, new_n11893, new_n11894, new_n11895,
    new_n11896, new_n11897, new_n11898_1, new_n11899, new_n11900,
    new_n11901, new_n11902, new_n11903, new_n11904, new_n11905_1,
    new_n11906, new_n11907, new_n11909, new_n11910, new_n11911, new_n11912,
    new_n11913, new_n11914, new_n11915, new_n11916, new_n11917, new_n11918,
    new_n11919, new_n11920, new_n11921, new_n11922, new_n11923, new_n11924,
    new_n11925, new_n11926_1, new_n11927, new_n11928, new_n11929,
    new_n11930, new_n11931, new_n11932, new_n11933, new_n11934, new_n11935,
    new_n11936, new_n11937, new_n11938, new_n11939, new_n11940, new_n11941,
    new_n11942, new_n11943, new_n11944, new_n11945, new_n11946, new_n11947,
    new_n11948, new_n11949, new_n11950, new_n11951, new_n11952, new_n11953,
    new_n11954, new_n11955, new_n11956, new_n11957, new_n11958, new_n11959,
    new_n11960, new_n11961, new_n11962, new_n11963, new_n11964,
    new_n11965_1, new_n11966, new_n11967, new_n11968, new_n11969,
    new_n11970, new_n11971, new_n11972, new_n11973, new_n11974, new_n11975,
    new_n11976, new_n11977, new_n11978, new_n11979, new_n11980_1,
    new_n11981, new_n11982, new_n11983, new_n11984, new_n11985, new_n11986,
    new_n11987, new_n11988, new_n11989, new_n11990, new_n11991, new_n11992,
    new_n11993, new_n11994, new_n11995, new_n11996, new_n11997, new_n11998,
    new_n11999, new_n12000_1, new_n12001, new_n12002, new_n12003_1,
    new_n12004, new_n12005, new_n12006, new_n12007, new_n12008, new_n12009,
    new_n12010, new_n12011_1, new_n12012, new_n12013, new_n12014,
    new_n12016, new_n12017, new_n12018, new_n12019, new_n12020, new_n12021,
    new_n12022, new_n12023, new_n12024, new_n12025, new_n12026, new_n12027,
    new_n12028, new_n12029, new_n12030, new_n12031, new_n12032, new_n12033,
    new_n12034, new_n12035, new_n12036, new_n12037, new_n12038, new_n12039,
    new_n12040, new_n12041, new_n12045, new_n12046, new_n12047, new_n12048,
    new_n12049, new_n12050, new_n12051, new_n12052, new_n12053, new_n12054,
    new_n12055, new_n12056, new_n12057, new_n12058, new_n12059, new_n12060,
    new_n12061, new_n12062, new_n12063, new_n12064, new_n12065, new_n12066,
    new_n12067, new_n12068, new_n12069, new_n12070, new_n12071,
    new_n12072_1, new_n12073, new_n12074, new_n12075, new_n12076,
    new_n12077, new_n12078, new_n12079, new_n12080, new_n12081, new_n12082,
    new_n12083, new_n12084, new_n12085, new_n12086, new_n12087, new_n12088,
    new_n12089, new_n12090, new_n12091, new_n12092, new_n12093, new_n12094,
    new_n12095, new_n12096, new_n12097, new_n12098, new_n12099, new_n12100,
    new_n12101, new_n12102, new_n12103, new_n12104, new_n12105, new_n12106,
    new_n12107, new_n12110, new_n12111, new_n12112, new_n12113_1,
    new_n12114, new_n12115, new_n12116, new_n12117, new_n12118, new_n12119,
    new_n12120, new_n12121_1, new_n12122, new_n12123, new_n12124,
    new_n12125, new_n12126, new_n12127, new_n12128, new_n12129, new_n12130,
    new_n12131_1, new_n12132, new_n12133, new_n12134, new_n12135,
    new_n12136, new_n12137, new_n12138, new_n12139, new_n12140, new_n12141,
    new_n12142, new_n12143, new_n12144, new_n12145, new_n12146_1,
    new_n12147, new_n12148, new_n12149, new_n12150, new_n12151,
    new_n12152_1, new_n12153_1, new_n12154, new_n12155, new_n12156,
    new_n12157_1, new_n12158_1, new_n12159, new_n12160, new_n12161_1,
    new_n12162, new_n12163, new_n12164, new_n12165, new_n12166, new_n12167,
    new_n12168, new_n12169, new_n12170, new_n12171, new_n12172, new_n12173,
    new_n12174, new_n12175, new_n12176, new_n12177, new_n12178,
    new_n12179_1, new_n12180, new_n12181, new_n12182, new_n12183,
    new_n12184, new_n12185, new_n12186, new_n12187, new_n12188, new_n12189,
    new_n12190, new_n12191, new_n12192_1, new_n12193, new_n12194,
    new_n12195, new_n12196, new_n12197, new_n12198, new_n12199, new_n12200,
    new_n12201, new_n12202, new_n12203, new_n12204, new_n12205, new_n12206,
    new_n12207, new_n12208, new_n12209_1, new_n12210, new_n12211,
    new_n12212, new_n12213, new_n12214, new_n12215, new_n12216, new_n12217,
    new_n12218, new_n12219, new_n12220, new_n12221, new_n12222,
    new_n12223_1, new_n12224, new_n12225_1, new_n12226, new_n12227,
    new_n12228_1, new_n12229, new_n12230, new_n12231, new_n12232,
    new_n12233, new_n12234, new_n12235_1, new_n12236, new_n12237,
    new_n12238, new_n12239, new_n12240, new_n12241, new_n12242, new_n12243,
    new_n12244, new_n12245, new_n12246, new_n12247, new_n12248, new_n12249,
    new_n12250, new_n12251, new_n12252, new_n12253, new_n12254, new_n12255,
    new_n12256, new_n12257, new_n12258, new_n12259, new_n12260, new_n12261,
    new_n12262, new_n12263, new_n12264, new_n12265, new_n12266, new_n12267,
    new_n12268, new_n12269, new_n12270, new_n12271, new_n12272, new_n12273,
    new_n12274, new_n12275, new_n12276, new_n12277, new_n12278, new_n12279,
    new_n12280, new_n12281, new_n12282, new_n12283, new_n12284, new_n12285,
    new_n12286, new_n12287, new_n12288, new_n12289, new_n12290, new_n12291,
    new_n12292, new_n12293, new_n12294, new_n12295, new_n12296, new_n12297,
    new_n12298, new_n12299, new_n12300, new_n12301, new_n12302_1,
    new_n12303, new_n12304_1, new_n12305, new_n12306, new_n12307,
    new_n12308, new_n12309, new_n12310, new_n12311, new_n12312, new_n12313,
    new_n12314, new_n12315_1, new_n12316, new_n12317, new_n12318,
    new_n12319, new_n12320, new_n12321, new_n12324_1, new_n12325_1,
    new_n12326, new_n12327, new_n12328, new_n12329_1, new_n12330_1,
    new_n12331, new_n12332, new_n12333, new_n12334, new_n12335, new_n12336,
    new_n12337, new_n12338, new_n12339, new_n12340, new_n12341_1,
    new_n12342, new_n12343, new_n12344, new_n12345, new_n12346_1,
    new_n12347, new_n12348, new_n12349_1, new_n12350, new_n12351,
    new_n12352, new_n12353, new_n12355, new_n12356, new_n12357, new_n12358,
    new_n12359, new_n12360, new_n12361, new_n12362, new_n12363,
    new_n12364_1, new_n12365, new_n12366, new_n12367, new_n12368,
    new_n12369, new_n12370, new_n12371, new_n12372, new_n12373, new_n12374,
    new_n12375, new_n12376, new_n12377, new_n12378, new_n12379,
    new_n12380_1, new_n12381, new_n12382, new_n12383_1, new_n12384_1,
    new_n12385, new_n12386, new_n12387, new_n12388, new_n12389, new_n12390,
    new_n12391, new_n12392, new_n12393, new_n12394, new_n12395, new_n12396,
    new_n12397_1, new_n12398_1, new_n12399, new_n12400, new_n12401,
    new_n12402, new_n12403, new_n12404, new_n12405, new_n12406, new_n12407,
    new_n12408_1, new_n12409, new_n12410, new_n12411, new_n12412,
    new_n12413, new_n12414, new_n12415, new_n12416, new_n12417, new_n12418,
    new_n12419, new_n12420, new_n12421, new_n12422, new_n12423, new_n12424,
    new_n12425, new_n12426, new_n12427, new_n12428, new_n12429, new_n12430,
    new_n12431, new_n12432, new_n12433, new_n12434, new_n12435, new_n12436,
    new_n12437, new_n12438, new_n12439, new_n12440, new_n12441, new_n12442,
    new_n12443, new_n12444, new_n12445, new_n12446_1, new_n12447,
    new_n12448, new_n12449_1, new_n12450, new_n12451, new_n12452,
    new_n12453, new_n12454, new_n12455, new_n12456, new_n12457, new_n12458,
    new_n12459, new_n12460, new_n12461_1, new_n12462_1, new_n12463,
    new_n12464, new_n12465, new_n12466, new_n12467_1, new_n12468,
    new_n12469_1, new_n12470, new_n12471, new_n12472, new_n12473,
    new_n12474, new_n12475, new_n12476, new_n12477, new_n12478, new_n12479,
    new_n12480, new_n12481, new_n12482, new_n12483, new_n12484, new_n12485,
    new_n12486, new_n12487, new_n12488, new_n12489, new_n12490, new_n12491,
    new_n12492, new_n12493, new_n12494, new_n12495_1, new_n12496,
    new_n12497, new_n12498, new_n12499, new_n12500, new_n12501, new_n12502,
    new_n12503, new_n12504, new_n12505, new_n12506, new_n12507_1,
    new_n12508, new_n12509, new_n12510, new_n12511, new_n12512, new_n12513,
    new_n12514, new_n12515_1, new_n12516_1, new_n12517, new_n12518,
    new_n12519, new_n12520, new_n12521, new_n12522, new_n12523, new_n12524,
    new_n12525, new_n12526, new_n12527, new_n12528, new_n12529, new_n12530,
    new_n12531, new_n12532, new_n12533, new_n12534, new_n12535, new_n12536,
    new_n12537, new_n12538, new_n12539, new_n12540_1, new_n12541,
    new_n12542, new_n12543, new_n12544, new_n12545_1, new_n12546_1,
    new_n12547, new_n12548, new_n12549, new_n12550, new_n12551,
    new_n12552_1, new_n12553, new_n12554, new_n12555, new_n12556,
    new_n12557, new_n12558, new_n12559, new_n12560, new_n12561,
    new_n12562_1, new_n12563, new_n12564, new_n12565, new_n12566_1,
    new_n12567, new_n12568, new_n12569_1, new_n12570, new_n12571,
    new_n12572, new_n12573, new_n12574, new_n12575, new_n12576, new_n12577,
    new_n12578, new_n12579, new_n12580, new_n12581, new_n12582, new_n12583,
    new_n12584, new_n12585, new_n12586, new_n12587_1, new_n12588,
    new_n12589, new_n12590, new_n12591, new_n12592, new_n12593_1,
    new_n12594, new_n12595, new_n12596, new_n12597, new_n12598, new_n12599,
    new_n12600, new_n12601, new_n12602, new_n12603, new_n12604, new_n12605,
    new_n12606, new_n12607_1, new_n12608, new_n12609, new_n12610,
    new_n12611, new_n12612, new_n12613, new_n12614, new_n12615, new_n12616,
    new_n12617, new_n12618, new_n12619, new_n12620_1, new_n12621_1,
    new_n12622, new_n12623, new_n12624, new_n12625, new_n12626_1,
    new_n12627, new_n12628, new_n12629, new_n12630, new_n12631, new_n12632,
    new_n12633, new_n12634, new_n12635, new_n12636, new_n12637, new_n12638,
    new_n12639, new_n12640, new_n12641, new_n12642, new_n12643, new_n12644,
    new_n12645, new_n12646, new_n12647, new_n12648, new_n12649,
    new_n12650_1, new_n12651, new_n12652, new_n12653, new_n12654_1,
    new_n12655, new_n12656, new_n12657_1, new_n12658, new_n12659,
    new_n12660, new_n12661, new_n12662, new_n12663, new_n12664,
    new_n12665_1, new_n12666, new_n12667, new_n12670_1, new_n12671,
    new_n12672, new_n12673, new_n12674, new_n12675, new_n12676, new_n12677,
    new_n12678, new_n12679, new_n12680, new_n12681, new_n12682, new_n12683,
    new_n12684, new_n12685, new_n12686, new_n12687, new_n12688, new_n12689,
    new_n12690, new_n12691, new_n12692, new_n12693, new_n12694, new_n12695,
    new_n12696, new_n12697, new_n12698, new_n12699, new_n12700, new_n12701,
    new_n12702_1, new_n12703, new_n12704, new_n12705, new_n12706,
    new_n12707_1, new_n12708, new_n12709, new_n12710, new_n12711,
    new_n12712, new_n12713, new_n12714, new_n12715, new_n12716, new_n12717,
    new_n12718, new_n12719, new_n12720, new_n12721, new_n12722, new_n12723,
    new_n12724, new_n12725_1, new_n12726, new_n12727_1, new_n12728,
    new_n12729, new_n12730, new_n12731, new_n12732, new_n12737, new_n12738,
    new_n12739, new_n12740_1, new_n12741, new_n12742_1, new_n12743,
    new_n12744, new_n12745, new_n12746_1, new_n12747, new_n12748,
    new_n12749, new_n12750, new_n12754, new_n12755, new_n12756_1,
    new_n12757, new_n12758, new_n12759, new_n12760, new_n12761, new_n12762,
    new_n12763, new_n12764, new_n12765, new_n12766, new_n12767, new_n12768,
    new_n12769, new_n12770, new_n12771, new_n12772, new_n12773, new_n12774,
    new_n12778, new_n12779, new_n12780, new_n12781, new_n12782,
    new_n12783_1, new_n12784, new_n12785, new_n12786, new_n12787,
    new_n12788, new_n12789, new_n12790, new_n12791, new_n12792, new_n12793,
    new_n12794, new_n12795, new_n12796, new_n12797, new_n12798, new_n12799,
    new_n12800, new_n12801_1, new_n12802, new_n12803, new_n12804,
    new_n12805, new_n12806, new_n12808, new_n12809, new_n12810,
    new_n12811_1, new_n12812_1, new_n12813, new_n12814, new_n12815,
    new_n12816_1, new_n12817, new_n12818, new_n12819, new_n12820,
    new_n12821_1, new_n12822, new_n12823, new_n12824, new_n12825,
    new_n12826, new_n12827, new_n12828, new_n12829, new_n12830, new_n12831,
    new_n12832, new_n12833, new_n12834, new_n12835, new_n12836, new_n12840,
    new_n12841, new_n12842, new_n12843_1, new_n12844, new_n12845,
    new_n12846, new_n12847, new_n12848, new_n12849, new_n12850, new_n12851,
    new_n12852, new_n12853, new_n12854, new_n12855, new_n12856, new_n12857,
    new_n12858, new_n12859, new_n12860, new_n12861_1, new_n12862,
    new_n12863, new_n12864_1, new_n12865_1, new_n12866, new_n12867,
    new_n12868, new_n12869, new_n12870_1, new_n12871_1, new_n12872,
    new_n12873_1, new_n12874, new_n12875_1, new_n12876, new_n12877,
    new_n12878, new_n12881, new_n12882, new_n12883, new_n12884, new_n12885,
    new_n12886, new_n12887, new_n12888, new_n12889, new_n12890, new_n12891,
    new_n12892_1, new_n12893, new_n12894, new_n12895, new_n12896,
    new_n12897, new_n12898, new_n12899, new_n12900_1, new_n12901,
    new_n12902, new_n12903, new_n12904_1, new_n12905, new_n12906,
    new_n12907, new_n12908, new_n12909, new_n12910, new_n12911, new_n12912,
    new_n12913, new_n12914, new_n12915, new_n12916, new_n12917_1,
    new_n12918, new_n12919, new_n12920, new_n12921, new_n12922, new_n12923,
    new_n12924, new_n12925, new_n12926, new_n12927, new_n12928, new_n12929,
    new_n12930, new_n12931, new_n12932, new_n12933, new_n12934, new_n12935,
    new_n12936, new_n12937, new_n12938, new_n12939, new_n12940,
    new_n12941_1, new_n12942_1, new_n12943, new_n12944, new_n12945,
    new_n12946, new_n12947, new_n12948, new_n12949, new_n12950, new_n12951,
    new_n12952, new_n12953, new_n12954, new_n12955, new_n12956_1,
    new_n12957, new_n12958, new_n12959, new_n12960, new_n12961, new_n12962,
    new_n12963, new_n12964, new_n12965, new_n12966, new_n12967, new_n12968,
    new_n12969, new_n12970, new_n12971, new_n12972, new_n12973, new_n12974,
    new_n12975, new_n12976, new_n12977, new_n12978_1, new_n12979,
    new_n12980_1, new_n12981, new_n12982, new_n12983, new_n12984,
    new_n12985_1, new_n12986, new_n12987_1, new_n12988, new_n12989,
    new_n12991, new_n12992_1, new_n12993, new_n12994, new_n12995,
    new_n12996, new_n12997, new_n12998, new_n12999, new_n13000, new_n13001,
    new_n13002, new_n13003, new_n13004, new_n13005_1, new_n13006,
    new_n13007, new_n13008, new_n13009, new_n13010, new_n13011, new_n13012,
    new_n13013, new_n13014, new_n13015, new_n13016, new_n13017, new_n13018,
    new_n13019, new_n13020, new_n13021, new_n13022, new_n13023, new_n13024,
    new_n13025, new_n13026_1, new_n13027, new_n13028, new_n13029,
    new_n13030, new_n13031, new_n13032, new_n13033, new_n13034, new_n13035,
    new_n13036, new_n13037, new_n13038, new_n13039, new_n13040, new_n13041,
    new_n13042, new_n13043_1, new_n13044_1, new_n13045, new_n13046,
    new_n13047, new_n13048_1, new_n13049, new_n13050, new_n13051,
    new_n13052, new_n13053, new_n13054_1, new_n13055, new_n13056,
    new_n13057, new_n13058, new_n13059, new_n13060, new_n13061, new_n13062,
    new_n13063, new_n13064, new_n13065, new_n13066, new_n13067, new_n13068,
    new_n13069, new_n13070, new_n13071, new_n13072, new_n13073,
    new_n13074_1, new_n13075, new_n13076, new_n13077, new_n13078,
    new_n13079, new_n13080, new_n13081, new_n13082_1, new_n13083,
    new_n13084, new_n13085, new_n13086, new_n13087, new_n13088, new_n13089,
    new_n13090, new_n13091, new_n13092, new_n13093, new_n13094, new_n13095,
    new_n13097, new_n13098, new_n13099, new_n13100, new_n13101, new_n13102,
    new_n13103, new_n13104, new_n13105, new_n13106, new_n13107, new_n13108,
    new_n13109, new_n13110_1, new_n13111, new_n13112, new_n13113,
    new_n13114, new_n13115, new_n13116_1, new_n13117, new_n13118,
    new_n13119, new_n13120, new_n13121, new_n13122_1, new_n13123,
    new_n13124, new_n13125, new_n13126, new_n13127, new_n13128, new_n13129,
    new_n13130, new_n13131, new_n13132, new_n13133, new_n13134, new_n13135,
    new_n13136, new_n13137_1, new_n13138, new_n13139, new_n13142,
    new_n13143, new_n13144_1, new_n13145, new_n13146, new_n13147,
    new_n13148, new_n13149, new_n13150, new_n13151, new_n13153, new_n13154,
    new_n13155, new_n13156, new_n13157, new_n13158, new_n13159, new_n13160,
    new_n13161, new_n13162, new_n13163, new_n13164, new_n13165, new_n13166,
    new_n13167, new_n13168_1, new_n13169, new_n13170, new_n13171,
    new_n13172, new_n13173, new_n13174, new_n13175, new_n13176, new_n13177,
    new_n13178, new_n13179, new_n13180, new_n13181, new_n13182, new_n13183,
    new_n13184, new_n13185, new_n13186, new_n13187, new_n13188, new_n13189,
    new_n13190_1, new_n13191, new_n13192, new_n13193, new_n13194,
    new_n13195, new_n13196, new_n13197, new_n13198_1, new_n13199_1,
    new_n13200, new_n13201, new_n13202, new_n13203, new_n13204_1,
    new_n13205, new_n13206, new_n13207, new_n13208, new_n13209_1,
    new_n13210, new_n13211, new_n13212, new_n13213, new_n13214, new_n13215,
    new_n13216, new_n13217, new_n13218, new_n13219, new_n13220, new_n13221,
    new_n13222, new_n13223, new_n13224, new_n13225, new_n13226, new_n13227,
    new_n13228, new_n13229, new_n13230, new_n13231, new_n13232, new_n13233,
    new_n13234, new_n13235, new_n13236, new_n13237, new_n13238, new_n13239,
    new_n13240, new_n13241, new_n13242, new_n13243, new_n13244, new_n13245,
    new_n13246, new_n13247, new_n13248, new_n13249, new_n13250, new_n13251,
    new_n13252, new_n13253, new_n13254, new_n13255, new_n13256, new_n13257,
    new_n13258, new_n13259, new_n13260, new_n13261, new_n13262,
    new_n13263_1, new_n13264, new_n13265, new_n13266, new_n13267,
    new_n13268, new_n13269, new_n13270_1, new_n13271, new_n13272,
    new_n13273_1, new_n13274, new_n13275, new_n13276, new_n13277,
    new_n13278, new_n13279, new_n13280, new_n13281, new_n13282, new_n13283,
    new_n13284, new_n13285_1, new_n13286, new_n13287, new_n13288,
    new_n13289, new_n13290, new_n13291, new_n13292, new_n13293, new_n13294,
    new_n13295, new_n13296, new_n13297, new_n13298, new_n13299, new_n13300,
    new_n13301, new_n13302, new_n13303, new_n13304, new_n13305, new_n13306,
    new_n13307, new_n13308, new_n13309, new_n13310, new_n13313, new_n13314,
    new_n13315, new_n13316, new_n13317, new_n13318, new_n13319_1,
    new_n13320, new_n13321, new_n13322, new_n13323, new_n13324, new_n13325,
    new_n13326, new_n13327, new_n13328, new_n13329, new_n13330, new_n13331,
    new_n13332, new_n13333_1, new_n13334, new_n13335, new_n13336,
    new_n13337, new_n13338_1, new_n13339, new_n13340, new_n13341,
    new_n13342, new_n13343, new_n13344, new_n13345, new_n13346, new_n13347,
    new_n13348, new_n13349, new_n13350, new_n13351, new_n13352, new_n13353,
    new_n13354, new_n13355, new_n13356, new_n13357, new_n13358, new_n13359,
    new_n13360, new_n13361, new_n13362, new_n13363, new_n13364, new_n13365,
    new_n13366, new_n13367_1, new_n13368, new_n13369, new_n13370,
    new_n13371, new_n13372, new_n13373, new_n13374, new_n13375, new_n13376,
    new_n13377, new_n13378, new_n13379, new_n13380, new_n13381, new_n13382,
    new_n13383, new_n13384, new_n13385, new_n13386, new_n13387, new_n13388,
    new_n13389, new_n13390, new_n13392, new_n13393, new_n13394, new_n13395,
    new_n13396, new_n13397, new_n13398, new_n13399, new_n13402, new_n13403,
    new_n13404, new_n13405, new_n13406, new_n13407_1, new_n13408,
    new_n13409_1, new_n13410, new_n13411, new_n13412, new_n13413,
    new_n13414, new_n13415, new_n13416, new_n13417, new_n13418,
    new_n13419_1, new_n13420, new_n13421, new_n13422, new_n13423,
    new_n13424_1, new_n13425, new_n13426, new_n13427, new_n13428,
    new_n13429, new_n13430, new_n13431, new_n13432, new_n13433, new_n13434,
    new_n13435, new_n13436, new_n13437, new_n13438, new_n13439, new_n13440,
    new_n13441, new_n13442, new_n13443, new_n13444, new_n13445, new_n13446,
    new_n13447, new_n13448, new_n13449, new_n13450, new_n13451, new_n13452,
    new_n13453_1, new_n13454, new_n13455, new_n13456_1, new_n13457_1,
    new_n13458, new_n13459, new_n13460_1, new_n13461, new_n13462,
    new_n13463, new_n13464, new_n13465, new_n13466, new_n13467, new_n13468,
    new_n13469, new_n13470, new_n13471, new_n13472, new_n13473, new_n13474,
    new_n13475, new_n13476, new_n13477_1, new_n13478, new_n13479,
    new_n13480, new_n13481, new_n13482, new_n13484_1, new_n13485,
    new_n13486_1, new_n13487_1, new_n13488, new_n13489, new_n13490_1,
    new_n13491, new_n13492, new_n13493, new_n13494_1, new_n13495,
    new_n13496, new_n13497, new_n13498, new_n13499, new_n13500_1,
    new_n13501_1, new_n13502, new_n13503, new_n13504, new_n13505,
    new_n13506_1, new_n13507, new_n13508, new_n13509, new_n13510,
    new_n13511, new_n13512, new_n13513, new_n13514, new_n13515, new_n13516,
    new_n13517, new_n13518, new_n13519, new_n13520, new_n13521, new_n13522,
    new_n13523, new_n13524, new_n13525, new_n13526, new_n13527, new_n13528,
    new_n13529, new_n13530, new_n13531, new_n13532, new_n13533, new_n13534,
    new_n13535, new_n13536, new_n13537, new_n13538, new_n13539, new_n13540,
    new_n13541, new_n13542, new_n13543, new_n13544, new_n13545, new_n13546,
    new_n13547, new_n13548_1, new_n13549_1, new_n13550, new_n13551_1,
    new_n13552, new_n13553, new_n13554, new_n13555, new_n13556, new_n13557,
    new_n13558, new_n13559, new_n13560, new_n13561, new_n13562, new_n13563,
    new_n13564, new_n13565, new_n13566, new_n13567, new_n13568, new_n13569,
    new_n13570, new_n13571, new_n13572, new_n13573, new_n13574, new_n13575,
    new_n13576, new_n13577, new_n13578, new_n13579, new_n13580, new_n13581,
    new_n13582, new_n13583, new_n13584, new_n13585, new_n13586, new_n13587,
    new_n13588, new_n13589, new_n13590, new_n13591, new_n13592, new_n13593,
    new_n13594, new_n13595, new_n13598, new_n13599, new_n13600, new_n13601,
    new_n13602_1, new_n13603, new_n13604, new_n13605, new_n13606,
    new_n13607, new_n13608, new_n13609, new_n13610, new_n13611, new_n13612,
    new_n13613, new_n13614, new_n13615, new_n13616, new_n13617, new_n13618,
    new_n13619, new_n13620, new_n13621, new_n13622, new_n13623, new_n13624,
    new_n13625, new_n13626_1, new_n13627, new_n13628, new_n13629,
    new_n13630, new_n13631, new_n13632, new_n13633, new_n13634, new_n13635,
    new_n13636, new_n13637, new_n13638, new_n13639, new_n13640, new_n13643,
    new_n13644, new_n13645, new_n13646, new_n13647, new_n13648, new_n13649,
    new_n13650, new_n13651, new_n13652, new_n13653, new_n13654, new_n13655,
    new_n13656, new_n13657, new_n13658, new_n13659, new_n13660, new_n13661,
    new_n13662, new_n13663, new_n13664, new_n13665, new_n13666, new_n13667,
    new_n13668_1, new_n13669, new_n13670, new_n13671, new_n13672,
    new_n13673, new_n13674, new_n13675, new_n13676, new_n13677_1,
    new_n13678, new_n13679, new_n13680, new_n13681, new_n13682,
    new_n13683_1, new_n13684, new_n13685, new_n13686, new_n13687,
    new_n13688, new_n13689, new_n13690, new_n13691, new_n13692, new_n13693,
    new_n13694, new_n13695, new_n13696, new_n13697, new_n13698, new_n13699,
    new_n13700, new_n13701, new_n13702, new_n13703, new_n13704, new_n13705,
    new_n13706, new_n13707, new_n13708_1, new_n13709, new_n13710_1,
    new_n13711, new_n13712, new_n13713, new_n13714_1, new_n13715,
    new_n13716, new_n13717, new_n13718, new_n13719_1, new_n13720,
    new_n13721, new_n13722_1, new_n13723, new_n13724, new_n13725,
    new_n13726, new_n13727, new_n13728, new_n13729, new_n13730, new_n13731,
    new_n13732, new_n13733, new_n13734, new_n13735, new_n13736, new_n13737,
    new_n13738, new_n13739, new_n13740, new_n13741, new_n13742, new_n13743,
    new_n13744, new_n13745, new_n13746, new_n13747, new_n13748, new_n13749,
    new_n13750, new_n13751, new_n13752, new_n13753, new_n13754_1,
    new_n13755, new_n13756, new_n13757, new_n13758, new_n13759, new_n13760,
    new_n13761, new_n13762, new_n13763, new_n13764_1, new_n13765,
    new_n13766, new_n13767, new_n13768, new_n13769, new_n13770, new_n13771,
    new_n13772, new_n13773, new_n13774, new_n13775_1, new_n13776,
    new_n13777, new_n13778, new_n13779, new_n13780, new_n13781_1,
    new_n13783_1, new_n13784, new_n13785, new_n13786, new_n13787,
    new_n13788, new_n13789, new_n13790, new_n13791, new_n13792, new_n13793,
    new_n13794, new_n13795, new_n13796, new_n13797, new_n13798_1,
    new_n13799, new_n13800, new_n13801, new_n13802, new_n13803, new_n13804,
    new_n13805, new_n13806, new_n13807, new_n13808, new_n13810, new_n13811,
    new_n13812, new_n13813, new_n13814, new_n13815, new_n13816, new_n13817,
    new_n13818, new_n13819, new_n13820, new_n13821, new_n13822, new_n13823,
    new_n13824, new_n13825, new_n13826, new_n13827, new_n13828, new_n13829,
    new_n13830, new_n13831, new_n13832, new_n13833, new_n13834,
    new_n13835_1, new_n13836, new_n13837, new_n13838, new_n13839,
    new_n13840, new_n13841, new_n13842, new_n13843, new_n13844, new_n13845,
    new_n13846, new_n13847, new_n13848, new_n13849, new_n13850_1,
    new_n13851_1, new_n13852, new_n13853, new_n13854, new_n13855,
    new_n13856, new_n13857, new_n13858, new_n13859, new_n13860, new_n13861,
    new_n13862, new_n13863, new_n13864, new_n13865, new_n13866, new_n13867,
    new_n13868, new_n13869, new_n13870, new_n13871, new_n13872, new_n13873,
    new_n13874, new_n13875, new_n13876, new_n13877, new_n13878, new_n13879,
    new_n13880, new_n13881, new_n13882, new_n13883, new_n13884, new_n13885,
    new_n13886, new_n13887, new_n13888, new_n13889, new_n13890, new_n13891,
    new_n13892, new_n13893, new_n13894, new_n13895, new_n13896, new_n13897,
    new_n13898, new_n13899, new_n13900, new_n13901, new_n13902, new_n13903,
    new_n13904, new_n13905, new_n13906, new_n13907, new_n13908, new_n13909,
    new_n13910, new_n13911, new_n13912_1, new_n13913, new_n13914_1,
    new_n13915, new_n13916, new_n13917, new_n13918, new_n13919, new_n13920,
    new_n13921, new_n13922_1, new_n13923_1, new_n13924, new_n13925,
    new_n13926, new_n13927, new_n13928, new_n13929, new_n13930, new_n13931,
    new_n13932, new_n13933, new_n13934, new_n13935, new_n13936, new_n13937,
    new_n13938, new_n13939, new_n13940, new_n13941, new_n13942, new_n13943,
    new_n13944, new_n13945, new_n13946, new_n13947, new_n13948, new_n13949,
    new_n13950, new_n13951_1, new_n13952, new_n13953, new_n13954,
    new_n13955, new_n13956, new_n13957, new_n13958, new_n13959, new_n13960,
    new_n13961, new_n13962, new_n13963, new_n13964, new_n13965, new_n13966,
    new_n13967, new_n13968, new_n13969, new_n13970, new_n13971, new_n13972,
    new_n13973, new_n13974, new_n13975, new_n13976, new_n13977, new_n13978,
    new_n13979, new_n13980, new_n13981, new_n13982, new_n13983, new_n13984,
    new_n13985, new_n13986, new_n13987, new_n13988, new_n13989, new_n13990,
    new_n13991, new_n13992, new_n13993, new_n13994, new_n13996, new_n13997,
    new_n13998, new_n13999, new_n14000, new_n14001, new_n14002, new_n14003,
    new_n14004_1, new_n14005, new_n14006, new_n14007, new_n14008,
    new_n14009, new_n14010, new_n14011, new_n14012, new_n14013, new_n14014,
    new_n14015, new_n14016, new_n14017, new_n14018, new_n14019, new_n14020,
    new_n14021, new_n14022, new_n14023, new_n14024, new_n14025, new_n14026,
    new_n14027, new_n14028, new_n14029, new_n14030, new_n14031, new_n14032,
    new_n14033, new_n14034, new_n14035, new_n14036_1, new_n14037,
    new_n14038, new_n14039, new_n14040, new_n14041, new_n14042, new_n14043,
    new_n14044, new_n14045, new_n14046, new_n14047, new_n14048, new_n14049,
    new_n14050, new_n14051, new_n14052, new_n14053, new_n14054, new_n14055,
    new_n14056, new_n14057, new_n14058, new_n14059_1, new_n14060,
    new_n14061, new_n14062, new_n14063, new_n14064, new_n14065, new_n14066,
    new_n14067, new_n14068, new_n14069, new_n14070, new_n14071_1,
    new_n14072, new_n14073, new_n14074, new_n14075, new_n14076, new_n14077,
    new_n14078, new_n14079, new_n14080, new_n14081_1, new_n14082,
    new_n14083, new_n14084, new_n14085, new_n14086, new_n14087, new_n14088,
    new_n14089, new_n14090_1, new_n14091, new_n14092, new_n14093,
    new_n14094, new_n14095_1, new_n14096, new_n14097, new_n14098,
    new_n14099, new_n14100, new_n14101, new_n14102, new_n14103, new_n14104,
    new_n14105, new_n14106, new_n14107_1, new_n14108, new_n14109,
    new_n14110, new_n14111, new_n14112, new_n14113, new_n14114, new_n14115,
    new_n14116, new_n14117, new_n14118, new_n14119, new_n14120,
    new_n14121_1, new_n14122, new_n14123, new_n14124, new_n14125,
    new_n14126_1, new_n14127, new_n14128, new_n14129, new_n14130_1,
    new_n14131, new_n14132, new_n14133, new_n14134, new_n14135,
    new_n14136_1, new_n14137, new_n14138, new_n14139, new_n14140,
    new_n14141, new_n14142, new_n14143, new_n14144, new_n14145, new_n14146,
    new_n14147_1, new_n14148_1, new_n14149, new_n14150, new_n14151,
    new_n14152, new_n14153, new_n14154, new_n14155, new_n14156, new_n14157,
    new_n14158, new_n14159, new_n14160, new_n14161, new_n14162, new_n14164,
    new_n14165, new_n14166, new_n14167, new_n14168, new_n14169, new_n14170,
    new_n14171, new_n14172, new_n14173, new_n14174_1, new_n14175,
    new_n14176, new_n14177, new_n14178, new_n14179, new_n14180, new_n14181,
    new_n14182, new_n14183, new_n14184, new_n14185, new_n14186, new_n14187,
    new_n14188, new_n14189, new_n14190_1, new_n14191, new_n14192,
    new_n14193, new_n14194, new_n14195, new_n14196, new_n14197, new_n14198,
    new_n14199, new_n14200, new_n14201, new_n14202, new_n14203, new_n14204,
    new_n14205, new_n14206, new_n14207, new_n14208, new_n14209, new_n14210,
    new_n14211_1, new_n14212, new_n14213, new_n14214, new_n14215,
    new_n14216, new_n14217, new_n14218, new_n14219, new_n14220, new_n14221,
    new_n14222_1, new_n14223, new_n14224, new_n14225, new_n14226,
    new_n14227, new_n14228, new_n14229, new_n14230_1, new_n14231,
    new_n14232, new_n14233, new_n14234, new_n14235, new_n14236, new_n14237,
    new_n14238, new_n14239, new_n14240, new_n14241, new_n14242, new_n14243,
    new_n14244, new_n14245, new_n14246, new_n14247, new_n14248, new_n14249,
    new_n14250, new_n14251, new_n14252, new_n14253, new_n14254, new_n14255,
    new_n14256, new_n14257, new_n14258, new_n14259, new_n14260, new_n14261,
    new_n14262, new_n14263, new_n14264, new_n14265, new_n14266,
    new_n14267_1, new_n14268, new_n14269, new_n14270, new_n14271_1,
    new_n14272, new_n14273, new_n14274, new_n14275_1, new_n14276,
    new_n14277_1, new_n14278, new_n14279, new_n14280, new_n14281,
    new_n14282, new_n14283, new_n14284, new_n14285, new_n14286, new_n14287,
    new_n14288, new_n14289, new_n14290, new_n14291, new_n14292, new_n14293,
    new_n14294_1, new_n14295, new_n14296, new_n14297, new_n14298,
    new_n14299, new_n14300, new_n14301, new_n14302, new_n14303, new_n14304,
    new_n14305, new_n14306, new_n14307, new_n14309, new_n14310_1,
    new_n14311, new_n14312, new_n14313, new_n14314, new_n14315, new_n14316,
    new_n14317, new_n14318, new_n14319, new_n14320, new_n14321, new_n14322,
    new_n14323_1, new_n14324, new_n14325, new_n14326_1, new_n14327,
    new_n14328, new_n14329, new_n14330, new_n14331, new_n14332, new_n14333,
    new_n14334, new_n14335, new_n14336, new_n14337, new_n14338, new_n14339,
    new_n14340, new_n14341, new_n14342_1, new_n14343, new_n14344,
    new_n14345_1, new_n14346, new_n14347, new_n14348, new_n14349,
    new_n14350, new_n14351, new_n14352, new_n14353_1, new_n14354,
    new_n14355, new_n14356, new_n14357, new_n14358, new_n14359, new_n14360,
    new_n14361, new_n14362, new_n14363, new_n14364_1, new_n14365,
    new_n14366, new_n14367, new_n14368, new_n14369, new_n14370, new_n14371,
    new_n14372, new_n14373, new_n14374, new_n14375_1, new_n14376,
    new_n14377, new_n14378, new_n14379, new_n14380, new_n14381, new_n14382,
    new_n14383, new_n14384, new_n14385, new_n14386, new_n14387, new_n14388,
    new_n14389, new_n14390, new_n14391, new_n14392, new_n14393, new_n14394,
    new_n14395, new_n14396, new_n14397, new_n14398, new_n14399, new_n14400,
    new_n14401, new_n14402, new_n14403, new_n14404, new_n14405, new_n14406,
    new_n14407, new_n14408, new_n14409, new_n14410, new_n14411,
    new_n14412_1, new_n14413, new_n14415, new_n14416, new_n14417,
    new_n14418, new_n14419, new_n14420, new_n14421, new_n14422, new_n14423,
    new_n14424, new_n14425, new_n14426, new_n14427, new_n14428, new_n14429,
    new_n14430, new_n14431, new_n14432, new_n14433, new_n14434, new_n14435,
    new_n14436, new_n14437, new_n14438, new_n14439, new_n14440_1,
    new_n14441, new_n14442, new_n14443, new_n14444, new_n14445, new_n14446,
    new_n14447, new_n14448, new_n14449, new_n14450, new_n14451, new_n14452,
    new_n14453, new_n14454, new_n14455, new_n14456, new_n14457_1,
    new_n14458, new_n14459, new_n14460, new_n14461, new_n14462, new_n14463,
    new_n14464_1, new_n14465, new_n14466, new_n14467, new_n14468,
    new_n14469, new_n14470, new_n14471_1, new_n14472, new_n14473,
    new_n14474, new_n14475_1, new_n14476, new_n14477, new_n14478,
    new_n14481, new_n14482, new_n14483, new_n14484, new_n14485, new_n14486,
    new_n14487, new_n14488, new_n14489, new_n14490, new_n14491, new_n14492,
    new_n14493, new_n14494, new_n14495, new_n14496, new_n14497, new_n14498,
    new_n14499, new_n14500, new_n14501, new_n14502, new_n14503, new_n14504,
    new_n14505, new_n14506, new_n14507, new_n14508, new_n14509,
    new_n14510_1, new_n14511, new_n14512, new_n14513, new_n14514,
    new_n14515, new_n14516, new_n14517, new_n14518, new_n14519, new_n14520,
    new_n14521, new_n14522, new_n14523, new_n14524, new_n14525, new_n14526,
    new_n14527, new_n14528, new_n14529, new_n14530, new_n14531, new_n14532,
    new_n14533, new_n14534, new_n14535, new_n14536, new_n14537, new_n14538,
    new_n14539, new_n14540, new_n14541_1, new_n14542, new_n14543,
    new_n14544, new_n14545, new_n14546_1, new_n14547_1, new_n14548,
    new_n14549, new_n14550, new_n14551, new_n14552, new_n14553, new_n14554,
    new_n14555, new_n14556, new_n14557, new_n14558, new_n14559, new_n14560,
    new_n14561, new_n14562, new_n14563, new_n14564, new_n14565, new_n14566,
    new_n14567, new_n14568, new_n14569, new_n14570_1, new_n14571,
    new_n14572, new_n14573, new_n14574, new_n14575_1, new_n14576_1,
    new_n14577, new_n14578, new_n14579, new_n14580, new_n14581, new_n14582,
    new_n14583, new_n14584, new_n14585, new_n14586, new_n14587, new_n14588,
    new_n14589, new_n14590, new_n14591, new_n14592, new_n14593_1,
    new_n14594, new_n14595, new_n14596, new_n14597, new_n14598, new_n14599,
    new_n14600, new_n14601, new_n14602, new_n14603_1, new_n14604,
    new_n14605, new_n14606, new_n14607, new_n14608, new_n14609, new_n14610,
    new_n14611, new_n14612, new_n14613, new_n14614, new_n14615, new_n14616,
    new_n14617, new_n14618, new_n14619, new_n14620, new_n14621, new_n14622,
    new_n14623, new_n14624, new_n14625, new_n14626, new_n14628, new_n14629,
    new_n14630, new_n14631, new_n14632, new_n14633_1, new_n14634,
    new_n14635, new_n14636_1, new_n14637, new_n14638, new_n14639,
    new_n14640, new_n14641, new_n14642, new_n14643, new_n14644, new_n14645,
    new_n14646, new_n14647, new_n14648, new_n14649, new_n14650, new_n14651,
    new_n14652, new_n14653, new_n14654, new_n14655, new_n14656, new_n14657,
    new_n14658, new_n14659, new_n14660, new_n14661, new_n14662, new_n14663,
    new_n14664, new_n14665, new_n14666, new_n14667, new_n14668, new_n14669,
    new_n14670, new_n14671, new_n14672, new_n14673, new_n14674, new_n14675,
    new_n14676, new_n14677, new_n14678, new_n14679, new_n14680_1,
    new_n14681, new_n14682, new_n14683, new_n14684_1, new_n14685,
    new_n14686, new_n14687, new_n14688, new_n14689, new_n14690, new_n14691,
    new_n14692_1, new_n14693, new_n14694, new_n14695, new_n14696,
    new_n14697, new_n14698, new_n14699, new_n14700, new_n14701_1,
    new_n14702_1, new_n14703, new_n14704_1, new_n14705, new_n14706,
    new_n14707, new_n14708, new_n14709, new_n14710, new_n14711, new_n14712,
    new_n14713, new_n14714, new_n14715, new_n14716, new_n14717, new_n14718,
    new_n14719, new_n14720, new_n14721, new_n14722, new_n14723, new_n14724,
    new_n14725, new_n14726, new_n14727, new_n14728, new_n14729, new_n14730,
    new_n14731, new_n14732, new_n14733, new_n14734_1, new_n14740,
    new_n14743, new_n14744, new_n14745, new_n14747, new_n14748, new_n14749,
    new_n14750, new_n14751, new_n14752, new_n14753, new_n14754, new_n14755,
    new_n14756, new_n14757, new_n14758, new_n14759, new_n14760, new_n14761,
    new_n14762, new_n14763_1, new_n14764, new_n14765, new_n14766,
    new_n14767, new_n14768, new_n14769, new_n14770, new_n14771,
    new_n14772_1, new_n14773, new_n14774, new_n14775, new_n14776,
    new_n14777, new_n14780, new_n14781, new_n14782, new_n14783, new_n14784,
    new_n14785, new_n14786, new_n14787, new_n14788, new_n14789,
    new_n14790_1, new_n14791, new_n14792, new_n14793, new_n14794,
    new_n14795, new_n14796, new_n14797, new_n14798, new_n14799, new_n14800,
    new_n14801_1, new_n14802, new_n14803, new_n14804, new_n14805,
    new_n14806, new_n14807, new_n14808, new_n14809, new_n14810, new_n14811,
    new_n14812, new_n14813, new_n14814, new_n14815, new_n14816, new_n14817,
    new_n14818, new_n14819_1, new_n14820, new_n14821, new_n14822,
    new_n14823, new_n14824, new_n14825, new_n14826_1, new_n14827_1,
    new_n14828, new_n14829, new_n14830, new_n14831, new_n14832, new_n14833,
    new_n14834, new_n14835, new_n14836, new_n14837, new_n14838,
    new_n14839_1, new_n14840, new_n14841, new_n14842, new_n14843,
    new_n14844, new_n14845, new_n14846, new_n14847, new_n14853, new_n14854,
    new_n14855, new_n14856, new_n14857, new_n14858, new_n14859, new_n14860,
    new_n14861, new_n14862, new_n14863, new_n14864, new_n14865, new_n14866,
    new_n14867, new_n14868, new_n14869, new_n14870, new_n14871, new_n14872,
    new_n14873, new_n14874, new_n14875, new_n14876, new_n14877, new_n14878,
    new_n14879, new_n14880, new_n14881, new_n14882, new_n14883, new_n14884,
    new_n14885, new_n14886, new_n14887, new_n14888, new_n14889, new_n14890,
    new_n14891_1, new_n14892, new_n14893, new_n14894, new_n14895,
    new_n14896, new_n14897, new_n14898, new_n14899_1, new_n14900,
    new_n14901, new_n14902, new_n14903, new_n14904, new_n14905, new_n14906,
    new_n14907, new_n14908, new_n14909, new_n14910, new_n14911, new_n14912,
    new_n14913, new_n14914, new_n14915, new_n14916, new_n14917, new_n14918,
    new_n14919, new_n14920, new_n14921, new_n14922, new_n14923, new_n14924,
    new_n14925, new_n14926, new_n14927, new_n14928, new_n14929, new_n14930,
    new_n14931_1, new_n14932, new_n14933, new_n14934, new_n14935,
    new_n14936, new_n14937, new_n14938, new_n14939, new_n14940, new_n14941,
    new_n14942, new_n14943, new_n14944_1, new_n14945, new_n14946,
    new_n14947, new_n14948, new_n14949, new_n14950, new_n14951, new_n14952,
    new_n14953, new_n14954_1, new_n14955, new_n14956, new_n14957,
    new_n14958, new_n14959, new_n14960, new_n14961, new_n14962, new_n14963,
    new_n14964, new_n14965, new_n14966, new_n14967, new_n14968, new_n14969,
    new_n14970, new_n14971, new_n14972, new_n14973, new_n14974, new_n14975,
    new_n14976, new_n14977_1, new_n14978, new_n14979, new_n14982,
    new_n14983, new_n14984, new_n14985, new_n14986, new_n14987, new_n14988,
    new_n14989_1, new_n14990, new_n14991, new_n14992, new_n14993,
    new_n14994, new_n14995, new_n14996, new_n14997, new_n14998, new_n14999,
    new_n15000, new_n15001, new_n15002_1, new_n15003, new_n15004_1,
    new_n15005, new_n15006, new_n15007, new_n15008, new_n15009, new_n15010,
    new_n15011_1, new_n15012, new_n15013, new_n15014, new_n15015,
    new_n15016, new_n15017, new_n15018, new_n15019_1, new_n15020,
    new_n15021, new_n15022, new_n15023, new_n15024, new_n15025, new_n15026,
    new_n15027, new_n15028, new_n15029, new_n15030, new_n15031_1,
    new_n15032, new_n15033_1, new_n15034, new_n15035, new_n15036,
    new_n15037, new_n15038, new_n15039, new_n15040, new_n15041, new_n15042,
    new_n15044, new_n15045, new_n15046, new_n15047, new_n15048, new_n15049,
    new_n15050, new_n15051, new_n15052_1, new_n15053_1, new_n15054,
    new_n15055, new_n15056, new_n15057, new_n15058, new_n15059, new_n15060,
    new_n15061, new_n15062, new_n15063, new_n15064, new_n15065, new_n15066,
    new_n15067, new_n15068, new_n15069, new_n15070, new_n15071, new_n15072,
    new_n15073, new_n15074, new_n15075, new_n15076, new_n15079, new_n15080,
    new_n15081, new_n15082_1, new_n15083, new_n15084, new_n15085,
    new_n15086, new_n15087, new_n15088, new_n15089, new_n15090, new_n15091,
    new_n15092, new_n15093, new_n15094_1, new_n15095, new_n15096,
    new_n15097, new_n15098, new_n15099, new_n15100, new_n15101, new_n15102,
    new_n15103, new_n15104, new_n15105, new_n15106, new_n15107, new_n15108,
    new_n15109, new_n15110, new_n15111, new_n15112, new_n15113, new_n15114,
    new_n15115, new_n15116, new_n15117, new_n15118_1, new_n15119,
    new_n15121, new_n15122, new_n15123, new_n15124, new_n15125, new_n15126,
    new_n15127, new_n15128_1, new_n15129, new_n15130, new_n15131,
    new_n15132, new_n15133, new_n15134, new_n15135, new_n15136, new_n15137,
    new_n15138, new_n15139_1, new_n15140, new_n15141, new_n15142,
    new_n15143, new_n15144, new_n15145_1, new_n15146_1, new_n15147,
    new_n15148, new_n15149, new_n15150, new_n15151, new_n15152, new_n15153,
    new_n15154, new_n15155, new_n15156, new_n15157, new_n15158, new_n15159,
    new_n15161, new_n15162, new_n15163, new_n15164, new_n15165_1,
    new_n15166, new_n15167_1, new_n15168, new_n15169, new_n15170,
    new_n15171, new_n15172, new_n15173, new_n15174, new_n15175,
    new_n15176_1, new_n15177, new_n15178, new_n15179, new_n15180_1,
    new_n15181, new_n15182_1, new_n15183, new_n15184, new_n15185,
    new_n15186, new_n15187, new_n15188, new_n15189, new_n15190, new_n15191,
    new_n15192, new_n15193, new_n15194, new_n15195, new_n15196, new_n15197,
    new_n15198, new_n15199, new_n15200, new_n15201, new_n15202, new_n15203,
    new_n15204, new_n15205_1, new_n15206, new_n15207, new_n15208,
    new_n15209, new_n15210, new_n15211, new_n15212, new_n15213, new_n15214,
    new_n15215, new_n15216, new_n15217, new_n15218, new_n15219, new_n15220,
    new_n15221, new_n15222, new_n15223, new_n15224, new_n15225, new_n15226,
    new_n15227, new_n15228, new_n15229, new_n15230_1, new_n15231,
    new_n15232, new_n15233, new_n15234, new_n15235, new_n15236, new_n15237,
    new_n15238, new_n15239, new_n15240, new_n15241_1, new_n15242,
    new_n15243, new_n15244, new_n15245, new_n15246, new_n15247, new_n15248,
    new_n15249, new_n15250, new_n15251, new_n15252, new_n15253, new_n15254,
    new_n15255_1, new_n15256, new_n15257, new_n15258_1, new_n15259,
    new_n15260, new_n15261, new_n15262, new_n15263, new_n15264, new_n15265,
    new_n15266, new_n15267, new_n15268, new_n15269, new_n15270,
    new_n15271_1, new_n15272, new_n15273, new_n15274, new_n15275_1,
    new_n15276, new_n15277, new_n15278, new_n15279, new_n15280, new_n15281,
    new_n15282, new_n15283, new_n15284, new_n15285, new_n15286, new_n15287,
    new_n15288, new_n15289_1, new_n15290, new_n15291, new_n15292,
    new_n15293, new_n15294, new_n15295, new_n15296, new_n15297, new_n15298,
    new_n15299, new_n15300_1, new_n15301, new_n15302, new_n15303,
    new_n15304, new_n15305, new_n15306, new_n15307_1, new_n15308,
    new_n15309, new_n15310, new_n15311, new_n15312, new_n15313, new_n15314,
    new_n15315, new_n15316, new_n15317, new_n15318, new_n15319, new_n15320,
    new_n15321, new_n15322, new_n15323, new_n15324, new_n15325, new_n15326,
    new_n15327_1, new_n15328, new_n15329, new_n15330, new_n15331,
    new_n15332_1, new_n15333, new_n15334, new_n15335, new_n15336,
    new_n15337, new_n15338, new_n15341, new_n15344, new_n15345_1,
    new_n15346, new_n15347, new_n15348, new_n15349, new_n15350, new_n15351,
    new_n15352, new_n15353_1, new_n15354, new_n15355, new_n15356,
    new_n15357, new_n15360, new_n15361, new_n15362, new_n15363, new_n15364,
    new_n15365, new_n15366_1, new_n15367, new_n15368, new_n15369,
    new_n15370, new_n15371, new_n15372, new_n15373, new_n15374, new_n15375,
    new_n15376, new_n15377, new_n15378_1, new_n15379, new_n15380,
    new_n15381, new_n15382_1, new_n15383, new_n15384, new_n15385,
    new_n15386, new_n15387, new_n15388, new_n15389, new_n15390, new_n15391,
    new_n15392, new_n15393, new_n15394, new_n15395, new_n15396, new_n15397,
    new_n15398, new_n15399, new_n15400, new_n15401, new_n15402, new_n15403,
    new_n15404, new_n15405, new_n15406, new_n15407_1, new_n15408,
    new_n15409, new_n15410, new_n15411, new_n15412, new_n15413, new_n15414,
    new_n15415, new_n15416, new_n15417, new_n15418, new_n15419, new_n15420,
    new_n15421, new_n15422, new_n15423, new_n15424_1, new_n15425,
    new_n15426, new_n15427, new_n15428_1, new_n15429, new_n15430,
    new_n15431, new_n15432, new_n15433, new_n15434, new_n15435_1,
    new_n15436, new_n15437, new_n15438_1, new_n15439, new_n15440,
    new_n15441, new_n15442, new_n15443, new_n15444, new_n15445, new_n15446,
    new_n15447, new_n15448, new_n15449, new_n15450, new_n15451, new_n15452,
    new_n15453, new_n15454, new_n15455, new_n15458, new_n15459, new_n15460,
    new_n15461, new_n15462, new_n15463, new_n15464, new_n15465_1,
    new_n15466, new_n15467_1, new_n15468, new_n15469, new_n15470_1,
    new_n15471, new_n15472, new_n15473, new_n15474, new_n15475, new_n15476,
    new_n15477_1, new_n15478, new_n15479, new_n15480, new_n15482,
    new_n15483, new_n15484, new_n15485, new_n15486, new_n15487, new_n15488,
    new_n15489, new_n15490_1, new_n15491, new_n15492, new_n15493,
    new_n15494, new_n15495, new_n15496_1, new_n15497, new_n15498,
    new_n15499, new_n15500, new_n15501_1, new_n15502, new_n15505,
    new_n15506_1, new_n15507, new_n15508_1, new_n15509, new_n15510,
    new_n15511, new_n15512, new_n15513, new_n15514, new_n15515, new_n15516,
    new_n15517, new_n15518, new_n15519, new_n15520, new_n15521, new_n15522,
    new_n15523, new_n15524, new_n15525, new_n15526, new_n15527, new_n15528,
    new_n15529, new_n15530, new_n15531, new_n15532, new_n15533, new_n15534,
    new_n15535, new_n15536, new_n15537, new_n15538, new_n15539_1,
    new_n15540, new_n15541, new_n15543, new_n15544, new_n15545,
    new_n15546_1, new_n15547, new_n15548, new_n15549, new_n15550,
    new_n15551, new_n15552, new_n15553, new_n15554, new_n15555_1,
    new_n15556, new_n15557, new_n15558_1, new_n15559_1, new_n15560,
    new_n15561, new_n15562, new_n15563, new_n15564, new_n15565, new_n15566,
    new_n15567, new_n15568, new_n15569, new_n15570_1, new_n15571,
    new_n15572, new_n15573_1, new_n15574, new_n15575, new_n15576,
    new_n15577, new_n15578, new_n15579, new_n15580, new_n15581, new_n15582,
    new_n15583, new_n15584, new_n15585, new_n15586, new_n15587,
    new_n15588_1, new_n15589, new_n15590_1, new_n15591, new_n15592,
    new_n15593, new_n15594, new_n15595, new_n15596, new_n15597,
    new_n15598_1, new_n15599, new_n15600, new_n15601, new_n15602_1,
    new_n15603, new_n15604, new_n15605, new_n15606, new_n15607, new_n15608,
    new_n15609, new_n15610, new_n15611, new_n15612, new_n15613,
    new_n15614_1, new_n15615, new_n15616, new_n15617, new_n15618,
    new_n15619, new_n15620, new_n15621, new_n15622, new_n15623, new_n15624,
    new_n15625, new_n15626, new_n15627, new_n15628, new_n15629, new_n15630,
    new_n15631, new_n15632, new_n15633, new_n15634, new_n15635,
    new_n15636_1, new_n15637, new_n15638, new_n15639, new_n15640,
    new_n15641, new_n15642, new_n15643, new_n15644, new_n15645, new_n15646,
    new_n15647, new_n15648, new_n15649, new_n15650, new_n15651,
    new_n15652_1, new_n15653, new_n15654, new_n15655, new_n15656,
    new_n15657, new_n15658, new_n15659, new_n15660, new_n15661,
    new_n15662_1, new_n15663, new_n15664, new_n15665, new_n15666,
    new_n15667, new_n15668, new_n15669, new_n15670, new_n15671, new_n15672,
    new_n15673, new_n15674, new_n15675, new_n15676, new_n15677, new_n15678,
    new_n15679, new_n15680, new_n15681, new_n15682, new_n15683, new_n15684,
    new_n15685, new_n15686, new_n15687, new_n15688, new_n15689, new_n15690,
    new_n15691, new_n15692, new_n15693, new_n15694, new_n15695, new_n15696,
    new_n15697, new_n15698, new_n15699, new_n15700, new_n15701, new_n15702,
    new_n15703, new_n15704, new_n15705, new_n15706, new_n15707, new_n15708,
    new_n15709, new_n15710, new_n15711, new_n15712, new_n15713, new_n15714,
    new_n15715, new_n15717, new_n15718, new_n15719, new_n15720, new_n15721,
    new_n15722, new_n15723, new_n15724, new_n15725, new_n15726, new_n15727,
    new_n15728, new_n15729, new_n15730, new_n15731, new_n15732, new_n15733,
    new_n15734, new_n15735, new_n15736, new_n15737, new_n15738, new_n15739,
    new_n15740, new_n15741, new_n15742, new_n15743_1, new_n15744,
    new_n15745, new_n15746, new_n15747, new_n15748, new_n15749_1,
    new_n15750, new_n15751, new_n15752, new_n15753, new_n15754, new_n15755,
    new_n15756, new_n15757, new_n15758, new_n15759, new_n15760,
    new_n15761_1, new_n15762_1, new_n15763, new_n15764, new_n15765,
    new_n15766_1, new_n15767, new_n15768, new_n15769, new_n15770,
    new_n15771, new_n15772, new_n15773, new_n15774, new_n15775, new_n15776,
    new_n15777, new_n15778, new_n15779, new_n15780_1, new_n15781,
    new_n15782, new_n15783, new_n15784, new_n15785, new_n15786, new_n15787,
    new_n15788, new_n15789, new_n15790, new_n15791, new_n15792,
    new_n15793_1, new_n15794, new_n15795, new_n15796, new_n15797,
    new_n15798, new_n15799, new_n15800, new_n15801, new_n15802, new_n15803,
    new_n15804, new_n15805, new_n15806, new_n15807, new_n15808, new_n15809,
    new_n15810, new_n15811, new_n15812_1, new_n15813, new_n15814,
    new_n15815_1, new_n15816_1, new_n15817, new_n15818, new_n15821,
    new_n15822, new_n15823, new_n15824, new_n15825, new_n15826, new_n15827,
    new_n15828, new_n15829, new_n15830, new_n15831_1, new_n15832,
    new_n15833, new_n15834, new_n15835, new_n15836, new_n15837, new_n15838,
    new_n15839, new_n15840, new_n15841, new_n15842, new_n15843, new_n15844,
    new_n15845, new_n15846_1, new_n15847, new_n15848, new_n15849,
    new_n15850, new_n15851, new_n15852, new_n15853, new_n15854, new_n15855,
    new_n15856, new_n15857, new_n15858, new_n15859_1, new_n15860,
    new_n15861, new_n15862, new_n15863, new_n15864, new_n15865, new_n15866,
    new_n15867, new_n15868, new_n15869_1, new_n15870, new_n15871,
    new_n15872, new_n15873, new_n15874, new_n15875, new_n15876, new_n15877,
    new_n15878, new_n15879, new_n15880, new_n15881, new_n15882, new_n15883,
    new_n15884_1, new_n15885_1, new_n15886, new_n15887, new_n15888,
    new_n15889_1, new_n15890, new_n15891, new_n15892, new_n15893,
    new_n15894, new_n15895, new_n15896, new_n15897, new_n15898, new_n15899,
    new_n15900, new_n15901, new_n15902, new_n15903, new_n15904, new_n15905,
    new_n15906, new_n15907, new_n15908, new_n15909, new_n15910, new_n15911,
    new_n15912, new_n15913, new_n15914, new_n15915, new_n15916,
    new_n15917_1, new_n15918_1, new_n15919, new_n15920, new_n15921,
    new_n15922_1, new_n15923, new_n15925, new_n15926, new_n15927,
    new_n15928, new_n15929, new_n15930, new_n15931, new_n15932, new_n15933,
    new_n15934, new_n15935, new_n15936_1, new_n15937, new_n15938,
    new_n15939, new_n15940, new_n15941, new_n15942, new_n15943, new_n15944,
    new_n15945, new_n15946, new_n15947_1, new_n15948, new_n15949,
    new_n15950, new_n15951, new_n15952, new_n15953, new_n15954, new_n15955,
    new_n15956_1, new_n15957, new_n15958_1, new_n15959, new_n15960,
    new_n15961, new_n15962, new_n15963, new_n15964, new_n15965, new_n15966,
    new_n15967_1, new_n15968, new_n15969, new_n15970, new_n15971,
    new_n15972, new_n15973, new_n15974, new_n15975, new_n15977, new_n15978,
    new_n15979_1, new_n15980, new_n15981, new_n15982, new_n15983,
    new_n15984, new_n15985, new_n15986_1, new_n15987, new_n15988,
    new_n15989, new_n15990, new_n15991, new_n15992, new_n15993, new_n15994,
    new_n15995, new_n15996, new_n15997, new_n15998, new_n16001, new_n16002,
    new_n16003, new_n16004, new_n16005, new_n16006, new_n16007, new_n16008,
    new_n16009, new_n16010, new_n16011, new_n16012, new_n16013_1,
    new_n16014, new_n16015, new_n16016, new_n16017, new_n16018, new_n16019,
    new_n16020, new_n16021, new_n16022, new_n16023, new_n16024, new_n16025,
    new_n16026, new_n16027, new_n16028, new_n16029_1, new_n16030,
    new_n16031, new_n16032, new_n16033, new_n16034, new_n16035, new_n16036,
    new_n16037, new_n16038, new_n16039, new_n16040, new_n16041, new_n16042,
    new_n16043, new_n16044, new_n16045, new_n16046, new_n16047, new_n16048,
    new_n16049, new_n16050, new_n16051, new_n16052, new_n16053, new_n16054,
    new_n16055, new_n16056, new_n16057, new_n16058, new_n16059,
    new_n16060_1, new_n16061, new_n16062_1, new_n16063, new_n16064,
    new_n16065, new_n16066, new_n16067, new_n16068_1, new_n16069,
    new_n16070, new_n16071, new_n16072, new_n16073, new_n16074, new_n16075,
    new_n16076, new_n16077, new_n16081, new_n16082, new_n16083, new_n16084,
    new_n16085, new_n16086, new_n16087, new_n16088, new_n16089, new_n16090,
    new_n16091, new_n16095, new_n16096, new_n16097, new_n16098_1,
    new_n16099, new_n16100, new_n16101, new_n16102, new_n16103, new_n16104,
    new_n16105, new_n16106, new_n16107, new_n16108, new_n16109,
    new_n16110_1, new_n16111, new_n16112, new_n16113, new_n16114,
    new_n16115, new_n16116, new_n16117, new_n16118, new_n16119, new_n16122,
    new_n16123, new_n16124, new_n16125, new_n16126, new_n16127, new_n16128,
    new_n16129, new_n16130, new_n16131, new_n16132, new_n16133, new_n16134,
    new_n16135, new_n16136, new_n16137, new_n16138, new_n16139, new_n16140,
    new_n16141, new_n16142_1, new_n16143, new_n16144, new_n16145,
    new_n16146, new_n16147, new_n16148, new_n16149, new_n16150, new_n16151,
    new_n16152, new_n16153, new_n16154, new_n16155, new_n16156, new_n16157,
    new_n16158_1, new_n16159, new_n16160, new_n16161, new_n16162,
    new_n16163, new_n16164, new_n16165, new_n16166, new_n16167_1,
    new_n16168, new_n16169, new_n16170, new_n16171, new_n16172, new_n16173,
    new_n16174, new_n16175, new_n16176, new_n16177, new_n16178, new_n16179,
    new_n16180, new_n16181, new_n16182, new_n16183, new_n16184,
    new_n16185_1, new_n16186, new_n16187, new_n16188, new_n16189,
    new_n16190, new_n16191, new_n16192, new_n16193, new_n16194, new_n16195,
    new_n16196_1, new_n16197, new_n16198, new_n16199, new_n16200,
    new_n16201, new_n16202, new_n16203, new_n16204, new_n16205,
    new_n16206_1, new_n16207, new_n16208, new_n16209, new_n16210,
    new_n16211, new_n16212, new_n16213, new_n16214, new_n16215_1,
    new_n16216, new_n16217_1, new_n16218_1, new_n16219_1, new_n16220,
    new_n16221, new_n16222, new_n16223_1, new_n16224, new_n16225,
    new_n16229, new_n16230_1, new_n16231, new_n16232, new_n16233,
    new_n16234, new_n16235, new_n16236, new_n16237, new_n16238, new_n16239,
    new_n16240, new_n16241, new_n16242, new_n16243_1, new_n16244,
    new_n16245, new_n16246, new_n16247_1, new_n16248, new_n16249,
    new_n16250, new_n16251, new_n16252, new_n16253, new_n16254, new_n16255,
    new_n16256, new_n16257, new_n16258, new_n16259, new_n16260, new_n16261,
    new_n16262, new_n16263, new_n16264, new_n16265, new_n16266, new_n16267,
    new_n16268, new_n16269, new_n16270, new_n16271, new_n16272, new_n16273,
    new_n16274, new_n16275_1, new_n16276, new_n16277, new_n16278,
    new_n16279_1, new_n16280, new_n16281, new_n16282, new_n16283,
    new_n16284, new_n16285, new_n16286, new_n16287, new_n16288, new_n16289,
    new_n16290, new_n16291, new_n16292, new_n16293, new_n16294, new_n16295,
    new_n16296, new_n16297, new_n16298, new_n16299, new_n16300, new_n16301,
    new_n16302, new_n16303, new_n16304, new_n16305, new_n16306, new_n16307,
    new_n16308, new_n16309, new_n16310, new_n16311, new_n16312, new_n16313,
    new_n16314, new_n16315, new_n16316, new_n16317, new_n16318, new_n16319,
    new_n16320, new_n16321, new_n16322_1, new_n16323, new_n16324,
    new_n16325, new_n16326, new_n16327_1, new_n16328, new_n16329,
    new_n16330, new_n16331, new_n16332, new_n16333, new_n16334, new_n16335,
    new_n16336, new_n16337, new_n16338, new_n16339, new_n16340, new_n16341,
    new_n16342, new_n16343, new_n16344, new_n16345, new_n16346, new_n16347,
    new_n16348, new_n16349, new_n16350_1, new_n16351, new_n16352,
    new_n16353, new_n16354, new_n16355, new_n16356, new_n16357, new_n16358,
    new_n16359, new_n16360, new_n16361, new_n16362, new_n16363, new_n16365,
    new_n16366, new_n16367_1, new_n16368, new_n16369, new_n16370,
    new_n16371, new_n16372, new_n16373, new_n16374, new_n16375, new_n16377,
    new_n16378, new_n16379_1, new_n16380, new_n16381, new_n16382,
    new_n16383, new_n16384, new_n16385, new_n16386, new_n16387, new_n16388,
    new_n16389, new_n16390, new_n16391, new_n16392, new_n16393, new_n16394,
    new_n16395, new_n16396_1, new_n16397, new_n16398_1, new_n16399,
    new_n16400, new_n16401, new_n16402, new_n16403, new_n16404, new_n16405,
    new_n16406_1, new_n16407_1, new_n16408, new_n16409, new_n16410,
    new_n16411, new_n16412, new_n16413, new_n16414, new_n16416, new_n16417,
    new_n16418, new_n16419_1, new_n16420, new_n16421, new_n16422,
    new_n16423, new_n16424_1, new_n16425, new_n16426, new_n16427,
    new_n16428_1, new_n16429, new_n16430, new_n16431, new_n16432,
    new_n16433_1, new_n16434, new_n16435, new_n16436, new_n16437,
    new_n16438, new_n16439_1, new_n16440_1, new_n16441, new_n16442,
    new_n16443, new_n16444, new_n16445_1, new_n16446, new_n16447,
    new_n16448, new_n16449, new_n16450, new_n16451, new_n16452, new_n16454,
    new_n16455, new_n16456, new_n16457, new_n16458, new_n16459,
    new_n16460_1, new_n16461, new_n16462, new_n16463, new_n16464,
    new_n16465, new_n16466, new_n16467, new_n16468, new_n16469, new_n16470,
    new_n16471, new_n16472, new_n16473, new_n16474, new_n16475,
    new_n16476_1, new_n16477, new_n16478, new_n16479, new_n16480,
    new_n16481_1, new_n16482_1, new_n16483, new_n16484, new_n16485,
    new_n16488, new_n16489, new_n16490, new_n16491, new_n16492,
    new_n16493_1, new_n16494, new_n16495, new_n16496, new_n16497,
    new_n16498, new_n16499, new_n16500, new_n16501, new_n16502_1,
    new_n16503, new_n16504, new_n16505, new_n16506_1, new_n16507_1,
    new_n16508, new_n16509, new_n16510, new_n16511, new_n16512, new_n16513,
    new_n16515, new_n16516_1, new_n16517_1, new_n16518, new_n16519,
    new_n16520, new_n16521_1, new_n16522, new_n16523, new_n16524_1,
    new_n16525, new_n16526, new_n16527_1, new_n16528, new_n16529,
    new_n16530, new_n16531, new_n16532, new_n16533, new_n16534, new_n16535,
    new_n16536, new_n16537, new_n16538, new_n16539, new_n16540, new_n16541,
    new_n16542, new_n16543, new_n16544_1, new_n16545, new_n16546,
    new_n16547, new_n16548, new_n16549, new_n16550, new_n16551, new_n16552,
    new_n16553, new_n16554_1, new_n16555, new_n16556, new_n16557,
    new_n16558, new_n16559, new_n16560, new_n16561, new_n16562, new_n16563,
    new_n16564, new_n16565, new_n16566, new_n16567, new_n16568, new_n16569,
    new_n16570, new_n16571, new_n16572, new_n16573, new_n16574, new_n16575,
    new_n16576, new_n16577, new_n16578, new_n16579, new_n16580, new_n16581,
    new_n16583_1, new_n16584_1, new_n16585, new_n16586, new_n16587,
    new_n16588, new_n16589_1, new_n16590, new_n16591, new_n16592,
    new_n16593, new_n16594, new_n16595, new_n16596_1, new_n16597,
    new_n16598, new_n16599, new_n16600, new_n16601, new_n16602, new_n16603,
    new_n16604, new_n16605, new_n16606, new_n16607, new_n16608_1,
    new_n16609, new_n16610, new_n16611, new_n16612, new_n16613, new_n16614,
    new_n16615, new_n16616, new_n16617_1, new_n16618, new_n16619,
    new_n16620, new_n16621, new_n16622, new_n16623, new_n16624, new_n16625,
    new_n16626, new_n16627, new_n16628, new_n16629, new_n16630_1,
    new_n16631, new_n16632, new_n16633, new_n16634, new_n16635, new_n16636,
    new_n16637, new_n16638, new_n16639, new_n16640_1, new_n16641,
    new_n16642, new_n16643, new_n16644, new_n16645, new_n16646, new_n16647,
    new_n16648, new_n16649, new_n16650, new_n16651, new_n16652, new_n16653,
    new_n16654, new_n16655, new_n16656_1, new_n16657, new_n16658,
    new_n16659, new_n16660, new_n16661, new_n16662, new_n16663, new_n16664,
    new_n16665, new_n16666, new_n16667, new_n16668, new_n16669, new_n16670,
    new_n16671, new_n16672, new_n16673, new_n16674_1, new_n16675,
    new_n16676, new_n16677, new_n16678, new_n16679, new_n16680, new_n16681,
    new_n16682_1, new_n16683, new_n16684_1, new_n16685, new_n16686,
    new_n16687, new_n16688_1, new_n16689, new_n16690, new_n16691,
    new_n16692, new_n16693, new_n16694, new_n16695, new_n16696, new_n16697,
    new_n16698, new_n16699, new_n16700, new_n16701, new_n16702, new_n16703,
    new_n16704, new_n16705, new_n16706, new_n16707, new_n16708, new_n16709,
    new_n16710, new_n16711, new_n16712, new_n16713, new_n16714, new_n16715,
    new_n16716, new_n16717, new_n16718, new_n16719, new_n16720, new_n16721,
    new_n16722_1, new_n16723, new_n16724, new_n16725, new_n16726,
    new_n16727, new_n16728, new_n16729, new_n16730, new_n16731, new_n16732,
    new_n16733_1, new_n16734, new_n16735, new_n16736, new_n16737,
    new_n16738, new_n16739, new_n16741, new_n16742, new_n16743_1,
    new_n16744, new_n16745, new_n16746, new_n16747, new_n16748, new_n16749,
    new_n16750, new_n16751, new_n16752, new_n16753, new_n16754, new_n16755,
    new_n16758, new_n16759, new_n16760, new_n16761, new_n16762, new_n16763,
    new_n16764, new_n16765, new_n16766, new_n16767, new_n16772, new_n16773,
    new_n16774, new_n16775, new_n16776, new_n16777, new_n16778, new_n16779,
    new_n16780, new_n16781, new_n16782, new_n16783, new_n16790, new_n16791,
    new_n16792, new_n16793, new_n16794, new_n16795, new_n16796, new_n16797,
    new_n16798_1, new_n16799, new_n16800, new_n16801, new_n16802,
    new_n16803, new_n16804, new_n16805, new_n16806, new_n16807, new_n16808,
    new_n16809, new_n16810, new_n16811, new_n16812_1, new_n16813,
    new_n16814, new_n16815, new_n16816, new_n16817, new_n16818_1,
    new_n16819, new_n16820, new_n16821, new_n16822, new_n16823,
    new_n16824_1, new_n16825, new_n16826, new_n16827, new_n16828,
    new_n16829, new_n16830, new_n16831, new_n16832, new_n16833,
    new_n16834_1, new_n16835, new_n16836, new_n16837_1, new_n16838,
    new_n16839, new_n16840, new_n16841_1, new_n16842, new_n16843,
    new_n16844, new_n16845, new_n16846, new_n16847, new_n16848, new_n16849,
    new_n16850, new_n16851, new_n16852, new_n16853, new_n16854, new_n16855,
    new_n16856, new_n16857, new_n16858, new_n16859, new_n16860, new_n16861,
    new_n16862, new_n16863, new_n16864, new_n16865, new_n16866, new_n16867,
    new_n16868, new_n16869, new_n16870, new_n16871, new_n16872, new_n16873,
    new_n16874, new_n16875, new_n16876, new_n16877, new_n16878, new_n16879,
    new_n16880, new_n16881, new_n16883, new_n16884, new_n16885_1,
    new_n16886, new_n16887, new_n16888, new_n16889, new_n16890, new_n16891,
    new_n16892, new_n16893, new_n16894, new_n16895, new_n16896, new_n16897,
    new_n16898, new_n16899, new_n16900, new_n16901, new_n16902, new_n16903,
    new_n16904, new_n16905_1, new_n16906, new_n16907, new_n16908,
    new_n16909, new_n16910, new_n16911_1, new_n16912, new_n16913,
    new_n16914, new_n16915, new_n16916, new_n16917, new_n16918, new_n16919,
    new_n16920, new_n16921, new_n16922, new_n16923, new_n16924, new_n16925,
    new_n16926, new_n16927, new_n16929, new_n16930, new_n16931, new_n16932,
    new_n16933, new_n16934, new_n16935, new_n16936, new_n16937, new_n16938,
    new_n16939, new_n16940, new_n16941, new_n16942, new_n16943, new_n16944,
    new_n16945, new_n16946, new_n16947, new_n16948, new_n16949, new_n16950,
    new_n16951_1, new_n16952, new_n16953, new_n16954_1, new_n16955,
    new_n16956, new_n16957, new_n16958, new_n16959, new_n16960, new_n16961,
    new_n16962, new_n16963, new_n16964, new_n16965, new_n16966, new_n16967,
    new_n16968_1, new_n16969, new_n16970, new_n16971_1, new_n16972,
    new_n16973, new_n16974, new_n16975, new_n16976, new_n16977, new_n16978,
    new_n16979, new_n16980, new_n16981, new_n16982, new_n16983, new_n16984,
    new_n16985, new_n16986, new_n16987, new_n16988_1, new_n16989_1,
    new_n16990, new_n16991, new_n16992, new_n16993, new_n16994_1,
    new_n16995, new_n16996, new_n16997, new_n16998, new_n16999, new_n17000,
    new_n17001, new_n17002, new_n17003, new_n17004, new_n17005,
    new_n17006_1, new_n17007, new_n17008, new_n17009, new_n17010,
    new_n17011, new_n17012, new_n17013, new_n17014, new_n17015, new_n17016,
    new_n17017, new_n17018, new_n17019, new_n17020, new_n17021, new_n17022,
    new_n17023, new_n17024, new_n17025, new_n17026, new_n17027, new_n17028,
    new_n17029, new_n17030, new_n17031, new_n17032, new_n17033, new_n17034,
    new_n17035_1, new_n17036, new_n17037_1, new_n17038, new_n17039,
    new_n17040, new_n17041, new_n17042, new_n17043, new_n17044, new_n17045,
    new_n17046, new_n17047, new_n17048, new_n17049, new_n17050, new_n17051,
    new_n17052, new_n17053, new_n17054, new_n17055, new_n17056, new_n17057,
    new_n17058, new_n17059, new_n17060, new_n17061, new_n17062, new_n17063,
    new_n17064, new_n17065, new_n17066, new_n17067, new_n17068_1,
    new_n17069_1, new_n17070_1, new_n17071, new_n17072, new_n17073,
    new_n17074, new_n17075_1, new_n17076, new_n17077_1, new_n17078,
    new_n17079, new_n17080, new_n17082, new_n17083, new_n17084_1,
    new_n17085, new_n17086, new_n17087, new_n17088, new_n17089,
    new_n17090_1, new_n17091, new_n17092, new_n17093, new_n17094,
    new_n17095_1, new_n17096, new_n17097, new_n17098, new_n17099,
    new_n17100, new_n17101, new_n17102, new_n17103, new_n17104_1,
    new_n17105, new_n17106_1, new_n17107, new_n17108, new_n17109,
    new_n17110, new_n17111, new_n17112, new_n17113, new_n17114, new_n17115,
    new_n17116, new_n17117, new_n17118, new_n17119_1, new_n17120,
    new_n17121, new_n17122, new_n17123, new_n17124, new_n17125, new_n17126,
    new_n17127, new_n17128, new_n17131, new_n17132, new_n17133, new_n17134,
    new_n17135, new_n17136, new_n17137, new_n17138_1, new_n17139,
    new_n17140, new_n17141, new_n17142, new_n17143, new_n17144, new_n17145,
    new_n17146, new_n17149, new_n17150, new_n17151, new_n17152, new_n17153,
    new_n17154, new_n17155, new_n17156, new_n17157, new_n17161, new_n17162,
    new_n17163_1, new_n17164, new_n17165, new_n17166, new_n17167,
    new_n17168_1, new_n17169, new_n17170, new_n17171, new_n17172,
    new_n17173, new_n17174, new_n17175, new_n17176, new_n17177, new_n17178,
    new_n17179, new_n17180, new_n17181, new_n17182, new_n17183, new_n17184,
    new_n17185, new_n17186, new_n17187, new_n17188, new_n17189, new_n17190,
    new_n17191, new_n17192, new_n17193, new_n17194, new_n17195, new_n17196,
    new_n17197, new_n17198, new_n17199, new_n17200, new_n17201,
    new_n17202_1, new_n17203, new_n17204, new_n17207, new_n17208,
    new_n17209, new_n17210, new_n17211, new_n17212, new_n17213, new_n17214,
    new_n17215, new_n17216, new_n17217, new_n17218, new_n17219_1,
    new_n17220, new_n17221, new_n17222, new_n17223, new_n17224, new_n17225,
    new_n17226, new_n17227, new_n17228, new_n17229, new_n17230, new_n17231,
    new_n17232_1, new_n17233, new_n17234, new_n17235, new_n17236_1,
    new_n17237, new_n17238, new_n17239, new_n17240, new_n17241, new_n17242,
    new_n17243_1, new_n17244, new_n17245, new_n17246, new_n17247,
    new_n17248, new_n17249, new_n17250_1, new_n17251_1, new_n17252,
    new_n17253, new_n17254, new_n17255, new_n17256, new_n17257, new_n17258,
    new_n17259, new_n17260, new_n17261, new_n17262, new_n17263_1,
    new_n17264, new_n17265, new_n17266, new_n17267, new_n17268, new_n17269,
    new_n17270, new_n17271, new_n17272, new_n17273, new_n17274, new_n17275,
    new_n17276, new_n17277, new_n17278, new_n17279, new_n17280, new_n17281,
    new_n17282, new_n17283, new_n17284, new_n17285_1, new_n17286,
    new_n17287, new_n17288, new_n17289, new_n17290, new_n17291, new_n17293,
    new_n17294, new_n17295, new_n17296, new_n17297, new_n17298, new_n17299,
    new_n17300, new_n17301, new_n17302_1, new_n17303, new_n17304,
    new_n17305, new_n17306, new_n17307, new_n17308, new_n17309, new_n17310,
    new_n17311, new_n17312, new_n17313, new_n17314, new_n17315, new_n17316,
    new_n17317, new_n17318, new_n17319, new_n17320_1, new_n17321,
    new_n17322, new_n17323, new_n17324, new_n17325, new_n17326, new_n17327,
    new_n17328, new_n17329, new_n17331, new_n17332, new_n17333, new_n17334,
    new_n17335, new_n17336, new_n17337_1, new_n17338, new_n17339,
    new_n17340, new_n17341, new_n17342, new_n17343, new_n17344_1,
    new_n17345, new_n17346, new_n17347, new_n17348, new_n17349, new_n17350,
    new_n17351_1, new_n17352, new_n17353, new_n17354, new_n17355,
    new_n17356, new_n17357, new_n17358, new_n17359_1, new_n17360,
    new_n17361, new_n17362, new_n17363, new_n17364, new_n17365, new_n17366,
    new_n17367, new_n17368, new_n17369, new_n17370, new_n17371, new_n17372,
    new_n17373, new_n17374, new_n17375, new_n17376, new_n17377, new_n17378,
    new_n17379, new_n17380, new_n17381, new_n17382, new_n17383, new_n17384,
    new_n17385, new_n17386, new_n17387_1, new_n17388, new_n17394,
    new_n17395, new_n17396, new_n17397, new_n17398, new_n17399, new_n17400,
    new_n17401, new_n17402, new_n17403, new_n17404, new_n17405, new_n17406,
    new_n17407, new_n17408, new_n17409, new_n17410, new_n17411, new_n17412,
    new_n17413, new_n17414, new_n17415, new_n17416, new_n17417, new_n17418,
    new_n17419, new_n17420, new_n17421_1, new_n17422, new_n17423,
    new_n17424, new_n17425, new_n17426, new_n17427, new_n17428, new_n17429,
    new_n17430, new_n17431, new_n17432_1, new_n17433, new_n17434,
    new_n17435, new_n17436_1, new_n17437, new_n17438, new_n17439,
    new_n17440_1, new_n17441, new_n17442, new_n17443, new_n17444,
    new_n17445, new_n17446, new_n17447, new_n17448, new_n17449,
    new_n17450_1, new_n17451, new_n17452, new_n17453, new_n17454,
    new_n17455, new_n17456, new_n17457, new_n17460, new_n17461_1,
    new_n17462, new_n17463, new_n17464, new_n17465, new_n17466_1,
    new_n17467, new_n17468, new_n17469, new_n17470, new_n17471, new_n17472,
    new_n17473, new_n17474, new_n17475, new_n17476, new_n17477, new_n17478,
    new_n17479, new_n17480, new_n17481, new_n17482, new_n17483, new_n17484,
    new_n17485, new_n17488, new_n17489, new_n17490, new_n17491, new_n17492,
    new_n17493_1, new_n17494, new_n17495, new_n17496, new_n17497,
    new_n17498, new_n17499, new_n17500_1, new_n17501, new_n17502,
    new_n17503, new_n17504, new_n17505, new_n17506, new_n17507, new_n17509,
    new_n17514, new_n17515, new_n17516, new_n17517, new_n17518, new_n17519,
    new_n17520, new_n17521, new_n17522, new_n17523, new_n17524_1,
    new_n17525, new_n17526, new_n17527, new_n17528, new_n17529_1,
    new_n17530, new_n17531, new_n17532, new_n17533, new_n17534, new_n17535,
    new_n17536, new_n17537, new_n17538, new_n17539, new_n17540, new_n17541,
    new_n17542, new_n17543, new_n17544, new_n17545, new_n17546, new_n17547,
    new_n17548, new_n17549, new_n17550, new_n17551, new_n17552, new_n17553,
    new_n17554, new_n17555, new_n17556, new_n17557_1, new_n17558,
    new_n17559, new_n17560, new_n17561, new_n17562, new_n17563, new_n17564,
    new_n17565, new_n17566, new_n17567, new_n17568, new_n17569, new_n17570,
    new_n17571, new_n17572, new_n17573, new_n17574, new_n17575, new_n17576,
    new_n17577, new_n17578, new_n17579, new_n17580, new_n17581, new_n17582,
    new_n17583_1, new_n17584, new_n17585, new_n17586, new_n17587,
    new_n17588, new_n17589, new_n17590, new_n17591, new_n17592_1,
    new_n17593, new_n17594, new_n17595, new_n17596, new_n17597, new_n17598,
    new_n17599, new_n17600, new_n17601, new_n17602, new_n17603, new_n17604,
    new_n17605, new_n17606, new_n17607, new_n17608, new_n17609, new_n17610,
    new_n17611, new_n17612, new_n17613, new_n17614, new_n17615, new_n17616,
    new_n17617, new_n17618, new_n17619, new_n17620, new_n17621, new_n17625,
    new_n17626, new_n17627, new_n17628, new_n17629, new_n17630, new_n17631,
    new_n17632, new_n17633, new_n17634, new_n17635, new_n17636, new_n17637,
    new_n17638_1, new_n17639, new_n17640, new_n17641, new_n17642,
    new_n17643, new_n17644, new_n17645, new_n17646, new_n17647, new_n17648,
    new_n17649, new_n17650, new_n17651, new_n17658, new_n17659, new_n17660,
    new_n17661, new_n17662, new_n17663, new_n17664_1, new_n17665,
    new_n17666, new_n17667, new_n17668, new_n17669, new_n17670, new_n17671,
    new_n17672, new_n17673, new_n17674, new_n17675, new_n17676, new_n17677,
    new_n17678, new_n17679, new_n17680, new_n17681, new_n17682, new_n17683,
    new_n17684, new_n17685, new_n17686, new_n17687_1, new_n17688,
    new_n17689, new_n17690, new_n17691, new_n17692, new_n17693, new_n17694,
    new_n17695, new_n17696, new_n17697, new_n17698, new_n17699, new_n17700,
    new_n17701, new_n17702, new_n17703, new_n17704, new_n17705, new_n17706,
    new_n17707, new_n17708, new_n17709, new_n17710, new_n17711, new_n17712,
    new_n17713, new_n17714, new_n17715, new_n17716, new_n17717, new_n17718,
    new_n17719, new_n17720, new_n17721_1, new_n17722, new_n17723,
    new_n17724, new_n17725, new_n17726, new_n17727, new_n17728, new_n17729,
    new_n17732, new_n17733, new_n17734, new_n17735_1, new_n17736,
    new_n17737, new_n17738_1, new_n17739, new_n17740, new_n17741,
    new_n17742, new_n17743, new_n17744, new_n17745, new_n17746_1,
    new_n17747, new_n17748, new_n17749_1, new_n17750, new_n17751,
    new_n17752, new_n17753, new_n17754, new_n17755, new_n17756, new_n17757,
    new_n17758, new_n17759, new_n17760, new_n17761, new_n17762, new_n17763,
    new_n17764, new_n17765, new_n17766, new_n17767, new_n17768, new_n17769,
    new_n17770, new_n17771, new_n17772, new_n17773, new_n17774, new_n17775,
    new_n17776, new_n17777, new_n17778, new_n17779, new_n17780, new_n17781,
    new_n17782, new_n17783, new_n17784_1, new_n17785, new_n17786,
    new_n17787, new_n17788, new_n17789, new_n17790, new_n17791, new_n17792,
    new_n17793, new_n17794, new_n17795, new_n17796, new_n17797, new_n17798,
    new_n17799, new_n17800, new_n17801, new_n17802, new_n17803, new_n17804,
    new_n17805, new_n17806, new_n17808, new_n17809, new_n17810, new_n17811,
    new_n17812, new_n17813, new_n17814, new_n17815, new_n17816, new_n17817,
    new_n17818, new_n17819, new_n17820_1, new_n17821, new_n17822,
    new_n17823, new_n17824, new_n17825, new_n17826, new_n17827, new_n17828,
    new_n17829, new_n17830, new_n17831, new_n17832, new_n17833, new_n17834,
    new_n17835, new_n17836, new_n17837, new_n17838, new_n17839, new_n17840,
    new_n17841, new_n17842, new_n17843, new_n17844, new_n17845, new_n17846,
    new_n17847, new_n17848, new_n17849, new_n17850, new_n17851, new_n17852,
    new_n17853, new_n17854, new_n17855_1, new_n17856, new_n17857,
    new_n17858, new_n17859, new_n17861, new_n17862, new_n17863, new_n17864,
    new_n17865, new_n17866, new_n17867, new_n17868, new_n17869, new_n17870,
    new_n17871, new_n17872, new_n17873, new_n17874, new_n17875, new_n17876,
    new_n17877_1, new_n17878, new_n17879, new_n17880, new_n17881,
    new_n17882, new_n17883, new_n17884, new_n17885, new_n17886, new_n17887,
    new_n17888, new_n17889_1, new_n17890, new_n17891, new_n17892,
    new_n17893, new_n17894, new_n17895, new_n17896, new_n17897, new_n17898,
    new_n17899, new_n17900, new_n17901, new_n17902, new_n17903, new_n17908,
    new_n17909, new_n17910, new_n17911_1, new_n17912_1, new_n17913,
    new_n17914, new_n17915, new_n17916, new_n17917, new_n17918, new_n17919,
    new_n17920, new_n17921, new_n17922, new_n17923, new_n17928, new_n17929,
    new_n17930, new_n17931_1, new_n17932, new_n17933, new_n17934,
    new_n17935, new_n17936, new_n17937, new_n17938, new_n17939, new_n17940,
    new_n17941, new_n17942, new_n17943, new_n17944, new_n17945, new_n17946,
    new_n17947, new_n17948_1, new_n17949, new_n17950, new_n17951,
    new_n17952, new_n17953, new_n17954_1, new_n17955, new_n17956_1,
    new_n17957, new_n17958, new_n17959_1, new_n17960, new_n17961,
    new_n17962, new_n17963_1, new_n17964, new_n17965, new_n17966,
    new_n17967, new_n17968_1, new_n17969, new_n17970, new_n17971,
    new_n17972, new_n17973, new_n17974, new_n17976_1, new_n17977,
    new_n17978, new_n17979, new_n17981, new_n17982, new_n17983, new_n17984,
    new_n17985, new_n17986, new_n17987, new_n17988, new_n17989, new_n17990,
    new_n17991, new_n17992, new_n17996, new_n17997, new_n17998_1,
    new_n17999, new_n18000, new_n18001, new_n18002, new_n18003, new_n18004,
    new_n18005, new_n18006, new_n18007, new_n18008, new_n18009, new_n18010,
    new_n18011, new_n18012, new_n18013, new_n18015, new_n18016, new_n18017,
    new_n18018, new_n18019, new_n18020, new_n18021, new_n18022, new_n18023,
    new_n18024, new_n18025_1, new_n18026, new_n18027, new_n18028,
    new_n18029, new_n18030, new_n18031, new_n18032, new_n18033, new_n18034,
    new_n18035_1, new_n18036, new_n18037, new_n18038, new_n18039,
    new_n18040, new_n18041, new_n18042, new_n18043_1, new_n18044,
    new_n18045_1, new_n18046, new_n18047, new_n18048, new_n18049,
    new_n18050, new_n18051, new_n18052, new_n18053, new_n18054, new_n18055,
    new_n18056, new_n18057, new_n18058, new_n18059_1, new_n18060,
    new_n18061_1, new_n18062, new_n18063, new_n18064, new_n18065,
    new_n18066, new_n18067, new_n18068, new_n18069, new_n18070,
    new_n18071_1, new_n18072, new_n18073, new_n18074, new_n18075,
    new_n18076, new_n18077, new_n18079, new_n18080, new_n18081, new_n18082,
    new_n18083, new_n18084, new_n18085, new_n18086, new_n18087, new_n18088,
    new_n18090, new_n18091, new_n18092, new_n18093, new_n18094, new_n18095,
    new_n18096, new_n18097, new_n18098, new_n18099, new_n18100, new_n18101,
    new_n18102, new_n18103, new_n18104, new_n18105_1, new_n18106,
    new_n18107, new_n18108, new_n18109, new_n18110, new_n18111, new_n18112,
    new_n18113, new_n18114, new_n18115, new_n18116, new_n18117, new_n18118,
    new_n18119, new_n18120, new_n18121, new_n18122, new_n18123, new_n18124,
    new_n18125, new_n18126, new_n18127, new_n18128, new_n18129, new_n18130,
    new_n18131, new_n18132, new_n18133, new_n18134, new_n18135, new_n18136,
    new_n18137, new_n18138, new_n18139, new_n18140, new_n18141, new_n18142,
    new_n18143_1, new_n18144, new_n18145_1, new_n18146, new_n18147,
    new_n18148, new_n18149, new_n18150, new_n18151_1, new_n18152_1,
    new_n18153, new_n18154, new_n18155, new_n18156, new_n18157_1,
    new_n18158, new_n18159, new_n18160, new_n18161, new_n18162, new_n18163,
    new_n18164, new_n18165, new_n18166, new_n18167, new_n18168, new_n18169,
    new_n18170, new_n18171_1, new_n18172, new_n18173, new_n18174,
    new_n18175, new_n18176, new_n18177, new_n18178, new_n18179, new_n18180,
    new_n18181, new_n18182, new_n18183, new_n18184, new_n18185, new_n18186,
    new_n18187, new_n18188, new_n18189, new_n18190, new_n18191, new_n18192,
    new_n18193_1, new_n18194, new_n18195, new_n18196, new_n18197,
    new_n18198, new_n18199, new_n18200, new_n18201, new_n18202, new_n18203,
    new_n18204, new_n18205, new_n18206, new_n18207, new_n18208, new_n18209,
    new_n18210, new_n18211, new_n18212, new_n18213, new_n18214, new_n18215,
    new_n18216, new_n18217, new_n18218, new_n18219, new_n18220, new_n18221,
    new_n18222, new_n18223, new_n18224, new_n18225, new_n18226,
    new_n18227_1, new_n18228, new_n18229, new_n18230, new_n18231,
    new_n18232_1, new_n18233, new_n18234, new_n18235, new_n18236,
    new_n18237, new_n18238_1, new_n18239, new_n18240, new_n18241_1,
    new_n18242, new_n18243, new_n18244, new_n18245, new_n18246, new_n18247,
    new_n18248, new_n18249, new_n18250, new_n18251, new_n18252, new_n18253,
    new_n18254_1, new_n18255, new_n18256, new_n18257, new_n18258,
    new_n18259, new_n18260, new_n18261, new_n18262, new_n18263, new_n18264,
    new_n18265, new_n18266, new_n18267, new_n18268, new_n18269, new_n18270,
    new_n18271, new_n18272, new_n18273, new_n18274_1, new_n18275,
    new_n18276, new_n18277, new_n18278, new_n18279, new_n18280, new_n18281,
    new_n18282, new_n18283, new_n18284, new_n18287, new_n18288_1,
    new_n18289, new_n18290_1, new_n18291, new_n18292, new_n18293,
    new_n18294, new_n18295_1, new_n18296, new_n18297, new_n18298,
    new_n18299, new_n18300, new_n18301_1, new_n18302, new_n18303,
    new_n18304_1, new_n18305, new_n18306, new_n18307, new_n18308,
    new_n18309, new_n18310_1, new_n18311_1, new_n18312, new_n18313,
    new_n18315, new_n18316, new_n18317, new_n18318, new_n18319, new_n18320,
    new_n18321, new_n18322, new_n18323_1, new_n18324, new_n18325,
    new_n18326, new_n18327, new_n18328, new_n18329, new_n18330, new_n18331,
    new_n18332_1, new_n18333, new_n18336, new_n18337, new_n18338,
    new_n18339, new_n18340, new_n18341, new_n18346, new_n18347, new_n18348,
    new_n18349, new_n18350_1, new_n18351, new_n18352, new_n18353,
    new_n18354, new_n18355, new_n18356, new_n18357, new_n18358, new_n18359,
    new_n18360, new_n18361, new_n18362_1, new_n18363, new_n18364,
    new_n18365, new_n18366, new_n18367, new_n18368, new_n18369, new_n18370,
    new_n18371, new_n18372, new_n18373, new_n18374, new_n18375, new_n18376,
    new_n18377_1, new_n18378, new_n18379, new_n18380, new_n18381,
    new_n18382, new_n18383, new_n18384, new_n18385, new_n18386, new_n18387,
    new_n18388, new_n18389, new_n18390, new_n18391, new_n18392, new_n18393,
    new_n18394, new_n18395, new_n18396, new_n18397, new_n18398, new_n18399,
    new_n18400, new_n18401, new_n18402, new_n18403, new_n18404,
    new_n18405_1, new_n18406, new_n18407, new_n18408, new_n18409_1,
    new_n18410, new_n18411, new_n18412, new_n18413, new_n18414_1,
    new_n18415, new_n18416, new_n18417, new_n18418_1, new_n18419,
    new_n18420, new_n18421, new_n18422, new_n18423, new_n18424, new_n18425,
    new_n18426, new_n18427, new_n18428, new_n18429, new_n18430, new_n18431,
    new_n18432, new_n18433, new_n18434, new_n18435, new_n18436,
    new_n18437_1, new_n18438, new_n18439_1, new_n18440, new_n18441,
    new_n18442, new_n18443, new_n18444_1, new_n18445_1, new_n18446,
    new_n18447, new_n18448, new_n18449, new_n18450, new_n18451, new_n18454,
    new_n18455, new_n18456, new_n18457, new_n18458, new_n18459, new_n18460,
    new_n18461, new_n18462, new_n18463, new_n18464, new_n18465, new_n18466,
    new_n18467_1, new_n18468, new_n18469, new_n18471, new_n18472,
    new_n18473, new_n18474, new_n18475, new_n18476, new_n18477, new_n18478,
    new_n18479, new_n18480, new_n18481, new_n18482_1, new_n18483_1,
    new_n18484, new_n18485, new_n18486, new_n18487, new_n18488, new_n18489,
    new_n18490, new_n18491, new_n18492, new_n18493, new_n18494, new_n18495,
    new_n18496_1, new_n18497, new_n18498, new_n18499, new_n18500,
    new_n18501, new_n18502, new_n18503, new_n18504, new_n18505, new_n18506,
    new_n18507, new_n18508, new_n18509_1, new_n18510, new_n18511,
    new_n18512, new_n18513_1, new_n18514, new_n18515_1, new_n18516,
    new_n18517, new_n18518, new_n18521, new_n18522, new_n18523, new_n18524,
    new_n18525, new_n18526, new_n18527, new_n18528, new_n18529, new_n18530,
    new_n18531, new_n18532, new_n18533, new_n18534, new_n18535, new_n18536,
    new_n18537_1, new_n18538, new_n18539, new_n18540, new_n18541,
    new_n18542, new_n18543, new_n18544, new_n18545, new_n18546, new_n18547,
    new_n18548, new_n18549, new_n18550, new_n18551, new_n18552, new_n18553,
    new_n18554, new_n18556, new_n18557, new_n18558_1, new_n18559,
    new_n18560, new_n18561, new_n18562, new_n18563, new_n18564, new_n18565,
    new_n18566, new_n18567, new_n18568, new_n18569, new_n18570, new_n18571,
    new_n18572_1, new_n18573, new_n18574_1, new_n18575, new_n18576_1,
    new_n18577, new_n18578_1, new_n18579, new_n18580, new_n18581,
    new_n18582_1, new_n18583_1, new_n18584_1, new_n18585, new_n18586,
    new_n18587, new_n18588, new_n18589, new_n18590, new_n18595, new_n18596,
    new_n18597, new_n18598, new_n18599, new_n18600, new_n18601, new_n18602,
    new_n18603, new_n18604, new_n18605, new_n18606, new_n18607, new_n18608,
    new_n18609, new_n18610_1, new_n18611, new_n18612, new_n18613,
    new_n18618, new_n18619, new_n18620, new_n18621, new_n18622, new_n18623,
    new_n18624, new_n18625, new_n18626, new_n18627, new_n18628, new_n18629,
    new_n18630, new_n18631, new_n18632, new_n18633, new_n18634,
    new_n18635_1, new_n18636, new_n18637, new_n18638, new_n18639,
    new_n18640, new_n18641, new_n18642, new_n18643, new_n18644, new_n18645,
    new_n18646, new_n18647, new_n18648, new_n18649_1, new_n18650,
    new_n18651, new_n18652, new_n18653_1, new_n18654, new_n18655,
    new_n18656, new_n18657, new_n18658, new_n18659, new_n18660, new_n18661,
    new_n18662, new_n18663, new_n18664, new_n18665, new_n18666, new_n18667,
    new_n18668, new_n18669, new_n18670, new_n18671, new_n18672, new_n18673,
    new_n18674, new_n18675, new_n18676, new_n18677, new_n18678,
    new_n18679_1, new_n18680, new_n18681, new_n18682, new_n18683,
    new_n18684, new_n18685, new_n18686, new_n18687, new_n18688, new_n18689,
    new_n18690_1, new_n18691, new_n18692, new_n18693_1, new_n18694,
    new_n18695, new_n18701, new_n18702, new_n18703, new_n18704, new_n18705,
    new_n18706, new_n18707, new_n18708_1, new_n18709, new_n18710,
    new_n18711, new_n18712, new_n18713, new_n18714, new_n18715, new_n18716,
    new_n18717, new_n18719, new_n18720, new_n18721_1, new_n18722,
    new_n18723, new_n18724, new_n18725_1, new_n18726, new_n18727,
    new_n18728, new_n18729, new_n18730, new_n18731, new_n18732, new_n18733,
    new_n18734, new_n18735, new_n18736, new_n18737_1, new_n18738,
    new_n18739, new_n18740, new_n18741, new_n18742, new_n18743, new_n18744,
    new_n18745_1, new_n18746, new_n18747, new_n18748, new_n18749,
    new_n18750, new_n18751_1, new_n18752, new_n18753, new_n18754,
    new_n18755, new_n18756, new_n18757, new_n18758, new_n18759, new_n18760,
    new_n18761, new_n18762, new_n18763, new_n18764, new_n18765, new_n18766,
    new_n18767, new_n18768, new_n18769, new_n18770, new_n18771, new_n18772,
    new_n18773, new_n18774, new_n18775, new_n18776, new_n18777, new_n18778,
    new_n18779, new_n18780_1, new_n18781, new_n18782_1, new_n18783,
    new_n18784, new_n18785, new_n18786, new_n18787, new_n18788, new_n18789,
    new_n18790, new_n18791, new_n18796, new_n18797, new_n18798, new_n18799,
    new_n18800, new_n18801, new_n18802_1, new_n18803, new_n18804,
    new_n18805, new_n18806, new_n18807, new_n18808, new_n18809, new_n18810,
    new_n18811, new_n18812, new_n18813, new_n18814, new_n18815, new_n18816,
    new_n18817, new_n18818, new_n18819, new_n18820, new_n18821, new_n18822,
    new_n18823, new_n18824, new_n18825, new_n18826, new_n18827, new_n18828,
    new_n18829, new_n18830_1, new_n18831_1, new_n18832, new_n18833,
    new_n18834, new_n18835, new_n18836, new_n18837, new_n18838, new_n18839,
    new_n18840, new_n18841, new_n18842, new_n18843_1, new_n18844,
    new_n18845, new_n18846, new_n18847, new_n18848, new_n18849, new_n18850,
    new_n18851, new_n18852, new_n18853, new_n18854, new_n18855, new_n18856,
    new_n18857, new_n18858_1, new_n18859_1, new_n18860, new_n18863,
    new_n18864_1, new_n18865_1, new_n18866, new_n18867, new_n18868,
    new_n18869, new_n18870, new_n18871, new_n18872, new_n18873, new_n18874,
    new_n18875, new_n18876, new_n18877, new_n18878, new_n18879,
    new_n18880_1, new_n18881, new_n18882, new_n18883, new_n18884,
    new_n18885, new_n18886_1, new_n18887_1, new_n18888, new_n18889,
    new_n18890, new_n18891, new_n18892, new_n18893, new_n18894, new_n18895,
    new_n18896, new_n18897, new_n18898, new_n18899, new_n18900,
    new_n18901_1, new_n18902, new_n18903, new_n18904, new_n18905,
    new_n18906, new_n18907_1, new_n18908, new_n18909, new_n18910,
    new_n18911, new_n18912, new_n18913, new_n18914, new_n18915, new_n18916,
    new_n18917, new_n18918, new_n18919_1, new_n18920, new_n18921,
    new_n18922, new_n18923, new_n18924, new_n18925, new_n18928, new_n18929,
    new_n18930, new_n18931, new_n18932, new_n18933, new_n18934, new_n18935,
    new_n18936, new_n18937, new_n18938, new_n18939, new_n18940_1,
    new_n18941, new_n18942, new_n18943, new_n18944, new_n18946, new_n18947,
    new_n18948, new_n18949, new_n18950, new_n18951, new_n18952, new_n18953,
    new_n18954, new_n18955, new_n18956, new_n18957, new_n18958, new_n18959,
    new_n18960, new_n18961, new_n18962_1, new_n18963, new_n18964,
    new_n18965, new_n18967, new_n18968, new_n18969, new_n18970_1,
    new_n18971, new_n18972, new_n18973, new_n18974, new_n18975, new_n18976,
    new_n18977_1, new_n18978, new_n18979, new_n18980, new_n18981,
    new_n18982_1, new_n18983, new_n18984, new_n18985, new_n18986,
    new_n18987, new_n18988, new_n18989, new_n18990, new_n18991, new_n18992,
    new_n18993, new_n18994, new_n18995, new_n18996, new_n18997, new_n18998,
    new_n18999_1, new_n19000, new_n19001, new_n19002, new_n19003,
    new_n19004, new_n19005_1, new_n19006, new_n19007, new_n19011,
    new_n19012, new_n19013, new_n19014, new_n19015, new_n19016, new_n19017,
    new_n19018, new_n19019, new_n19020, new_n19021, new_n19022, new_n19023,
    new_n19024, new_n19025, new_n19026, new_n19027, new_n19028, new_n19029,
    new_n19030, new_n19031, new_n19032, new_n19033_1, new_n19034,
    new_n19035, new_n19036, new_n19037, new_n19038, new_n19039, new_n19040,
    new_n19041, new_n19042_1, new_n19043, new_n19044_1, new_n19045,
    new_n19046, new_n19047, new_n19048, new_n19049, new_n19050, new_n19051,
    new_n19052, new_n19053, new_n19054, new_n19055, new_n19056, new_n19057,
    new_n19058, new_n19059, new_n19061, new_n19062, new_n19063, new_n19064,
    new_n19065, new_n19066, new_n19067, new_n19068, new_n19069, new_n19070,
    new_n19071, new_n19072, new_n19073, new_n19074, new_n19075, new_n19076,
    new_n19077, new_n19078, new_n19079, new_n19080, new_n19081_1,
    new_n19082, new_n19083, new_n19084, new_n19085, new_n19086, new_n19087,
    new_n19088, new_n19090, new_n19091, new_n19092, new_n19093, new_n19094,
    new_n19095, new_n19096, new_n19097, new_n19098, new_n19099, new_n19100,
    new_n19101, new_n19102, new_n19103, new_n19104, new_n19105, new_n19110,
    new_n19111, new_n19112, new_n19113, new_n19114, new_n19115,
    new_n19116_1, new_n19117, new_n19118, new_n19121, new_n19122,
    new_n19123, new_n19124, new_n19125_1, new_n19126, new_n19127,
    new_n19128, new_n19129, new_n19130, new_n19131, new_n19132, new_n19133,
    new_n19134, new_n19135, new_n19136, new_n19137, new_n19138, new_n19139,
    new_n19140, new_n19141_1, new_n19142, new_n19143, new_n19144_1,
    new_n19145, new_n19146, new_n19147, new_n19148, new_n19149, new_n19150,
    new_n19151, new_n19152, new_n19153, new_n19154, new_n19155, new_n19156,
    new_n19157, new_n19158, new_n19159, new_n19160, new_n19161, new_n19162,
    new_n19163_1, new_n19164_1, new_n19165, new_n19166, new_n19167,
    new_n19168, new_n19169, new_n19170, new_n19171, new_n19172, new_n19173,
    new_n19174_1, new_n19175, new_n19176_1, new_n19177, new_n19178,
    new_n19179, new_n19180, new_n19181, new_n19182, new_n19183, new_n19184,
    new_n19185, new_n19186, new_n19191, new_n19192, new_n19193, new_n19194,
    new_n19195, new_n19196_1, new_n19197, new_n19198, new_n19199,
    new_n19200, new_n19201, new_n19202_1, new_n19203, new_n19204,
    new_n19205, new_n19206, new_n19207, new_n19208, new_n19209, new_n19210,
    new_n19211, new_n19212, new_n19216, new_n19217, new_n19218, new_n19219,
    new_n19220_1, new_n19221_1, new_n19222, new_n19223_1, new_n19224_1,
    new_n19225, new_n19226, new_n19227, new_n19228_1, new_n19229,
    new_n19230, new_n19231, new_n19232, new_n19233_1, new_n19234_1,
    new_n19235, new_n19236, new_n19237, new_n19238, new_n19239, new_n19240,
    new_n19241, new_n19242, new_n19243, new_n19244_1, new_n19245,
    new_n19246, new_n19247, new_n19248, new_n19249, new_n19250, new_n19251,
    new_n19252, new_n19253, new_n19254, new_n19255, new_n19256, new_n19257,
    new_n19258, new_n19259, new_n19260, new_n19261, new_n19262, new_n19263,
    new_n19264, new_n19265, new_n19266, new_n19267, new_n19268, new_n19269,
    new_n19270_1, new_n19271, new_n19272, new_n19273, new_n19274,
    new_n19275, new_n19276, new_n19277, new_n19278, new_n19279, new_n19280,
    new_n19281, new_n19282_1, new_n19283, new_n19284, new_n19285,
    new_n19286, new_n19287, new_n19288, new_n19289, new_n19290, new_n19291,
    new_n19292, new_n19293, new_n19294, new_n19295, new_n19296, new_n19297,
    new_n19298, new_n19299, new_n19300, new_n19301, new_n19302, new_n19303,
    new_n19304, new_n19305, new_n19306, new_n19307, new_n19308, new_n19309,
    new_n19310, new_n19318, new_n19319, new_n19320, new_n19321, new_n19322,
    new_n19323_1, new_n19324, new_n19325, new_n19326, new_n19327_1,
    new_n19328, new_n19329, new_n19330, new_n19331, new_n19332,
    new_n19333_1, new_n19334, new_n19335, new_n19336, new_n19337,
    new_n19338, new_n19339, new_n19340, new_n19341, new_n19342, new_n19343,
    new_n19344, new_n19345, new_n19346, new_n19347, new_n19348_1,
    new_n19349, new_n19350, new_n19351, new_n19352, new_n19353,
    new_n19354_1, new_n19355, new_n19356, new_n19357_1, new_n19358,
    new_n19359, new_n19363, new_n19364, new_n19365, new_n19366,
    new_n19367_1, new_n19368, new_n19369, new_n19370, new_n19371,
    new_n19372, new_n19373, new_n19374, new_n19375, new_n19376, new_n19377,
    new_n19378, new_n19379, new_n19380, new_n19381, new_n19382, new_n19383,
    new_n19384, new_n19385_1, new_n19386, new_n19387, new_n19388,
    new_n19389_1, new_n19390, new_n19391, new_n19392, new_n19393,
    new_n19394, new_n19395, new_n19396, new_n19397, new_n19398, new_n19399,
    new_n19400, new_n19401_1, new_n19402, new_n19403, new_n19404,
    new_n19405, new_n19406, new_n19407, new_n19408, new_n19409, new_n19410,
    new_n19411, new_n19412, new_n19413, new_n19414_1, new_n19415,
    new_n19416, new_n19417, new_n19418, new_n19419, new_n19420, new_n19421,
    new_n19422, new_n19423, new_n19424_1, new_n19425, new_n19426,
    new_n19427, new_n19428, new_n19429, new_n19430, new_n19431, new_n19432,
    new_n19433, new_n19434, new_n19435, new_n19436, new_n19437, new_n19438,
    new_n19439, new_n19440, new_n19441, new_n19442, new_n19443, new_n19444,
    new_n19445, new_n19446, new_n19447, new_n19448, new_n19449,
    new_n19450_1, new_n19451, new_n19452, new_n19453, new_n19454_1,
    new_n19455, new_n19457, new_n19458_1, new_n19459, new_n19460,
    new_n19461, new_n19462, new_n19463, new_n19464, new_n19465, new_n19466,
    new_n19470, new_n19471, new_n19472_1, new_n19473, new_n19474,
    new_n19475, new_n19476, new_n19477_1, new_n19478, new_n19479,
    new_n19480, new_n19481, new_n19482, new_n19483, new_n19484, new_n19485,
    new_n19486, new_n19487, new_n19488, new_n19489, new_n19490, new_n19491,
    new_n19492, new_n19494_1, new_n19495, new_n19496_1, new_n19497,
    new_n19498, new_n19499, new_n19500, new_n19501, new_n19502, new_n19503,
    new_n19504, new_n19505, new_n19506, new_n19507, new_n19508, new_n19509,
    new_n19510, new_n19511, new_n19512, new_n19513, new_n19514_1,
    new_n19515_1, new_n19516, new_n19517, new_n19518, new_n19519,
    new_n19520, new_n19521, new_n19522, new_n19523_1, new_n19524,
    new_n19525, new_n19526, new_n19527, new_n19528, new_n19529, new_n19530,
    new_n19531_1, new_n19532, new_n19533, new_n19534, new_n19535,
    new_n19536, new_n19537, new_n19538, new_n19539_1, new_n19540,
    new_n19541, new_n19542, new_n19543, new_n19544, new_n19545, new_n19546,
    new_n19547, new_n19548, new_n19549, new_n19550, new_n19551, new_n19552,
    new_n19553, new_n19554, new_n19555, new_n19556, new_n19557, new_n19558,
    new_n19559, new_n19560, new_n19561, new_n19562, new_n19564, new_n19567,
    new_n19568, new_n19569, new_n19570_1, new_n19571, new_n19572,
    new_n19573, new_n19574, new_n19575_1, new_n19576, new_n19577,
    new_n19578, new_n19579, new_n19580, new_n19581, new_n19582, new_n19583,
    new_n19584_1, new_n19585, new_n19586, new_n19587, new_n19588,
    new_n19589, new_n19590, new_n19591, new_n19592, new_n19593, new_n19594,
    new_n19595, new_n19596, new_n19597, new_n19598, new_n19599, new_n19600,
    new_n19601, new_n19602_1, new_n19603, new_n19604, new_n19605,
    new_n19606, new_n19607, new_n19608_1, new_n19609, new_n19610,
    new_n19611, new_n19612, new_n19613, new_n19614, new_n19615, new_n19616,
    new_n19617_1, new_n19618_1, new_n19619, new_n19620, new_n19621,
    new_n19622, new_n19623_1, new_n19624, new_n19625, new_n19626,
    new_n19627, new_n19628, new_n19629, new_n19630, new_n19631, new_n19632,
    new_n19633, new_n19634, new_n19635, new_n19636, new_n19637, new_n19638,
    new_n19639, new_n19640, new_n19641_1, new_n19642, new_n19643,
    new_n19644, new_n19645, new_n19646, new_n19647, new_n19648_1,
    new_n19649, new_n19650, new_n19651, new_n19652_1, new_n19653,
    new_n19654, new_n19655, new_n19656, new_n19657, new_n19658, new_n19659,
    new_n19660, new_n19661, new_n19662, new_n19663, new_n19664_1,
    new_n19665, new_n19668, new_n19669, new_n19670, new_n19671, new_n19672,
    new_n19673, new_n19674, new_n19675, new_n19676, new_n19677, new_n19678,
    new_n19679, new_n19680_1, new_n19681, new_n19682, new_n19683,
    new_n19684, new_n19685, new_n19686, new_n19687, new_n19688, new_n19689,
    new_n19690, new_n19691, new_n19692, new_n19693, new_n19694, new_n19695,
    new_n19696, new_n19697, new_n19698, new_n19699, new_n19700,
    new_n19701_1, new_n19702, new_n19703, new_n19704, new_n19705,
    new_n19706, new_n19707, new_n19708, new_n19709, new_n19710, new_n19711,
    new_n19712, new_n19713, new_n19714, new_n19715, new_n19716, new_n19717,
    new_n19718, new_n19719, new_n19720, new_n19721, new_n19722, new_n19723,
    new_n19724, new_n19725, new_n19726, new_n19727, new_n19728, new_n19729,
    new_n19730, new_n19731, new_n19732, new_n19733, new_n19740, new_n19741,
    new_n19742, new_n19746, new_n19747, new_n19748, new_n19749_1,
    new_n19750, new_n19751, new_n19752, new_n19753, new_n19754, new_n19755,
    new_n19756_1, new_n19757, new_n19758, new_n19759, new_n19760,
    new_n19761, new_n19762, new_n19763, new_n19764, new_n19765, new_n19766,
    new_n19767_1, new_n19768, new_n19769, new_n19770_1, new_n19771,
    new_n19772, new_n19773, new_n19774, new_n19775, new_n19776, new_n19777,
    new_n19778, new_n19779, new_n19780_1, new_n19781, new_n19782,
    new_n19783, new_n19784, new_n19785, new_n19786, new_n19787, new_n19788,
    new_n19789_1, new_n19790, new_n19791, new_n19792_1, new_n19793,
    new_n19794, new_n19795, new_n19796, new_n19797, new_n19798_1,
    new_n19799, new_n19800, new_n19801, new_n19802, new_n19803_1,
    new_n19804, new_n19805, new_n19806, new_n19807, new_n19808, new_n19809,
    new_n19810, new_n19811, new_n19812, new_n19813, new_n19814, new_n19815,
    new_n19816, new_n19817, new_n19818, new_n19819, new_n19820, new_n19821,
    new_n19822, new_n19823, new_n19824, new_n19825, new_n19826, new_n19827,
    new_n19828, new_n19829, new_n19830, new_n19831, new_n19832, new_n19833,
    new_n19834, new_n19835, new_n19836, new_n19837, new_n19838, new_n19839,
    new_n19840, new_n19841, new_n19842, new_n19843, new_n19844, new_n19845,
    new_n19846, new_n19847, new_n19848, new_n19849, new_n19850, new_n19851,
    new_n19852, new_n19853, new_n19854, new_n19855, new_n19856, new_n19857,
    new_n19858, new_n19859, new_n19860, new_n19861, new_n19862, new_n19863,
    new_n19864, new_n19865, new_n19866, new_n19867, new_n19868, new_n19869,
    new_n19870, new_n19871, new_n19872, new_n19873_1, new_n19874,
    new_n19875, new_n19876, new_n19877, new_n19878, new_n19879, new_n19882,
    new_n19883, new_n19884, new_n19885, new_n19886, new_n19887, new_n19888,
    new_n19889, new_n19890, new_n19891, new_n19892, new_n19893, new_n19894,
    new_n19895, new_n19896, new_n19897, new_n19898, new_n19899, new_n19900,
    new_n19901, new_n19902, new_n19903, new_n19904, new_n19905_1,
    new_n19906, new_n19907, new_n19908, new_n19909_1, new_n19910,
    new_n19911_1, new_n19912, new_n19913, new_n19914, new_n19915,
    new_n19916_1, new_n19917, new_n19918, new_n19919, new_n19920,
    new_n19921, new_n19922_1, new_n19923_1, new_n19924, new_n19925,
    new_n19926, new_n19927, new_n19928, new_n19929, new_n19930_1,
    new_n19931, new_n19932, new_n19933, new_n19934, new_n19935, new_n19936,
    new_n19937, new_n19938, new_n19939, new_n19940, new_n19941_1,
    new_n19942, new_n19943, new_n19944, new_n19945, new_n19946, new_n19947,
    new_n19948, new_n19949, new_n19950, new_n19951, new_n19952, new_n19953,
    new_n19954, new_n19955, new_n19956, new_n19957, new_n19958, new_n19959,
    new_n19960, new_n19961, new_n19962, new_n19963, new_n19964, new_n19965,
    new_n19966, new_n19967, new_n19968_1, new_n19969, new_n19970,
    new_n19971, new_n19972, new_n19977, new_n19978, new_n19979, new_n19980,
    new_n19981, new_n19982, new_n19983, new_n19984, new_n19985, new_n19986,
    new_n19987, new_n19988_1, new_n19989, new_n19990, new_n19991,
    new_n19992, new_n19993, new_n19994, new_n19995, new_n19996, new_n19997,
    new_n19998, new_n19999, new_n20000, new_n20001, new_n20002, new_n20003,
    new_n20004_1, new_n20005, new_n20006, new_n20007, new_n20008,
    new_n20009, new_n20010, new_n20011, new_n20012, new_n20013_1,
    new_n20014, new_n20015, new_n20016, new_n20017_1, new_n20018,
    new_n20019, new_n20020, new_n20021, new_n20022, new_n20023, new_n20024,
    new_n20025, new_n20026, new_n20027, new_n20028, new_n20029, new_n20030,
    new_n20031, new_n20032, new_n20033_1, new_n20034, new_n20035,
    new_n20036_1, new_n20037, new_n20038, new_n20039, new_n20040_1,
    new_n20041, new_n20042, new_n20043, new_n20044, new_n20045, new_n20046,
    new_n20047, new_n20048, new_n20049, new_n20050, new_n20051, new_n20052,
    new_n20053, new_n20054, new_n20055, new_n20056, new_n20057, new_n20058,
    new_n20059, new_n20060, new_n20061_1, new_n20062, new_n20063,
    new_n20064, new_n20065, new_n20066, new_n20067, new_n20068,
    new_n20069_1, new_n20071, new_n20072, new_n20073, new_n20074,
    new_n20075, new_n20076, new_n20077_1, new_n20078, new_n20080,
    new_n20081, new_n20082, new_n20083, new_n20084, new_n20085,
    new_n20086_1, new_n20087, new_n20088, new_n20089, new_n20090,
    new_n20091, new_n20092, new_n20093, new_n20094, new_n20095,
    new_n20096_1, new_n20097, new_n20098, new_n20099, new_n20100,
    new_n20101, new_n20102, new_n20103_1, new_n20104, new_n20105,
    new_n20106, new_n20113, new_n20114, new_n20115, new_n20116, new_n20117,
    new_n20118, new_n20119, new_n20120, new_n20121, new_n20122, new_n20123,
    new_n20124, new_n20125, new_n20126_1, new_n20127, new_n20128,
    new_n20129, new_n20132, new_n20142, new_n20143, new_n20144, new_n20145,
    new_n20146, new_n20147, new_n20148, new_n20149_1, new_n20150,
    new_n20151_1, new_n20152, new_n20153, new_n20154, new_n20155,
    new_n20156, new_n20157, new_n20158, new_n20159, new_n20160, new_n20161,
    new_n20162, new_n20163, new_n20164, new_n20165, new_n20166, new_n20167,
    new_n20168, new_n20169_1, new_n20170, new_n20171, new_n20172,
    new_n20173, new_n20174, new_n20175, new_n20176, new_n20177, new_n20178,
    new_n20179_1, new_n20180, new_n20181, new_n20182, new_n20183,
    new_n20185, new_n20186, new_n20187_1, new_n20188, new_n20189,
    new_n20190, new_n20191, new_n20192, new_n20193, new_n20194, new_n20195,
    new_n20196, new_n20197, new_n20198, new_n20199, new_n20200, new_n20201,
    new_n20202, new_n20203, new_n20204, new_n20205, new_n20206, new_n20207,
    new_n20208, new_n20209, new_n20210, new_n20211, new_n20212, new_n20214,
    new_n20215, new_n20216, new_n20217, new_n20218, new_n20219, new_n20220,
    new_n20221, new_n20222, new_n20223, new_n20224, new_n20225, new_n20226,
    new_n20227, new_n20228, new_n20229, new_n20230, new_n20231, new_n20232,
    new_n20233, new_n20234, new_n20235_1, new_n20236, new_n20237,
    new_n20238, new_n20239, new_n20240, new_n20241, new_n20242, new_n20243,
    new_n20244, new_n20245, new_n20246, new_n20247, new_n20248, new_n20249,
    new_n20250_1, new_n20251, new_n20252, new_n20253, new_n20254,
    new_n20255, new_n20256, new_n20257, new_n20258, new_n20259_1,
    new_n20260, new_n20261, new_n20262, new_n20263, new_n20264, new_n20265,
    new_n20266, new_n20267, new_n20268, new_n20269, new_n20270, new_n20271,
    new_n20272, new_n20273, new_n20274, new_n20275, new_n20276, new_n20277,
    new_n20278, new_n20279_1, new_n20280, new_n20281, new_n20282,
    new_n20283, new_n20284, new_n20285, new_n20286, new_n20287_1,
    new_n20288, new_n20289, new_n20290, new_n20291, new_n20292, new_n20293,
    new_n20294, new_n20295, new_n20296, new_n20297, new_n20298, new_n20299,
    new_n20300, new_n20301_1, new_n20302, new_n20303, new_n20304,
    new_n20305, new_n20306, new_n20307, new_n20308, new_n20309, new_n20310,
    new_n20311, new_n20312, new_n20313, new_n20314, new_n20315, new_n20316,
    new_n20317, new_n20318, new_n20319, new_n20320, new_n20321, new_n20322,
    new_n20323, new_n20324, new_n20325, new_n20326, new_n20327, new_n20328,
    new_n20329, new_n20330_1, new_n20331, new_n20332, new_n20333_1,
    new_n20334, new_n20335, new_n20336, new_n20337, new_n20338, new_n20339,
    new_n20340, new_n20341, new_n20342, new_n20343, new_n20344, new_n20345,
    new_n20346, new_n20347, new_n20348, new_n20349_1, new_n20350,
    new_n20351, new_n20352, new_n20353, new_n20354, new_n20355_1,
    new_n20356, new_n20357, new_n20358, new_n20359_1, new_n20360,
    new_n20361, new_n20362, new_n20363, new_n20364, new_n20365,
    new_n20366_1, new_n20367, new_n20368, new_n20369, new_n20370,
    new_n20371, new_n20372, new_n20373, new_n20374, new_n20375, new_n20376,
    new_n20377, new_n20378, new_n20379, new_n20380, new_n20381, new_n20382,
    new_n20383, new_n20384, new_n20385_1, new_n20386, new_n20387,
    new_n20392, new_n20393, new_n20394, new_n20395, new_n20396, new_n20397,
    new_n20398, new_n20399, new_n20400, new_n20401, new_n20402_1,
    new_n20403_1, new_n20404, new_n20405, new_n20406, new_n20407,
    new_n20408, new_n20409_1, new_n20410, new_n20411_1, new_n20414,
    new_n20415, new_n20416, new_n20417, new_n20418, new_n20419, new_n20420,
    new_n20421, new_n20422, new_n20423, new_n20424_1, new_n20425,
    new_n20426, new_n20427, new_n20428, new_n20429_1, new_n20430,
    new_n20431, new_n20432, new_n20433, new_n20436_1, new_n20437,
    new_n20438, new_n20439, new_n20440, new_n20441_1, new_n20442,
    new_n20447, new_n20448, new_n20452, new_n20453, new_n20454,
    new_n20455_1, new_n20456, new_n20457, new_n20458, new_n20459,
    new_n20460, new_n20461, new_n20462, new_n20463, new_n20464, new_n20465,
    new_n20466, new_n20467, new_n20468, new_n20472, new_n20473, new_n20474,
    new_n20475, new_n20476, new_n20477, new_n20478_1, new_n20479,
    new_n20480, new_n20482, new_n20483, new_n20484, new_n20485, new_n20486,
    new_n20487, new_n20488, new_n20489_1, new_n20490_1, new_n20491,
    new_n20492, new_n20493, new_n20494, new_n20495_1, new_n20496,
    new_n20497, new_n20498, new_n20499, new_n20501, new_n20502, new_n20503,
    new_n20504, new_n20505, new_n20506, new_n20507, new_n20508, new_n20509,
    new_n20510, new_n20511, new_n20512, new_n20513, new_n20514,
    new_n20515_1, new_n20516, new_n20517, new_n20518, new_n20519,
    new_n20520, new_n20521, new_n20522, new_n20523, new_n20524, new_n20525,
    new_n20526, new_n20527, new_n20528, new_n20529, new_n20530, new_n20531,
    new_n20532, new_n20533_1, new_n20534, new_n20535, new_n20536,
    new_n20538, new_n20539, new_n20540, new_n20541, new_n20542, new_n20543,
    new_n20544, new_n20545, new_n20546, new_n20547, new_n20548, new_n20549,
    new_n20550, new_n20551, new_n20552, new_n20553, new_n20554, new_n20555,
    new_n20556, new_n20557, new_n20558, new_n20559, new_n20560, new_n20561,
    new_n20562, new_n20563, new_n20564, new_n20565, new_n20566, new_n20567,
    new_n20568, new_n20569, new_n20570, new_n20571, new_n20572, new_n20573,
    new_n20574, new_n20575, new_n20576, new_n20577, new_n20578, new_n20579,
    new_n20580, new_n20581, new_n20582_1, new_n20583, new_n20584,
    new_n20585, new_n20586, new_n20587, new_n20588, new_n20589,
    new_n20590_1, new_n20591, new_n20592, new_n20593, new_n20594,
    new_n20595, new_n20596, new_n20597, new_n20598, new_n20599, new_n20600,
    new_n20601, new_n20602_1, new_n20603, new_n20604_1, new_n20605,
    new_n20606, new_n20607, new_n20608, new_n20609_1, new_n20610,
    new_n20611, new_n20612, new_n20613, new_n20614, new_n20615, new_n20616,
    new_n20617, new_n20618, new_n20619, new_n20620, new_n20621, new_n20626,
    new_n20627, new_n20628, new_n20629_1, new_n20630, new_n20631,
    new_n20632, new_n20633, new_n20634, new_n20635, new_n20636, new_n20637,
    new_n20638, new_n20639, new_n20640, new_n20641, new_n20642, new_n20643,
    new_n20644, new_n20645, new_n20646, new_n20647, new_n20648, new_n20649,
    new_n20650, new_n20651, new_n20652, new_n20653, new_n20654, new_n20655,
    new_n20656, new_n20657, new_n20658_1, new_n20659, new_n20660,
    new_n20661_1, new_n20662, new_n20663, new_n20664, new_n20665,
    new_n20666, new_n20667, new_n20668, new_n20669, new_n20670, new_n20671,
    new_n20672, new_n20673_1, new_n20674, new_n20675, new_n20676,
    new_n20677, new_n20678_1, new_n20679, new_n20680_1, new_n20681,
    new_n20682, new_n20683, new_n20684, new_n20685_1, new_n20686,
    new_n20687, new_n20688, new_n20689, new_n20690, new_n20691_1,
    new_n20692, new_n20693, new_n20694, new_n20695, new_n20696_1,
    new_n20697, new_n20698, new_n20699, new_n20700_1, new_n20701,
    new_n20702, new_n20703, new_n20704_1, new_n20705_1, new_n20706,
    new_n20707, new_n20708, new_n20709_1, new_n20710, new_n20711,
    new_n20712, new_n20713_1, new_n20714, new_n20715, new_n20716,
    new_n20717, new_n20718, new_n20719, new_n20720, new_n20721,
    new_n20722_1, new_n20723_1, new_n20724, new_n20725, new_n20726,
    new_n20727, new_n20728, new_n20729, new_n20730, new_n20731, new_n20732,
    new_n20733, new_n20734, new_n20735, new_n20736, new_n20737, new_n20738,
    new_n20739, new_n20740, new_n20742, new_n20743, new_n20748_1,
    new_n20751, new_n20752, new_n20753, new_n20754, new_n20755, new_n20756,
    new_n20757, new_n20758, new_n20759, new_n20760, new_n20761_1,
    new_n20762, new_n20763, new_n20764, new_n20765, new_n20766, new_n20767,
    new_n20768, new_n20769, new_n20770, new_n20771, new_n20772, new_n20773,
    new_n20774_1, new_n20775, new_n20776, new_n20777, new_n20778,
    new_n20779, new_n20780, new_n20781, new_n20782, new_n20783, new_n20784,
    new_n20786, new_n20787, new_n20788_1, new_n20789, new_n20790,
    new_n20791, new_n20792, new_n20793, new_n20794_1, new_n20795_1,
    new_n20796, new_n20797, new_n20798, new_n20799, new_n20800, new_n20801,
    new_n20802, new_n20803_1, new_n20804, new_n20805, new_n20806,
    new_n20807, new_n20808, new_n20809, new_n20810, new_n20811, new_n20812,
    new_n20813, new_n20814, new_n20815, new_n20824, new_n20825,
    new_n20826_1, new_n20827, new_n20828, new_n20829, new_n20830,
    new_n20831, new_n20832, new_n20833, new_n20834, new_n20835, new_n20839,
    new_n20840, new_n20841, new_n20842, new_n20843, new_n20844, new_n20845,
    new_n20846, new_n20847, new_n20848, new_n20849, new_n20850, new_n20851,
    new_n20852, new_n20853, new_n20854, new_n20855, new_n20856, new_n20857,
    new_n20858, new_n20859, new_n20860, new_n20861, new_n20862, new_n20863,
    new_n20864, new_n20865, new_n20866, new_n20867, new_n20868,
    new_n20869_1, new_n20872, new_n20873, new_n20874, new_n20875,
    new_n20876, new_n20877, new_n20878, new_n20879_1, new_n20880,
    new_n20881, new_n20882, new_n20883, new_n20884, new_n20885, new_n20886,
    new_n20887, new_n20888, new_n20889, new_n20890, new_n20891, new_n20892,
    new_n20893, new_n20894, new_n20895, new_n20896, new_n20897, new_n20898,
    new_n20899, new_n20900, new_n20901, new_n20902, new_n20903, new_n20904,
    new_n20905, new_n20906, new_n20907, new_n20908, new_n20909, new_n20910,
    new_n20911, new_n20912, new_n20913, new_n20914, new_n20915_1,
    new_n20916, new_n20917, new_n20918, new_n20919, new_n20920, new_n20921,
    new_n20922, new_n20923_1, new_n20924, new_n20925, new_n20926,
    new_n20927, new_n20928, new_n20929_1, new_n20930, new_n20931,
    new_n20932, new_n20933, new_n20934, new_n20936_1, new_n20937,
    new_n20938, new_n20939, new_n20940, new_n20941, new_n20942, new_n20943,
    new_n20944, new_n20945, new_n20946_1, new_n20947, new_n20948,
    new_n20949, new_n20950, new_n20951, new_n20952, new_n20953, new_n20954,
    new_n20955, new_n20956, new_n20957, new_n20958, new_n20959, new_n20960,
    new_n20961, new_n20962, new_n20963, new_n20964, new_n20965, new_n20966,
    new_n20967, new_n20968, new_n20970, new_n20971, new_n20973, new_n20974,
    new_n20975, new_n20976, new_n20977, new_n20978, new_n20979, new_n20980,
    new_n20981, new_n20982, new_n20983, new_n20984, new_n20985,
    new_n20986_1, new_n20987, new_n20988, new_n20989, new_n20990,
    new_n20991, new_n20992, new_n20993, new_n20994, new_n20995, new_n20996,
    new_n20997, new_n20998, new_n20999, new_n21000, new_n21001, new_n21002,
    new_n21003, new_n21004, new_n21005, new_n21006, new_n21007, new_n21010,
    new_n21011, new_n21014, new_n21015, new_n21016, new_n21017_1,
    new_n21018, new_n21019, new_n21020, new_n21021, new_n21022, new_n21023,
    new_n21024, new_n21025, new_n21026, new_n21027, new_n21028, new_n21029,
    new_n21030, new_n21031, new_n21032, new_n21033, new_n21034_1,
    new_n21035, new_n21036, new_n21037, new_n21038, new_n21039, new_n21040,
    new_n21041, new_n21042, new_n21043, new_n21044, new_n21045,
    new_n21046_1, new_n21047, new_n21048, new_n21049, new_n21050,
    new_n21051, new_n21052, new_n21055, new_n21056, new_n21057, new_n21058,
    new_n21059, new_n21060, new_n21061, new_n21062_1, new_n21063,
    new_n21064, new_n21065, new_n21066, new_n21067, new_n21068, new_n21069,
    new_n21070, new_n21071, new_n21072, new_n21073, new_n21074, new_n21075,
    new_n21076, new_n21077, new_n21078_1, new_n21086, new_n21087,
    new_n21088, new_n21089, new_n21090, new_n21091, new_n21092,
    new_n21093_1, new_n21094_1, new_n21095_1, new_n21096, new_n21097,
    new_n21098, new_n21099, new_n21100, new_n21101, new_n21102, new_n21103,
    new_n21104, new_n21105, new_n21106, new_n21107, new_n21108, new_n21109,
    new_n21110, new_n21111, new_n21112, new_n21113, new_n21114, new_n21115,
    new_n21116, new_n21117, new_n21118, new_n21119, new_n21120, new_n21121,
    new_n21122, new_n21123_1, new_n21124, new_n21125, new_n21126,
    new_n21127, new_n21128, new_n21129, new_n21130, new_n21131, new_n21132,
    new_n21133, new_n21134_1, new_n21135, new_n21136, new_n21137,
    new_n21138_1, new_n21139, new_n21140, new_n21141, new_n21142,
    new_n21143, new_n21150, new_n21154_1, new_n21155, new_n21156,
    new_n21157_1, new_n21158, new_n21159, new_n21160, new_n21161,
    new_n21162, new_n21163, new_n21164, new_n21180, new_n21182_1,
    new_n21183, new_n21184, new_n21185, new_n21186, new_n21187, new_n21188,
    new_n21189, new_n21190, new_n21191, new_n21192, new_n21193_1,
    new_n21194, new_n21195, new_n21196, new_n21197, new_n21198, new_n21199,
    new_n21200, new_n21201, new_n21202, new_n21203_1, new_n21204,
    new_n21206, new_n21207, new_n21208, new_n21209, new_n21210, new_n21211,
    new_n21212, new_n21213, new_n21214, new_n21215, new_n21216, new_n21217,
    new_n21218, new_n21219, new_n21220, new_n21221, new_n21222_1,
    new_n21223, new_n21224, new_n21226_1, new_n21227, new_n21228,
    new_n21229, new_n21230, new_n21231, new_n21232, new_n21233, new_n21234,
    new_n21235, new_n21236, new_n21237, new_n21238_1, new_n21239,
    new_n21240, new_n21241, new_n21246, new_n21247, new_n21248, new_n21249,
    new_n21250, new_n21251, new_n21252, new_n21253, new_n21254_1,
    new_n21255, new_n21256, new_n21257, new_n21258, new_n21259, new_n21260,
    new_n21261, new_n21262, new_n21263, new_n21264, new_n21267, new_n21274,
    new_n21275, new_n21276_1, new_n21277, new_n21278, new_n21279,
    new_n21280, new_n21286, new_n21287_1, new_n21288, new_n21289,
    new_n21290, new_n21291, new_n21292, new_n21293, new_n21294, new_n21295,
    new_n21300, new_n21306, new_n21307, new_n21308, new_n21309, new_n21310,
    new_n21311, new_n21312, new_n21313, new_n21314, new_n21315, new_n21316,
    new_n21317_1, new_n21318, new_n21319, new_n21320, new_n21321,
    new_n21322, new_n21327, new_n21328, new_n21329, new_n21330, new_n21331,
    new_n21332, new_n21339, new_n21340, new_n21341, new_n21342, new_n21343,
    new_n21344, new_n21345, new_n21346, new_n21347, new_n21348,
    new_n21349_1, new_n21350, new_n21351, new_n21352, new_n21353,
    new_n21354, new_n21355, new_n21356, new_n21357, new_n21358, new_n21359,
    new_n21360, new_n21361, new_n21362, new_n21363, new_n21364,
    new_n21365_1, new_n21366, new_n21367_1, new_n21368, new_n21369,
    new_n21370, new_n21371, new_n21372, new_n21373, new_n21374, new_n21375,
    new_n21376, new_n21377, new_n21378, new_n21379, new_n21380, new_n21381,
    new_n21382, new_n21385, new_n21386, new_n21387, new_n21388, new_n21389,
    new_n21390, new_n21391, new_n21392, new_n21393, new_n21395,
    new_n21396_1, new_n21397, new_n21398_1, new_n21399_1, new_n21400,
    new_n21401, new_n21402, new_n21403, new_n21404_1, new_n21405,
    new_n21406, new_n21407, new_n21408, new_n21409, new_n21410, new_n21411,
    new_n21421, new_n21422, new_n21423, new_n21424, new_n21425, new_n21426,
    new_n21427, new_n21428, new_n21429, new_n21430, new_n21431, new_n21432,
    new_n21433, new_n21434, new_n21435, new_n21436, new_n21437, new_n21438,
    new_n21439, new_n21440, new_n21441, new_n21442, new_n21443, new_n21444,
    new_n21445, new_n21446_1, new_n21447, new_n21448, new_n21449,
    new_n21450, new_n21451, new_n21452, new_n21453, new_n21459, new_n21460,
    new_n21461, new_n21462, new_n21472_1, new_n21473, new_n21474,
    new_n21475, new_n21476, new_n21477, new_n21478, new_n21479, new_n21480,
    new_n21481, new_n21482, new_n21483, new_n21484, new_n21485, new_n21486,
    new_n21487, new_n21488, new_n21489_1, new_n21490, new_n21491,
    new_n21492, new_n21493, new_n21494, new_n21495, new_n21496, new_n21497,
    new_n21498, new_n21499, new_n21500, new_n21501, new_n21502, new_n21503,
    new_n21504, new_n21505, new_n21506, new_n21507, new_n21508, new_n21509,
    new_n21510, new_n21511, new_n21512, new_n21513, new_n21514, new_n21515,
    new_n21516, new_n21517, new_n21518, new_n21519, new_n21520, new_n21521,
    new_n21522, new_n21523, new_n21524, new_n21525_1, new_n21526,
    new_n21527, new_n21528, new_n21529, new_n21530, new_n21531, new_n21532,
    new_n21533, new_n21534, new_n21535, new_n21536, new_n21537,
    new_n21538_1, new_n21539, new_n21540, new_n21541, new_n21542,
    new_n21543, new_n21544, new_n21546, new_n21547, new_n21548,
    new_n21549_1, new_n21550, new_n21551, new_n21552, new_n21553,
    new_n21554, new_n21555, new_n21556, new_n21557, new_n21558, new_n21559,
    new_n21560, new_n21561, new_n21562, new_n21563, new_n21564, new_n21565,
    new_n21566, new_n21567, new_n21568, new_n21569, new_n21570, new_n21571,
    new_n21572, new_n21573, new_n21574, new_n21575, new_n21576, new_n21577,
    new_n21578, new_n21579, new_n21580, new_n21581, new_n21582, new_n21583,
    new_n21584, new_n21585, new_n21586, new_n21587, new_n21588, new_n21589,
    new_n21590, new_n21591, new_n21592, new_n21593, new_n21594, new_n21595,
    new_n21596, new_n21597, new_n21598, new_n21599_1, new_n21600,
    new_n21601, new_n21602, new_n21603, new_n21604, new_n21605, new_n21606,
    new_n21607, new_n21608, new_n21609, new_n21610, new_n21611, new_n21612,
    new_n21613, new_n21614, new_n21617, new_n21618, new_n21619, new_n21620,
    new_n21621, new_n21622, new_n21623, new_n21624, new_n21625, new_n21626,
    new_n21627, new_n21628_1, new_n21629, new_n21635, new_n21636,
    new_n21637_1, new_n21638, new_n21639, new_n21640, new_n21641,
    new_n21642, new_n21643, new_n21644, new_n21645_1, new_n21646,
    new_n21647, new_n21648, new_n21649_1, new_n21650, new_n21651,
    new_n21652, new_n21653, new_n21654_1, new_n21655, new_n21656,
    new_n21657, new_n21658, new_n21659, new_n21660, new_n21661, new_n21662,
    new_n21663, new_n21664, new_n21665_1, new_n21666, new_n21667,
    new_n21668, new_n21669, new_n21670, new_n21671, new_n21672, new_n21673,
    new_n21674_1, new_n21675, new_n21676, new_n21677, new_n21678,
    new_n21679, new_n21680_1, new_n21681, new_n21682, new_n21683,
    new_n21684, new_n21685_1, new_n21686, new_n21687_1, new_n21688,
    new_n21689, new_n21690, new_n21691, new_n21692, new_n21693, new_n21694,
    new_n21695, new_n21696, new_n21697, new_n21698, new_n21699, new_n21700,
    new_n21701, new_n21702, new_n21703, new_n21704, new_n21705, new_n21706,
    new_n21708, new_n21709, new_n21710, new_n21711, new_n21712, new_n21713,
    new_n21714, new_n21715, new_n21716, new_n21717_1, new_n21720,
    new_n21721, new_n21722, new_n21723, new_n21724, new_n21725, new_n21726,
    new_n21727, new_n21728, new_n21729, new_n21735_1, new_n21736,
    new_n21737, new_n21738, new_n21739, new_n21740, new_n21741, new_n21742,
    new_n21743, new_n21744, new_n21745, new_n21746, new_n21747, new_n21748,
    new_n21749_1, new_n21750_1, new_n21751, new_n21752, new_n21753_1,
    new_n21754, new_n21755, new_n21756, new_n21757, new_n21758, new_n21759,
    new_n21760, new_n21761, new_n21762, new_n21763, new_n21764,
    new_n21765_1, new_n21766, new_n21767, new_n21768, new_n21769,
    new_n21770, new_n21771, new_n21772, new_n21773, new_n21774, new_n21775,
    new_n21776, new_n21777, new_n21778, new_n21779_1, new_n21780,
    new_n21781, new_n21782, new_n21783, new_n21784_1, new_n21785,
    new_n21786, new_n21787, new_n21788, new_n21789, new_n21790, new_n21791,
    new_n21792, new_n21793, new_n21794, new_n21795, new_n21796, new_n21797,
    new_n21798, new_n21799, new_n21800_1, new_n21801, new_n21802,
    new_n21810, new_n21811, new_n21812, new_n21813, new_n21814, new_n21819,
    new_n21822, new_n21824, new_n21825, new_n21826, new_n21827, new_n21828,
    new_n21829, new_n21830, new_n21831, new_n21832_1, new_n21833,
    new_n21834, new_n21835, new_n21836, new_n21837, new_n21838,
    new_n21839_1, new_n21840, new_n21841, new_n21842, new_n21843,
    new_n21844, new_n21845, new_n21846, new_n21847, new_n21848, new_n21849,
    new_n21850, new_n21851, new_n21852, new_n21853, new_n21854, new_n21855,
    new_n21856, new_n21857, new_n21858, new_n21859, new_n21860, new_n21861,
    new_n21862, new_n21863, new_n21864, new_n21865, new_n21866, new_n21867,
    new_n21868, new_n21869, new_n21872, new_n21873, new_n21874_1,
    new_n21875, new_n21883, new_n21884, new_n21885, new_n21886, new_n21887,
    new_n21888, new_n21889, new_n21890, new_n21891, new_n21895, new_n21903,
    new_n21904, new_n21905_1, new_n21906, new_n21907, new_n21908,
    new_n21909, new_n21910, new_n21911, new_n21912, new_n21913, new_n21914,
    new_n21915_1, new_n21916, new_n21918, new_n21919, new_n21920,
    new_n21921, new_n21922, new_n21923, new_n21924, new_n21925, new_n21926,
    new_n21927, new_n21928, new_n21929, new_n21930, new_n21931, new_n21932,
    new_n21933, new_n21934_1, new_n21940, new_n21941, new_n21942,
    new_n21943_1, new_n21944, new_n21945, new_n21946, new_n21947,
    new_n21948, new_n21949, new_n21950, new_n21951, new_n21952, new_n21953,
    new_n21954, new_n21955, new_n21956, new_n21957_1, new_n21958,
    new_n21959, new_n21960_1, new_n21961, new_n21962, new_n21963,
    new_n21964, new_n21965, new_n21966, new_n21967, new_n21968, new_n21969,
    new_n21972, new_n21973, new_n21974, new_n21975, new_n21976_1,
    new_n21977, new_n21978, new_n21979, new_n21980, new_n21981_1,
    new_n21982, new_n21983, new_n21984, new_n21985, new_n21986_1,
    new_n21987, new_n21988, new_n21989, new_n21990, new_n21991, new_n21992,
    new_n21993_1, new_n21994, new_n21996, new_n21997_1, new_n21998,
    new_n21999, new_n22000, new_n22001, new_n22002, new_n22003, new_n22004,
    new_n22005, new_n22006, new_n22007, new_n22008, new_n22009, new_n22013,
    new_n22015, new_n22016_1, new_n22021, new_n22022, new_n22023,
    new_n22024, new_n22025, new_n22026, new_n22027_1, new_n22028,
    new_n22029, new_n22030, new_n22031, new_n22032, new_n22033, new_n22034,
    new_n22035, new_n22036, new_n22037, new_n22038, new_n22039, new_n22040,
    new_n22041, new_n22042, new_n22043_1, new_n22044, new_n22045,
    new_n22046, new_n22047, new_n22048, new_n22049, new_n22050_1,
    new_n22051, new_n22052, new_n22053, new_n22054, new_n22055, new_n22056,
    new_n22057, new_n22058, new_n22059, new_n22060, new_n22061, new_n22062,
    new_n22063_1, new_n22064, new_n22065, new_n22067, new_n22068_1,
    new_n22069, new_n22070, new_n22071, new_n22072_1, new_n22073,
    new_n22074, new_n22075, new_n22076_1, new_n22077, new_n22078,
    new_n22079, new_n22080, new_n22081, new_n22082, new_n22083, new_n22084,
    new_n22085, new_n22086, new_n22087, new_n22088, new_n22089,
    new_n22090_1, new_n22091, new_n22092, new_n22093, new_n22094,
    new_n22095, new_n22096, new_n22097, new_n22098, new_n22099, new_n22100,
    new_n22101, new_n22102, new_n22103, new_n22104, new_n22105, new_n22106,
    new_n22107_1, new_n22108, new_n22109, new_n22110, new_n22111,
    new_n22112, new_n22113_1, new_n22114, new_n22115, new_n22116,
    new_n22117, new_n22123, new_n22132, new_n22133, new_n22134, new_n22135,
    new_n22141, new_n22148, new_n22149, new_n22150_1, new_n22151,
    new_n22152, new_n22153, new_n22154, new_n22155, new_n22156,
    new_n22157_1, new_n22158, new_n22159, new_n22160, new_n22161,
    new_n22162, new_n22163, new_n22164, new_n22165, new_n22166, new_n22167,
    new_n22168, new_n22169, new_n22170, new_n22171, new_n22172,
    new_n22173_1, new_n22174, new_n22175, new_n22176, new_n22177,
    new_n22178, new_n22179, new_n22180, new_n22181, new_n22182, new_n22183,
    new_n22184, new_n22187, new_n22188, new_n22189, new_n22190, new_n22191,
    new_n22192, new_n22193, new_n22194, new_n22195, new_n22196, new_n22197,
    new_n22198_1, new_n22205, new_n22206, new_n22207, new_n22208,
    new_n22209, new_n22210, new_n22211, new_n22212, new_n22213_1,
    new_n22214, new_n22215, new_n22216, new_n22217, new_n22218, new_n22219,
    new_n22220, new_n22221, new_n22222, new_n22223, new_n22224, new_n22225,
    new_n22226, new_n22227, new_n22228, new_n22229, new_n22230, new_n22231,
    new_n22232, new_n22233, new_n22234, new_n22235, new_n22236, new_n22237,
    new_n22238, new_n22239, new_n22240, new_n22241, new_n22242, new_n22243,
    new_n22244, new_n22245, new_n22246, new_n22247, new_n22248, new_n22249,
    new_n22250, new_n22251, new_n22252, new_n22253_1, new_n22254,
    new_n22255, new_n22256, new_n22257, new_n22258, new_n22259, new_n22260,
    new_n22261, new_n22262, new_n22263, new_n22264, new_n22265, new_n22266,
    new_n22267, new_n22268, new_n22269, new_n22270_1, new_n22271,
    new_n22272, new_n22273, new_n22274_1, new_n22275, new_n22276,
    new_n22277, new_n22278, new_n22279, new_n22280, new_n22281, new_n22282,
    new_n22283_1, new_n22284, new_n22285, new_n22286, new_n22287,
    new_n22288, new_n22289, new_n22290_1, new_n22291, new_n22292,
    new_n22293, new_n22294, new_n22295, new_n22296, new_n22297, new_n22298,
    new_n22299, new_n22300, new_n22301, new_n22302, new_n22303, new_n22304,
    new_n22305, new_n22306, new_n22307, new_n22308, new_n22309_1,
    new_n22310, new_n22311_1, new_n22312, new_n22313, new_n22314,
    new_n22315, new_n22316, new_n22317_1, new_n22318, new_n22319,
    new_n22320, new_n22321, new_n22322, new_n22323, new_n22324, new_n22325,
    new_n22326, new_n22327, new_n22328, new_n22329, new_n22330, new_n22331,
    new_n22332_1, new_n22333, new_n22337, new_n22340, new_n22341_1,
    new_n22342, new_n22343, new_n22344, new_n22345, new_n22346, new_n22347,
    new_n22348, new_n22349, new_n22350, new_n22351, new_n22352,
    new_n22353_1, new_n22354, new_n22355, new_n22360, new_n22361,
    new_n22362, new_n22363, new_n22364, new_n22365, new_n22366, new_n22367,
    new_n22368, new_n22369, new_n22370, new_n22371, new_n22372, new_n22373,
    new_n22374, new_n22375, new_n22376, new_n22377, new_n22378,
    new_n22379_1, new_n22380, new_n22381, new_n22382, new_n22383,
    new_n22384, new_n22386, new_n22387, new_n22388, new_n22389, new_n22390,
    new_n22391, new_n22395, new_n22396, new_n22397, new_n22398, new_n22404,
    new_n22409, new_n22410, new_n22411, new_n22412, new_n22413, new_n22414,
    new_n22415, new_n22416, new_n22417, new_n22418, new_n22419, new_n22420,
    new_n22421, new_n22422, new_n22423, new_n22424, new_n22425, new_n22426,
    new_n22427, new_n22428, new_n22429, new_n22430, new_n22431, new_n22452,
    new_n22453, new_n22454, new_n22455, new_n22456, new_n22457, new_n22458,
    new_n22459, new_n22460, new_n22461, new_n22462, new_n22463, new_n22464,
    new_n22465, new_n22466, new_n22467_1, new_n22468, new_n22469,
    new_n22470_1, new_n22471, new_n22472, new_n22473, new_n22474,
    new_n22475, new_n22476, new_n22477, new_n22478, new_n22479, new_n22480,
    new_n22481, new_n22482, new_n22483, new_n22484_1, new_n22485,
    new_n22486, new_n22487, new_n22495, new_n22496, new_n22497, new_n22498,
    new_n22499, new_n22500, new_n22501, new_n22502, new_n22503, new_n22504,
    new_n22505, new_n22506, new_n22507, new_n22508, new_n22512, new_n22513,
    new_n22516, new_n22517, new_n22518, new_n22519, new_n22520, new_n22521,
    new_n22522, new_n22523, new_n22526, new_n22527, new_n22528, new_n22529,
    new_n22530, new_n22531, new_n22532, new_n22533_1, new_n22534,
    new_n22535, new_n22536, new_n22537, new_n22538, new_n22539, new_n22540,
    new_n22541, new_n22542, new_n22543, new_n22544, new_n22545, new_n22546,
    new_n22547, new_n22550, new_n22551, new_n22552, new_n22553,
    new_n22554_1, new_n22555, new_n22556, new_n22557, new_n22558,
    new_n22559, new_n22560, new_n22561, new_n22562, new_n22563, new_n22564,
    new_n22565, new_n22566, new_n22567, new_n22568, new_n22569, new_n22570,
    new_n22571, new_n22572, new_n22573, new_n22574, new_n22575, new_n22576,
    new_n22577, new_n22578, new_n22579, new_n22580, new_n22581, new_n22582,
    new_n22583, new_n22584_1, new_n22585, new_n22586, new_n22587,
    new_n22608, new_n22612, new_n22613, new_n22614, new_n22615, new_n22616,
    new_n22617, new_n22618, new_n22619_1, new_n22620_1, new_n22621,
    new_n22622, new_n22623_1, new_n22624, new_n22625, new_n22628,
    new_n22629, new_n22630, new_n22631_1, new_n22632, new_n22633,
    new_n22634, new_n22635, new_n22636, new_n22637, new_n22638, new_n22639,
    new_n22640, new_n22641, new_n22642, new_n22643, new_n22644, new_n22645,
    new_n22646, new_n22647, new_n22651, new_n22652, new_n22653, new_n22654,
    new_n22655, new_n22656, new_n22657, new_n22661, new_n22664, new_n22667,
    new_n22668, new_n22669, new_n22670, new_n22671, new_n22672, new_n22673,
    new_n22675, new_n22676, new_n22677, new_n22678, new_n22679, new_n22680,
    new_n22681, new_n22682, new_n22683, new_n22684, new_n22685, new_n22686,
    new_n22687, new_n22688, new_n22689, new_n22690, new_n22691, new_n22692,
    new_n22693, new_n22714_1, new_n22717, new_n22718, new_n22719,
    new_n22720, new_n22721, new_n22722, new_n22723, new_n22724, new_n22725,
    new_n22726, new_n22727, new_n22728, new_n22729, new_n22730, new_n22731,
    new_n22732, new_n22733, new_n22734, new_n22735, new_n22736, new_n22737,
    new_n22742, new_n22743, new_n22744, new_n22745, new_n22757, new_n22760,
    new_n22775, new_n22776, new_n22777, new_n22778, new_n22779_1,
    new_n22780, new_n22794, new_n22795, new_n22796, new_n22797, new_n22798,
    new_n22799, new_n22800, new_n22804, new_n22805, new_n22806, new_n22807,
    new_n22808, new_n22809, new_n22810, new_n22815, new_n22816, new_n22817,
    new_n22818, new_n22819_1, new_n22820, new_n22821, new_n22822,
    new_n22823, new_n22826, new_n22827, new_n22842, new_n22843_1,
    new_n22844, new_n22847, new_n22848, new_n22849, new_n22850,
    new_n22858_1, new_n22859, new_n22868, new_n22874, new_n22879_1,
    new_n22880, new_n22881, new_n22882, new_n22883, new_n22884, new_n22885,
    new_n22886, new_n22887, new_n22888, new_n22896, new_n22898, new_n22899,
    new_n22900, new_n22901, new_n22902, new_n22903_1, new_n22904,
    new_n22905, new_n22906, new_n22907_1, new_n22909, new_n22910_1,
    new_n22911, new_n22912, new_n22923, new_n22924, new_n22926, new_n22927,
    new_n22928, new_n22929, new_n22930, new_n22931, new_n22932, new_n22933,
    new_n22934, new_n22935, new_n22936, new_n22937, new_n22938,
    new_n22939_1, new_n22957, new_n22958, new_n22959, new_n22960,
    new_n22961, new_n22962, new_n22963, new_n22964, new_n22965, new_n22966,
    new_n22967, new_n22968, new_n22969, new_n22972, new_n22973, new_n22974,
    new_n22975, new_n22979, new_n22981, new_n22982, new_n22983, new_n22984,
    new_n22985, new_n22986, new_n22987, new_n22988, new_n22991, new_n22992,
    new_n22993, new_n22994, new_n22995, new_n22998_1, new_n22999,
    new_n23000, new_n23001, new_n23002, new_n23004, new_n23005,
    new_n23006_1, new_n23007_1, new_n23008, new_n23009_1, new_n23010,
    new_n23011, new_n23012, new_n23013, new_n23014_1, new_n23015,
    new_n23016, new_n23017, new_n23018, new_n23019, new_n23020, new_n23021,
    new_n23022, new_n23023, new_n23024, new_n23025, new_n23026, new_n23030,
    new_n23031, new_n23032, new_n23033, new_n23034, new_n23035_1,
    new_n23049, new_n23050, new_n23061, new_n23068_1, new_n23069,
    new_n23070, new_n23071, new_n23072, new_n23073, new_n23081, new_n23100,
    new_n23122, new_n23123, new_n23137, new_n23138, new_n23139, new_n23140,
    new_n23141, new_n23142, new_n23143, new_n23144, new_n23151, new_n23159,
    new_n23160_1, new_n23161, new_n23162, new_n23163, new_n23164,
    new_n23165, new_n23166_1, new_n23167, new_n23168, new_n23169,
    new_n23170, new_n23176, new_n23177, new_n23178, new_n23179, new_n23180,
    new_n23181, new_n23182, new_n23183, new_n23184, new_n23187, new_n23188,
    new_n23189, new_n23190, new_n23196, new_n23197, new_n23198, new_n23199,
    new_n23201, new_n23202, new_n23203, new_n23204, new_n23205, new_n23206,
    new_n23207, new_n23208, new_n23209, new_n23210, new_n23211, new_n23212,
    new_n23213, new_n23214, new_n23215, new_n23227, new_n23255, new_n23256,
    new_n23257, new_n23258, new_n23269, new_n23275, new_n23276, new_n23277,
    new_n23278, new_n23279, new_n23294, new_n23301, new_n23302, new_n23303,
    new_n23304_1, new_n23305_1, new_n23306, new_n23307, new_n23308,
    new_n23323, new_n23324, new_n23325, new_n23326, new_n23327, new_n23328,
    new_n23329, new_n23330, new_n23335, new_n23341_1, new_n23342_1,
    new_n23343, new_n23344, new_n23345, new_n23346, new_n23347, new_n23348,
    new_n23349, new_n23350, new_n23363, new_n23364, new_n23365,
    new_n23369_1, new_n23374, new_n23375, new_n23376, new_n23377,
    new_n23384, new_n23385, new_n23386, new_n23387, new_n23388, new_n23389,
    new_n23390, new_n23396, new_n23397, new_n23405, new_n23406, new_n23407,
    new_n23408, new_n23409, new_n23412, new_n23415, new_n23416, new_n23417,
    new_n23418, new_n23431, new_n23432, new_n23433_1, new_n23434_1,
    new_n23436, new_n23447, new_n23448, new_n23449, new_n23450_1,
    new_n23453, new_n23461, new_n23462, new_n23463_1, new_n23464,
    new_n23465, new_n23466, new_n23467, new_n23468, new_n23469,
    new_n23471_1, new_n23476, new_n23477, new_n23478, new_n23479,
    new_n23481, new_n23482, new_n23483, new_n23484, new_n23489, new_n23490,
    new_n23491, new_n23492, new_n23493_1, new_n23494, new_n23495,
    new_n23496, new_n23497, new_n23498, new_n23499, new_n23500, new_n23501,
    new_n23502, new_n23503, new_n23504, new_n23505, new_n23506, new_n23507,
    new_n23508, new_n23509, new_n23510, new_n23515, new_n23516, new_n23517,
    new_n23518, new_n23522, new_n23532, new_n23533, new_n23534, new_n23535,
    new_n23536, new_n23555, new_n23556, new_n23557, new_n23558, new_n23559,
    new_n23560, new_n23562, new_n23563, new_n23564, new_n23565, new_n23566,
    new_n23567, new_n23578, new_n23590, new_n23591, new_n23595, new_n23596,
    new_n23597, new_n23598, new_n23600, new_n23601, new_n23603, new_n23613,
    new_n23614, new_n23615, new_n23616, new_n23617, new_n23626,
    new_n23637_1, new_n23646, new_n23655, new_n23656, new_n23666,
    new_n23667, new_n23668, new_n23669_1, new_n23675, new_n23676,
    new_n23677, new_n23678, new_n23681, new_n23682, new_n23683,
    new_n23684_1, new_n23705, new_n23725, new_n23735, new_n23736,
    new_n23737, new_n23751, new_n23752, new_n23767, new_n23783, new_n23788,
    new_n23791, new_n23792, new_n23798, new_n23799, new_n23800, new_n23804,
    new_n23805, new_n23806, new_n23807, new_n23809, new_n23822, new_n23825,
    new_n23826, new_n23827, new_n23828, new_n23831_1, new_n23834,
    new_n23835, new_n23836, new_n23837, new_n23851, new_n23852, new_n23855,
    new_n23867, new_n23869, new_n23870, new_n23871, new_n23872, new_n23875,
    new_n23876, new_n23886, new_n23888_1, new_n23893, new_n23894,
    new_n23895_1, new_n23896, new_n23902, new_n23903_1, new_n23913_1,
    new_n23927, new_n23936, new_n23937, new_n23940;
  xnor_4 g00000(.A(n10739), .B(n9942), .Y(new_n2349));
  not_8  g00001(.A(n21753), .Y(new_n2350));
  nor_5  g00002(.A(n25643), .B(new_n2350), .Y(new_n2351));
  xnor_4 g00003(.A(n25643), .B(n21753), .Y(new_n2352));
  not_8  g00004(.A(n21832), .Y(new_n2353));
  nor_5  g00005(.A(new_n2353), .B(n9557), .Y(new_n2354));
  xnor_4 g00006(.A(n21832), .B(n9557), .Y(new_n2355_1));
  not_8  g00007(.A(n26913), .Y(new_n2356));
  nor_5  g00008(.A(new_n2356), .B(n3136), .Y(new_n2357));
  xnor_4 g00009(.A(n26913), .B(n3136), .Y(new_n2358));
  not_8  g00010(.A(n6385), .Y(new_n2359));
  nor_5  g00011(.A(n16223), .B(new_n2359), .Y(new_n2360));
  not_8  g00012(.A(n16223), .Y(new_n2361_1));
  nor_5  g00013(.A(new_n2361_1), .B(n6385), .Y(new_n2362));
  not_8  g00014(.A(n20138), .Y(new_n2363_1));
  nor_5  g00015(.A(new_n2363_1), .B(n19494), .Y(new_n2364));
  not_8  g00016(.A(n19494), .Y(new_n2365));
  nor_5  g00017(.A(n20138), .B(new_n2365), .Y(new_n2366));
  not_8  g00018(.A(n9251), .Y(new_n2367));
  nor_5  g00019(.A(new_n2367), .B(n2387), .Y(new_n2368));
  not_8  g00020(.A(new_n2368), .Y(new_n2369));
  nor_5  g00021(.A(new_n2369), .B(new_n2366), .Y(new_n2370));
  nor_5  g00022(.A(new_n2370), .B(new_n2364), .Y(new_n2371));
  nor_5  g00023(.A(new_n2371), .B(new_n2362), .Y(new_n2372));
  nor_5  g00024(.A(new_n2372), .B(new_n2360), .Y(new_n2373));
  and_5  g00025(.A(new_n2373), .B(new_n2358), .Y(new_n2374_1));
  or_5   g00026(.A(new_n2374_1), .B(new_n2357), .Y(new_n2375));
  and_5  g00027(.A(new_n2375), .B(new_n2355_1), .Y(new_n2376));
  or_5   g00028(.A(new_n2376), .B(new_n2354), .Y(new_n2377));
  and_5  g00029(.A(new_n2377), .B(new_n2352), .Y(new_n2378));
  or_5   g00030(.A(new_n2378), .B(new_n2351), .Y(new_n2379));
  xor_4  g00031(.A(new_n2379), .B(new_n2349), .Y(new_n2380));
  not_8  g00032(.A(n5704), .Y(new_n2381));
  xnor_4 g00033(.A(n13781), .B(new_n2381), .Y(new_n2382));
  not_8  g00034(.A(n13781), .Y(new_n2383));
  nor_5  g00035(.A(new_n2383), .B(new_n2381), .Y(new_n2384));
  xnor_4 g00036(.A(n18409), .B(n11486), .Y(new_n2385));
  xnor_4 g00037(.A(new_n2385), .B(new_n2384), .Y(new_n2386));
  nor_5  g00038(.A(new_n2386), .B(new_n2382), .Y(new_n2387_1));
  not_8  g00039(.A(new_n2387_1), .Y(new_n2388_1));
  not_8  g00040(.A(n13708), .Y(new_n2389));
  xnor_4 g00041(.A(n16722), .B(new_n2389), .Y(new_n2390));
  nor_5  g00042(.A(n18409), .B(n11486), .Y(new_n2391));
  nor_5  g00043(.A(new_n2385), .B(new_n2384), .Y(new_n2392));
  nor_5  g00044(.A(new_n2392), .B(new_n2391), .Y(new_n2393));
  xnor_4 g00045(.A(new_n2393), .B(new_n2390), .Y(new_n2394));
  not_8  g00046(.A(new_n2394), .Y(new_n2395));
  nor_5  g00047(.A(new_n2395), .B(new_n2388_1), .Y(new_n2396));
  not_8  g00048(.A(new_n2396), .Y(new_n2397));
  not_8  g00049(.A(n3480), .Y(new_n2398));
  xnor_4 g00050(.A(n19911), .B(new_n2398), .Y(new_n2399));
  nor_5  g00051(.A(n16722), .B(n13708), .Y(new_n2400));
  or_5   g00052(.A(new_n2392), .B(new_n2391), .Y(new_n2401));
  and_5  g00053(.A(new_n2401), .B(new_n2390), .Y(new_n2402));
  nor_5  g00054(.A(new_n2402), .B(new_n2400), .Y(new_n2403));
  xnor_4 g00055(.A(new_n2403), .B(new_n2399), .Y(new_n2404));
  not_8  g00056(.A(new_n2404), .Y(new_n2405));
  nor_5  g00057(.A(new_n2405), .B(new_n2397), .Y(new_n2406));
  not_8  g00058(.A(new_n2406), .Y(new_n2407));
  not_8  g00059(.A(n2731), .Y(new_n2408));
  xnor_4 g00060(.A(n3018), .B(new_n2408), .Y(new_n2409_1));
  nor_5  g00061(.A(n19911), .B(n3480), .Y(new_n2410));
  or_5   g00062(.A(new_n2402), .B(new_n2400), .Y(new_n2411));
  and_5  g00063(.A(new_n2411), .B(new_n2399), .Y(new_n2412));
  nor_5  g00064(.A(new_n2412), .B(new_n2410), .Y(new_n2413));
  xnor_4 g00065(.A(new_n2413), .B(new_n2409_1), .Y(new_n2414));
  not_8  g00066(.A(new_n2414), .Y(new_n2415));
  nor_5  g00067(.A(new_n2415), .B(new_n2407), .Y(new_n2416_1));
  not_8  g00068(.A(new_n2416_1), .Y(new_n2417));
  xnor_4 g00069(.A(n26660), .B(n18907), .Y(new_n2418));
  nor_5  g00070(.A(n3018), .B(n2731), .Y(new_n2419));
  or_5   g00071(.A(new_n2412), .B(new_n2410), .Y(new_n2420_1));
  and_5  g00072(.A(new_n2420_1), .B(new_n2409_1), .Y(new_n2421_1));
  nor_5  g00073(.A(new_n2421_1), .B(new_n2419), .Y(new_n2422));
  xnor_4 g00074(.A(new_n2422), .B(new_n2418), .Y(new_n2423));
  nor_5  g00075(.A(new_n2423), .B(new_n2417), .Y(new_n2424));
  not_8  g00076(.A(n13783), .Y(new_n2425));
  xnor_4 g00077(.A(n22332), .B(new_n2425), .Y(new_n2426));
  nor_5  g00078(.A(n26660), .B(n18907), .Y(new_n2427));
  nor_5  g00079(.A(new_n2422), .B(new_n2418), .Y(new_n2428));
  nor_5  g00080(.A(new_n2428), .B(new_n2427), .Y(new_n2429));
  xnor_4 g00081(.A(new_n2429), .B(new_n2426), .Y(new_n2430));
  not_8  g00082(.A(new_n2430), .Y(new_n2431));
  xnor_4 g00083(.A(new_n2431), .B(new_n2424), .Y(new_n2432));
  xnor_4 g00084(.A(n13490), .B(n7751), .Y(new_n2433));
  nor_5  g00085(.A(n26823), .B(n22660), .Y(new_n2434));
  xnor_4 g00086(.A(n26823), .B(n22660), .Y(new_n2435));
  nor_5  g00087(.A(n4812), .B(n1777), .Y(new_n2436));
  xnor_4 g00088(.A(n4812), .B(n1777), .Y(new_n2437));
  nor_5  g00089(.A(n24278), .B(n8745), .Y(new_n2438));
  xnor_4 g00090(.A(n24278), .B(n8745), .Y(new_n2439));
  nor_5  g00091(.A(n24618), .B(n15636), .Y(new_n2440_1));
  not_8  g00092(.A(n15636), .Y(new_n2441));
  xnor_4 g00093(.A(n24618), .B(new_n2441), .Y(new_n2442));
  not_8  g00094(.A(n3952), .Y(new_n2443));
  not_8  g00095(.A(n20077), .Y(new_n2444_1));
  nor_5  g00096(.A(new_n2444_1), .B(new_n2443), .Y(new_n2445));
  or_5   g00097(.A(n20077), .B(n3952), .Y(new_n2446));
  not_8  g00098(.A(n6794), .Y(new_n2447));
  not_8  g00099(.A(n12315), .Y(new_n2448));
  nor_5  g00100(.A(new_n2448), .B(new_n2447), .Y(new_n2449));
  and_5  g00101(.A(new_n2449), .B(new_n2446), .Y(new_n2450));
  nor_5  g00102(.A(new_n2450), .B(new_n2445), .Y(new_n2451));
  and_5  g00103(.A(new_n2451), .B(new_n2442), .Y(new_n2452));
  nor_5  g00104(.A(new_n2452), .B(new_n2440_1), .Y(new_n2453));
  nor_5  g00105(.A(new_n2453), .B(new_n2439), .Y(new_n2454));
  nor_5  g00106(.A(new_n2454), .B(new_n2438), .Y(new_n2455));
  nor_5  g00107(.A(new_n2455), .B(new_n2437), .Y(new_n2456));
  nor_5  g00108(.A(new_n2456), .B(new_n2436), .Y(new_n2457));
  nor_5  g00109(.A(new_n2457), .B(new_n2435), .Y(new_n2458));
  nor_5  g00110(.A(new_n2458), .B(new_n2434), .Y(new_n2459));
  xnor_4 g00111(.A(new_n2459), .B(new_n2433), .Y(new_n2460));
  xnor_4 g00112(.A(new_n2460), .B(new_n2432), .Y(new_n2461));
  xnor_4 g00113(.A(new_n2423), .B(new_n2416_1), .Y(new_n2462));
  xnor_4 g00114(.A(new_n2457), .B(new_n2435), .Y(new_n2463));
  nor_5  g00115(.A(new_n2463), .B(new_n2462), .Y(new_n2464));
  xnor_4 g00116(.A(new_n2415), .B(new_n2406), .Y(new_n2465));
  xnor_4 g00117(.A(new_n2455), .B(new_n2437), .Y(new_n2466));
  nor_5  g00118(.A(new_n2466), .B(new_n2465), .Y(new_n2467));
  xnor_4 g00119(.A(new_n2466), .B(new_n2465), .Y(new_n2468));
  xnor_4 g00120(.A(new_n2405), .B(new_n2396), .Y(new_n2469));
  xnor_4 g00121(.A(new_n2453), .B(new_n2439), .Y(new_n2470));
  nor_5  g00122(.A(new_n2470), .B(new_n2469), .Y(new_n2471));
  xnor_4 g00123(.A(new_n2395), .B(new_n2387_1), .Y(new_n2472));
  xnor_4 g00124(.A(new_n2451), .B(new_n2442), .Y(new_n2473));
  nor_5  g00125(.A(new_n2473), .B(new_n2472), .Y(new_n2474));
  not_8  g00126(.A(new_n2473), .Y(new_n2475));
  xnor_4 g00127(.A(new_n2475), .B(new_n2472), .Y(new_n2476));
  not_8  g00128(.A(new_n2382), .Y(new_n2477));
  xnor_4 g00129(.A(n12315), .B(n6794), .Y(new_n2478));
  nor_5  g00130(.A(new_n2478), .B(new_n2477), .Y(new_n2479_1));
  xnor_4 g00131(.A(n20077), .B(n3952), .Y(new_n2480));
  xnor_4 g00132(.A(new_n2480), .B(new_n2449), .Y(new_n2481));
  nor_5  g00133(.A(new_n2481), .B(new_n2479_1), .Y(new_n2482));
  or_5   g00134(.A(n13781), .B(n5704), .Y(new_n2483));
  and_5  g00135(.A(new_n2392), .B(new_n2483), .Y(new_n2484));
  or_5   g00136(.A(new_n2484), .B(new_n2387_1), .Y(new_n2485));
  not_8  g00137(.A(new_n2479_1), .Y(new_n2486));
  nor_5  g00138(.A(new_n2480), .B(new_n2486), .Y(new_n2487));
  nor_5  g00139(.A(new_n2487), .B(new_n2482), .Y(new_n2488));
  and_5  g00140(.A(new_n2488), .B(new_n2485), .Y(new_n2489));
  or_5   g00141(.A(new_n2489), .B(new_n2482), .Y(new_n2490));
  and_5  g00142(.A(new_n2490), .B(new_n2476), .Y(new_n2491));
  nor_5  g00143(.A(new_n2491), .B(new_n2474), .Y(new_n2492));
  xnor_4 g00144(.A(new_n2470), .B(new_n2469), .Y(new_n2493));
  nor_5  g00145(.A(new_n2493), .B(new_n2492), .Y(new_n2494));
  nor_5  g00146(.A(new_n2494), .B(new_n2471), .Y(new_n2495));
  nor_5  g00147(.A(new_n2495), .B(new_n2468), .Y(new_n2496));
  nor_5  g00148(.A(new_n2496), .B(new_n2467), .Y(new_n2497));
  xnor_4 g00149(.A(new_n2463), .B(new_n2462), .Y(new_n2498));
  nor_5  g00150(.A(new_n2498), .B(new_n2497), .Y(new_n2499));
  nor_5  g00151(.A(new_n2499), .B(new_n2464), .Y(new_n2500));
  xnor_4 g00152(.A(new_n2500), .B(new_n2461), .Y(new_n2501));
  xor_4  g00153(.A(new_n2501), .B(new_n2380), .Y(new_n2502));
  xor_4  g00154(.A(new_n2377), .B(new_n2352), .Y(new_n2503));
  xnor_4 g00155(.A(new_n2498), .B(new_n2497), .Y(new_n2504));
  nor_5  g00156(.A(new_n2504), .B(new_n2503), .Y(new_n2505));
  xnor_4 g00157(.A(new_n2504), .B(new_n2503), .Y(new_n2506));
  xor_4  g00158(.A(new_n2375), .B(new_n2355_1), .Y(new_n2507));
  xnor_4 g00159(.A(new_n2495), .B(new_n2468), .Y(new_n2508));
  nor_5  g00160(.A(new_n2508), .B(new_n2507), .Y(new_n2509));
  xnor_4 g00161(.A(new_n2508), .B(new_n2507), .Y(new_n2510));
  xnor_4 g00162(.A(new_n2373), .B(new_n2358), .Y(new_n2511));
  xnor_4 g00163(.A(new_n2493), .B(new_n2492), .Y(new_n2512));
  not_8  g00164(.A(new_n2512), .Y(new_n2513_1));
  and_5  g00165(.A(new_n2513_1), .B(new_n2511), .Y(new_n2514));
  xnor_4 g00166(.A(new_n2513_1), .B(new_n2511), .Y(new_n2515_1));
  xor_4  g00167(.A(new_n2490), .B(new_n2476), .Y(new_n2516));
  xnor_4 g00168(.A(n16223), .B(n6385), .Y(new_n2517));
  xnor_4 g00169(.A(new_n2517), .B(new_n2371), .Y(new_n2518));
  and_5  g00170(.A(new_n2518), .B(new_n2516), .Y(new_n2519));
  xnor_4 g00171(.A(new_n2518), .B(new_n2516), .Y(new_n2520));
  xnor_4 g00172(.A(n9251), .B(n2387), .Y(new_n2521));
  xnor_4 g00173(.A(new_n2478), .B(new_n2382), .Y(new_n2522));
  not_8  g00174(.A(new_n2522), .Y(new_n2523));
  or_5   g00175(.A(new_n2523), .B(new_n2521), .Y(new_n2524));
  xnor_4 g00176(.A(n20138), .B(n19494), .Y(new_n2525));
  xnor_4 g00177(.A(new_n2525), .B(new_n2369), .Y(new_n2526));
  and_5  g00178(.A(new_n2526), .B(new_n2524), .Y(new_n2527));
  xnor_4 g00179(.A(new_n2488), .B(new_n2485), .Y(new_n2528));
  not_8  g00180(.A(new_n2528), .Y(new_n2529));
  xor_4  g00181(.A(new_n2526), .B(new_n2524), .Y(new_n2530));
  and_5  g00182(.A(new_n2530), .B(new_n2529), .Y(new_n2531));
  nor_5  g00183(.A(new_n2531), .B(new_n2527), .Y(new_n2532));
  nor_5  g00184(.A(new_n2532), .B(new_n2520), .Y(new_n2533_1));
  nor_5  g00185(.A(new_n2533_1), .B(new_n2519), .Y(new_n2534));
  nor_5  g00186(.A(new_n2534), .B(new_n2515_1), .Y(new_n2535_1));
  nor_5  g00187(.A(new_n2535_1), .B(new_n2514), .Y(new_n2536));
  nor_5  g00188(.A(new_n2536), .B(new_n2510), .Y(new_n2537_1));
  nor_5  g00189(.A(new_n2537_1), .B(new_n2509), .Y(new_n2538));
  nor_5  g00190(.A(new_n2538), .B(new_n2506), .Y(new_n2539));
  nor_5  g00191(.A(new_n2539), .B(new_n2505), .Y(new_n2540));
  xor_4  g00192(.A(new_n2540), .B(new_n2502), .Y(n7));
  not_8  g00193(.A(n4588), .Y(new_n2542));
  xnor_4 g00194(.A(n3618), .B(n1681), .Y(new_n2543));
  xnor_4 g00195(.A(new_n2543), .B(new_n2542), .Y(new_n2544));
  xnor_4 g00196(.A(n22843), .B(n583), .Y(new_n2545));
  xnor_4 g00197(.A(new_n2545), .B(n22201), .Y(new_n2546));
  xnor_4 g00198(.A(new_n2546), .B(new_n2544), .Y(n50));
  not_8  g00199(.A(n21687), .Y(new_n2548));
  xnor_4 g00200(.A(n19922), .B(n6773), .Y(new_n2549));
  xnor_4 g00201(.A(new_n2549), .B(new_n2548), .Y(new_n2550));
  xnor_4 g00202(.A(n21398), .B(n14090), .Y(new_n2551));
  xnor_4 g00203(.A(new_n2551), .B(n25926), .Y(new_n2552));
  xnor_4 g00204(.A(new_n2552), .B(new_n2550), .Y(n55));
  not_8  g00205(.A(n9396), .Y(new_n2554));
  xnor_4 g00206(.A(n20040), .B(new_n2554), .Y(new_n2555_1));
  not_8  g00207(.A(new_n2555_1), .Y(new_n2556));
  nor_5  g00208(.A(n19531), .B(n1999), .Y(new_n2557));
  not_8  g00209(.A(n19531), .Y(new_n2558));
  xnor_4 g00210(.A(new_n2558), .B(n1999), .Y(new_n2559));
  not_8  g00211(.A(new_n2559), .Y(new_n2560_1));
  nor_5  g00212(.A(n25168), .B(n18345), .Y(new_n2561_1));
  not_8  g00213(.A(n18345), .Y(new_n2562));
  xnor_4 g00214(.A(n25168), .B(new_n2562), .Y(new_n2563));
  not_8  g00215(.A(new_n2563), .Y(new_n2564));
  nor_5  g00216(.A(n13190), .B(n9318), .Y(new_n2565));
  not_8  g00217(.A(n13190), .Y(new_n2566));
  xnor_4 g00218(.A(new_n2566), .B(n9318), .Y(new_n2567));
  not_8  g00219(.A(new_n2567), .Y(new_n2568));
  nor_5  g00220(.A(n19477), .B(n3460), .Y(new_n2569));
  xnor_4 g00221(.A(n19477), .B(n3460), .Y(new_n2570_1));
  nor_5  g00222(.A(n11223), .B(n5226), .Y(new_n2571));
  xnor_4 g00223(.A(n11223), .B(n5226), .Y(new_n2572));
  nor_5  g00224(.A(n17664), .B(n5115), .Y(new_n2573_1));
  not_8  g00225(.A(n17664), .Y(new_n2574));
  xnor_4 g00226(.A(new_n2574), .B(n5115), .Y(new_n2575));
  not_8  g00227(.A(new_n2575), .Y(new_n2576));
  nor_5  g00228(.A(n26572), .B(n23369), .Y(new_n2577));
  not_8  g00229(.A(n23369), .Y(new_n2578_1));
  xnor_4 g00230(.A(n26572), .B(new_n2578_1), .Y(new_n2579));
  not_8  g00231(.A(new_n2579), .Y(new_n2580));
  nor_5  g00232(.A(n11667), .B(n1136), .Y(new_n2581));
  not_8  g00233(.A(n19234), .Y(new_n2582_1));
  not_8  g00234(.A(n21398), .Y(new_n2583));
  nor_5  g00235(.A(new_n2583), .B(new_n2582_1), .Y(new_n2584));
  xnor_4 g00236(.A(n11667), .B(n1136), .Y(new_n2585));
  nor_5  g00237(.A(new_n2585), .B(new_n2584), .Y(new_n2586));
  nor_5  g00238(.A(new_n2586), .B(new_n2581), .Y(new_n2587));
  nor_5  g00239(.A(new_n2587), .B(new_n2580), .Y(new_n2588));
  nor_5  g00240(.A(new_n2588), .B(new_n2577), .Y(new_n2589));
  nor_5  g00241(.A(new_n2589), .B(new_n2576), .Y(new_n2590));
  nor_5  g00242(.A(new_n2590), .B(new_n2573_1), .Y(new_n2591));
  nor_5  g00243(.A(new_n2591), .B(new_n2572), .Y(new_n2592));
  nor_5  g00244(.A(new_n2592), .B(new_n2571), .Y(new_n2593));
  nor_5  g00245(.A(new_n2593), .B(new_n2570_1), .Y(new_n2594));
  nor_5  g00246(.A(new_n2594), .B(new_n2569), .Y(new_n2595));
  nor_5  g00247(.A(new_n2595), .B(new_n2568), .Y(new_n2596));
  nor_5  g00248(.A(new_n2596), .B(new_n2565), .Y(new_n2597));
  nor_5  g00249(.A(new_n2597), .B(new_n2564), .Y(new_n2598));
  nor_5  g00250(.A(new_n2598), .B(new_n2561_1), .Y(new_n2599));
  nor_5  g00251(.A(new_n2599), .B(new_n2560_1), .Y(new_n2600));
  nor_5  g00252(.A(new_n2600), .B(new_n2557), .Y(new_n2601));
  xnor_4 g00253(.A(new_n2601), .B(new_n2556), .Y(new_n2602_1));
  not_8  g00254(.A(new_n2602_1), .Y(new_n2603));
  xnor_4 g00255(.A(new_n2603), .B(n25365), .Y(new_n2604));
  xnor_4 g00256(.A(new_n2599), .B(new_n2560_1), .Y(new_n2605));
  and_5  g00257(.A(new_n2605), .B(n14704), .Y(new_n2606));
  not_8  g00258(.A(new_n2605), .Y(new_n2607));
  xnor_4 g00259(.A(new_n2607), .B(n14704), .Y(new_n2608));
  xnor_4 g00260(.A(new_n2597), .B(new_n2564), .Y(new_n2609));
  and_5  g00261(.A(new_n2609), .B(n19270), .Y(new_n2610));
  not_8  g00262(.A(new_n2609), .Y(new_n2611));
  xnor_4 g00263(.A(new_n2611), .B(n19270), .Y(new_n2612));
  xnor_4 g00264(.A(new_n2595), .B(new_n2568), .Y(new_n2613));
  and_5  g00265(.A(new_n2613), .B(n8687), .Y(new_n2614));
  xnor_4 g00266(.A(new_n2593), .B(new_n2570_1), .Y(new_n2615));
  nor_5  g00267(.A(new_n2615), .B(n24768), .Y(new_n2616));
  xnor_4 g00268(.A(new_n2615), .B(n24768), .Y(new_n2617));
  xnor_4 g00269(.A(new_n2591), .B(new_n2572), .Y(new_n2618));
  nor_5  g00270(.A(new_n2618), .B(n26483), .Y(new_n2619_1));
  xnor_4 g00271(.A(new_n2618), .B(n26483), .Y(new_n2620));
  xnor_4 g00272(.A(new_n2589), .B(new_n2576), .Y(new_n2621));
  and_5  g00273(.A(new_n2621), .B(n15979), .Y(new_n2622));
  not_8  g00274(.A(new_n2621), .Y(new_n2623));
  xnor_4 g00275(.A(new_n2623), .B(n15979), .Y(new_n2624));
  xnor_4 g00276(.A(new_n2587), .B(new_n2580), .Y(new_n2625));
  and_5  g00277(.A(new_n2625), .B(n8638), .Y(new_n2626));
  xnor_4 g00278(.A(new_n2585), .B(new_n2584), .Y(new_n2627));
  nor_5  g00279(.A(new_n2627), .B(n16247), .Y(new_n2628));
  not_8  g00280(.A(n23541), .Y(new_n2629));
  xnor_4 g00281(.A(n21398), .B(n19234), .Y(new_n2630));
  or_5   g00282(.A(new_n2630), .B(new_n2629), .Y(new_n2631));
  not_8  g00283(.A(n16247), .Y(new_n2632));
  xnor_4 g00284(.A(new_n2627), .B(new_n2632), .Y(new_n2633));
  and_5  g00285(.A(new_n2633), .B(new_n2631), .Y(new_n2634));
  nor_5  g00286(.A(new_n2634), .B(new_n2628), .Y(new_n2635));
  not_8  g00287(.A(new_n2625), .Y(new_n2636));
  xnor_4 g00288(.A(new_n2636), .B(n8638), .Y(new_n2637));
  and_5  g00289(.A(new_n2637), .B(new_n2635), .Y(new_n2638));
  or_5   g00290(.A(new_n2638), .B(new_n2626), .Y(new_n2639));
  and_5  g00291(.A(new_n2639), .B(new_n2624), .Y(new_n2640));
  nor_5  g00292(.A(new_n2640), .B(new_n2622), .Y(new_n2641));
  not_8  g00293(.A(new_n2641), .Y(new_n2642));
  nor_5  g00294(.A(new_n2642), .B(new_n2620), .Y(new_n2643));
  nor_5  g00295(.A(new_n2643), .B(new_n2619_1), .Y(new_n2644));
  nor_5  g00296(.A(new_n2644), .B(new_n2617), .Y(new_n2645));
  nor_5  g00297(.A(new_n2645), .B(new_n2616), .Y(new_n2646_1));
  not_8  g00298(.A(new_n2613), .Y(new_n2647));
  xnor_4 g00299(.A(new_n2647), .B(n8687), .Y(new_n2648));
  and_5  g00300(.A(new_n2648), .B(new_n2646_1), .Y(new_n2649));
  or_5   g00301(.A(new_n2649), .B(new_n2614), .Y(new_n2650));
  and_5  g00302(.A(new_n2650), .B(new_n2612), .Y(new_n2651));
  or_5   g00303(.A(new_n2651), .B(new_n2610), .Y(new_n2652));
  and_5  g00304(.A(new_n2652), .B(new_n2608), .Y(new_n2653));
  nor_5  g00305(.A(new_n2653), .B(new_n2606), .Y(new_n2654));
  xnor_4 g00306(.A(new_n2654), .B(new_n2604), .Y(new_n2655));
  not_8  g00307(.A(new_n2655), .Y(new_n2656));
  nor_5  g00308(.A(n18151), .B(n11503), .Y(new_n2657));
  not_8  g00309(.A(new_n2657), .Y(new_n2658));
  nor_5  g00310(.A(new_n2658), .B(n16971), .Y(new_n2659_1));
  not_8  g00311(.A(new_n2659_1), .Y(new_n2660));
  nor_5  g00312(.A(new_n2660), .B(n10411), .Y(new_n2661_1));
  not_8  g00313(.A(new_n2661_1), .Y(new_n2662));
  nor_5  g00314(.A(new_n2662), .B(n23430), .Y(new_n2663));
  not_8  g00315(.A(new_n2663), .Y(new_n2664));
  nor_5  g00316(.A(new_n2664), .B(n5579), .Y(new_n2665));
  not_8  g00317(.A(new_n2665), .Y(new_n2666));
  nor_5  g00318(.A(new_n2666), .B(n25523), .Y(new_n2667));
  not_8  g00319(.A(new_n2667), .Y(new_n2668));
  nor_5  g00320(.A(new_n2668), .B(n8439), .Y(new_n2669));
  not_8  g00321(.A(new_n2669), .Y(new_n2670));
  nor_5  g00322(.A(new_n2670), .B(n22793), .Y(new_n2671));
  not_8  g00323(.A(new_n2671), .Y(new_n2672));
  xnor_4 g00324(.A(new_n2672), .B(n13951), .Y(new_n2673));
  not_8  g00325(.A(n2944), .Y(new_n2674));
  xnor_4 g00326(.A(n22270), .B(new_n2674), .Y(new_n2675));
  nor_5  g00327(.A(n8806), .B(n767), .Y(new_n2676));
  not_8  g00328(.A(n767), .Y(new_n2677));
  xnor_4 g00329(.A(n8806), .B(new_n2677), .Y(new_n2678));
  nor_5  g00330(.A(n7330), .B(n2479), .Y(new_n2679));
  not_8  g00331(.A(n2479), .Y(new_n2680_1));
  xnor_4 g00332(.A(n7330), .B(new_n2680_1), .Y(new_n2681));
  nor_5  g00333(.A(n22492), .B(n9372), .Y(new_n2682));
  not_8  g00334(.A(n22492), .Y(new_n2683));
  xnor_4 g00335(.A(new_n2683), .B(n9372), .Y(new_n2684));
  nor_5  g00336(.A(n12821), .B(n6596), .Y(new_n2685));
  not_8  g00337(.A(n6596), .Y(new_n2686));
  xnor_4 g00338(.A(n12821), .B(new_n2686), .Y(new_n2687));
  nor_5  g00339(.A(n15289), .B(n3468), .Y(new_n2688));
  not_8  g00340(.A(n3468), .Y(new_n2689));
  xnor_4 g00341(.A(n15289), .B(new_n2689), .Y(new_n2690));
  nor_5  g00342(.A(n18558), .B(n6556), .Y(new_n2691));
  not_8  g00343(.A(n6556), .Y(new_n2692));
  xnor_4 g00344(.A(n18558), .B(new_n2692), .Y(new_n2693_1));
  nor_5  g00345(.A(n22871), .B(n7149), .Y(new_n2694));
  not_8  g00346(.A(n7149), .Y(new_n2695));
  xnor_4 g00347(.A(n22871), .B(new_n2695), .Y(new_n2696));
  nor_5  g00348(.A(n14275), .B(n14148), .Y(new_n2697));
  not_8  g00349(.A(n1152), .Y(new_n2698));
  not_8  g00350(.A(n25023), .Y(new_n2699));
  or_5   g00351(.A(new_n2699), .B(new_n2698), .Y(new_n2700));
  not_8  g00352(.A(n14148), .Y(new_n2701));
  xnor_4 g00353(.A(n14275), .B(new_n2701), .Y(new_n2702));
  and_5  g00354(.A(new_n2702), .B(new_n2700), .Y(new_n2703_1));
  or_5   g00355(.A(new_n2703_1), .B(new_n2697), .Y(new_n2704));
  and_5  g00356(.A(new_n2704), .B(new_n2696), .Y(new_n2705));
  or_5   g00357(.A(new_n2705), .B(new_n2694), .Y(new_n2706_1));
  and_5  g00358(.A(new_n2706_1), .B(new_n2693_1), .Y(new_n2707));
  or_5   g00359(.A(new_n2707), .B(new_n2691), .Y(new_n2708));
  and_5  g00360(.A(new_n2708), .B(new_n2690), .Y(new_n2709));
  or_5   g00361(.A(new_n2709), .B(new_n2688), .Y(new_n2710));
  and_5  g00362(.A(new_n2710), .B(new_n2687), .Y(new_n2711_1));
  or_5   g00363(.A(new_n2711_1), .B(new_n2685), .Y(new_n2712));
  and_5  g00364(.A(new_n2712), .B(new_n2684), .Y(new_n2713));
  or_5   g00365(.A(new_n2713), .B(new_n2682), .Y(new_n2714));
  and_5  g00366(.A(new_n2714), .B(new_n2681), .Y(new_n2715));
  or_5   g00367(.A(new_n2715), .B(new_n2679), .Y(new_n2716));
  and_5  g00368(.A(new_n2716), .B(new_n2678), .Y(new_n2717));
  nor_5  g00369(.A(new_n2717), .B(new_n2676), .Y(new_n2718));
  xnor_4 g00370(.A(new_n2718), .B(new_n2675), .Y(new_n2719));
  xnor_4 g00371(.A(new_n2719), .B(new_n2673), .Y(new_n2720));
  xnor_4 g00372(.A(new_n2669), .B(n22793), .Y(new_n2721));
  nor_5  g00373(.A(new_n2715), .B(new_n2679), .Y(new_n2722));
  xnor_4 g00374(.A(new_n2722), .B(new_n2678), .Y(new_n2723));
  and_5  g00375(.A(new_n2723), .B(new_n2721), .Y(new_n2724));
  not_8  g00376(.A(new_n2723), .Y(new_n2725));
  xnor_4 g00377(.A(new_n2725), .B(new_n2721), .Y(new_n2726));
  xnor_4 g00378(.A(new_n2667), .B(n8439), .Y(new_n2727));
  nor_5  g00379(.A(new_n2713), .B(new_n2682), .Y(new_n2728));
  xnor_4 g00380(.A(new_n2728), .B(new_n2681), .Y(new_n2729));
  nor_5  g00381(.A(new_n2729), .B(new_n2727), .Y(new_n2730));
  xnor_4 g00382(.A(new_n2729), .B(new_n2727), .Y(new_n2731_1));
  xnor_4 g00383(.A(new_n2665), .B(n25523), .Y(new_n2732));
  xor_4  g00384(.A(new_n2712), .B(new_n2684), .Y(new_n2733));
  nor_5  g00385(.A(new_n2733), .B(new_n2732), .Y(new_n2734));
  xnor_4 g00386(.A(new_n2733), .B(new_n2732), .Y(new_n2735));
  xnor_4 g00387(.A(new_n2663), .B(n5579), .Y(new_n2736));
  nor_5  g00388(.A(new_n2709), .B(new_n2688), .Y(new_n2737));
  xnor_4 g00389(.A(new_n2737), .B(new_n2687), .Y(new_n2738));
  nor_5  g00390(.A(new_n2738), .B(new_n2736), .Y(new_n2739));
  not_8  g00391(.A(new_n2738), .Y(new_n2740));
  xnor_4 g00392(.A(new_n2740), .B(new_n2736), .Y(new_n2741));
  xnor_4 g00393(.A(new_n2661_1), .B(n23430), .Y(new_n2742));
  nor_5  g00394(.A(new_n2707), .B(new_n2691), .Y(new_n2743_1));
  xnor_4 g00395(.A(new_n2743_1), .B(new_n2690), .Y(new_n2744));
  nor_5  g00396(.A(new_n2744), .B(new_n2742), .Y(new_n2745));
  xnor_4 g00397(.A(new_n2659_1), .B(n10411), .Y(new_n2746));
  nor_5  g00398(.A(new_n2705), .B(new_n2694), .Y(new_n2747));
  xnor_4 g00399(.A(new_n2747), .B(new_n2693_1), .Y(new_n2748));
  nor_5  g00400(.A(new_n2748), .B(new_n2746), .Y(new_n2749));
  xnor_4 g00401(.A(new_n2748), .B(new_n2746), .Y(new_n2750));
  xnor_4 g00402(.A(new_n2657), .B(n16971), .Y(new_n2751));
  nor_5  g00403(.A(new_n2703_1), .B(new_n2697), .Y(new_n2752));
  xnor_4 g00404(.A(new_n2752), .B(new_n2696), .Y(new_n2753));
  nor_5  g00405(.A(new_n2753), .B(new_n2751), .Y(new_n2754));
  xnor_4 g00406(.A(new_n2753), .B(new_n2751), .Y(new_n2755));
  not_8  g00407(.A(n11503), .Y(new_n2756));
  xnor_4 g00408(.A(n18151), .B(new_n2756), .Y(new_n2757));
  nor_5  g00409(.A(new_n2699), .B(new_n2698), .Y(new_n2758));
  xnor_4 g00410(.A(new_n2702), .B(new_n2758), .Y(new_n2759));
  nor_5  g00411(.A(new_n2759), .B(new_n2757), .Y(new_n2760));
  xnor_4 g00412(.A(n25023), .B(n1152), .Y(new_n2761_1));
  nor_5  g00413(.A(new_n2761_1), .B(n18151), .Y(new_n2762));
  not_8  g00414(.A(new_n2759), .Y(new_n2763));
  xnor_4 g00415(.A(new_n2763), .B(new_n2757), .Y(new_n2764));
  and_5  g00416(.A(new_n2764), .B(new_n2762), .Y(new_n2765));
  nor_5  g00417(.A(new_n2765), .B(new_n2760), .Y(new_n2766));
  nor_5  g00418(.A(new_n2766), .B(new_n2755), .Y(new_n2767));
  nor_5  g00419(.A(new_n2767), .B(new_n2754), .Y(new_n2768));
  nor_5  g00420(.A(new_n2768), .B(new_n2750), .Y(new_n2769));
  or_5   g00421(.A(new_n2769), .B(new_n2749), .Y(new_n2770));
  not_8  g00422(.A(new_n2744), .Y(new_n2771));
  xnor_4 g00423(.A(new_n2771), .B(new_n2742), .Y(new_n2772));
  and_5  g00424(.A(new_n2772), .B(new_n2770), .Y(new_n2773));
  or_5   g00425(.A(new_n2773), .B(new_n2745), .Y(new_n2774_1));
  and_5  g00426(.A(new_n2774_1), .B(new_n2741), .Y(new_n2775));
  nor_5  g00427(.A(new_n2775), .B(new_n2739), .Y(new_n2776));
  nor_5  g00428(.A(new_n2776), .B(new_n2735), .Y(new_n2777));
  nor_5  g00429(.A(new_n2777), .B(new_n2734), .Y(new_n2778));
  nor_5  g00430(.A(new_n2778), .B(new_n2731_1), .Y(new_n2779_1));
  nor_5  g00431(.A(new_n2779_1), .B(new_n2730), .Y(new_n2780));
  and_5  g00432(.A(new_n2780), .B(new_n2726), .Y(new_n2781));
  or_5   g00433(.A(new_n2781), .B(new_n2724), .Y(new_n2782));
  xor_4  g00434(.A(new_n2782), .B(new_n2720), .Y(new_n2783_1));
  xnor_4 g00435(.A(new_n2783_1), .B(new_n2656), .Y(new_n2784));
  nor_5  g00436(.A(new_n2651), .B(new_n2610), .Y(new_n2785));
  xnor_4 g00437(.A(new_n2785), .B(new_n2608), .Y(new_n2786));
  not_8  g00438(.A(new_n2786), .Y(new_n2787));
  xnor_4 g00439(.A(new_n2780), .B(new_n2726), .Y(new_n2788));
  nor_5  g00440(.A(new_n2788), .B(new_n2787), .Y(new_n2789));
  xnor_4 g00441(.A(new_n2788), .B(new_n2786), .Y(new_n2790));
  nor_5  g00442(.A(new_n2649), .B(new_n2614), .Y(new_n2791));
  xnor_4 g00443(.A(new_n2791), .B(new_n2612), .Y(new_n2792));
  xnor_4 g00444(.A(new_n2778), .B(new_n2731_1), .Y(new_n2793));
  nor_5  g00445(.A(new_n2793), .B(new_n2792), .Y(new_n2794));
  xnor_4 g00446(.A(new_n2793), .B(new_n2792), .Y(new_n2795));
  xnor_4 g00447(.A(new_n2648), .B(new_n2646_1), .Y(new_n2796));
  not_8  g00448(.A(new_n2796), .Y(new_n2797));
  xnor_4 g00449(.A(new_n2776), .B(new_n2735), .Y(new_n2798));
  nor_5  g00450(.A(new_n2798), .B(new_n2797), .Y(new_n2799));
  xnor_4 g00451(.A(new_n2798), .B(new_n2796), .Y(new_n2800));
  xnor_4 g00452(.A(new_n2644), .B(new_n2617), .Y(new_n2801));
  not_8  g00453(.A(new_n2801), .Y(new_n2802));
  xor_4  g00454(.A(new_n2774_1), .B(new_n2741), .Y(new_n2803));
  nor_5  g00455(.A(new_n2803), .B(new_n2802), .Y(new_n2804));
  xnor_4 g00456(.A(new_n2803), .B(new_n2801), .Y(new_n2805));
  xnor_4 g00457(.A(new_n2641), .B(new_n2620), .Y(new_n2806));
  xor_4  g00458(.A(new_n2772), .B(new_n2770), .Y(new_n2807));
  and_5  g00459(.A(new_n2807), .B(new_n2806), .Y(new_n2808));
  xnor_4 g00460(.A(new_n2807), .B(new_n2806), .Y(new_n2809_1));
  xnor_4 g00461(.A(new_n2768), .B(new_n2750), .Y(new_n2810));
  nor_5  g00462(.A(new_n2638), .B(new_n2626), .Y(new_n2811));
  xnor_4 g00463(.A(new_n2811), .B(new_n2624), .Y(new_n2812));
  nor_5  g00464(.A(new_n2812), .B(new_n2810), .Y(new_n2813));
  not_8  g00465(.A(new_n2812), .Y(new_n2814));
  xnor_4 g00466(.A(new_n2814), .B(new_n2810), .Y(new_n2815));
  xnor_4 g00467(.A(new_n2766), .B(new_n2755), .Y(new_n2816_1));
  xnor_4 g00468(.A(new_n2637), .B(new_n2635), .Y(new_n2817));
  not_8  g00469(.A(new_n2817), .Y(new_n2818));
  and_5  g00470(.A(new_n2818), .B(new_n2816_1), .Y(new_n2819));
  xnor_4 g00471(.A(new_n2817), .B(new_n2816_1), .Y(new_n2820));
  xnor_4 g00472(.A(new_n2764), .B(new_n2762), .Y(new_n2821));
  nor_5  g00473(.A(new_n2630), .B(new_n2629), .Y(new_n2822));
  xnor_4 g00474(.A(new_n2633), .B(new_n2822), .Y(new_n2823));
  not_8  g00475(.A(new_n2823), .Y(new_n2824));
  nor_5  g00476(.A(new_n2824), .B(new_n2821), .Y(new_n2825));
  xnor_4 g00477(.A(new_n2630), .B(n23541), .Y(new_n2826_1));
  not_8  g00478(.A(new_n2826_1), .Y(new_n2827));
  not_8  g00479(.A(n18151), .Y(new_n2828));
  xnor_4 g00480(.A(new_n2761_1), .B(new_n2828), .Y(new_n2829));
  nor_5  g00481(.A(new_n2829), .B(new_n2827), .Y(new_n2830));
  xnor_4 g00482(.A(new_n2824), .B(new_n2821), .Y(new_n2831));
  nor_5  g00483(.A(new_n2831), .B(new_n2830), .Y(new_n2832));
  nor_5  g00484(.A(new_n2832), .B(new_n2825), .Y(new_n2833));
  and_5  g00485(.A(new_n2833), .B(new_n2820), .Y(new_n2834));
  nor_5  g00486(.A(new_n2834), .B(new_n2819), .Y(new_n2835));
  and_5  g00487(.A(new_n2835), .B(new_n2815), .Y(new_n2836));
  nor_5  g00488(.A(new_n2836), .B(new_n2813), .Y(new_n2837));
  nor_5  g00489(.A(new_n2837), .B(new_n2809_1), .Y(new_n2838));
  nor_5  g00490(.A(new_n2838), .B(new_n2808), .Y(new_n2839));
  and_5  g00491(.A(new_n2839), .B(new_n2805), .Y(new_n2840));
  nor_5  g00492(.A(new_n2840), .B(new_n2804), .Y(new_n2841));
  and_5  g00493(.A(new_n2841), .B(new_n2800), .Y(new_n2842));
  nor_5  g00494(.A(new_n2842), .B(new_n2799), .Y(new_n2843));
  nor_5  g00495(.A(new_n2843), .B(new_n2795), .Y(new_n2844));
  nor_5  g00496(.A(new_n2844), .B(new_n2794), .Y(new_n2845));
  and_5  g00497(.A(new_n2845), .B(new_n2790), .Y(new_n2846));
  nor_5  g00498(.A(new_n2846), .B(new_n2789), .Y(new_n2847));
  xnor_4 g00499(.A(new_n2847), .B(new_n2784), .Y(n108));
  xnor_4 g00500(.A(n22379), .B(n767), .Y(new_n2849));
  not_8  g00501(.A(n1662), .Y(new_n2850));
  nor_5  g00502(.A(n7330), .B(new_n2850), .Y(new_n2851));
  xnor_4 g00503(.A(n7330), .B(n1662), .Y(new_n2852));
  not_8  g00504(.A(n12875), .Y(new_n2853_1));
  nor_5  g00505(.A(n22492), .B(new_n2853_1), .Y(new_n2854));
  xnor_4 g00506(.A(n22492), .B(n12875), .Y(new_n2855));
  not_8  g00507(.A(n2035), .Y(new_n2856));
  nor_5  g00508(.A(n12821), .B(new_n2856), .Y(new_n2857));
  xnor_4 g00509(.A(n12821), .B(n2035), .Y(new_n2858_1));
  not_8  g00510(.A(n5213), .Y(new_n2859));
  nor_5  g00511(.A(new_n2859), .B(n3468), .Y(new_n2860_1));
  xnor_4 g00512(.A(n5213), .B(n3468), .Y(new_n2861));
  not_8  g00513(.A(n4665), .Y(new_n2862));
  nor_5  g00514(.A(n18558), .B(new_n2862), .Y(new_n2863));
  xnor_4 g00515(.A(n18558), .B(n4665), .Y(new_n2864));
  nor_5  g00516(.A(n19005), .B(new_n2695), .Y(new_n2865));
  not_8  g00517(.A(n19005), .Y(new_n2866));
  nor_5  g00518(.A(new_n2866), .B(n7149), .Y(new_n2867));
  nor_5  g00519(.A(new_n2701), .B(n4326), .Y(new_n2868));
  not_8  g00520(.A(n4326), .Y(new_n2869));
  or_5   g00521(.A(n14148), .B(new_n2869), .Y(new_n2870));
  nor_5  g00522(.A(n5438), .B(new_n2698), .Y(new_n2871));
  and_5  g00523(.A(new_n2871), .B(new_n2870), .Y(new_n2872));
  nor_5  g00524(.A(new_n2872), .B(new_n2868), .Y(new_n2873));
  nor_5  g00525(.A(new_n2873), .B(new_n2867), .Y(new_n2874));
  nor_5  g00526(.A(new_n2874), .B(new_n2865), .Y(new_n2875));
  and_5  g00527(.A(new_n2875), .B(new_n2864), .Y(new_n2876));
  or_5   g00528(.A(new_n2876), .B(new_n2863), .Y(new_n2877));
  and_5  g00529(.A(new_n2877), .B(new_n2861), .Y(new_n2878));
  or_5   g00530(.A(new_n2878), .B(new_n2860_1), .Y(new_n2879));
  and_5  g00531(.A(new_n2879), .B(new_n2858_1), .Y(new_n2880));
  or_5   g00532(.A(new_n2880), .B(new_n2857), .Y(new_n2881));
  and_5  g00533(.A(new_n2881), .B(new_n2855), .Y(new_n2882));
  or_5   g00534(.A(new_n2882), .B(new_n2854), .Y(new_n2883));
  and_5  g00535(.A(new_n2883), .B(new_n2852), .Y(new_n2884));
  or_5   g00536(.A(new_n2884), .B(new_n2851), .Y(new_n2885));
  xor_4  g00537(.A(new_n2885), .B(new_n2849), .Y(new_n2886_1));
  not_8  g00538(.A(n6814), .Y(new_n2887_1));
  xnor_4 g00539(.A(n10763), .B(new_n2887_1), .Y(new_n2888));
  nor_5  g00540(.A(n19701), .B(n7437), .Y(new_n2889));
  not_8  g00541(.A(n7437), .Y(new_n2890));
  xnor_4 g00542(.A(n19701), .B(new_n2890), .Y(new_n2891));
  nor_5  g00543(.A(n23529), .B(n20700), .Y(new_n2892));
  not_8  g00544(.A(n20700), .Y(new_n2893));
  xnor_4 g00545(.A(n23529), .B(new_n2893), .Y(new_n2894));
  nor_5  g00546(.A(n24620), .B(n7099), .Y(new_n2895));
  not_8  g00547(.A(n7099), .Y(new_n2896));
  xnor_4 g00548(.A(n24620), .B(new_n2896), .Y(new_n2897));
  nor_5  g00549(.A(n12811), .B(n5211), .Y(new_n2898));
  xnor_4 g00550(.A(n12811), .B(n5211), .Y(new_n2899));
  nor_5  g00551(.A(n12956), .B(n1118), .Y(new_n2900));
  xnor_4 g00552(.A(n12956), .B(n1118), .Y(new_n2901));
  nor_5  g00553(.A(n25974), .B(n18295), .Y(new_n2902));
  not_8  g00554(.A(n18295), .Y(new_n2903));
  xnor_4 g00555(.A(n25974), .B(new_n2903), .Y(new_n2904));
  nor_5  g00556(.A(n6502), .B(n1630), .Y(new_n2905));
  not_8  g00557(.A(n1451), .Y(new_n2906));
  not_8  g00558(.A(n15780), .Y(new_n2907));
  or_5   g00559(.A(new_n2907), .B(new_n2906), .Y(new_n2908));
  not_8  g00560(.A(n1630), .Y(new_n2909));
  xnor_4 g00561(.A(n6502), .B(new_n2909), .Y(new_n2910));
  and_5  g00562(.A(new_n2910), .B(new_n2908), .Y(new_n2911));
  or_5   g00563(.A(new_n2911), .B(new_n2905), .Y(new_n2912));
  and_5  g00564(.A(new_n2912), .B(new_n2904), .Y(new_n2913));
  nor_5  g00565(.A(new_n2913), .B(new_n2902), .Y(new_n2914));
  nor_5  g00566(.A(new_n2914), .B(new_n2901), .Y(new_n2915));
  nor_5  g00567(.A(new_n2915), .B(new_n2900), .Y(new_n2916));
  nor_5  g00568(.A(new_n2916), .B(new_n2899), .Y(new_n2917));
  or_5   g00569(.A(new_n2917), .B(new_n2898), .Y(new_n2918));
  and_5  g00570(.A(new_n2918), .B(new_n2897), .Y(new_n2919));
  or_5   g00571(.A(new_n2919), .B(new_n2895), .Y(new_n2920));
  and_5  g00572(.A(new_n2920), .B(new_n2894), .Y(new_n2921));
  or_5   g00573(.A(new_n2921), .B(new_n2892), .Y(new_n2922));
  and_5  g00574(.A(new_n2922), .B(new_n2891), .Y(new_n2923));
  or_5   g00575(.A(new_n2923), .B(new_n2889), .Y(new_n2924));
  xor_4  g00576(.A(new_n2924), .B(new_n2888), .Y(new_n2925));
  not_8  g00577(.A(n12657), .Y(new_n2926));
  xnor_4 g00578(.A(n27089), .B(new_n2926), .Y(new_n2927));
  nor_5  g00579(.A(n17077), .B(n11841), .Y(new_n2928));
  not_8  g00580(.A(n11841), .Y(new_n2929_1));
  xnor_4 g00581(.A(n17077), .B(new_n2929_1), .Y(new_n2930));
  not_8  g00582(.A(new_n2930), .Y(new_n2931));
  nor_5  g00583(.A(n26510), .B(n10710), .Y(new_n2932));
  not_8  g00584(.A(n10710), .Y(new_n2933));
  xnor_4 g00585(.A(n26510), .B(new_n2933), .Y(new_n2934));
  not_8  g00586(.A(new_n2934), .Y(new_n2935));
  nor_5  g00587(.A(n23068), .B(n20929), .Y(new_n2936));
  not_8  g00588(.A(n20929), .Y(new_n2937));
  xnor_4 g00589(.A(n23068), .B(new_n2937), .Y(new_n2938));
  not_8  g00590(.A(new_n2938), .Y(new_n2939));
  nor_5  g00591(.A(n19514), .B(n8006), .Y(new_n2940));
  not_8  g00592(.A(n8006), .Y(new_n2941));
  xnor_4 g00593(.A(n19514), .B(new_n2941), .Y(new_n2942));
  nor_5  g00594(.A(n25074), .B(n10053), .Y(new_n2943));
  not_8  g00595(.A(n10053), .Y(new_n2944_1));
  xnor_4 g00596(.A(n25074), .B(new_n2944_1), .Y(new_n2945));
  nor_5  g00597(.A(n16396), .B(n8399), .Y(new_n2946));
  not_8  g00598(.A(n8399), .Y(new_n2947));
  xnor_4 g00599(.A(n16396), .B(new_n2947), .Y(new_n2948_1));
  not_8  g00600(.A(new_n2948_1), .Y(new_n2949));
  nor_5  g00601(.A(n9507), .B(n9399), .Y(new_n2950));
  not_8  g00602(.A(n2088), .Y(new_n2951));
  not_8  g00603(.A(n26979), .Y(new_n2952));
  nor_5  g00604(.A(new_n2952), .B(new_n2951), .Y(new_n2953));
  xnor_4 g00605(.A(n9507), .B(n9399), .Y(new_n2954));
  nor_5  g00606(.A(new_n2954), .B(new_n2953), .Y(new_n2955));
  nor_5  g00607(.A(new_n2955), .B(new_n2950), .Y(new_n2956));
  nor_5  g00608(.A(new_n2956), .B(new_n2949), .Y(new_n2957));
  or_5   g00609(.A(new_n2957), .B(new_n2946), .Y(new_n2958));
  and_5  g00610(.A(new_n2958), .B(new_n2945), .Y(new_n2959));
  or_5   g00611(.A(new_n2959), .B(new_n2943), .Y(new_n2960));
  and_5  g00612(.A(new_n2960), .B(new_n2942), .Y(new_n2961_1));
  nor_5  g00613(.A(new_n2961_1), .B(new_n2940), .Y(new_n2962));
  nor_5  g00614(.A(new_n2962), .B(new_n2939), .Y(new_n2963));
  nor_5  g00615(.A(new_n2963), .B(new_n2936), .Y(new_n2964));
  nor_5  g00616(.A(new_n2964), .B(new_n2935), .Y(new_n2965));
  nor_5  g00617(.A(new_n2965), .B(new_n2932), .Y(new_n2966));
  nor_5  g00618(.A(new_n2966), .B(new_n2931), .Y(new_n2967));
  nor_5  g00619(.A(new_n2967), .B(new_n2928), .Y(new_n2968));
  xnor_4 g00620(.A(new_n2968), .B(new_n2927), .Y(new_n2969));
  xnor_4 g00621(.A(new_n2969), .B(new_n2925), .Y(new_n2970));
  nor_5  g00622(.A(new_n2921), .B(new_n2892), .Y(new_n2971_1));
  xnor_4 g00623(.A(new_n2971_1), .B(new_n2891), .Y(new_n2972));
  xnor_4 g00624(.A(new_n2966), .B(new_n2930), .Y(new_n2973));
  not_8  g00625(.A(new_n2973), .Y(new_n2974));
  nor_5  g00626(.A(new_n2974), .B(new_n2972), .Y(new_n2975));
  not_8  g00627(.A(new_n2972), .Y(new_n2976));
  xnor_4 g00628(.A(new_n2974), .B(new_n2976), .Y(new_n2977));
  nor_5  g00629(.A(new_n2919), .B(new_n2895), .Y(new_n2978_1));
  xnor_4 g00630(.A(new_n2978_1), .B(new_n2894), .Y(new_n2979_1));
  not_8  g00631(.A(new_n2979_1), .Y(new_n2980));
  xnor_4 g00632(.A(new_n2964), .B(new_n2934), .Y(new_n2981));
  nor_5  g00633(.A(new_n2981), .B(new_n2980), .Y(new_n2982));
  xnor_4 g00634(.A(new_n2981), .B(new_n2980), .Y(new_n2983));
  nor_5  g00635(.A(new_n2917), .B(new_n2898), .Y(new_n2984));
  xnor_4 g00636(.A(new_n2984), .B(new_n2897), .Y(new_n2985_1));
  not_8  g00637(.A(new_n2985_1), .Y(new_n2986));
  xnor_4 g00638(.A(new_n2962), .B(new_n2938), .Y(new_n2987));
  nor_5  g00639(.A(new_n2987), .B(new_n2986), .Y(new_n2988));
  xnor_4 g00640(.A(new_n2987), .B(new_n2986), .Y(new_n2989));
  xnor_4 g00641(.A(new_n2916), .B(new_n2899), .Y(new_n2990));
  nor_5  g00642(.A(new_n2959), .B(new_n2943), .Y(new_n2991));
  xnor_4 g00643(.A(new_n2991), .B(new_n2942), .Y(new_n2992));
  nor_5  g00644(.A(new_n2992), .B(new_n2990), .Y(new_n2993));
  not_8  g00645(.A(new_n2992), .Y(new_n2994));
  xnor_4 g00646(.A(new_n2994), .B(new_n2990), .Y(new_n2995));
  xnor_4 g00647(.A(new_n2914), .B(new_n2901), .Y(new_n2996));
  nor_5  g00648(.A(new_n2957), .B(new_n2946), .Y(new_n2997));
  xnor_4 g00649(.A(new_n2997), .B(new_n2945), .Y(new_n2998));
  nor_5  g00650(.A(new_n2998), .B(new_n2996), .Y(new_n2999_1));
  not_8  g00651(.A(new_n2998), .Y(new_n3000));
  xnor_4 g00652(.A(new_n3000), .B(new_n2996), .Y(new_n3001));
  xor_4  g00653(.A(new_n2912), .B(new_n2904), .Y(new_n3002));
  xnor_4 g00654(.A(new_n2956), .B(new_n2948_1), .Y(new_n3003));
  not_8  g00655(.A(new_n3003), .Y(new_n3004));
  nor_5  g00656(.A(new_n3004), .B(new_n3002), .Y(new_n3005));
  xnor_4 g00657(.A(new_n3003), .B(new_n3002), .Y(new_n3006));
  nor_5  g00658(.A(new_n2907), .B(new_n2906), .Y(new_n3007));
  xnor_4 g00659(.A(new_n2910), .B(new_n3007), .Y(new_n3008));
  not_8  g00660(.A(new_n3008), .Y(new_n3009));
  xnor_4 g00661(.A(new_n2954), .B(new_n2953), .Y(new_n3010_1));
  not_8  g00662(.A(new_n3010_1), .Y(new_n3011));
  nor_5  g00663(.A(new_n3011), .B(new_n3009), .Y(new_n3012));
  xnor_4 g00664(.A(n15780), .B(new_n2906), .Y(new_n3013));
  xnor_4 g00665(.A(n26979), .B(new_n2951), .Y(new_n3014));
  not_8  g00666(.A(new_n3014), .Y(new_n3015));
  nor_5  g00667(.A(new_n3015), .B(new_n3013), .Y(new_n3016));
  xnor_4 g00668(.A(new_n3010_1), .B(new_n3009), .Y(new_n3017_1));
  and_5  g00669(.A(new_n3017_1), .B(new_n3016), .Y(new_n3018_1));
  nor_5  g00670(.A(new_n3018_1), .B(new_n3012), .Y(new_n3019));
  and_5  g00671(.A(new_n3019), .B(new_n3006), .Y(new_n3020_1));
  nor_5  g00672(.A(new_n3020_1), .B(new_n3005), .Y(new_n3021));
  and_5  g00673(.A(new_n3021), .B(new_n3001), .Y(new_n3022));
  or_5   g00674(.A(new_n3022), .B(new_n2999_1), .Y(new_n3023));
  and_5  g00675(.A(new_n3023), .B(new_n2995), .Y(new_n3024));
  nor_5  g00676(.A(new_n3024), .B(new_n2993), .Y(new_n3025));
  nor_5  g00677(.A(new_n3025), .B(new_n2989), .Y(new_n3026));
  nor_5  g00678(.A(new_n3026), .B(new_n2988), .Y(new_n3027));
  nor_5  g00679(.A(new_n3027), .B(new_n2983), .Y(new_n3028));
  nor_5  g00680(.A(new_n3028), .B(new_n2982), .Y(new_n3029));
  and_5  g00681(.A(new_n3029), .B(new_n2977), .Y(new_n3030_1));
  or_5   g00682(.A(new_n3030_1), .B(new_n2975), .Y(new_n3031));
  xor_4  g00683(.A(new_n3031), .B(new_n2970), .Y(new_n3032));
  xnor_4 g00684(.A(new_n3032), .B(new_n2886_1), .Y(new_n3033));
  xor_4  g00685(.A(new_n2883), .B(new_n2852), .Y(new_n3034));
  xor_4  g00686(.A(new_n3029), .B(new_n2977), .Y(new_n3035));
  nor_5  g00687(.A(new_n3035), .B(new_n3034), .Y(new_n3036));
  xnor_4 g00688(.A(new_n3035), .B(new_n3034), .Y(new_n3037));
  xor_4  g00689(.A(new_n2881), .B(new_n2855), .Y(new_n3038));
  xnor_4 g00690(.A(new_n3027), .B(new_n2983), .Y(new_n3039));
  nor_5  g00691(.A(new_n3039), .B(new_n3038), .Y(new_n3040));
  xnor_4 g00692(.A(new_n3039), .B(new_n3038), .Y(new_n3041));
  xor_4  g00693(.A(new_n2879), .B(new_n2858_1), .Y(new_n3042));
  xnor_4 g00694(.A(new_n3025), .B(new_n2989), .Y(new_n3043));
  nor_5  g00695(.A(new_n3043), .B(new_n3042), .Y(new_n3044));
  xnor_4 g00696(.A(new_n3043), .B(new_n3042), .Y(new_n3045));
  xor_4  g00697(.A(new_n2877), .B(new_n2861), .Y(new_n3046));
  nor_5  g00698(.A(new_n3022), .B(new_n2999_1), .Y(new_n3047));
  xnor_4 g00699(.A(new_n3047), .B(new_n2995), .Y(new_n3048));
  not_8  g00700(.A(new_n3048), .Y(new_n3049));
  nor_5  g00701(.A(new_n3049), .B(new_n3046), .Y(new_n3050));
  xnor_4 g00702(.A(new_n3049), .B(new_n3046), .Y(new_n3051));
  xnor_4 g00703(.A(new_n3021), .B(new_n3001), .Y(new_n3052));
  not_8  g00704(.A(new_n3052), .Y(new_n3053));
  xnor_4 g00705(.A(new_n2875), .B(new_n2864), .Y(new_n3054));
  and_5  g00706(.A(new_n3054), .B(new_n3053), .Y(new_n3055));
  xnor_4 g00707(.A(new_n3054), .B(new_n3053), .Y(new_n3056));
  xnor_4 g00708(.A(new_n3019), .B(new_n3006), .Y(new_n3057));
  xnor_4 g00709(.A(n19005), .B(n7149), .Y(new_n3058));
  xnor_4 g00710(.A(new_n3058), .B(new_n2873), .Y(new_n3059));
  and_5  g00711(.A(new_n3059), .B(new_n3057), .Y(new_n3060));
  xnor_4 g00712(.A(new_n3059), .B(new_n3057), .Y(new_n3061));
  xnor_4 g00713(.A(n5438), .B(n1152), .Y(new_n3062));
  not_8  g00714(.A(new_n3013), .Y(new_n3063));
  xnor_4 g00715(.A(new_n3015), .B(new_n3063), .Y(new_n3064));
  nor_5  g00716(.A(new_n3064), .B(new_n3062), .Y(new_n3065));
  xnor_4 g00717(.A(n14148), .B(n4326), .Y(new_n3066));
  xnor_4 g00718(.A(new_n3066), .B(new_n2871), .Y(new_n3067_1));
  nor_5  g00719(.A(new_n3067_1), .B(new_n3065), .Y(new_n3068));
  xnor_4 g00720(.A(new_n3017_1), .B(new_n3016), .Y(new_n3069));
  xnor_4 g00721(.A(new_n3067_1), .B(new_n3065), .Y(new_n3070));
  nor_5  g00722(.A(new_n3070), .B(new_n3069), .Y(new_n3071));
  nor_5  g00723(.A(new_n3071), .B(new_n3068), .Y(new_n3072));
  nor_5  g00724(.A(new_n3072), .B(new_n3061), .Y(new_n3073));
  nor_5  g00725(.A(new_n3073), .B(new_n3060), .Y(new_n3074));
  nor_5  g00726(.A(new_n3074), .B(new_n3056), .Y(new_n3075));
  nor_5  g00727(.A(new_n3075), .B(new_n3055), .Y(new_n3076_1));
  nor_5  g00728(.A(new_n3076_1), .B(new_n3051), .Y(new_n3077));
  nor_5  g00729(.A(new_n3077), .B(new_n3050), .Y(new_n3078));
  nor_5  g00730(.A(new_n3078), .B(new_n3045), .Y(new_n3079));
  nor_5  g00731(.A(new_n3079), .B(new_n3044), .Y(new_n3080));
  nor_5  g00732(.A(new_n3080), .B(new_n3041), .Y(new_n3081));
  nor_5  g00733(.A(new_n3081), .B(new_n3040), .Y(new_n3082));
  nor_5  g00734(.A(new_n3082), .B(new_n3037), .Y(new_n3083));
  nor_5  g00735(.A(new_n3083), .B(new_n3036), .Y(new_n3084));
  xnor_4 g00736(.A(new_n3084), .B(new_n3033), .Y(n142));
  not_8  g00737(.A(n5025), .Y(new_n3086));
  not_8  g00738(.A(n4319), .Y(new_n3087));
  xnor_4 g00739(.A(n7335), .B(new_n3087), .Y(new_n3088));
  not_8  g00740(.A(new_n3088), .Y(new_n3089_1));
  nor_5  g00741(.A(n23463), .B(n5696), .Y(new_n3090));
  not_8  g00742(.A(n5696), .Y(new_n3091));
  xnor_4 g00743(.A(n23463), .B(new_n3091), .Y(new_n3092));
  not_8  g00744(.A(new_n3092), .Y(new_n3093));
  nor_5  g00745(.A(n13367), .B(n13074), .Y(new_n3094));
  not_8  g00746(.A(n13074), .Y(new_n3095));
  xnor_4 g00747(.A(n13367), .B(new_n3095), .Y(new_n3096));
  not_8  g00748(.A(new_n3096), .Y(new_n3097));
  nor_5  g00749(.A(n10739), .B(n932), .Y(new_n3098));
  not_8  g00750(.A(n10739), .Y(new_n3099));
  xnor_4 g00751(.A(new_n3099), .B(n932), .Y(new_n3100));
  not_8  g00752(.A(new_n3100), .Y(new_n3101));
  nor_5  g00753(.A(n21753), .B(n6691), .Y(new_n3102));
  xnor_4 g00754(.A(new_n2350), .B(n6691), .Y(new_n3103));
  not_8  g00755(.A(new_n3103), .Y(new_n3104));
  nor_5  g00756(.A(n21832), .B(n3260), .Y(new_n3105));
  not_8  g00757(.A(n3260), .Y(new_n3106));
  xnor_4 g00758(.A(n21832), .B(new_n3106), .Y(new_n3107));
  not_8  g00759(.A(new_n3107), .Y(new_n3108));
  nor_5  g00760(.A(n26913), .B(n20489), .Y(new_n3109));
  not_8  g00761(.A(n20489), .Y(new_n3110));
  xnor_4 g00762(.A(n26913), .B(new_n3110), .Y(new_n3111));
  not_8  g00763(.A(new_n3111), .Y(new_n3112));
  nor_5  g00764(.A(n16223), .B(n2355), .Y(new_n3113));
  xnor_4 g00765(.A(n16223), .B(n2355), .Y(new_n3114));
  nor_5  g00766(.A(n19494), .B(n11121), .Y(new_n3115));
  not_8  g00767(.A(n2387), .Y(new_n3116));
  not_8  g00768(.A(n16217), .Y(new_n3117));
  nor_5  g00769(.A(new_n3117), .B(new_n3116), .Y(new_n3118));
  xnor_4 g00770(.A(new_n2365), .B(n11121), .Y(new_n3119));
  not_8  g00771(.A(new_n3119), .Y(new_n3120));
  nor_5  g00772(.A(new_n3120), .B(new_n3118), .Y(new_n3121));
  nor_5  g00773(.A(new_n3121), .B(new_n3115), .Y(new_n3122));
  nor_5  g00774(.A(new_n3122), .B(new_n3114), .Y(new_n3123));
  nor_5  g00775(.A(new_n3123), .B(new_n3113), .Y(new_n3124));
  nor_5  g00776(.A(new_n3124), .B(new_n3112), .Y(new_n3125_1));
  nor_5  g00777(.A(new_n3125_1), .B(new_n3109), .Y(new_n3126_1));
  nor_5  g00778(.A(new_n3126_1), .B(new_n3108), .Y(new_n3127));
  nor_5  g00779(.A(new_n3127), .B(new_n3105), .Y(new_n3128));
  nor_5  g00780(.A(new_n3128), .B(new_n3104), .Y(new_n3129));
  nor_5  g00781(.A(new_n3129), .B(new_n3102), .Y(new_n3130));
  nor_5  g00782(.A(new_n3130), .B(new_n3101), .Y(new_n3131));
  nor_5  g00783(.A(new_n3131), .B(new_n3098), .Y(new_n3132));
  nor_5  g00784(.A(new_n3132), .B(new_n3097), .Y(new_n3133));
  nor_5  g00785(.A(new_n3133), .B(new_n3094), .Y(new_n3134));
  nor_5  g00786(.A(new_n3134), .B(new_n3093), .Y(new_n3135));
  nor_5  g00787(.A(new_n3135), .B(new_n3090), .Y(new_n3136_1));
  xnor_4 g00788(.A(new_n3136_1), .B(new_n3089_1), .Y(new_n3137));
  and_5  g00789(.A(new_n3137), .B(new_n3086), .Y(new_n3138));
  xnor_4 g00790(.A(new_n3137), .B(new_n3086), .Y(new_n3139));
  not_8  g00791(.A(n6485), .Y(new_n3140));
  xnor_4 g00792(.A(new_n3134), .B(new_n3093), .Y(new_n3141));
  and_5  g00793(.A(new_n3141), .B(new_n3140), .Y(new_n3142));
  xnor_4 g00794(.A(new_n3141), .B(new_n3140), .Y(new_n3143));
  not_8  g00795(.A(n26036), .Y(new_n3144));
  xnor_4 g00796(.A(new_n3132), .B(new_n3097), .Y(new_n3145));
  and_5  g00797(.A(new_n3145), .B(new_n3144), .Y(new_n3146));
  xnor_4 g00798(.A(new_n3145), .B(new_n3144), .Y(new_n3147));
  not_8  g00799(.A(n19770), .Y(new_n3148));
  xnor_4 g00800(.A(new_n3130), .B(new_n3101), .Y(new_n3149));
  and_5  g00801(.A(new_n3149), .B(new_n3148), .Y(new_n3150));
  xnor_4 g00802(.A(new_n3149), .B(new_n3148), .Y(new_n3151));
  not_8  g00803(.A(n8782), .Y(new_n3152));
  xnor_4 g00804(.A(new_n3128), .B(new_n3104), .Y(new_n3153));
  and_5  g00805(.A(new_n3153), .B(new_n3152), .Y(new_n3154));
  xnor_4 g00806(.A(new_n3153), .B(new_n3152), .Y(new_n3155));
  not_8  g00807(.A(n8678), .Y(new_n3156));
  xnor_4 g00808(.A(new_n3126_1), .B(new_n3108), .Y(new_n3157));
  and_5  g00809(.A(new_n3157), .B(new_n3156), .Y(new_n3158));
  xnor_4 g00810(.A(new_n3157), .B(new_n3156), .Y(new_n3159));
  xnor_4 g00811(.A(new_n3124), .B(new_n3111), .Y(new_n3160));
  nor_5  g00812(.A(new_n3160), .B(n1432), .Y(new_n3161_1));
  not_8  g00813(.A(n1432), .Y(new_n3162));
  not_8  g00814(.A(new_n3160), .Y(new_n3163));
  xnor_4 g00815(.A(new_n3163), .B(new_n3162), .Y(new_n3164_1));
  xnor_4 g00816(.A(new_n3122), .B(new_n3114), .Y(new_n3165));
  not_8  g00817(.A(new_n3165), .Y(new_n3166));
  nor_5  g00818(.A(new_n3166), .B(n21599), .Y(new_n3167));
  xnor_4 g00819(.A(new_n3166), .B(n21599), .Y(new_n3168));
  not_8  g00820(.A(n25336), .Y(new_n3169));
  xnor_4 g00821(.A(n16217), .B(n2387), .Y(new_n3170));
  nor_5  g00822(.A(new_n3170), .B(n11424), .Y(new_n3171));
  and_5  g00823(.A(new_n3171), .B(new_n3169), .Y(new_n3172));
  xnor_4 g00824(.A(new_n3171), .B(new_n3169), .Y(new_n3173));
  xnor_4 g00825(.A(new_n3119), .B(new_n3118), .Y(new_n3174));
  nor_5  g00826(.A(new_n3174), .B(new_n3173), .Y(new_n3175));
  nor_5  g00827(.A(new_n3175), .B(new_n3172), .Y(new_n3176));
  nor_5  g00828(.A(new_n3176), .B(new_n3168), .Y(new_n3177));
  nor_5  g00829(.A(new_n3177), .B(new_n3167), .Y(new_n3178));
  nor_5  g00830(.A(new_n3178), .B(new_n3164_1), .Y(new_n3179));
  nor_5  g00831(.A(new_n3179), .B(new_n3161_1), .Y(new_n3180));
  nor_5  g00832(.A(new_n3180), .B(new_n3159), .Y(new_n3181));
  nor_5  g00833(.A(new_n3181), .B(new_n3158), .Y(new_n3182));
  nor_5  g00834(.A(new_n3182), .B(new_n3155), .Y(new_n3183));
  nor_5  g00835(.A(new_n3183), .B(new_n3154), .Y(new_n3184));
  nor_5  g00836(.A(new_n3184), .B(new_n3151), .Y(new_n3185));
  nor_5  g00837(.A(new_n3185), .B(new_n3150), .Y(new_n3186));
  nor_5  g00838(.A(new_n3186), .B(new_n3147), .Y(new_n3187));
  nor_5  g00839(.A(new_n3187), .B(new_n3146), .Y(new_n3188));
  nor_5  g00840(.A(new_n3188), .B(new_n3143), .Y(new_n3189));
  nor_5  g00841(.A(new_n3189), .B(new_n3142), .Y(new_n3190));
  nor_5  g00842(.A(new_n3190), .B(new_n3139), .Y(new_n3191));
  nor_5  g00843(.A(new_n3191), .B(new_n3138), .Y(new_n3192));
  nor_5  g00844(.A(n7335), .B(n4319), .Y(new_n3193));
  nor_5  g00845(.A(new_n3136_1), .B(new_n3089_1), .Y(new_n3194));
  nor_5  g00846(.A(new_n3194), .B(new_n3193), .Y(new_n3195));
  not_8  g00847(.A(new_n3195), .Y(new_n3196));
  nand_5 g00848(.A(new_n3196), .B(new_n3192), .Y(new_n3197));
  not_8  g00849(.A(n9967), .Y(new_n3198));
  nor_5  g00850(.A(n12315), .B(n3952), .Y(new_n3199));
  not_8  g00851(.A(new_n3199), .Y(new_n3200));
  nor_5  g00852(.A(new_n3200), .B(n24618), .Y(new_n3201));
  not_8  g00853(.A(new_n3201), .Y(new_n3202));
  nor_5  g00854(.A(new_n3202), .B(n24278), .Y(new_n3203));
  not_8  g00855(.A(new_n3203), .Y(new_n3204));
  nor_5  g00856(.A(new_n3204), .B(n4812), .Y(new_n3205));
  not_8  g00857(.A(new_n3205), .Y(new_n3206));
  nor_5  g00858(.A(new_n3206), .B(n26823), .Y(new_n3207));
  not_8  g00859(.A(new_n3207), .Y(new_n3208_1));
  nor_5  g00860(.A(new_n3208_1), .B(n7751), .Y(new_n3209));
  not_8  g00861(.A(new_n3209), .Y(new_n3210));
  nor_5  g00862(.A(new_n3210), .B(n20946), .Y(new_n3211));
  and_5  g00863(.A(new_n3211), .B(new_n3198), .Y(new_n3212));
  xnor_4 g00864(.A(new_n3212), .B(n3425), .Y(new_n3213));
  not_8  g00865(.A(new_n3213), .Y(new_n3214));
  xor_4  g00866(.A(new_n3190), .B(new_n3139), .Y(new_n3215));
  nor_5  g00867(.A(new_n3215), .B(new_n3214), .Y(new_n3216));
  not_8  g00868(.A(n3425), .Y(new_n3217));
  and_5  g00869(.A(new_n3212), .B(new_n3217), .Y(new_n3218));
  xnor_4 g00870(.A(new_n3215), .B(new_n3214), .Y(new_n3219_1));
  xnor_4 g00871(.A(new_n3211), .B(n9967), .Y(new_n3220));
  not_8  g00872(.A(new_n3220), .Y(new_n3221));
  xor_4  g00873(.A(new_n3188), .B(new_n3143), .Y(new_n3222));
  nor_5  g00874(.A(new_n3222), .B(new_n3221), .Y(new_n3223));
  not_8  g00875(.A(new_n3222), .Y(new_n3224));
  xnor_4 g00876(.A(new_n3224), .B(new_n3220), .Y(new_n3225));
  xnor_4 g00877(.A(new_n3209), .B(n20946), .Y(new_n3226));
  not_8  g00878(.A(new_n3226), .Y(new_n3227));
  xor_4  g00879(.A(new_n3186), .B(new_n3147), .Y(new_n3228_1));
  nor_5  g00880(.A(new_n3228_1), .B(new_n3227), .Y(new_n3229));
  xnor_4 g00881(.A(new_n3228_1), .B(new_n3227), .Y(new_n3230));
  xnor_4 g00882(.A(new_n3207), .B(n7751), .Y(new_n3231));
  not_8  g00883(.A(new_n3231), .Y(new_n3232));
  xor_4  g00884(.A(new_n3184), .B(new_n3151), .Y(new_n3233));
  nor_5  g00885(.A(new_n3233), .B(new_n3232), .Y(new_n3234));
  xnor_4 g00886(.A(new_n3233), .B(new_n3232), .Y(new_n3235_1));
  xnor_4 g00887(.A(new_n3205), .B(n26823), .Y(new_n3236));
  not_8  g00888(.A(new_n3236), .Y(new_n3237));
  xor_4  g00889(.A(new_n3182), .B(new_n3155), .Y(new_n3238));
  nor_5  g00890(.A(new_n3238), .B(new_n3237), .Y(new_n3239));
  xnor_4 g00891(.A(new_n3238), .B(new_n3237), .Y(new_n3240));
  xnor_4 g00892(.A(new_n3203), .B(n4812), .Y(new_n3241));
  not_8  g00893(.A(new_n3241), .Y(new_n3242));
  xor_4  g00894(.A(new_n3180), .B(new_n3159), .Y(new_n3243));
  nor_5  g00895(.A(new_n3243), .B(new_n3242), .Y(new_n3244_1));
  xnor_4 g00896(.A(new_n3243), .B(new_n3242), .Y(new_n3245));
  xnor_4 g00897(.A(new_n3201), .B(n24278), .Y(new_n3246));
  not_8  g00898(.A(new_n3246), .Y(new_n3247));
  xor_4  g00899(.A(new_n3178), .B(new_n3164_1), .Y(new_n3248));
  nor_5  g00900(.A(new_n3248), .B(new_n3247), .Y(new_n3249));
  xnor_4 g00901(.A(new_n3248), .B(new_n3247), .Y(new_n3250));
  xnor_4 g00902(.A(new_n3199), .B(n24618), .Y(new_n3251));
  not_8  g00903(.A(new_n3251), .Y(new_n3252));
  xor_4  g00904(.A(new_n3176), .B(new_n3168), .Y(new_n3253_1));
  nor_5  g00905(.A(new_n3253_1), .B(new_n3252), .Y(new_n3254));
  xnor_4 g00906(.A(new_n3253_1), .B(new_n3252), .Y(new_n3255));
  not_8  g00907(.A(n11424), .Y(new_n3256));
  xnor_4 g00908(.A(new_n3170), .B(new_n3256), .Y(new_n3257));
  nor_5  g00909(.A(new_n3257), .B(new_n2448), .Y(new_n3258));
  and_5  g00910(.A(new_n3258), .B(new_n2443), .Y(new_n3259));
  xnor_4 g00911(.A(new_n3120), .B(new_n3118), .Y(new_n3260_1));
  xnor_4 g00912(.A(new_n3260_1), .B(new_n3173), .Y(new_n3261));
  xnor_4 g00913(.A(n12315), .B(new_n2443), .Y(new_n3262));
  nor_5  g00914(.A(new_n3262), .B(new_n3258), .Y(new_n3263_1));
  or_5   g00915(.A(new_n3263_1), .B(new_n3259), .Y(new_n3264));
  nor_5  g00916(.A(new_n3264), .B(new_n3261), .Y(new_n3265));
  nor_5  g00917(.A(new_n3265), .B(new_n3259), .Y(new_n3266));
  nor_5  g00918(.A(new_n3266), .B(new_n3255), .Y(new_n3267));
  nor_5  g00919(.A(new_n3267), .B(new_n3254), .Y(new_n3268));
  nor_5  g00920(.A(new_n3268), .B(new_n3250), .Y(new_n3269));
  nor_5  g00921(.A(new_n3269), .B(new_n3249), .Y(new_n3270));
  nor_5  g00922(.A(new_n3270), .B(new_n3245), .Y(new_n3271));
  nor_5  g00923(.A(new_n3271), .B(new_n3244_1), .Y(new_n3272));
  nor_5  g00924(.A(new_n3272), .B(new_n3240), .Y(new_n3273));
  nor_5  g00925(.A(new_n3273), .B(new_n3239), .Y(new_n3274));
  nor_5  g00926(.A(new_n3274), .B(new_n3235_1), .Y(new_n3275));
  nor_5  g00927(.A(new_n3275), .B(new_n3234), .Y(new_n3276));
  nor_5  g00928(.A(new_n3276), .B(new_n3230), .Y(new_n3277));
  nor_5  g00929(.A(new_n3277), .B(new_n3229), .Y(new_n3278));
  nor_5  g00930(.A(new_n3278), .B(new_n3225), .Y(new_n3279_1));
  nor_5  g00931(.A(new_n3279_1), .B(new_n3223), .Y(new_n3280));
  nor_5  g00932(.A(new_n3280), .B(new_n3219_1), .Y(new_n3281));
  or_5   g00933(.A(new_n3281), .B(new_n3218), .Y(new_n3282));
  nor_5  g00934(.A(new_n3282), .B(new_n3216), .Y(new_n3283));
  not_8  g00935(.A(new_n3283), .Y(new_n3284));
  nor_5  g00936(.A(new_n3284), .B(new_n3197), .Y(new_n3285));
  nor_5  g00937(.A(n7593), .B(n5101), .Y(new_n3286));
  xnor_4 g00938(.A(n7593), .B(n5101), .Y(new_n3287));
  nor_5  g00939(.A(n16507), .B(n337), .Y(new_n3288));
  xnor_4 g00940(.A(n16507), .B(n337), .Y(new_n3289_1));
  nor_5  g00941(.A(n22470), .B(n3228), .Y(new_n3290));
  xnor_4 g00942(.A(n22470), .B(n3228), .Y(new_n3291));
  nor_5  g00943(.A(n19116), .B(n5302), .Y(new_n3292));
  xnor_4 g00944(.A(n19116), .B(n5302), .Y(new_n3293));
  nor_5  g00945(.A(n25738), .B(n6861), .Y(new_n3294));
  xnor_4 g00946(.A(n25738), .B(n6861), .Y(new_n3295));
  nor_5  g00947(.A(n21471), .B(n19357), .Y(new_n3296));
  xnor_4 g00948(.A(n21471), .B(n19357), .Y(new_n3297));
  nor_5  g00949(.A(n18737), .B(n2328), .Y(new_n3298));
  xnor_4 g00950(.A(n18737), .B(n2328), .Y(new_n3299));
  nor_5  g00951(.A(n15053), .B(n14603), .Y(new_n3300));
  not_8  g00952(.A(n14603), .Y(new_n3301_1));
  xnor_4 g00953(.A(n15053), .B(new_n3301_1), .Y(new_n3302));
  nor_5  g00954(.A(n25471), .B(n20794), .Y(new_n3303));
  not_8  g00955(.A(n16502), .Y(new_n3304));
  not_8  g00956(.A(n23333), .Y(new_n3305));
  nor_5  g00957(.A(new_n3305), .B(new_n3304), .Y(new_n3306_1));
  not_8  g00958(.A(n20794), .Y(new_n3307));
  xnor_4 g00959(.A(n25471), .B(new_n3307), .Y(new_n3308));
  not_8  g00960(.A(new_n3308), .Y(new_n3309));
  nor_5  g00961(.A(new_n3309), .B(new_n3306_1), .Y(new_n3310));
  or_5   g00962(.A(new_n3310), .B(new_n3303), .Y(new_n3311));
  and_5  g00963(.A(new_n3311), .B(new_n3302), .Y(new_n3312));
  nor_5  g00964(.A(new_n3312), .B(new_n3300), .Y(new_n3313));
  nor_5  g00965(.A(new_n3313), .B(new_n3299), .Y(new_n3314));
  nor_5  g00966(.A(new_n3314), .B(new_n3298), .Y(new_n3315));
  nor_5  g00967(.A(new_n3315), .B(new_n3297), .Y(new_n3316_1));
  nor_5  g00968(.A(new_n3316_1), .B(new_n3296), .Y(new_n3317));
  nor_5  g00969(.A(new_n3317), .B(new_n3295), .Y(new_n3318));
  nor_5  g00970(.A(new_n3318), .B(new_n3294), .Y(new_n3319));
  nor_5  g00971(.A(new_n3319), .B(new_n3293), .Y(new_n3320_1));
  nor_5  g00972(.A(new_n3320_1), .B(new_n3292), .Y(new_n3321));
  nor_5  g00973(.A(new_n3321), .B(new_n3291), .Y(new_n3322));
  nor_5  g00974(.A(new_n3322), .B(new_n3290), .Y(new_n3323));
  nor_5  g00975(.A(new_n3323), .B(new_n3289_1), .Y(new_n3324_1));
  nor_5  g00976(.A(new_n3324_1), .B(new_n3288), .Y(new_n3325));
  nor_5  g00977(.A(new_n3325), .B(new_n3287), .Y(new_n3326));
  nor_5  g00978(.A(new_n3326), .B(new_n3286), .Y(new_n3327));
  xnor_4 g00979(.A(new_n3196), .B(new_n3192), .Y(new_n3328));
  not_8  g00980(.A(new_n3328), .Y(new_n3329));
  xnor_4 g00981(.A(new_n3329), .B(new_n3284), .Y(new_n3330));
  and_5  g00982(.A(new_n3330), .B(new_n3327), .Y(new_n3331));
  nor_5  g00983(.A(new_n3330), .B(new_n3327), .Y(new_n3332_1));
  xor_4  g00984(.A(new_n3280), .B(new_n3219_1), .Y(new_n3333));
  xnor_4 g00985(.A(new_n3325), .B(new_n3287), .Y(new_n3334));
  nor_5  g00986(.A(new_n3334), .B(new_n3333), .Y(new_n3335));
  xnor_4 g00987(.A(new_n3334), .B(new_n3333), .Y(new_n3336));
  xor_4  g00988(.A(new_n3278), .B(new_n3225), .Y(new_n3337));
  xnor_4 g00989(.A(new_n3323), .B(new_n3289_1), .Y(new_n3338));
  nor_5  g00990(.A(new_n3338), .B(new_n3337), .Y(new_n3339));
  xnor_4 g00991(.A(new_n3338), .B(new_n3337), .Y(new_n3340_1));
  xor_4  g00992(.A(new_n3276), .B(new_n3230), .Y(new_n3341));
  xnor_4 g00993(.A(new_n3321), .B(new_n3291), .Y(new_n3342));
  nor_5  g00994(.A(new_n3342), .B(new_n3341), .Y(new_n3343_1));
  xnor_4 g00995(.A(new_n3342), .B(new_n3341), .Y(new_n3344));
  xor_4  g00996(.A(new_n3274), .B(new_n3235_1), .Y(new_n3345));
  xnor_4 g00997(.A(new_n3319), .B(new_n3293), .Y(new_n3346));
  nor_5  g00998(.A(new_n3346), .B(new_n3345), .Y(new_n3347));
  xnor_4 g00999(.A(new_n3346), .B(new_n3345), .Y(new_n3348));
  xor_4  g01000(.A(new_n3272), .B(new_n3240), .Y(new_n3349_1));
  xnor_4 g01001(.A(new_n3317), .B(new_n3295), .Y(new_n3350));
  nor_5  g01002(.A(new_n3350), .B(new_n3349_1), .Y(new_n3351));
  xnor_4 g01003(.A(new_n3350), .B(new_n3349_1), .Y(new_n3352));
  xor_4  g01004(.A(new_n3270), .B(new_n3245), .Y(new_n3353));
  xnor_4 g01005(.A(new_n3315), .B(new_n3297), .Y(new_n3354));
  nor_5  g01006(.A(new_n3354), .B(new_n3353), .Y(new_n3355));
  xnor_4 g01007(.A(new_n3354), .B(new_n3353), .Y(new_n3356));
  xor_4  g01008(.A(new_n3268), .B(new_n3250), .Y(new_n3357));
  xnor_4 g01009(.A(new_n3313), .B(new_n3299), .Y(new_n3358));
  nor_5  g01010(.A(new_n3358), .B(new_n3357), .Y(new_n3359));
  xnor_4 g01011(.A(new_n3358), .B(new_n3357), .Y(new_n3360));
  xor_4  g01012(.A(new_n3266), .B(new_n3255), .Y(new_n3361));
  nor_5  g01013(.A(new_n3310), .B(new_n3303), .Y(new_n3362));
  xnor_4 g01014(.A(new_n3362), .B(new_n3302), .Y(new_n3363));
  not_8  g01015(.A(new_n3363), .Y(new_n3364));
  nor_5  g01016(.A(new_n3364), .B(new_n3361), .Y(new_n3365));
  xnor_4 g01017(.A(new_n3364), .B(new_n3361), .Y(new_n3366_1));
  xnor_4 g01018(.A(n23333), .B(new_n3304), .Y(new_n3367));
  xnor_4 g01019(.A(new_n3257), .B(n12315), .Y(new_n3368));
  and_5  g01020(.A(new_n3368), .B(new_n3367), .Y(new_n3369));
  xnor_4 g01021(.A(new_n3309), .B(new_n3306_1), .Y(new_n3370));
  nor_5  g01022(.A(new_n3370), .B(new_n3369), .Y(new_n3371));
  xor_4  g01023(.A(new_n3264), .B(new_n3261), .Y(new_n3372));
  not_8  g01024(.A(new_n3372), .Y(new_n3373));
  and_5  g01025(.A(new_n3369), .B(new_n3308), .Y(new_n3374));
  nor_5  g01026(.A(new_n3374), .B(new_n3371), .Y(new_n3375));
  and_5  g01027(.A(new_n3375), .B(new_n3373), .Y(new_n3376));
  nor_5  g01028(.A(new_n3376), .B(new_n3371), .Y(new_n3377));
  nor_5  g01029(.A(new_n3377), .B(new_n3366_1), .Y(new_n3378));
  nor_5  g01030(.A(new_n3378), .B(new_n3365), .Y(new_n3379));
  nor_5  g01031(.A(new_n3379), .B(new_n3360), .Y(new_n3380));
  nor_5  g01032(.A(new_n3380), .B(new_n3359), .Y(new_n3381));
  nor_5  g01033(.A(new_n3381), .B(new_n3356), .Y(new_n3382));
  nor_5  g01034(.A(new_n3382), .B(new_n3355), .Y(new_n3383));
  nor_5  g01035(.A(new_n3383), .B(new_n3352), .Y(new_n3384));
  nor_5  g01036(.A(new_n3384), .B(new_n3351), .Y(new_n3385));
  nor_5  g01037(.A(new_n3385), .B(new_n3348), .Y(new_n3386));
  nor_5  g01038(.A(new_n3386), .B(new_n3347), .Y(new_n3387));
  nor_5  g01039(.A(new_n3387), .B(new_n3344), .Y(new_n3388));
  nor_5  g01040(.A(new_n3388), .B(new_n3343_1), .Y(new_n3389));
  nor_5  g01041(.A(new_n3389), .B(new_n3340_1), .Y(new_n3390_1));
  nor_5  g01042(.A(new_n3390_1), .B(new_n3339), .Y(new_n3391));
  nor_5  g01043(.A(new_n3391), .B(new_n3336), .Y(new_n3392));
  or_5   g01044(.A(new_n3392), .B(new_n3335), .Y(new_n3393));
  nor_5  g01045(.A(new_n3393), .B(new_n3332_1), .Y(new_n3394));
  nor_5  g01046(.A(new_n3394), .B(new_n3331), .Y(new_n3395));
  not_8  g01047(.A(new_n3395), .Y(new_n3396));
  and_5  g01048(.A(new_n3396), .B(new_n3285), .Y(new_n3397));
  nor_5  g01049(.A(new_n3283), .B(new_n3197), .Y(new_n3398));
  or_5   g01050(.A(new_n3196), .B(new_n3192), .Y(new_n3399));
  nor_5  g01051(.A(new_n3399), .B(new_n3284), .Y(new_n3400));
  or_5   g01052(.A(new_n3400), .B(new_n3398), .Y(new_n3401));
  nor_5  g01053(.A(new_n3401), .B(new_n3395), .Y(new_n3402));
  nor_5  g01054(.A(new_n3402), .B(new_n3285), .Y(new_n3403));
  nor_5  g01055(.A(new_n3403), .B(new_n3397), .Y(n175));
  not_8  g01056(.A(n14130), .Y(new_n3405));
  nor_5  g01057(.A(n20138), .B(n9251), .Y(new_n3406));
  not_8  g01058(.A(new_n3406), .Y(new_n3407));
  nor_5  g01059(.A(new_n3407), .B(n6385), .Y(new_n3408));
  not_8  g01060(.A(new_n3408), .Y(new_n3409));
  nor_5  g01061(.A(new_n3409), .B(n3136), .Y(new_n3410));
  not_8  g01062(.A(new_n3410), .Y(new_n3411));
  nor_5  g01063(.A(new_n3411), .B(n9557), .Y(new_n3412));
  not_8  g01064(.A(new_n3412), .Y(new_n3413));
  nor_5  g01065(.A(new_n3413), .B(n25643), .Y(new_n3414));
  not_8  g01066(.A(new_n3414), .Y(new_n3415));
  nor_5  g01067(.A(new_n3415), .B(n9942), .Y(new_n3416));
  not_8  g01068(.A(new_n3416), .Y(new_n3417));
  nor_5  g01069(.A(new_n3417), .B(n16482), .Y(new_n3418));
  and_5  g01070(.A(new_n3418), .B(new_n3405), .Y(new_n3419));
  xnor_4 g01071(.A(new_n3419), .B(n8856), .Y(new_n3420));
  xnor_4 g01072(.A(new_n3420), .B(n25494), .Y(new_n3421));
  xnor_4 g01073(.A(new_n3418), .B(n14130), .Y(new_n3422));
  nor_5  g01074(.A(new_n3422), .B(n10117), .Y(new_n3423));
  not_8  g01075(.A(n10117), .Y(new_n3424));
  xnor_4 g01076(.A(new_n3422), .B(new_n3424), .Y(new_n3425_1));
  xnor_4 g01077(.A(new_n3416), .B(n16482), .Y(new_n3426_1));
  nor_5  g01078(.A(new_n3426_1), .B(n13460), .Y(new_n3427));
  not_8  g01079(.A(n13460), .Y(new_n3428));
  xnor_4 g01080(.A(new_n3426_1), .B(new_n3428), .Y(new_n3429));
  xnor_4 g01081(.A(new_n3414), .B(n9942), .Y(new_n3430));
  nor_5  g01082(.A(new_n3430), .B(n6104), .Y(new_n3431));
  not_8  g01083(.A(n6104), .Y(new_n3432));
  xnor_4 g01084(.A(new_n3430), .B(new_n3432), .Y(new_n3433));
  xnor_4 g01085(.A(new_n3412), .B(n25643), .Y(new_n3434));
  nor_5  g01086(.A(new_n3434), .B(n4119), .Y(new_n3435));
  not_8  g01087(.A(n4119), .Y(new_n3436));
  xnor_4 g01088(.A(new_n3434), .B(new_n3436), .Y(new_n3437));
  xnor_4 g01089(.A(new_n3410), .B(n9557), .Y(new_n3438));
  nor_5  g01090(.A(new_n3438), .B(n14510), .Y(new_n3439));
  not_8  g01091(.A(n14510), .Y(new_n3440));
  xnor_4 g01092(.A(new_n3438), .B(new_n3440), .Y(new_n3441));
  xnor_4 g01093(.A(new_n3408), .B(n3136), .Y(new_n3442));
  nor_5  g01094(.A(new_n3442), .B(n13263), .Y(new_n3443));
  xnor_4 g01095(.A(new_n3406), .B(n6385), .Y(new_n3444));
  nor_5  g01096(.A(new_n3444), .B(n20455), .Y(new_n3445));
  not_8  g01097(.A(n20455), .Y(new_n3446));
  xnor_4 g01098(.A(new_n3444), .B(new_n3446), .Y(new_n3447));
  not_8  g01099(.A(n1639), .Y(new_n3448));
  xnor_4 g01100(.A(n20138), .B(n9251), .Y(new_n3449));
  and_5  g01101(.A(new_n3449), .B(new_n3448), .Y(new_n3450));
  not_8  g01102(.A(n16968), .Y(new_n3451_1));
  or_5   g01103(.A(new_n3451_1), .B(new_n2367), .Y(new_n3452));
  xnor_4 g01104(.A(new_n3449), .B(n1639), .Y(new_n3453));
  and_5  g01105(.A(new_n3453), .B(new_n3452), .Y(new_n3454));
  or_5   g01106(.A(new_n3454), .B(new_n3450), .Y(new_n3455));
  and_5  g01107(.A(new_n3455), .B(new_n3447), .Y(new_n3456));
  or_5   g01108(.A(new_n3456), .B(new_n3445), .Y(new_n3457));
  not_8  g01109(.A(n13263), .Y(new_n3458));
  xnor_4 g01110(.A(new_n3442), .B(new_n3458), .Y(new_n3459_1));
  and_5  g01111(.A(new_n3459_1), .B(new_n3457), .Y(new_n3460_1));
  or_5   g01112(.A(new_n3460_1), .B(new_n3443), .Y(new_n3461));
  and_5  g01113(.A(new_n3461), .B(new_n3441), .Y(new_n3462));
  or_5   g01114(.A(new_n3462), .B(new_n3439), .Y(new_n3463));
  and_5  g01115(.A(new_n3463), .B(new_n3437), .Y(new_n3464));
  or_5   g01116(.A(new_n3464), .B(new_n3435), .Y(new_n3465));
  and_5  g01117(.A(new_n3465), .B(new_n3433), .Y(new_n3466));
  or_5   g01118(.A(new_n3466), .B(new_n3431), .Y(new_n3467));
  and_5  g01119(.A(new_n3467), .B(new_n3429), .Y(new_n3468_1));
  or_5   g01120(.A(new_n3468_1), .B(new_n3427), .Y(new_n3469));
  and_5  g01121(.A(new_n3469), .B(new_n3425_1), .Y(new_n3470));
  nor_5  g01122(.A(new_n3470), .B(new_n3423), .Y(new_n3471));
  xnor_4 g01123(.A(new_n3471), .B(new_n3421), .Y(new_n3472));
  xnor_4 g01124(.A(new_n3472), .B(n26180), .Y(new_n3473));
  nor_5  g01125(.A(new_n3468_1), .B(new_n3427), .Y(new_n3474));
  xnor_4 g01126(.A(new_n3474), .B(new_n3425_1), .Y(new_n3475));
  not_8  g01127(.A(new_n3475), .Y(new_n3476));
  nor_5  g01128(.A(new_n3476), .B(n24004), .Y(new_n3477));
  xnor_4 g01129(.A(new_n3475), .B(n24004), .Y(new_n3478));
  nor_5  g01130(.A(new_n3466), .B(new_n3431), .Y(new_n3479));
  xnor_4 g01131(.A(new_n3479), .B(new_n3429), .Y(new_n3480_1));
  not_8  g01132(.A(new_n3480_1), .Y(new_n3481));
  nor_5  g01133(.A(new_n3481), .B(n12871), .Y(new_n3482));
  xnor_4 g01134(.A(new_n3480_1), .B(n12871), .Y(new_n3483));
  nor_5  g01135(.A(new_n3464), .B(new_n3435), .Y(new_n3484));
  xnor_4 g01136(.A(new_n3484), .B(new_n3433), .Y(new_n3485));
  not_8  g01137(.A(new_n3485), .Y(new_n3486));
  nor_5  g01138(.A(new_n3486), .B(n23304), .Y(new_n3487));
  xnor_4 g01139(.A(new_n3485), .B(n23304), .Y(new_n3488));
  nor_5  g01140(.A(new_n3462), .B(new_n3439), .Y(new_n3489));
  xnor_4 g01141(.A(new_n3489), .B(new_n3437), .Y(new_n3490));
  not_8  g01142(.A(new_n3490), .Y(new_n3491));
  nor_5  g01143(.A(new_n3491), .B(n19361), .Y(new_n3492));
  xnor_4 g01144(.A(new_n3490), .B(n19361), .Y(new_n3493));
  xor_4  g01145(.A(new_n3461), .B(new_n3441), .Y(new_n3494));
  not_8  g01146(.A(new_n3494), .Y(new_n3495));
  nor_5  g01147(.A(new_n3495), .B(n1437), .Y(new_n3496));
  not_8  g01148(.A(n1437), .Y(new_n3497));
  xnor_4 g01149(.A(new_n3495), .B(new_n3497), .Y(new_n3498));
  nor_5  g01150(.A(new_n3456), .B(new_n3445), .Y(new_n3499));
  xnor_4 g01151(.A(new_n3459_1), .B(new_n3499), .Y(new_n3500));
  not_8  g01152(.A(new_n3500), .Y(new_n3501));
  nor_5  g01153(.A(new_n3501), .B(n4722), .Y(new_n3502_1));
  not_8  g01154(.A(n4722), .Y(new_n3503));
  xnor_4 g01155(.A(new_n3501), .B(new_n3503), .Y(new_n3504));
  not_8  g01156(.A(n14633), .Y(new_n3505));
  nor_5  g01157(.A(new_n3454), .B(new_n3450), .Y(new_n3506_1));
  xnor_4 g01158(.A(new_n3506_1), .B(new_n3447), .Y(new_n3507));
  nor_5  g01159(.A(new_n3507), .B(new_n3505), .Y(new_n3508));
  not_8  g01160(.A(new_n3507), .Y(new_n3509));
  xnor_4 g01161(.A(new_n3509), .B(new_n3505), .Y(new_n3510));
  not_8  g01162(.A(n8721), .Y(new_n3511));
  nor_5  g01163(.A(new_n3451_1), .B(new_n2367), .Y(new_n3512));
  xnor_4 g01164(.A(new_n3453), .B(new_n3512), .Y(new_n3513));
  nor_5  g01165(.A(new_n3513), .B(new_n3511), .Y(new_n3514));
  not_8  g01166(.A(n18578), .Y(new_n3515));
  xnor_4 g01167(.A(n16968), .B(n9251), .Y(new_n3516_1));
  nor_5  g01168(.A(new_n3516_1), .B(new_n3515), .Y(new_n3517));
  xnor_4 g01169(.A(new_n3513), .B(n8721), .Y(new_n3518));
  and_5  g01170(.A(new_n3518), .B(new_n3517), .Y(new_n3519));
  or_5   g01171(.A(new_n3519), .B(new_n3514), .Y(new_n3520));
  and_5  g01172(.A(new_n3520), .B(new_n3510), .Y(new_n3521));
  nor_5  g01173(.A(new_n3521), .B(new_n3508), .Y(new_n3522));
  and_5  g01174(.A(new_n3522), .B(new_n3504), .Y(new_n3523));
  or_5   g01175(.A(new_n3523), .B(new_n3502_1), .Y(new_n3524));
  and_5  g01176(.A(new_n3524), .B(new_n3498), .Y(new_n3525));
  or_5   g01177(.A(new_n3525), .B(new_n3496), .Y(new_n3526));
  and_5  g01178(.A(new_n3526), .B(new_n3493), .Y(new_n3527));
  or_5   g01179(.A(new_n3527), .B(new_n3492), .Y(new_n3528_1));
  and_5  g01180(.A(new_n3528_1), .B(new_n3488), .Y(new_n3529));
  or_5   g01181(.A(new_n3529), .B(new_n3487), .Y(new_n3530));
  and_5  g01182(.A(new_n3530), .B(new_n3483), .Y(new_n3531));
  or_5   g01183(.A(new_n3531), .B(new_n3482), .Y(new_n3532));
  and_5  g01184(.A(new_n3532), .B(new_n3478), .Y(new_n3533));
  nor_5  g01185(.A(new_n3533), .B(new_n3477), .Y(new_n3534));
  xnor_4 g01186(.A(new_n3534), .B(new_n3473), .Y(new_n3535));
  xnor_4 g01187(.A(n3506), .B(n2743), .Y(new_n3536));
  not_8  g01188(.A(n7026), .Y(new_n3537));
  nor_5  g01189(.A(n14899), .B(new_n3537), .Y(new_n3538));
  xnor_4 g01190(.A(n14899), .B(n7026), .Y(new_n3539));
  not_8  g01191(.A(n13719), .Y(new_n3540));
  nor_5  g01192(.A(n18444), .B(new_n3540), .Y(new_n3541_1));
  xnor_4 g01193(.A(n18444), .B(n13719), .Y(new_n3542));
  not_8  g01194(.A(n442), .Y(new_n3543));
  nor_5  g01195(.A(n24638), .B(new_n3543), .Y(new_n3544));
  xnor_4 g01196(.A(n24638), .B(n442), .Y(new_n3545));
  not_8  g01197(.A(n9172), .Y(new_n3546));
  nor_5  g01198(.A(n21674), .B(new_n3546), .Y(new_n3547));
  xnor_4 g01199(.A(n21674), .B(n9172), .Y(new_n3548));
  not_8  g01200(.A(n4913), .Y(new_n3549));
  nor_5  g01201(.A(n17251), .B(new_n3549), .Y(new_n3550));
  xnor_4 g01202(.A(n17251), .B(n4913), .Y(new_n3551));
  not_8  g01203(.A(n604), .Y(new_n3552));
  nor_5  g01204(.A(n14790), .B(new_n3552), .Y(new_n3553));
  xnor_4 g01205(.A(n14790), .B(n604), .Y(new_n3554));
  not_8  g01206(.A(n10096), .Y(new_n3555_1));
  nor_5  g01207(.A(n16824), .B(new_n3555_1), .Y(new_n3556));
  and_5  g01208(.A(n16824), .B(new_n3555_1), .Y(new_n3557));
  not_8  g01209(.A(n16994), .Y(new_n3558));
  nor_5  g01210(.A(new_n3558), .B(n16521), .Y(new_n3559));
  not_8  g01211(.A(n16521), .Y(new_n3560));
  nor_5  g01212(.A(n16994), .B(new_n3560), .Y(new_n3561_1));
  not_8  g01213(.A(n9246), .Y(new_n3562));
  nor_5  g01214(.A(new_n3562), .B(n7139), .Y(new_n3563_1));
  not_8  g01215(.A(new_n3563_1), .Y(new_n3564));
  nor_5  g01216(.A(new_n3564), .B(new_n3561_1), .Y(new_n3565));
  nor_5  g01217(.A(new_n3565), .B(new_n3559), .Y(new_n3566));
  nor_5  g01218(.A(new_n3566), .B(new_n3557), .Y(new_n3567));
  nor_5  g01219(.A(new_n3567), .B(new_n3556), .Y(new_n3568));
  and_5  g01220(.A(new_n3568), .B(new_n3554), .Y(new_n3569));
  or_5   g01221(.A(new_n3569), .B(new_n3553), .Y(new_n3570_1));
  and_5  g01222(.A(new_n3570_1), .B(new_n3551), .Y(new_n3571));
  or_5   g01223(.A(new_n3571), .B(new_n3550), .Y(new_n3572));
  and_5  g01224(.A(new_n3572), .B(new_n3548), .Y(new_n3573));
  or_5   g01225(.A(new_n3573), .B(new_n3547), .Y(new_n3574));
  and_5  g01226(.A(new_n3574), .B(new_n3545), .Y(new_n3575));
  or_5   g01227(.A(new_n3575), .B(new_n3544), .Y(new_n3576));
  and_5  g01228(.A(new_n3576), .B(new_n3542), .Y(new_n3577));
  or_5   g01229(.A(new_n3577), .B(new_n3541_1), .Y(new_n3578));
  and_5  g01230(.A(new_n3578), .B(new_n3539), .Y(new_n3579));
  or_5   g01231(.A(new_n3579), .B(new_n3538), .Y(new_n3580));
  xor_4  g01232(.A(new_n3580), .B(new_n3536), .Y(new_n3581));
  not_8  g01233(.A(new_n3581), .Y(new_n3582_1));
  not_8  g01234(.A(n21489), .Y(new_n3583));
  nor_5  g01235(.A(n25565), .B(n21993), .Y(new_n3584));
  not_8  g01236(.A(new_n3584), .Y(new_n3585));
  nor_5  g01237(.A(new_n3585), .B(n11273), .Y(new_n3586));
  not_8  g01238(.A(new_n3586), .Y(new_n3587));
  nor_5  g01239(.A(new_n3587), .B(n22290), .Y(new_n3588));
  not_8  g01240(.A(new_n3588), .Y(new_n3589));
  nor_5  g01241(.A(new_n3589), .B(n9598), .Y(new_n3590));
  not_8  g01242(.A(new_n3590), .Y(new_n3591));
  nor_5  g01243(.A(new_n3591), .B(n7670), .Y(new_n3592));
  not_8  g01244(.A(new_n3592), .Y(new_n3593));
  nor_5  g01245(.A(new_n3593), .B(n13912), .Y(new_n3594));
  not_8  g01246(.A(new_n3594), .Y(new_n3595));
  nor_5  g01247(.A(new_n3595), .B(n20213), .Y(new_n3596));
  and_5  g01248(.A(new_n3596), .B(new_n3583), .Y(new_n3597));
  xnor_4 g01249(.A(new_n3597), .B(n9259), .Y(new_n3598));
  xnor_4 g01250(.A(new_n3598), .B(new_n3582_1), .Y(new_n3599));
  xor_4  g01251(.A(new_n3578), .B(new_n3539), .Y(new_n3600));
  not_8  g01252(.A(new_n3600), .Y(new_n3601));
  xnor_4 g01253(.A(new_n3596), .B(n21489), .Y(new_n3602));
  not_8  g01254(.A(new_n3602), .Y(new_n3603));
  nor_5  g01255(.A(new_n3603), .B(new_n3601), .Y(new_n3604));
  xnor_4 g01256(.A(new_n3602), .B(new_n3601), .Y(new_n3605));
  nor_5  g01257(.A(new_n3575), .B(new_n3544), .Y(new_n3606));
  xnor_4 g01258(.A(new_n3606), .B(new_n3542), .Y(new_n3607));
  xnor_4 g01259(.A(new_n3594), .B(n20213), .Y(new_n3608));
  nor_5  g01260(.A(new_n3608), .B(new_n3607), .Y(new_n3609));
  not_8  g01261(.A(new_n3607), .Y(new_n3610));
  not_8  g01262(.A(new_n3608), .Y(new_n3611));
  xnor_4 g01263(.A(new_n3611), .B(new_n3610), .Y(new_n3612));
  xor_4  g01264(.A(new_n3574), .B(new_n3545), .Y(new_n3613));
  xnor_4 g01265(.A(new_n3592), .B(n13912), .Y(new_n3614));
  nor_5  g01266(.A(new_n3614), .B(new_n3613), .Y(new_n3615));
  xnor_4 g01267(.A(new_n3614), .B(new_n3613), .Y(new_n3616));
  xor_4  g01268(.A(new_n3572), .B(new_n3548), .Y(new_n3617_1));
  xnor_4 g01269(.A(new_n3590), .B(n7670), .Y(new_n3618_1));
  nor_5  g01270(.A(new_n3618_1), .B(new_n3617_1), .Y(new_n3619));
  xnor_4 g01271(.A(new_n3618_1), .B(new_n3617_1), .Y(new_n3620));
  xnor_4 g01272(.A(new_n3588), .B(n9598), .Y(new_n3621));
  xor_4  g01273(.A(new_n3570_1), .B(new_n3551), .Y(new_n3622));
  nor_5  g01274(.A(new_n3622), .B(new_n3621), .Y(new_n3623));
  xnor_4 g01275(.A(new_n3622), .B(new_n3621), .Y(new_n3624));
  xnor_4 g01276(.A(new_n3586), .B(n22290), .Y(new_n3625));
  not_8  g01277(.A(new_n3625), .Y(new_n3626));
  xnor_4 g01278(.A(new_n3568), .B(new_n3554), .Y(new_n3627));
  and_5  g01279(.A(new_n3627), .B(new_n3626), .Y(new_n3628));
  xnor_4 g01280(.A(new_n3584), .B(n11273), .Y(new_n3629));
  not_8  g01281(.A(new_n3629), .Y(new_n3630));
  xnor_4 g01282(.A(n16824), .B(n10096), .Y(new_n3631));
  xnor_4 g01283(.A(new_n3631), .B(new_n3566), .Y(new_n3632));
  and_5  g01284(.A(new_n3632), .B(new_n3630), .Y(new_n3633));
  xnor_4 g01285(.A(new_n3632), .B(new_n3629), .Y(new_n3634));
  not_8  g01286(.A(n21993), .Y(new_n3635));
  xnor_4 g01287(.A(n25565), .B(new_n3635), .Y(new_n3636));
  xnor_4 g01288(.A(n16994), .B(n16521), .Y(new_n3637));
  xnor_4 g01289(.A(new_n3637), .B(new_n3564), .Y(new_n3638));
  not_8  g01290(.A(new_n3638), .Y(new_n3639));
  nor_5  g01291(.A(new_n3639), .B(new_n3636), .Y(new_n3640));
  xnor_4 g01292(.A(n9246), .B(n7139), .Y(new_n3641));
  nor_5  g01293(.A(new_n3641), .B(new_n3635), .Y(new_n3642_1));
  not_8  g01294(.A(new_n3636), .Y(new_n3643));
  xnor_4 g01295(.A(new_n3638), .B(new_n3643), .Y(new_n3644));
  nor_5  g01296(.A(new_n3644), .B(new_n3642_1), .Y(new_n3645));
  or_5   g01297(.A(new_n3645), .B(new_n3640), .Y(new_n3646));
  and_5  g01298(.A(new_n3646), .B(new_n3634), .Y(new_n3647));
  or_5   g01299(.A(new_n3647), .B(new_n3633), .Y(new_n3648));
  xnor_4 g01300(.A(new_n3627), .B(new_n3625), .Y(new_n3649_1));
  and_5  g01301(.A(new_n3649_1), .B(new_n3648), .Y(new_n3650));
  nor_5  g01302(.A(new_n3650), .B(new_n3628), .Y(new_n3651));
  nor_5  g01303(.A(new_n3651), .B(new_n3624), .Y(new_n3652));
  nor_5  g01304(.A(new_n3652), .B(new_n3623), .Y(new_n3653));
  nor_5  g01305(.A(new_n3653), .B(new_n3620), .Y(new_n3654));
  nor_5  g01306(.A(new_n3654), .B(new_n3619), .Y(new_n3655));
  nor_5  g01307(.A(new_n3655), .B(new_n3616), .Y(new_n3656));
  nor_5  g01308(.A(new_n3656), .B(new_n3615), .Y(new_n3657));
  nor_5  g01309(.A(new_n3657), .B(new_n3612), .Y(new_n3658));
  nor_5  g01310(.A(new_n3658), .B(new_n3609), .Y(new_n3659));
  and_5  g01311(.A(new_n3659), .B(new_n3605), .Y(new_n3660));
  or_5   g01312(.A(new_n3660), .B(new_n3604), .Y(new_n3661));
  xor_4  g01313(.A(new_n3661), .B(new_n3599), .Y(new_n3662));
  xnor_4 g01314(.A(new_n3662), .B(new_n3535), .Y(new_n3663));
  nor_5  g01315(.A(new_n3531), .B(new_n3482), .Y(new_n3664));
  xnor_4 g01316(.A(new_n3664), .B(new_n3478), .Y(new_n3665_1));
  not_8  g01317(.A(new_n3665_1), .Y(new_n3666));
  xor_4  g01318(.A(new_n3659), .B(new_n3605), .Y(new_n3667));
  nor_5  g01319(.A(new_n3667), .B(new_n3666), .Y(new_n3668));
  xnor_4 g01320(.A(new_n3667), .B(new_n3666), .Y(new_n3669));
  xor_4  g01321(.A(new_n3530), .B(new_n3483), .Y(new_n3670));
  not_8  g01322(.A(new_n3670), .Y(new_n3671));
  xnor_4 g01323(.A(new_n3657), .B(new_n3612), .Y(new_n3672));
  nor_5  g01324(.A(new_n3672), .B(new_n3671), .Y(new_n3673));
  xnor_4 g01325(.A(new_n3672), .B(new_n3671), .Y(new_n3674));
  xor_4  g01326(.A(new_n3528_1), .B(new_n3488), .Y(new_n3675));
  not_8  g01327(.A(new_n3675), .Y(new_n3676));
  xnor_4 g01328(.A(new_n3655), .B(new_n3616), .Y(new_n3677));
  nor_5  g01329(.A(new_n3677), .B(new_n3676), .Y(new_n3678));
  xnor_4 g01330(.A(new_n3677), .B(new_n3676), .Y(new_n3679_1));
  xor_4  g01331(.A(new_n3526), .B(new_n3493), .Y(new_n3680));
  not_8  g01332(.A(new_n3680), .Y(new_n3681));
  xnor_4 g01333(.A(new_n3653), .B(new_n3620), .Y(new_n3682));
  nor_5  g01334(.A(new_n3682), .B(new_n3681), .Y(new_n3683));
  xnor_4 g01335(.A(new_n3682), .B(new_n3681), .Y(new_n3684));
  xor_4  g01336(.A(new_n3524), .B(new_n3498), .Y(new_n3685));
  not_8  g01337(.A(new_n3685), .Y(new_n3686));
  xnor_4 g01338(.A(new_n3651), .B(new_n3624), .Y(new_n3687));
  nor_5  g01339(.A(new_n3687), .B(new_n3686), .Y(new_n3688));
  xnor_4 g01340(.A(new_n3687), .B(new_n3686), .Y(new_n3689));
  xnor_4 g01341(.A(new_n3522), .B(new_n3504), .Y(new_n3690));
  not_8  g01342(.A(new_n3690), .Y(new_n3691));
  xor_4  g01343(.A(new_n3649_1), .B(new_n3648), .Y(new_n3692));
  and_5  g01344(.A(new_n3692), .B(new_n3691), .Y(new_n3693));
  xnor_4 g01345(.A(new_n3692), .B(new_n3691), .Y(new_n3694));
  nor_5  g01346(.A(new_n3519), .B(new_n3514), .Y(new_n3695));
  xnor_4 g01347(.A(new_n3695), .B(new_n3510), .Y(new_n3696));
  not_8  g01348(.A(new_n3696), .Y(new_n3697));
  xor_4  g01349(.A(new_n3646), .B(new_n3634), .Y(new_n3698));
  and_5  g01350(.A(new_n3698), .B(new_n3697), .Y(new_n3699));
  xnor_4 g01351(.A(new_n3698), .B(new_n3697), .Y(new_n3700));
  xnor_4 g01352(.A(new_n3644), .B(new_n3642_1), .Y(new_n3701));
  xor_4  g01353(.A(new_n3518), .B(new_n3517), .Y(new_n3702));
  nor_5  g01354(.A(new_n3702), .B(new_n3701), .Y(new_n3703));
  xnor_4 g01355(.A(new_n3516_1), .B(n18578), .Y(new_n3704));
  xnor_4 g01356(.A(new_n3641), .B(n21993), .Y(new_n3705));
  and_5  g01357(.A(new_n3705), .B(new_n3704), .Y(new_n3706));
  xnor_4 g01358(.A(new_n3702), .B(new_n3701), .Y(new_n3707));
  nor_5  g01359(.A(new_n3707), .B(new_n3706), .Y(new_n3708));
  nor_5  g01360(.A(new_n3708), .B(new_n3703), .Y(new_n3709));
  nor_5  g01361(.A(new_n3709), .B(new_n3700), .Y(new_n3710_1));
  nor_5  g01362(.A(new_n3710_1), .B(new_n3699), .Y(new_n3711));
  nor_5  g01363(.A(new_n3711), .B(new_n3694), .Y(new_n3712));
  nor_5  g01364(.A(new_n3712), .B(new_n3693), .Y(new_n3713));
  nor_5  g01365(.A(new_n3713), .B(new_n3689), .Y(new_n3714));
  nor_5  g01366(.A(new_n3714), .B(new_n3688), .Y(new_n3715));
  nor_5  g01367(.A(new_n3715), .B(new_n3684), .Y(new_n3716));
  nor_5  g01368(.A(new_n3716), .B(new_n3683), .Y(new_n3717));
  nor_5  g01369(.A(new_n3717), .B(new_n3679_1), .Y(new_n3718));
  nor_5  g01370(.A(new_n3718), .B(new_n3678), .Y(new_n3719));
  nor_5  g01371(.A(new_n3719), .B(new_n3674), .Y(new_n3720));
  nor_5  g01372(.A(new_n3720), .B(new_n3673), .Y(new_n3721));
  nor_5  g01373(.A(new_n3721), .B(new_n3669), .Y(new_n3722));
  nor_5  g01374(.A(new_n3722), .B(new_n3668), .Y(new_n3723));
  xnor_4 g01375(.A(new_n3723), .B(new_n3663), .Y(n235));
  not_8  g01376(.A(n25749), .Y(new_n3725_1));
  not_8  g01377(.A(n19327), .Y(new_n3726));
  nor_5  g01378(.A(n25435), .B(n13319), .Y(new_n3727));
  not_8  g01379(.A(new_n3727), .Y(new_n3728));
  nor_5  g01380(.A(new_n3728), .B(n15967), .Y(new_n3729));
  not_8  g01381(.A(new_n3729), .Y(new_n3730));
  nor_5  g01382(.A(new_n3730), .B(n25797), .Y(new_n3731));
  not_8  g01383(.A(new_n3731), .Y(new_n3732));
  nor_5  g01384(.A(new_n3732), .B(n6369), .Y(new_n3733_1));
  not_8  g01385(.A(new_n3733_1), .Y(new_n3734));
  nor_5  g01386(.A(new_n3734), .B(n21134), .Y(new_n3735));
  xnor_4 g01387(.A(new_n3735), .B(n2113), .Y(new_n3736));
  xnor_4 g01388(.A(new_n3736), .B(new_n3726), .Y(new_n3737));
  xnor_4 g01389(.A(new_n3733_1), .B(n21134), .Y(new_n3738));
  nor_5  g01390(.A(new_n3738), .B(n22597), .Y(new_n3739));
  not_8  g01391(.A(n22597), .Y(new_n3740_1));
  xnor_4 g01392(.A(new_n3738), .B(new_n3740_1), .Y(new_n3741));
  xnor_4 g01393(.A(new_n3731), .B(n6369), .Y(new_n3742));
  nor_5  g01394(.A(new_n3742), .B(n26107), .Y(new_n3743));
  not_8  g01395(.A(n26107), .Y(new_n3744));
  xnor_4 g01396(.A(new_n3742), .B(new_n3744), .Y(new_n3745));
  xnor_4 g01397(.A(new_n3729), .B(n25797), .Y(new_n3746));
  nor_5  g01398(.A(new_n3746), .B(n342), .Y(new_n3747));
  xnor_4 g01399(.A(new_n3727), .B(n15967), .Y(new_n3748));
  nor_5  g01400(.A(new_n3748), .B(n26553), .Y(new_n3749));
  not_8  g01401(.A(new_n3748), .Y(new_n3750));
  xnor_4 g01402(.A(new_n3750), .B(n26553), .Y(new_n3751));
  not_8  g01403(.A(n13319), .Y(new_n3752));
  xnor_4 g01404(.A(n25435), .B(new_n3752), .Y(new_n3753));
  nor_5  g01405(.A(new_n3753), .B(n4964), .Y(new_n3754));
  not_8  g01406(.A(n7876), .Y(new_n3755_1));
  not_8  g01407(.A(n25435), .Y(new_n3756));
  or_5   g01408(.A(new_n3756), .B(new_n3755_1), .Y(new_n3757));
  not_8  g01409(.A(new_n3753), .Y(new_n3758_1));
  xnor_4 g01410(.A(new_n3758_1), .B(n4964), .Y(new_n3759));
  and_5  g01411(.A(new_n3759), .B(new_n3757), .Y(new_n3760_1));
  or_5   g01412(.A(new_n3760_1), .B(new_n3754), .Y(new_n3761));
  and_5  g01413(.A(new_n3761), .B(new_n3751), .Y(new_n3762));
  or_5   g01414(.A(new_n3762), .B(new_n3749), .Y(new_n3763));
  xor_4  g01415(.A(new_n3746), .B(n342), .Y(new_n3764));
  and_5  g01416(.A(new_n3764), .B(new_n3763), .Y(new_n3765));
  or_5   g01417(.A(new_n3765), .B(new_n3747), .Y(new_n3766));
  and_5  g01418(.A(new_n3766), .B(new_n3745), .Y(new_n3767));
  or_5   g01419(.A(new_n3767), .B(new_n3743), .Y(new_n3768));
  and_5  g01420(.A(new_n3768), .B(new_n3741), .Y(new_n3769));
  nor_5  g01421(.A(new_n3769), .B(new_n3739), .Y(new_n3770));
  xnor_4 g01422(.A(new_n3770), .B(new_n3737), .Y(new_n3771));
  not_8  g01423(.A(new_n3771), .Y(new_n3772));
  xnor_4 g01424(.A(new_n3772), .B(new_n3725_1), .Y(new_n3773));
  not_8  g01425(.A(n3161), .Y(new_n3774));
  xor_4  g01426(.A(new_n3768), .B(new_n3741), .Y(new_n3775));
  nor_5  g01427(.A(new_n3775), .B(new_n3774), .Y(new_n3776));
  xnor_4 g01428(.A(new_n3775), .B(n3161), .Y(new_n3777));
  not_8  g01429(.A(n9003), .Y(new_n3778));
  nor_5  g01430(.A(new_n3765), .B(new_n3747), .Y(new_n3779));
  xnor_4 g01431(.A(new_n3779), .B(new_n3745), .Y(new_n3780));
  nor_5  g01432(.A(new_n3780), .B(new_n3778), .Y(new_n3781_1));
  not_8  g01433(.A(new_n3780), .Y(new_n3782));
  xnor_4 g01434(.A(new_n3782), .B(new_n3778), .Y(new_n3783));
  not_8  g01435(.A(n4957), .Y(new_n3784));
  xor_4  g01436(.A(new_n3764), .B(new_n3763), .Y(new_n3785_1));
  nor_5  g01437(.A(new_n3785_1), .B(new_n3784), .Y(new_n3786));
  xnor_4 g01438(.A(new_n3785_1), .B(n4957), .Y(new_n3787));
  not_8  g01439(.A(n7524), .Y(new_n3788));
  nor_5  g01440(.A(new_n3760_1), .B(new_n3754), .Y(new_n3789));
  xnor_4 g01441(.A(new_n3789), .B(new_n3751), .Y(new_n3790));
  nor_5  g01442(.A(new_n3790), .B(new_n3788), .Y(new_n3791));
  not_8  g01443(.A(new_n3790), .Y(new_n3792));
  xnor_4 g01444(.A(new_n3792), .B(new_n3788), .Y(new_n3793));
  not_8  g01445(.A(n15743), .Y(new_n3794_1));
  nor_5  g01446(.A(new_n3756), .B(new_n3755_1), .Y(new_n3795_1));
  xnor_4 g01447(.A(new_n3759), .B(new_n3795_1), .Y(new_n3796));
  nor_5  g01448(.A(new_n3796), .B(new_n3794_1), .Y(new_n3797));
  not_8  g01449(.A(n20658), .Y(new_n3798));
  xnor_4 g01450(.A(n25435), .B(new_n3755_1), .Y(new_n3799));
  not_8  g01451(.A(new_n3799), .Y(new_n3800));
  nor_5  g01452(.A(new_n3800), .B(new_n3798), .Y(new_n3801));
  xnor_4 g01453(.A(new_n3796), .B(n15743), .Y(new_n3802));
  and_5  g01454(.A(new_n3802), .B(new_n3801), .Y(new_n3803));
  or_5   g01455(.A(new_n3803), .B(new_n3797), .Y(new_n3804));
  and_5  g01456(.A(new_n3804), .B(new_n3793), .Y(new_n3805));
  or_5   g01457(.A(new_n3805), .B(new_n3791), .Y(new_n3806));
  and_5  g01458(.A(new_n3806), .B(new_n3787), .Y(new_n3807));
  or_5   g01459(.A(new_n3807), .B(new_n3786), .Y(new_n3808));
  and_5  g01460(.A(new_n3808), .B(new_n3783), .Y(new_n3809));
  or_5   g01461(.A(new_n3809), .B(new_n3781_1), .Y(new_n3810));
  and_5  g01462(.A(new_n3810), .B(new_n3777), .Y(new_n3811));
  or_5   g01463(.A(new_n3811), .B(new_n3776), .Y(new_n3812));
  xor_4  g01464(.A(new_n3812), .B(new_n3773), .Y(new_n3813));
  xnor_4 g01465(.A(n26510), .B(n22332), .Y(new_n3814));
  not_8  g01466(.A(n23068), .Y(new_n3815));
  and_5  g01467(.A(new_n3815), .B(n18907), .Y(new_n3816));
  xnor_4 g01468(.A(n23068), .B(n18907), .Y(new_n3817));
  nor_5  g01469(.A(n19514), .B(new_n2408), .Y(new_n3818));
  xnor_4 g01470(.A(n19514), .B(n2731), .Y(new_n3819));
  and_5  g01471(.A(n19911), .B(new_n2944_1), .Y(new_n3820));
  xnor_4 g01472(.A(n19911), .B(n10053), .Y(new_n3821));
  nor_5  g01473(.A(n13708), .B(new_n2947), .Y(new_n3822));
  nor_5  g01474(.A(new_n2389), .B(n8399), .Y(new_n3823));
  not_8  g01475(.A(n9507), .Y(new_n3824));
  nor_5  g01476(.A(n18409), .B(new_n3824), .Y(new_n3825));
  not_8  g01477(.A(n18409), .Y(new_n3826));
  nor_5  g01478(.A(new_n3826), .B(n9507), .Y(new_n3827));
  nor_5  g01479(.A(new_n2952), .B(n5704), .Y(new_n3828_1));
  not_8  g01480(.A(new_n3828_1), .Y(new_n3829));
  nor_5  g01481(.A(new_n3829), .B(new_n3827), .Y(new_n3830));
  nor_5  g01482(.A(new_n3830), .B(new_n3825), .Y(new_n3831));
  nor_5  g01483(.A(new_n3831), .B(new_n3823), .Y(new_n3832));
  nor_5  g01484(.A(new_n3832), .B(new_n3822), .Y(new_n3833));
  and_5  g01485(.A(new_n3833), .B(new_n3821), .Y(new_n3834));
  or_5   g01486(.A(new_n3834), .B(new_n3820), .Y(new_n3835));
  and_5  g01487(.A(new_n3835), .B(new_n3819), .Y(new_n3836));
  or_5   g01488(.A(new_n3836), .B(new_n3818), .Y(new_n3837));
  and_5  g01489(.A(new_n3837), .B(new_n3817), .Y(new_n3838));
  or_5   g01490(.A(new_n3838), .B(new_n3816), .Y(new_n3839));
  xor_4  g01491(.A(new_n3839), .B(new_n3814), .Y(new_n3840));
  nor_5  g01492(.A(n22043), .B(n12121), .Y(new_n3841));
  not_8  g01493(.A(new_n3841), .Y(new_n3842_1));
  nor_5  g01494(.A(new_n3842_1), .B(n19618), .Y(new_n3843));
  not_8  g01495(.A(new_n3843), .Y(new_n3844));
  nor_5  g01496(.A(new_n3844), .B(n1204), .Y(new_n3845));
  not_8  g01497(.A(new_n3845), .Y(new_n3846));
  nor_5  g01498(.A(new_n3846), .B(n626), .Y(new_n3847));
  not_8  g01499(.A(new_n3847), .Y(new_n3848));
  nor_5  g01500(.A(new_n3848), .B(n5337), .Y(new_n3849));
  xnor_4 g01501(.A(new_n3849), .B(n4325), .Y(new_n3850_1));
  xnor_4 g01502(.A(new_n3850_1), .B(new_n3840), .Y(new_n3851));
  xor_4  g01503(.A(new_n3837), .B(new_n3817), .Y(new_n3852));
  xnor_4 g01504(.A(new_n3847), .B(n5337), .Y(new_n3853));
  nor_5  g01505(.A(new_n3853), .B(new_n3852), .Y(new_n3854));
  xnor_4 g01506(.A(new_n3853), .B(new_n3852), .Y(new_n3855));
  xor_4  g01507(.A(new_n3835), .B(new_n3819), .Y(new_n3856));
  xnor_4 g01508(.A(new_n3845), .B(n626), .Y(new_n3857));
  nor_5  g01509(.A(new_n3857), .B(new_n3856), .Y(new_n3858));
  xnor_4 g01510(.A(new_n3857), .B(new_n3856), .Y(new_n3859));
  xnor_4 g01511(.A(new_n3843), .B(n1204), .Y(new_n3860));
  xnor_4 g01512(.A(new_n3833), .B(new_n3821), .Y(new_n3861));
  not_8  g01513(.A(new_n3861), .Y(new_n3862));
  nor_5  g01514(.A(new_n3862), .B(new_n3860), .Y(new_n3863));
  xnor_4 g01515(.A(new_n3861), .B(new_n3860), .Y(new_n3864));
  xnor_4 g01516(.A(new_n3841), .B(n19618), .Y(new_n3865));
  xnor_4 g01517(.A(n13708), .B(n8399), .Y(new_n3866));
  xnor_4 g01518(.A(new_n3866), .B(new_n3831), .Y(new_n3867));
  not_8  g01519(.A(new_n3867), .Y(new_n3868));
  nor_5  g01520(.A(new_n3868), .B(new_n3865), .Y(new_n3869_1));
  xnor_4 g01521(.A(new_n3867), .B(new_n3865), .Y(new_n3870));
  xnor_4 g01522(.A(n22043), .B(n12121), .Y(new_n3871_1));
  xnor_4 g01523(.A(n18409), .B(n9507), .Y(new_n3872));
  xnor_4 g01524(.A(new_n3872), .B(new_n3829), .Y(new_n3873));
  nor_5  g01525(.A(new_n3873), .B(new_n3871_1), .Y(new_n3874));
  not_8  g01526(.A(n12121), .Y(new_n3875));
  xnor_4 g01527(.A(n26979), .B(n5704), .Y(new_n3876));
  nor_5  g01528(.A(new_n3876), .B(new_n3875), .Y(new_n3877));
  xor_4  g01529(.A(new_n3873), .B(new_n3871_1), .Y(new_n3878));
  and_5  g01530(.A(new_n3878), .B(new_n3877), .Y(new_n3879));
  nor_5  g01531(.A(new_n3879), .B(new_n3874), .Y(new_n3880));
  and_5  g01532(.A(new_n3880), .B(new_n3870), .Y(new_n3881));
  or_5   g01533(.A(new_n3881), .B(new_n3869_1), .Y(new_n3882));
  and_5  g01534(.A(new_n3882), .B(new_n3864), .Y(new_n3883));
  nor_5  g01535(.A(new_n3883), .B(new_n3863), .Y(new_n3884));
  nor_5  g01536(.A(new_n3884), .B(new_n3859), .Y(new_n3885));
  nor_5  g01537(.A(new_n3885), .B(new_n3858), .Y(new_n3886));
  nor_5  g01538(.A(new_n3886), .B(new_n3855), .Y(new_n3887));
  nor_5  g01539(.A(new_n3887), .B(new_n3854), .Y(new_n3888));
  xnor_4 g01540(.A(new_n3888), .B(new_n3851), .Y(new_n3889));
  xnor_4 g01541(.A(new_n3889), .B(new_n3813), .Y(new_n3890));
  xnor_4 g01542(.A(new_n3886), .B(new_n3855), .Y(new_n3891_1));
  xor_4  g01543(.A(new_n3810), .B(new_n3777), .Y(new_n3892));
  nor_5  g01544(.A(new_n3892), .B(new_n3891_1), .Y(new_n3893));
  xnor_4 g01545(.A(new_n3892), .B(new_n3891_1), .Y(new_n3894));
  xnor_4 g01546(.A(new_n3884), .B(new_n3859), .Y(new_n3895));
  xor_4  g01547(.A(new_n3808), .B(new_n3783), .Y(new_n3896));
  nor_5  g01548(.A(new_n3896), .B(new_n3895), .Y(new_n3897));
  xnor_4 g01549(.A(new_n3896), .B(new_n3895), .Y(new_n3898));
  xor_4  g01550(.A(new_n3882), .B(new_n3864), .Y(new_n3899));
  not_8  g01551(.A(new_n3899), .Y(new_n3900));
  xor_4  g01552(.A(new_n3806), .B(new_n3787), .Y(new_n3901));
  nor_5  g01553(.A(new_n3901), .B(new_n3900), .Y(new_n3902));
  xnor_4 g01554(.A(new_n3901), .B(new_n3900), .Y(new_n3903));
  xnor_4 g01555(.A(new_n3880), .B(new_n3870), .Y(new_n3904));
  xor_4  g01556(.A(new_n3804), .B(new_n3793), .Y(new_n3905));
  nor_5  g01557(.A(new_n3905), .B(new_n3904), .Y(new_n3906));
  xnor_4 g01558(.A(new_n3905), .B(new_n3904), .Y(new_n3907));
  xnor_4 g01559(.A(new_n3878), .B(new_n3877), .Y(new_n3908));
  not_8  g01560(.A(new_n3908), .Y(new_n3909_1));
  xor_4  g01561(.A(new_n3802), .B(new_n3801), .Y(new_n3910));
  nor_5  g01562(.A(new_n3910), .B(new_n3909_1), .Y(new_n3911));
  xnor_4 g01563(.A(new_n3800), .B(new_n3798), .Y(new_n3912));
  xnor_4 g01564(.A(new_n3876), .B(n12121), .Y(new_n3913));
  not_8  g01565(.A(new_n3913), .Y(new_n3914));
  nor_5  g01566(.A(new_n3914), .B(new_n3912), .Y(new_n3915));
  xnor_4 g01567(.A(new_n3910), .B(new_n3909_1), .Y(new_n3916));
  nor_5  g01568(.A(new_n3916), .B(new_n3915), .Y(new_n3917));
  nor_5  g01569(.A(new_n3917), .B(new_n3911), .Y(new_n3918_1));
  nor_5  g01570(.A(new_n3918_1), .B(new_n3907), .Y(new_n3919));
  nor_5  g01571(.A(new_n3919), .B(new_n3906), .Y(new_n3920));
  nor_5  g01572(.A(new_n3920), .B(new_n3903), .Y(new_n3921));
  nor_5  g01573(.A(new_n3921), .B(new_n3902), .Y(new_n3922));
  nor_5  g01574(.A(new_n3922), .B(new_n3898), .Y(new_n3923));
  nor_5  g01575(.A(new_n3923), .B(new_n3897), .Y(new_n3924));
  nor_5  g01576(.A(new_n3924), .B(new_n3894), .Y(new_n3925_1));
  nor_5  g01577(.A(new_n3925_1), .B(new_n3893), .Y(new_n3926));
  xnor_4 g01578(.A(new_n3926), .B(new_n3890), .Y(n242));
  nor_5  g01579(.A(n21398), .B(n11667), .Y(new_n3928));
  not_8  g01580(.A(new_n3928), .Y(new_n3929));
  nor_5  g01581(.A(new_n3929), .B(n26572), .Y(new_n3930));
  not_8  g01582(.A(new_n3930), .Y(new_n3931));
  nor_5  g01583(.A(new_n3931), .B(n5115), .Y(new_n3932_1));
  not_8  g01584(.A(new_n3932_1), .Y(new_n3933));
  nor_5  g01585(.A(new_n3933), .B(n11223), .Y(new_n3934_1));
  xnor_4 g01586(.A(new_n3934_1), .B(n19477), .Y(new_n3935));
  xnor_4 g01587(.A(new_n3935), .B(n11011), .Y(new_n3936));
  xnor_4 g01588(.A(new_n3932_1), .B(n11223), .Y(new_n3937));
  nor_5  g01589(.A(new_n3937), .B(n16029), .Y(new_n3938));
  not_8  g01590(.A(n16029), .Y(new_n3939));
  xnor_4 g01591(.A(new_n3937), .B(new_n3939), .Y(new_n3940));
  xnor_4 g01592(.A(new_n3930), .B(n5115), .Y(new_n3941));
  and_5  g01593(.A(new_n3941), .B(n16476), .Y(new_n3942));
  not_8  g01594(.A(n16476), .Y(new_n3943));
  xnor_4 g01595(.A(new_n3941), .B(new_n3943), .Y(new_n3944));
  xnor_4 g01596(.A(new_n3928), .B(n26572), .Y(new_n3945_1));
  nor_5  g01597(.A(new_n3945_1), .B(n11615), .Y(new_n3946));
  not_8  g01598(.A(n11615), .Y(new_n3947));
  xnor_4 g01599(.A(new_n3945_1), .B(new_n3947), .Y(new_n3948));
  not_8  g01600(.A(n22433), .Y(new_n3949));
  xnor_4 g01601(.A(n21398), .B(n11667), .Y(new_n3950));
  and_5  g01602(.A(new_n3950), .B(new_n3949), .Y(new_n3951));
  not_8  g01603(.A(n14090), .Y(new_n3952_1));
  or_5   g01604(.A(new_n2583), .B(new_n3952_1), .Y(new_n3953));
  xnor_4 g01605(.A(new_n3950), .B(n22433), .Y(new_n3954));
  and_5  g01606(.A(new_n3954), .B(new_n3953), .Y(new_n3955));
  or_5   g01607(.A(new_n3955), .B(new_n3951), .Y(new_n3956));
  and_5  g01608(.A(new_n3956), .B(new_n3948), .Y(new_n3957));
  nor_5  g01609(.A(new_n3957), .B(new_n3946), .Y(new_n3958));
  and_5  g01610(.A(new_n3958), .B(new_n3944), .Y(new_n3959_1));
  nor_5  g01611(.A(new_n3959_1), .B(new_n3942), .Y(new_n3960));
  and_5  g01612(.A(new_n3960), .B(new_n3940), .Y(new_n3961));
  nor_5  g01613(.A(new_n3961), .B(new_n3938), .Y(new_n3962_1));
  xnor_4 g01614(.A(new_n3962_1), .B(new_n3936), .Y(new_n3963));
  xnor_4 g01615(.A(new_n3963), .B(n13677), .Y(new_n3964));
  xnor_4 g01616(.A(new_n3960), .B(new_n3940), .Y(new_n3965));
  nor_5  g01617(.A(new_n3965), .B(n18926), .Y(new_n3966));
  not_8  g01618(.A(n5451), .Y(new_n3967));
  xnor_4 g01619(.A(new_n3958), .B(new_n3944), .Y(new_n3968));
  nor_5  g01620(.A(new_n3968), .B(new_n3967), .Y(new_n3969));
  not_8  g01621(.A(new_n3968), .Y(new_n3970));
  xnor_4 g01622(.A(new_n3970), .B(new_n3967), .Y(new_n3971_1));
  not_8  g01623(.A(n5330), .Y(new_n3972));
  nor_5  g01624(.A(new_n3955), .B(new_n3951), .Y(new_n3973));
  xnor_4 g01625(.A(new_n3973), .B(new_n3948), .Y(new_n3974));
  nor_5  g01626(.A(new_n3974), .B(new_n3972), .Y(new_n3975));
  not_8  g01627(.A(new_n3974), .Y(new_n3976));
  xnor_4 g01628(.A(new_n3976), .B(new_n3972), .Y(new_n3977));
  not_8  g01629(.A(n7657), .Y(new_n3978));
  nor_5  g01630(.A(new_n2583), .B(new_n3952_1), .Y(new_n3979));
  xnor_4 g01631(.A(new_n3954), .B(new_n3979), .Y(new_n3980));
  nor_5  g01632(.A(new_n3980), .B(new_n3978), .Y(new_n3981));
  not_8  g01633(.A(n25926), .Y(new_n3982));
  nor_5  g01634(.A(new_n2551), .B(new_n3982), .Y(new_n3983_1));
  not_8  g01635(.A(new_n3980), .Y(new_n3984_1));
  xnor_4 g01636(.A(new_n3984_1), .B(new_n3978), .Y(new_n3985));
  and_5  g01637(.A(new_n3985), .B(new_n3983_1), .Y(new_n3986));
  or_5   g01638(.A(new_n3986), .B(new_n3981), .Y(new_n3987));
  and_5  g01639(.A(new_n3987), .B(new_n3977), .Y(new_n3988));
  or_5   g01640(.A(new_n3988), .B(new_n3975), .Y(new_n3989));
  and_5  g01641(.A(new_n3989), .B(new_n3971_1), .Y(new_n3990));
  nor_5  g01642(.A(new_n3990), .B(new_n3969), .Y(new_n3991));
  not_8  g01643(.A(new_n3991), .Y(new_n3992));
  xnor_4 g01644(.A(new_n3965), .B(n18926), .Y(new_n3993));
  nor_5  g01645(.A(new_n3993), .B(new_n3992), .Y(new_n3994));
  nor_5  g01646(.A(new_n3994), .B(new_n3966), .Y(new_n3995));
  xnor_4 g01647(.A(new_n3995), .B(new_n3964), .Y(new_n3996));
  nor_5  g01648(.A(n21687), .B(n6729), .Y(new_n3997));
  not_8  g01649(.A(new_n3997), .Y(new_n3998));
  nor_5  g01650(.A(new_n3998), .B(n8285), .Y(new_n3999));
  not_8  g01651(.A(new_n3999), .Y(new_n4000_1));
  nor_5  g01652(.A(new_n4000_1), .B(n20169), .Y(new_n4001));
  not_8  g01653(.A(new_n4001), .Y(new_n4002));
  nor_5  g01654(.A(new_n4002), .B(n19789), .Y(new_n4003));
  xnor_4 g01655(.A(new_n4003), .B(n12398), .Y(new_n4004));
  nor_5  g01656(.A(n19922), .B(n10792), .Y(new_n4005));
  not_8  g01657(.A(new_n4005), .Y(new_n4006));
  nor_5  g01658(.A(new_n4006), .B(n9323), .Y(new_n4007));
  not_8  g01659(.A(new_n4007), .Y(new_n4008));
  nor_5  g01660(.A(new_n4008), .B(n1949), .Y(new_n4009));
  not_8  g01661(.A(new_n4009), .Y(new_n4010_1));
  nor_5  g01662(.A(new_n4010_1), .B(n15424), .Y(new_n4011));
  xnor_4 g01663(.A(new_n4011), .B(n25694), .Y(new_n4012));
  not_8  g01664(.A(new_n4012), .Y(new_n4013));
  xnor_4 g01665(.A(new_n4013), .B(n20151), .Y(new_n4014_1));
  not_8  g01666(.A(n7693), .Y(new_n4015));
  xnor_4 g01667(.A(new_n4009), .B(n15424), .Y(new_n4016));
  not_8  g01668(.A(new_n4016), .Y(new_n4017));
  nor_5  g01669(.A(new_n4017), .B(new_n4015), .Y(new_n4018));
  xnor_4 g01670(.A(new_n4007), .B(n1949), .Y(new_n4019));
  and_5  g01671(.A(new_n4019), .B(n10405), .Y(new_n4020));
  not_8  g01672(.A(n10405), .Y(new_n4021));
  xnor_4 g01673(.A(new_n4019), .B(new_n4021), .Y(new_n4022));
  xnor_4 g01674(.A(new_n4005), .B(n9323), .Y(new_n4023));
  nor_5  g01675(.A(new_n4023), .B(n11302), .Y(new_n4024));
  not_8  g01676(.A(new_n4023), .Y(new_n4025));
  xnor_4 g01677(.A(new_n4025), .B(n11302), .Y(new_n4026));
  xnor_4 g01678(.A(n19922), .B(n10792), .Y(new_n4027));
  not_8  g01679(.A(new_n4027), .Y(new_n4028));
  nor_5  g01680(.A(new_n4028), .B(n17090), .Y(new_n4029));
  not_8  g01681(.A(n6773), .Y(new_n4030));
  not_8  g01682(.A(n19922), .Y(new_n4031));
  or_5   g01683(.A(new_n4031), .B(new_n4030), .Y(new_n4032));
  xnor_4 g01684(.A(new_n4027), .B(n17090), .Y(new_n4033));
  and_5  g01685(.A(new_n4033), .B(new_n4032), .Y(new_n4034));
  or_5   g01686(.A(new_n4034), .B(new_n4029), .Y(new_n4035));
  and_5  g01687(.A(new_n4035), .B(new_n4026), .Y(new_n4036));
  nor_5  g01688(.A(new_n4036), .B(new_n4024), .Y(new_n4037));
  and_5  g01689(.A(new_n4037), .B(new_n4022), .Y(new_n4038));
  or_5   g01690(.A(new_n4038), .B(new_n4020), .Y(new_n4039));
  xnor_4 g01691(.A(new_n4017), .B(n7693), .Y(new_n4040));
  and_5  g01692(.A(new_n4040), .B(new_n4039), .Y(new_n4041));
  nor_5  g01693(.A(new_n4041), .B(new_n4018), .Y(new_n4042));
  xnor_4 g01694(.A(new_n4042), .B(new_n4014_1), .Y(new_n4043));
  not_8  g01695(.A(new_n4043), .Y(new_n4044));
  xnor_4 g01696(.A(new_n4044), .B(new_n4004), .Y(new_n4045));
  xnor_4 g01697(.A(new_n4001), .B(n19789), .Y(new_n4046));
  xor_4  g01698(.A(new_n4040), .B(new_n4039), .Y(new_n4047));
  and_5  g01699(.A(new_n4047), .B(new_n4046), .Y(new_n4048));
  not_8  g01700(.A(new_n4047), .Y(new_n4049));
  xnor_4 g01701(.A(new_n4049), .B(new_n4046), .Y(new_n4050));
  xnor_4 g01702(.A(new_n4037), .B(new_n4022), .Y(new_n4051));
  not_8  g01703(.A(new_n4051), .Y(new_n4052));
  xnor_4 g01704(.A(new_n3999), .B(n20169), .Y(new_n4053));
  nor_5  g01705(.A(new_n4053), .B(new_n4052), .Y(new_n4054));
  xnor_4 g01706(.A(new_n4053), .B(new_n4051), .Y(new_n4055));
  nor_5  g01707(.A(new_n4034), .B(new_n4029), .Y(new_n4056));
  xnor_4 g01708(.A(new_n4056), .B(new_n4026), .Y(new_n4057));
  not_8  g01709(.A(new_n4057), .Y(new_n4058));
  xnor_4 g01710(.A(new_n3997), .B(n8285), .Y(new_n4059));
  and_5  g01711(.A(new_n4059), .B(new_n4058), .Y(new_n4060));
  xnor_4 g01712(.A(new_n4059), .B(new_n4057), .Y(new_n4061));
  xnor_4 g01713(.A(n21687), .B(n6729), .Y(new_n4062));
  nor_5  g01714(.A(new_n4031), .B(new_n4030), .Y(new_n4063));
  xnor_4 g01715(.A(new_n4033), .B(new_n4063), .Y(new_n4064));
  nor_5  g01716(.A(new_n4064), .B(new_n4062), .Y(new_n4065));
  nor_5  g01717(.A(new_n2549), .B(new_n2548), .Y(new_n4066));
  not_8  g01718(.A(new_n4064), .Y(new_n4067));
  xnor_4 g01719(.A(new_n4067), .B(new_n4062), .Y(new_n4068));
  and_5  g01720(.A(new_n4068), .B(new_n4066), .Y(new_n4069));
  or_5   g01721(.A(new_n4069), .B(new_n4065), .Y(new_n4070));
  and_5  g01722(.A(new_n4070), .B(new_n4061), .Y(new_n4071_1));
  nor_5  g01723(.A(new_n4071_1), .B(new_n4060), .Y(new_n4072));
  and_5  g01724(.A(new_n4072), .B(new_n4055), .Y(new_n4073));
  nor_5  g01725(.A(new_n4073), .B(new_n4054), .Y(new_n4074));
  and_5  g01726(.A(new_n4074), .B(new_n4050), .Y(new_n4075));
  or_5   g01727(.A(new_n4075), .B(new_n4048), .Y(new_n4076));
  xor_4  g01728(.A(new_n4076), .B(new_n4045), .Y(new_n4077));
  xnor_4 g01729(.A(new_n4077), .B(new_n3996), .Y(new_n4078));
  xnor_4 g01730(.A(new_n4074), .B(new_n4050), .Y(new_n4079));
  xnor_4 g01731(.A(new_n3993), .B(new_n3991), .Y(new_n4080));
  and_5  g01732(.A(new_n4080), .B(new_n4079), .Y(new_n4081));
  xnor_4 g01733(.A(new_n4080), .B(new_n4079), .Y(new_n4082));
  xnor_4 g01734(.A(new_n4072), .B(new_n4055), .Y(new_n4083));
  xor_4  g01735(.A(new_n3989), .B(new_n3971_1), .Y(new_n4084));
  nor_5  g01736(.A(new_n4084), .B(new_n4083), .Y(new_n4085_1));
  xnor_4 g01737(.A(new_n4084), .B(new_n4083), .Y(new_n4086));
  xor_4  g01738(.A(new_n3987), .B(new_n3977), .Y(new_n4087));
  xor_4  g01739(.A(new_n4070), .B(new_n4061), .Y(new_n4088_1));
  nor_5  g01740(.A(new_n4088_1), .B(new_n4087), .Y(new_n4089_1));
  xnor_4 g01741(.A(new_n4088_1), .B(new_n4087), .Y(new_n4090));
  xor_4  g01742(.A(new_n4068), .B(new_n4066), .Y(new_n4091));
  xor_4  g01743(.A(new_n3985), .B(new_n3983_1), .Y(new_n4092));
  nor_5  g01744(.A(new_n4092), .B(new_n4091), .Y(new_n4093));
  not_8  g01745(.A(new_n2552), .Y(new_n4094));
  nor_5  g01746(.A(new_n4094), .B(new_n2550), .Y(new_n4095));
  xnor_4 g01747(.A(new_n4092), .B(new_n4091), .Y(new_n4096));
  nor_5  g01748(.A(new_n4096), .B(new_n4095), .Y(new_n4097));
  nor_5  g01749(.A(new_n4097), .B(new_n4093), .Y(new_n4098));
  nor_5  g01750(.A(new_n4098), .B(new_n4090), .Y(new_n4099));
  nor_5  g01751(.A(new_n4099), .B(new_n4089_1), .Y(new_n4100_1));
  nor_5  g01752(.A(new_n4100_1), .B(new_n4086), .Y(new_n4101));
  nor_5  g01753(.A(new_n4101), .B(new_n4085_1), .Y(new_n4102));
  nor_5  g01754(.A(new_n4102), .B(new_n4082), .Y(new_n4103_1));
  nor_5  g01755(.A(new_n4103_1), .B(new_n4081), .Y(new_n4104));
  xnor_4 g01756(.A(new_n4104), .B(new_n4078), .Y(n243));
  not_8  g01757(.A(n11302), .Y(new_n4106));
  xnor_4 g01758(.A(n24786), .B(new_n4106), .Y(new_n4107));
  nor_5  g01759(.A(n27120), .B(n17090), .Y(new_n4108));
  not_8  g01760(.A(n23065), .Y(new_n4109));
  or_5   g01761(.A(new_n4109), .B(new_n4030), .Y(new_n4110));
  not_8  g01762(.A(n17090), .Y(new_n4111));
  xnor_4 g01763(.A(n27120), .B(new_n4111), .Y(new_n4112));
  and_5  g01764(.A(new_n4112), .B(new_n4110), .Y(new_n4113));
  nor_5  g01765(.A(new_n4113), .B(new_n4108), .Y(new_n4114));
  xnor_4 g01766(.A(new_n4114), .B(new_n4107), .Y(new_n4115));
  not_8  g01767(.A(new_n4115), .Y(new_n4116));
  xnor_4 g01768(.A(n20036), .B(n1689), .Y(new_n4117));
  not_8  g01769(.A(n22274), .Y(new_n4118));
  nor_5  g01770(.A(new_n4118), .B(n11192), .Y(new_n4119_1));
  not_8  g01771(.A(n11192), .Y(new_n4120));
  nor_5  g01772(.A(n22274), .B(new_n4120), .Y(new_n4121));
  not_8  g01773(.A(n24129), .Y(new_n4122));
  nor_5  g01774(.A(new_n4122), .B(n9380), .Y(new_n4123_1));
  not_8  g01775(.A(new_n4123_1), .Y(new_n4124));
  nor_5  g01776(.A(new_n4124), .B(new_n4121), .Y(new_n4125));
  nor_5  g01777(.A(new_n4125), .B(new_n4119_1), .Y(new_n4126));
  xnor_4 g01778(.A(new_n4126), .B(new_n4117), .Y(new_n4127));
  xnor_4 g01779(.A(new_n4127), .B(new_n4116), .Y(new_n4128));
  nor_5  g01780(.A(new_n4109), .B(new_n4030), .Y(new_n4129));
  xnor_4 g01781(.A(new_n4112), .B(new_n4129), .Y(new_n4130));
  xnor_4 g01782(.A(n22274), .B(n11192), .Y(new_n4131));
  xnor_4 g01783(.A(new_n4131), .B(new_n4124), .Y(new_n4132));
  nor_5  g01784(.A(new_n4132), .B(new_n4130), .Y(new_n4133));
  xnor_4 g01785(.A(n23065), .B(new_n4030), .Y(new_n4134_1));
  not_8  g01786(.A(new_n4134_1), .Y(new_n4135));
  xnor_4 g01787(.A(n24129), .B(n9380), .Y(new_n4136));
  nor_5  g01788(.A(new_n4136), .B(new_n4135), .Y(new_n4137));
  not_8  g01789(.A(new_n4130), .Y(new_n4138));
  xnor_4 g01790(.A(new_n4132), .B(new_n4138), .Y(new_n4139));
  and_5  g01791(.A(new_n4139), .B(new_n4137), .Y(new_n4140));
  nor_5  g01792(.A(new_n4140), .B(new_n4133), .Y(new_n4141));
  xnor_4 g01793(.A(new_n4141), .B(new_n4128), .Y(new_n4142));
  not_8  g01794(.A(n919), .Y(new_n4143));
  xnor_4 g01795(.A(n5330), .B(new_n4143), .Y(new_n4144));
  nor_5  g01796(.A(n25316), .B(n7657), .Y(new_n4145));
  not_8  g01797(.A(n20385), .Y(new_n4146_1));
  or_5   g01798(.A(new_n3982), .B(new_n4146_1), .Y(new_n4147));
  xnor_4 g01799(.A(n25316), .B(new_n3978), .Y(new_n4148));
  and_5  g01800(.A(new_n4148), .B(new_n4147), .Y(new_n4149));
  nor_5  g01801(.A(new_n4149), .B(new_n4145), .Y(new_n4150_1));
  xnor_4 g01802(.A(new_n4150_1), .B(new_n4144), .Y(new_n4151_1));
  xnor_4 g01803(.A(new_n4151_1), .B(new_n4142), .Y(new_n4152_1));
  xor_4  g01804(.A(new_n4139), .B(new_n4137), .Y(new_n4153_1));
  nor_5  g01805(.A(new_n3982), .B(new_n4146_1), .Y(new_n4154));
  xnor_4 g01806(.A(new_n4148), .B(new_n4154), .Y(new_n4155));
  nor_5  g01807(.A(new_n4155), .B(new_n4153_1), .Y(new_n4156));
  xnor_4 g01808(.A(n25926), .B(n20385), .Y(new_n4157));
  xnor_4 g01809(.A(new_n4136), .B(new_n4134_1), .Y(new_n4158));
  nor_5  g01810(.A(new_n4158), .B(new_n4157), .Y(new_n4159));
  not_8  g01811(.A(new_n4155), .Y(new_n4160));
  xnor_4 g01812(.A(new_n4160), .B(new_n4153_1), .Y(new_n4161));
  and_5  g01813(.A(new_n4161), .B(new_n4159), .Y(new_n4162));
  nor_5  g01814(.A(new_n4162), .B(new_n4156), .Y(new_n4163));
  xnor_4 g01815(.A(new_n4163), .B(new_n4152_1), .Y(n248));
  not_8  g01816(.A(n6369), .Y(new_n4165_1));
  nor_5  g01817(.A(n24732), .B(n6631), .Y(new_n4166));
  not_8  g01818(.A(new_n4166), .Y(new_n4167));
  nor_5  g01819(.A(new_n4167), .B(n14684), .Y(new_n4168));
  not_8  g01820(.A(new_n4168), .Y(new_n4169));
  nor_5  g01821(.A(new_n4169), .B(n17035), .Y(new_n4170));
  xnor_4 g01822(.A(new_n4170), .B(n19905), .Y(new_n4171));
  xnor_4 g01823(.A(new_n4171), .B(new_n4165_1), .Y(new_n4172_1));
  xnor_4 g01824(.A(new_n4168), .B(n17035), .Y(new_n4173_1));
  and_5  g01825(.A(new_n4173_1), .B(n25797), .Y(new_n4174));
  xnor_4 g01826(.A(new_n4173_1), .B(n25797), .Y(new_n4175));
  xnor_4 g01827(.A(new_n4166), .B(n14684), .Y(new_n4176_1));
  nor_5  g01828(.A(new_n4176_1), .B(n15967), .Y(new_n4177));
  not_8  g01829(.A(n15967), .Y(new_n4178));
  xnor_4 g01830(.A(new_n4176_1), .B(new_n4178), .Y(new_n4179));
  not_8  g01831(.A(n6631), .Y(new_n4180));
  xnor_4 g01832(.A(n24732), .B(new_n4180), .Y(new_n4181));
  nor_5  g01833(.A(new_n4181), .B(n13319), .Y(new_n4182));
  not_8  g01834(.A(n24732), .Y(new_n4183));
  or_5   g01835(.A(new_n3756), .B(new_n4183), .Y(new_n4184));
  not_8  g01836(.A(new_n4181), .Y(new_n4185));
  xnor_4 g01837(.A(new_n4185), .B(n13319), .Y(new_n4186_1));
  and_5  g01838(.A(new_n4186_1), .B(new_n4184), .Y(new_n4187));
  or_5   g01839(.A(new_n4187), .B(new_n4182), .Y(new_n4188));
  and_5  g01840(.A(new_n4188), .B(new_n4179), .Y(new_n4189));
  nor_5  g01841(.A(new_n4189), .B(new_n4177), .Y(new_n4190));
  not_8  g01842(.A(new_n4190), .Y(new_n4191));
  nor_5  g01843(.A(new_n4191), .B(new_n4175), .Y(new_n4192));
  nor_5  g01844(.A(new_n4192), .B(new_n4174), .Y(new_n4193));
  xnor_4 g01845(.A(new_n4193), .B(new_n4172_1), .Y(new_n4194));
  not_8  g01846(.A(new_n4194), .Y(new_n4195));
  nor_5  g01847(.A(n14148), .B(n1152), .Y(new_n4196));
  not_8  g01848(.A(new_n4196), .Y(new_n4197));
  nor_5  g01849(.A(new_n4197), .B(n7149), .Y(new_n4198));
  not_8  g01850(.A(new_n4198), .Y(new_n4199));
  nor_5  g01851(.A(new_n4199), .B(n18558), .Y(new_n4200));
  xnor_4 g01852(.A(new_n4200), .B(n3468), .Y(new_n4201));
  not_8  g01853(.A(new_n4201), .Y(new_n4202));
  xnor_4 g01854(.A(new_n4202), .B(n19514), .Y(new_n4203));
  xnor_4 g01855(.A(new_n4198), .B(n18558), .Y(new_n4204_1));
  and_5  g01856(.A(new_n4204_1), .B(n10053), .Y(new_n4205_1));
  xnor_4 g01857(.A(new_n4204_1), .B(new_n2944_1), .Y(new_n4206));
  xnor_4 g01858(.A(new_n4196), .B(n7149), .Y(new_n4207));
  not_8  g01859(.A(new_n4207), .Y(new_n4208));
  nor_5  g01860(.A(new_n4208), .B(new_n2947), .Y(new_n4209));
  xnor_4 g01861(.A(new_n4208), .B(n8399), .Y(new_n4210));
  xnor_4 g01862(.A(n14148), .B(n1152), .Y(new_n4211));
  nor_5  g01863(.A(new_n4211), .B(new_n3824), .Y(new_n4212));
  nor_5  g01864(.A(new_n2952), .B(new_n2698), .Y(new_n4213));
  xnor_4 g01865(.A(new_n4211), .B(n9507), .Y(new_n4214));
  and_5  g01866(.A(new_n4214), .B(new_n4213), .Y(new_n4215_1));
  or_5   g01867(.A(new_n4215_1), .B(new_n4212), .Y(new_n4216));
  and_5  g01868(.A(new_n4216), .B(new_n4210), .Y(new_n4217));
  or_5   g01869(.A(new_n4217), .B(new_n4209), .Y(new_n4218));
  and_5  g01870(.A(new_n4218), .B(new_n4206), .Y(new_n4219));
  nor_5  g01871(.A(new_n4219), .B(new_n4205_1), .Y(new_n4220));
  xnor_4 g01872(.A(new_n4220), .B(new_n4203), .Y(new_n4221_1));
  not_8  g01873(.A(new_n4221_1), .Y(new_n4222));
  not_8  g01874(.A(n626), .Y(new_n4223));
  nor_5  g01875(.A(n10057), .B(n8920), .Y(new_n4224_1));
  not_8  g01876(.A(new_n4224_1), .Y(new_n4225));
  nor_5  g01877(.A(new_n4225), .B(n26748), .Y(new_n4226));
  not_8  g01878(.A(new_n4226), .Y(new_n4227));
  nor_5  g01879(.A(new_n4227), .B(n21276), .Y(new_n4228));
  xnor_4 g01880(.A(new_n4228), .B(n13668), .Y(new_n4229));
  xnor_4 g01881(.A(new_n4229), .B(new_n4223), .Y(new_n4230));
  xnor_4 g01882(.A(new_n4226), .B(n21276), .Y(new_n4231_1));
  and_5  g01883(.A(new_n4231_1), .B(n1204), .Y(new_n4232));
  not_8  g01884(.A(n1204), .Y(new_n4233));
  xnor_4 g01885(.A(new_n4231_1), .B(new_n4233), .Y(new_n4234));
  xnor_4 g01886(.A(new_n4224_1), .B(n26748), .Y(new_n4235));
  and_5  g01887(.A(new_n4235), .B(n19618), .Y(new_n4236));
  not_8  g01888(.A(n19618), .Y(new_n4237));
  xnor_4 g01889(.A(new_n4235), .B(new_n4237), .Y(new_n4238));
  xnor_4 g01890(.A(n10057), .B(n8920), .Y(new_n4239));
  not_8  g01891(.A(new_n4239), .Y(new_n4240));
  nor_5  g01892(.A(new_n4240), .B(n22043), .Y(new_n4241));
  not_8  g01893(.A(n8920), .Y(new_n4242));
  or_5   g01894(.A(new_n3875), .B(new_n4242), .Y(new_n4243));
  xnor_4 g01895(.A(new_n4239), .B(n22043), .Y(new_n4244));
  and_5  g01896(.A(new_n4244), .B(new_n4243), .Y(new_n4245));
  nor_5  g01897(.A(new_n4245), .B(new_n4241), .Y(new_n4246));
  and_5  g01898(.A(new_n4246), .B(new_n4238), .Y(new_n4247));
  or_5   g01899(.A(new_n4247), .B(new_n4236), .Y(new_n4248));
  and_5  g01900(.A(new_n4248), .B(new_n4234), .Y(new_n4249));
  nor_5  g01901(.A(new_n4249), .B(new_n4232), .Y(new_n4250));
  xnor_4 g01902(.A(new_n4250), .B(new_n4230), .Y(new_n4251));
  xnor_4 g01903(.A(new_n4251), .B(new_n4222), .Y(new_n4252));
  nor_5  g01904(.A(new_n4217), .B(new_n4209), .Y(new_n4253));
  xnor_4 g01905(.A(new_n4253), .B(new_n4206), .Y(new_n4254));
  not_8  g01906(.A(new_n4254), .Y(new_n4255));
  nor_5  g01907(.A(new_n4247), .B(new_n4236), .Y(new_n4256_1));
  xnor_4 g01908(.A(new_n4256_1), .B(new_n4234), .Y(new_n4257));
  not_8  g01909(.A(new_n4257), .Y(new_n4258));
  nor_5  g01910(.A(new_n4258), .B(new_n4255), .Y(new_n4259));
  xnor_4 g01911(.A(new_n4258), .B(new_n4255), .Y(new_n4260));
  xnor_4 g01912(.A(new_n4246), .B(new_n4238), .Y(new_n4261));
  xnor_4 g01913(.A(new_n4214), .B(new_n4213), .Y(new_n4262));
  nor_5  g01914(.A(new_n3875), .B(new_n4242), .Y(new_n4263));
  xnor_4 g01915(.A(new_n4244), .B(new_n4263), .Y(new_n4264));
  nor_5  g01916(.A(new_n4264), .B(new_n4262), .Y(new_n4265));
  xnor_4 g01917(.A(n12121), .B(n8920), .Y(new_n4266_1));
  xnor_4 g01918(.A(n26979), .B(new_n2698), .Y(new_n4267));
  not_8  g01919(.A(new_n4267), .Y(new_n4268));
  nor_5  g01920(.A(new_n4268), .B(new_n4266_1), .Y(new_n4269));
  not_8  g01921(.A(new_n4262), .Y(new_n4270));
  xnor_4 g01922(.A(new_n4264), .B(new_n4270), .Y(new_n4271));
  and_5  g01923(.A(new_n4271), .B(new_n4269), .Y(new_n4272_1));
  nor_5  g01924(.A(new_n4272_1), .B(new_n4265), .Y(new_n4273));
  nor_5  g01925(.A(new_n4273), .B(new_n4261), .Y(new_n4274));
  nor_5  g01926(.A(new_n4215_1), .B(new_n4212), .Y(new_n4275));
  xnor_4 g01927(.A(new_n4275), .B(new_n4210), .Y(new_n4276));
  not_8  g01928(.A(new_n4261), .Y(new_n4277));
  xnor_4 g01929(.A(new_n4273), .B(new_n4277), .Y(new_n4278));
  and_5  g01930(.A(new_n4278), .B(new_n4276), .Y(new_n4279));
  nor_5  g01931(.A(new_n4279), .B(new_n4274), .Y(new_n4280));
  nor_5  g01932(.A(new_n4280), .B(new_n4260), .Y(new_n4281));
  or_5   g01933(.A(new_n4281), .B(new_n4259), .Y(new_n4282));
  xor_4  g01934(.A(new_n4282), .B(new_n4252), .Y(new_n4283));
  xnor_4 g01935(.A(new_n4283), .B(new_n4195), .Y(new_n4284));
  xnor_4 g01936(.A(new_n4190), .B(new_n4175), .Y(new_n4285));
  not_8  g01937(.A(new_n4285), .Y(new_n4286));
  xnor_4 g01938(.A(new_n4280), .B(new_n4260), .Y(new_n4287));
  nor_5  g01939(.A(new_n4287), .B(new_n4286), .Y(new_n4288));
  xnor_4 g01940(.A(new_n4287), .B(new_n4285), .Y(new_n4289));
  not_8  g01941(.A(new_n4276), .Y(new_n4290));
  xnor_4 g01942(.A(new_n4278), .B(new_n4290), .Y(new_n4291));
  not_8  g01943(.A(new_n4291), .Y(new_n4292));
  xor_4  g01944(.A(new_n4188), .B(new_n4179), .Y(new_n4293));
  nor_5  g01945(.A(new_n4293), .B(new_n4292), .Y(new_n4294));
  xnor_4 g01946(.A(new_n4293), .B(new_n4291), .Y(new_n4295));
  xnor_4 g01947(.A(new_n4271), .B(new_n4269), .Y(new_n4296));
  not_8  g01948(.A(new_n4296), .Y(new_n4297));
  nor_5  g01949(.A(new_n4297), .B(new_n4186_1), .Y(new_n4298));
  xor_4  g01950(.A(new_n4186_1), .B(new_n4184), .Y(new_n4299));
  nor_5  g01951(.A(new_n4299), .B(new_n4296), .Y(new_n4300));
  xnor_4 g01952(.A(n25435), .B(n24732), .Y(new_n4301));
  xnor_4 g01953(.A(new_n4267), .B(new_n4266_1), .Y(new_n4302));
  not_8  g01954(.A(new_n4302), .Y(new_n4303));
  nor_5  g01955(.A(new_n4303), .B(new_n4301), .Y(new_n4304));
  nor_5  g01956(.A(new_n4304), .B(new_n4300), .Y(new_n4305));
  nor_5  g01957(.A(new_n4305), .B(new_n4298), .Y(new_n4306_1));
  and_5  g01958(.A(new_n4306_1), .B(new_n4295), .Y(new_n4307));
  or_5   g01959(.A(new_n4307), .B(new_n4294), .Y(new_n4308));
  and_5  g01960(.A(new_n4308), .B(new_n4289), .Y(new_n4309));
  nor_5  g01961(.A(new_n4309), .B(new_n4288), .Y(new_n4310));
  xnor_4 g01962(.A(new_n4310), .B(new_n4284), .Y(n266));
  not_8  g01963(.A(n21839), .Y(new_n4312));
  nor_5  g01964(.A(n22270), .B(new_n4312), .Y(new_n4313));
  xnor_4 g01965(.A(n22270), .B(n21839), .Y(new_n4314));
  not_8  g01966(.A(n27089), .Y(new_n4315));
  nor_5  g01967(.A(new_n4315), .B(n8806), .Y(new_n4316));
  xnor_4 g01968(.A(n27089), .B(n8806), .Y(new_n4317));
  nor_5  g01969(.A(new_n2929_1), .B(n2479), .Y(new_n4318));
  xnor_4 g01970(.A(n11841), .B(n2479), .Y(new_n4319_1));
  nor_5  g01971(.A(new_n2933), .B(n9372), .Y(new_n4320));
  xnor_4 g01972(.A(n10710), .B(n9372), .Y(new_n4321));
  nor_5  g01973(.A(new_n2937), .B(n6596), .Y(new_n4322));
  xnor_4 g01974(.A(n20929), .B(n6596), .Y(new_n4323));
  nor_5  g01975(.A(n15289), .B(new_n2941), .Y(new_n4324));
  xnor_4 g01976(.A(n15289), .B(n8006), .Y(new_n4325_1));
  and_5  g01977(.A(n25074), .B(new_n2692), .Y(new_n4326_1));
  xnor_4 g01978(.A(n25074), .B(n6556), .Y(new_n4327));
  not_8  g01979(.A(n16396), .Y(new_n4328));
  and_5  g01980(.A(n22871), .B(new_n4328), .Y(new_n4329));
  nor_5  g01981(.A(n22871), .B(new_n4328), .Y(new_n4330));
  not_8  g01982(.A(n9399), .Y(new_n4331));
  and_5  g01983(.A(n14275), .B(new_n4331), .Y(new_n4332));
  nor_5  g01984(.A(n14275), .B(new_n4331), .Y(new_n4333));
  nor_5  g01985(.A(new_n2699), .B(n2088), .Y(new_n4334));
  not_8  g01986(.A(new_n4334), .Y(new_n4335));
  nor_5  g01987(.A(new_n4335), .B(new_n4333), .Y(new_n4336));
  nor_5  g01988(.A(new_n4336), .B(new_n4332), .Y(new_n4337));
  nor_5  g01989(.A(new_n4337), .B(new_n4330), .Y(new_n4338));
  nor_5  g01990(.A(new_n4338), .B(new_n4329), .Y(new_n4339));
  and_5  g01991(.A(new_n4339), .B(new_n4327), .Y(new_n4340_1));
  or_5   g01992(.A(new_n4340_1), .B(new_n4326_1), .Y(new_n4341));
  and_5  g01993(.A(new_n4341), .B(new_n4325_1), .Y(new_n4342));
  or_5   g01994(.A(new_n4342), .B(new_n4324), .Y(new_n4343));
  and_5  g01995(.A(new_n4343), .B(new_n4323), .Y(new_n4344));
  or_5   g01996(.A(new_n4344), .B(new_n4322), .Y(new_n4345));
  and_5  g01997(.A(new_n4345), .B(new_n4321), .Y(new_n4346));
  or_5   g01998(.A(new_n4346), .B(new_n4320), .Y(new_n4347));
  and_5  g01999(.A(new_n4347), .B(new_n4319_1), .Y(new_n4348));
  or_5   g02000(.A(new_n4348), .B(new_n4318), .Y(new_n4349));
  and_5  g02001(.A(new_n4349), .B(new_n4317), .Y(new_n4350));
  or_5   g02002(.A(new_n4350), .B(new_n4316), .Y(new_n4351));
  and_5  g02003(.A(new_n4351), .B(new_n4314), .Y(new_n4352));
  nor_5  g02004(.A(new_n4352), .B(new_n4313), .Y(new_n4353));
  nor_5  g02005(.A(new_n4350), .B(new_n4316), .Y(new_n4354));
  xnor_4 g02006(.A(new_n4354), .B(new_n4314), .Y(new_n4355));
  nor_5  g02007(.A(new_n4355), .B(n23272), .Y(new_n4356));
  not_8  g02008(.A(new_n4355), .Y(new_n4357));
  xnor_4 g02009(.A(new_n4357), .B(n23272), .Y(new_n4358));
  xor_4  g02010(.A(new_n4349), .B(new_n4317), .Y(new_n4359));
  nor_5  g02011(.A(new_n4359), .B(n11481), .Y(new_n4360));
  not_8  g02012(.A(n11481), .Y(new_n4361));
  xnor_4 g02013(.A(new_n4359), .B(new_n4361), .Y(new_n4362));
  xor_4  g02014(.A(new_n4347), .B(new_n4319_1), .Y(new_n4363));
  nor_5  g02015(.A(new_n4363), .B(n16439), .Y(new_n4364));
  not_8  g02016(.A(n16439), .Y(new_n4365));
  xnor_4 g02017(.A(new_n4363), .B(new_n4365), .Y(new_n4366));
  xor_4  g02018(.A(new_n4345), .B(new_n4321), .Y(new_n4367));
  nor_5  g02019(.A(new_n4367), .B(n15241), .Y(new_n4368));
  not_8  g02020(.A(n15241), .Y(new_n4369));
  xnor_4 g02021(.A(new_n4367), .B(new_n4369), .Y(new_n4370));
  xor_4  g02022(.A(new_n4343), .B(new_n4323), .Y(new_n4371));
  nor_5  g02023(.A(new_n4371), .B(n7678), .Y(new_n4372));
  not_8  g02024(.A(n7678), .Y(new_n4373));
  xnor_4 g02025(.A(new_n4371), .B(new_n4373), .Y(new_n4374_1));
  xor_4  g02026(.A(new_n4341), .B(new_n4325_1), .Y(new_n4375));
  nor_5  g02027(.A(new_n4375), .B(n3785), .Y(new_n4376_1));
  not_8  g02028(.A(n3785), .Y(new_n4377));
  xnor_4 g02029(.A(new_n4375), .B(new_n4377), .Y(new_n4378));
  xnor_4 g02030(.A(new_n4339), .B(new_n4327), .Y(new_n4379));
  not_8  g02031(.A(new_n4379), .Y(new_n4380));
  nor_5  g02032(.A(new_n4380), .B(n20250), .Y(new_n4381));
  not_8  g02033(.A(n20250), .Y(new_n4382));
  xnor_4 g02034(.A(new_n4380), .B(new_n4382), .Y(new_n4383));
  not_8  g02035(.A(n5822), .Y(new_n4384));
  xnor_4 g02036(.A(n22871), .B(n16396), .Y(new_n4385));
  xnor_4 g02037(.A(new_n4385), .B(new_n4337), .Y(new_n4386));
  nor_5  g02038(.A(new_n4386), .B(new_n4384), .Y(new_n4387));
  not_8  g02039(.A(new_n4386), .Y(new_n4388));
  or_5   g02040(.A(new_n4388), .B(n5822), .Y(new_n4389));
  xnor_4 g02041(.A(n14275), .B(n9399), .Y(new_n4390));
  xnor_4 g02042(.A(new_n4390), .B(new_n4335), .Y(new_n4391));
  not_8  g02043(.A(new_n4391), .Y(new_n4392));
  nor_5  g02044(.A(new_n4392), .B(n26443), .Y(new_n4393));
  not_8  g02045(.A(n1681), .Y(new_n4394));
  xnor_4 g02046(.A(n25023), .B(n2088), .Y(new_n4395));
  or_5   g02047(.A(new_n4395), .B(new_n4394), .Y(new_n4396));
  xnor_4 g02048(.A(new_n4391), .B(n26443), .Y(new_n4397));
  and_5  g02049(.A(new_n4397), .B(new_n4396), .Y(new_n4398));
  nor_5  g02050(.A(new_n4398), .B(new_n4393), .Y(new_n4399));
  and_5  g02051(.A(new_n4399), .B(new_n4389), .Y(new_n4400));
  nor_5  g02052(.A(new_n4400), .B(new_n4387), .Y(new_n4401_1));
  and_5  g02053(.A(new_n4401_1), .B(new_n4383), .Y(new_n4402));
  or_5   g02054(.A(new_n4402), .B(new_n4381), .Y(new_n4403));
  and_5  g02055(.A(new_n4403), .B(new_n4378), .Y(new_n4404));
  or_5   g02056(.A(new_n4404), .B(new_n4376_1), .Y(new_n4405));
  and_5  g02057(.A(new_n4405), .B(new_n4374_1), .Y(new_n4406));
  or_5   g02058(.A(new_n4406), .B(new_n4372), .Y(new_n4407));
  and_5  g02059(.A(new_n4407), .B(new_n4370), .Y(new_n4408));
  or_5   g02060(.A(new_n4408), .B(new_n4368), .Y(new_n4409_1));
  and_5  g02061(.A(new_n4409_1), .B(new_n4366), .Y(new_n4410));
  or_5   g02062(.A(new_n4410), .B(new_n4364), .Y(new_n4411));
  and_5  g02063(.A(new_n4411), .B(new_n4362), .Y(new_n4412));
  or_5   g02064(.A(new_n4412), .B(new_n4360), .Y(new_n4413));
  and_5  g02065(.A(new_n4413), .B(new_n4358), .Y(new_n4414));
  nor_5  g02066(.A(new_n4414), .B(new_n4356), .Y(new_n4415));
  and_5  g02067(.A(new_n4415), .B(new_n4353), .Y(new_n4416));
  not_8  g02068(.A(new_n4416), .Y(new_n4417));
  not_8  g02069(.A(new_n3934_1), .Y(new_n4418));
  nor_5  g02070(.A(new_n4418), .B(n19477), .Y(new_n4419));
  not_8  g02071(.A(new_n4419), .Y(new_n4420));
  nor_5  g02072(.A(new_n4420), .B(n9318), .Y(new_n4421));
  not_8  g02073(.A(new_n4421), .Y(new_n4422));
  nor_5  g02074(.A(new_n4422), .B(n25168), .Y(new_n4423));
  not_8  g02075(.A(new_n4423), .Y(new_n4424_1));
  nor_5  g02076(.A(new_n4424_1), .B(n1999), .Y(new_n4425));
  and_5  g02077(.A(new_n4425), .B(new_n2554), .Y(new_n4426_1));
  xnor_4 g02078(.A(new_n4425), .B(n9396), .Y(new_n4427));
  nor_5  g02079(.A(new_n4427), .B(n18880), .Y(new_n4428));
  xnor_4 g02080(.A(new_n4423), .B(n1999), .Y(new_n4429));
  nor_5  g02081(.A(new_n4429), .B(n25475), .Y(new_n4430));
  not_8  g02082(.A(n25475), .Y(new_n4431));
  xnor_4 g02083(.A(new_n4429), .B(new_n4431), .Y(new_n4432_1));
  xnor_4 g02084(.A(new_n4421), .B(n25168), .Y(new_n4433));
  nor_5  g02085(.A(new_n4433), .B(n23849), .Y(new_n4434));
  not_8  g02086(.A(n23849), .Y(new_n4435));
  xnor_4 g02087(.A(new_n4433), .B(new_n4435), .Y(new_n4436));
  xnor_4 g02088(.A(new_n4419), .B(n9318), .Y(new_n4437));
  nor_5  g02089(.A(new_n4437), .B(n12446), .Y(new_n4438));
  nor_5  g02090(.A(new_n3935), .B(n11011), .Y(new_n4439));
  nor_5  g02091(.A(new_n3962_1), .B(new_n3936), .Y(new_n4440));
  or_5   g02092(.A(new_n4440), .B(new_n4439), .Y(new_n4441_1));
  not_8  g02093(.A(n12446), .Y(new_n4442));
  xnor_4 g02094(.A(new_n4437), .B(new_n4442), .Y(new_n4443));
  and_5  g02095(.A(new_n4443), .B(new_n4441_1), .Y(new_n4444));
  or_5   g02096(.A(new_n4444), .B(new_n4438), .Y(new_n4445));
  and_5  g02097(.A(new_n4445), .B(new_n4436), .Y(new_n4446));
  or_5   g02098(.A(new_n4446), .B(new_n4434), .Y(new_n4447));
  and_5  g02099(.A(new_n4447), .B(new_n4432_1), .Y(new_n4448));
  nor_5  g02100(.A(new_n4448), .B(new_n4430), .Y(new_n4449));
  and_5  g02101(.A(new_n4427), .B(n18880), .Y(new_n4450));
  nor_5  g02102(.A(new_n4450), .B(new_n4449), .Y(new_n4451_1));
  nor_5  g02103(.A(new_n4451_1), .B(new_n4428), .Y(new_n4452));
  nor_5  g02104(.A(new_n4452), .B(new_n4426_1), .Y(new_n4453));
  nor_5  g02105(.A(n24032), .B(n22843), .Y(new_n4454));
  not_8  g02106(.A(new_n4454), .Y(new_n4455));
  nor_5  g02107(.A(new_n4455), .B(n6785), .Y(new_n4456));
  not_8  g02108(.A(new_n4456), .Y(new_n4457));
  nor_5  g02109(.A(new_n4457), .B(n24879), .Y(new_n4458));
  not_8  g02110(.A(new_n4458), .Y(new_n4459));
  nor_5  g02111(.A(new_n4459), .B(n268), .Y(new_n4460));
  not_8  g02112(.A(new_n4460), .Y(new_n4461));
  nor_5  g02113(.A(new_n4461), .B(n12587), .Y(new_n4462));
  not_8  g02114(.A(new_n4462), .Y(new_n4463));
  nor_5  g02115(.A(new_n4463), .B(n25381), .Y(new_n4464));
  not_8  g02116(.A(new_n4464), .Y(new_n4465));
  nor_5  g02117(.A(new_n4465), .B(n16376), .Y(new_n4466));
  not_8  g02118(.A(new_n4466), .Y(new_n4467));
  nor_5  g02119(.A(new_n4467), .B(n24196), .Y(new_n4468));
  xnor_4 g02120(.A(new_n4468), .B(n18105), .Y(new_n4469));
  not_8  g02121(.A(new_n4469), .Y(new_n4470));
  not_8  g02122(.A(n18880), .Y(new_n4471));
  xnor_4 g02123(.A(new_n4427), .B(new_n4471), .Y(new_n4472));
  xnor_4 g02124(.A(new_n4472), .B(new_n4449), .Y(new_n4473));
  nor_5  g02125(.A(new_n4473), .B(new_n4470), .Y(new_n4474));
  not_8  g02126(.A(new_n4468), .Y(new_n4475));
  nor_5  g02127(.A(new_n4475), .B(n18105), .Y(new_n4476_1));
  not_8  g02128(.A(new_n4473), .Y(new_n4477));
  xnor_4 g02129(.A(new_n4477), .B(new_n4470), .Y(new_n4478_1));
  xnor_4 g02130(.A(new_n4466), .B(n24196), .Y(new_n4479));
  nor_5  g02131(.A(new_n4446), .B(new_n4434), .Y(new_n4480));
  xnor_4 g02132(.A(new_n4480), .B(new_n4432_1), .Y(new_n4481));
  not_8  g02133(.A(new_n4481), .Y(new_n4482));
  nor_5  g02134(.A(new_n4482), .B(new_n4479), .Y(new_n4483));
  xnor_4 g02135(.A(new_n4482), .B(new_n4479), .Y(new_n4484));
  xnor_4 g02136(.A(new_n4464), .B(n16376), .Y(new_n4485));
  nor_5  g02137(.A(new_n4444), .B(new_n4438), .Y(new_n4486));
  xnor_4 g02138(.A(new_n4486), .B(new_n4436), .Y(new_n4487));
  not_8  g02139(.A(new_n4487), .Y(new_n4488));
  nor_5  g02140(.A(new_n4488), .B(new_n4485), .Y(new_n4489));
  xnor_4 g02141(.A(new_n4488), .B(new_n4485), .Y(new_n4490));
  xnor_4 g02142(.A(new_n4462), .B(n25381), .Y(new_n4491));
  xor_4  g02143(.A(new_n4443), .B(new_n4441_1), .Y(new_n4492));
  not_8  g02144(.A(new_n4492), .Y(new_n4493));
  nor_5  g02145(.A(new_n4493), .B(new_n4491), .Y(new_n4494));
  xnor_4 g02146(.A(new_n4493), .B(new_n4491), .Y(new_n4495));
  xnor_4 g02147(.A(new_n4460), .B(n12587), .Y(new_n4496));
  nor_5  g02148(.A(new_n4496), .B(new_n3963), .Y(new_n4497));
  xnor_4 g02149(.A(new_n4496), .B(new_n3963), .Y(new_n4498));
  xnor_4 g02150(.A(new_n4458), .B(n268), .Y(new_n4499));
  nor_5  g02151(.A(new_n4499), .B(new_n3965), .Y(new_n4500));
  xnor_4 g02152(.A(new_n4456), .B(n24879), .Y(new_n4501));
  nor_5  g02153(.A(new_n4501), .B(new_n3970), .Y(new_n4502));
  xnor_4 g02154(.A(new_n4501), .B(new_n3968), .Y(new_n4503));
  xnor_4 g02155(.A(new_n4454), .B(n6785), .Y(new_n4504));
  and_5  g02156(.A(new_n4504), .B(new_n3976), .Y(new_n4505));
  xnor_4 g02157(.A(new_n4504), .B(new_n3974), .Y(new_n4506));
  not_8  g02158(.A(n22843), .Y(new_n4507));
  xnor_4 g02159(.A(n24032), .B(new_n4507), .Y(new_n4508));
  nor_5  g02160(.A(new_n4508), .B(new_n3984_1), .Y(new_n4509));
  or_5   g02161(.A(new_n2551), .B(new_n4507), .Y(new_n4510));
  xnor_4 g02162(.A(new_n4508), .B(new_n3980), .Y(new_n4511));
  and_5  g02163(.A(new_n4511), .B(new_n4510), .Y(new_n4512));
  nor_5  g02164(.A(new_n4512), .B(new_n4509), .Y(new_n4513));
  and_5  g02165(.A(new_n4513), .B(new_n4506), .Y(new_n4514_1));
  nor_5  g02166(.A(new_n4514_1), .B(new_n4505), .Y(new_n4515));
  and_5  g02167(.A(new_n4515), .B(new_n4503), .Y(new_n4516));
  nor_5  g02168(.A(new_n4516), .B(new_n4502), .Y(new_n4517));
  xnor_4 g02169(.A(new_n4499), .B(new_n3965), .Y(new_n4518));
  nor_5  g02170(.A(new_n4518), .B(new_n4517), .Y(new_n4519));
  nor_5  g02171(.A(new_n4519), .B(new_n4500), .Y(new_n4520));
  nor_5  g02172(.A(new_n4520), .B(new_n4498), .Y(new_n4521));
  nor_5  g02173(.A(new_n4521), .B(new_n4497), .Y(new_n4522));
  nor_5  g02174(.A(new_n4522), .B(new_n4495), .Y(new_n4523));
  nor_5  g02175(.A(new_n4523), .B(new_n4494), .Y(new_n4524));
  nor_5  g02176(.A(new_n4524), .B(new_n4490), .Y(new_n4525));
  nor_5  g02177(.A(new_n4525), .B(new_n4489), .Y(new_n4526));
  nor_5  g02178(.A(new_n4526), .B(new_n4484), .Y(new_n4527));
  nor_5  g02179(.A(new_n4527), .B(new_n4483), .Y(new_n4528));
  and_5  g02180(.A(new_n4528), .B(new_n4478_1), .Y(new_n4529_1));
  or_5   g02181(.A(new_n4529_1), .B(new_n4476_1), .Y(new_n4530));
  nor_5  g02182(.A(new_n4530), .B(new_n4474), .Y(new_n4531));
  not_8  g02183(.A(new_n4531), .Y(new_n4532));
  nor_5  g02184(.A(new_n4532), .B(new_n4453), .Y(new_n4533));
  xnor_4 g02185(.A(new_n4533), .B(new_n4417), .Y(new_n4534));
  not_8  g02186(.A(new_n4415), .Y(new_n4535));
  xnor_4 g02187(.A(new_n4535), .B(new_n4353), .Y(new_n4536));
  not_8  g02188(.A(new_n4536), .Y(new_n4537));
  not_8  g02189(.A(new_n4453), .Y(new_n4538));
  xnor_4 g02190(.A(new_n4532), .B(new_n4538), .Y(new_n4539));
  and_5  g02191(.A(new_n4539), .B(new_n4537), .Y(new_n4540));
  xnor_4 g02192(.A(new_n4539), .B(new_n4537), .Y(new_n4541));
  xnor_4 g02193(.A(new_n4528), .B(new_n4478_1), .Y(new_n4542));
  nor_5  g02194(.A(new_n4412), .B(new_n4360), .Y(new_n4543));
  xnor_4 g02195(.A(new_n4543), .B(new_n4358), .Y(new_n4544));
  and_5  g02196(.A(new_n4544), .B(new_n4542), .Y(new_n4545));
  xnor_4 g02197(.A(new_n4544), .B(new_n4542), .Y(new_n4546));
  xnor_4 g02198(.A(new_n4526), .B(new_n4484), .Y(new_n4547));
  xor_4  g02199(.A(new_n4411), .B(new_n4362), .Y(new_n4548));
  not_8  g02200(.A(new_n4548), .Y(new_n4549));
  nor_5  g02201(.A(new_n4549), .B(new_n4547), .Y(new_n4550));
  xnor_4 g02202(.A(new_n4549), .B(new_n4547), .Y(new_n4551));
  xnor_4 g02203(.A(new_n4524), .B(new_n4490), .Y(new_n4552_1));
  xor_4  g02204(.A(new_n4409_1), .B(new_n4366), .Y(new_n4553));
  not_8  g02205(.A(new_n4553), .Y(new_n4554));
  nor_5  g02206(.A(new_n4554), .B(new_n4552_1), .Y(new_n4555));
  xnor_4 g02207(.A(new_n4554), .B(new_n4552_1), .Y(new_n4556));
  xnor_4 g02208(.A(new_n4522), .B(new_n4495), .Y(new_n4557));
  xor_4  g02209(.A(new_n4407), .B(new_n4370), .Y(new_n4558));
  not_8  g02210(.A(new_n4558), .Y(new_n4559));
  nor_5  g02211(.A(new_n4559), .B(new_n4557), .Y(new_n4560));
  xnor_4 g02212(.A(new_n4559), .B(new_n4557), .Y(new_n4561));
  xnor_4 g02213(.A(new_n4520), .B(new_n4498), .Y(new_n4562));
  xor_4  g02214(.A(new_n4405), .B(new_n4374_1), .Y(new_n4563));
  not_8  g02215(.A(new_n4563), .Y(new_n4564));
  nor_5  g02216(.A(new_n4564), .B(new_n4562), .Y(new_n4565));
  xnor_4 g02217(.A(new_n4564), .B(new_n4562), .Y(new_n4566));
  xor_4  g02218(.A(new_n4403), .B(new_n4378), .Y(new_n4567));
  not_8  g02219(.A(new_n4567), .Y(new_n4568));
  xnor_4 g02220(.A(new_n4518), .B(new_n4517), .Y(new_n4569));
  nor_5  g02221(.A(new_n4569), .B(new_n4568), .Y(new_n4570));
  xnor_4 g02222(.A(new_n4569), .B(new_n4568), .Y(new_n4571));
  xnor_4 g02223(.A(new_n4515), .B(new_n4503), .Y(new_n4572));
  xnor_4 g02224(.A(new_n4401_1), .B(new_n4383), .Y(new_n4573));
  nor_5  g02225(.A(new_n4573), .B(new_n4572), .Y(new_n4574));
  not_8  g02226(.A(new_n4573), .Y(new_n4575));
  xnor_4 g02227(.A(new_n4575), .B(new_n4572), .Y(new_n4576));
  xnor_4 g02228(.A(new_n4513), .B(new_n4506), .Y(new_n4577));
  xnor_4 g02229(.A(new_n4388), .B(new_n4384), .Y(new_n4578));
  xnor_4 g02230(.A(new_n4578), .B(new_n4399), .Y(new_n4579));
  nor_5  g02231(.A(new_n4579), .B(new_n4577), .Y(new_n4580));
  xor_4  g02232(.A(new_n4397), .B(new_n4396), .Y(new_n4581));
  xor_4  g02233(.A(new_n4511), .B(new_n4510), .Y(new_n4582));
  and_5  g02234(.A(new_n4582), .B(new_n4581), .Y(new_n4583));
  xnor_4 g02235(.A(new_n2551), .B(new_n4507), .Y(new_n4584));
  xnor_4 g02236(.A(new_n4395), .B(n1681), .Y(new_n4585));
  not_8  g02237(.A(new_n4585), .Y(new_n4586));
  nor_5  g02238(.A(new_n4586), .B(new_n4584), .Y(new_n4587));
  xnor_4 g02239(.A(new_n4582), .B(new_n4581), .Y(new_n4588_1));
  nor_5  g02240(.A(new_n4588_1), .B(new_n4587), .Y(new_n4589));
  nor_5  g02241(.A(new_n4589), .B(new_n4583), .Y(new_n4590_1));
  not_8  g02242(.A(new_n4579), .Y(new_n4591));
  xnor_4 g02243(.A(new_n4591), .B(new_n4577), .Y(new_n4592));
  and_5  g02244(.A(new_n4592), .B(new_n4590_1), .Y(new_n4593));
  nor_5  g02245(.A(new_n4593), .B(new_n4580), .Y(new_n4594));
  and_5  g02246(.A(new_n4594), .B(new_n4576), .Y(new_n4595_1));
  nor_5  g02247(.A(new_n4595_1), .B(new_n4574), .Y(new_n4596));
  nor_5  g02248(.A(new_n4596), .B(new_n4571), .Y(new_n4597));
  nor_5  g02249(.A(new_n4597), .B(new_n4570), .Y(new_n4598));
  nor_5  g02250(.A(new_n4598), .B(new_n4566), .Y(new_n4599));
  nor_5  g02251(.A(new_n4599), .B(new_n4565), .Y(new_n4600));
  nor_5  g02252(.A(new_n4600), .B(new_n4561), .Y(new_n4601));
  nor_5  g02253(.A(new_n4601), .B(new_n4560), .Y(new_n4602));
  nor_5  g02254(.A(new_n4602), .B(new_n4556), .Y(new_n4603));
  nor_5  g02255(.A(new_n4603), .B(new_n4555), .Y(new_n4604));
  nor_5  g02256(.A(new_n4604), .B(new_n4551), .Y(new_n4605));
  nor_5  g02257(.A(new_n4605), .B(new_n4550), .Y(new_n4606));
  nor_5  g02258(.A(new_n4606), .B(new_n4546), .Y(new_n4607));
  nor_5  g02259(.A(new_n4607), .B(new_n4545), .Y(new_n4608));
  nor_5  g02260(.A(new_n4608), .B(new_n4541), .Y(new_n4609));
  nor_5  g02261(.A(new_n4609), .B(new_n4540), .Y(new_n4610));
  not_8  g02262(.A(new_n4610), .Y(new_n4611));
  xnor_4 g02263(.A(new_n4611), .B(new_n4534), .Y(n298));
  xnor_4 g02264(.A(n21735), .B(n20604), .Y(new_n4613));
  not_8  g02265(.A(n16158), .Y(new_n4614));
  and_5  g02266(.A(n24085), .B(new_n4614), .Y(new_n4615));
  xnor_4 g02267(.A(n24085), .B(n16158), .Y(new_n4616));
  not_8  g02268(.A(n5752), .Y(new_n4617));
  and_5  g02269(.A(n14071), .B(new_n4617), .Y(new_n4618));
  xnor_4 g02270(.A(n14071), .B(n5752), .Y(new_n4619));
  not_8  g02271(.A(n18171), .Y(new_n4620));
  nor_5  g02272(.A(new_n4620), .B(n1738), .Y(new_n4621));
  and_5  g02273(.A(new_n4620), .B(n1738), .Y(new_n4622));
  not_8  g02274(.A(n25073), .Y(new_n4623));
  nor_5  g02275(.A(new_n4623), .B(n12152), .Y(new_n4624_1));
  nand_5 g02276(.A(new_n4623), .B(n12152), .Y(new_n4625));
  not_8  g02277(.A(n22309), .Y(new_n4626));
  nor_5  g02278(.A(new_n4626), .B(n19107), .Y(new_n4627));
  and_5  g02279(.A(new_n4627), .B(new_n4625), .Y(new_n4628));
  nor_5  g02280(.A(new_n4628), .B(new_n4624_1), .Y(new_n4629));
  nor_5  g02281(.A(new_n4629), .B(new_n4622), .Y(new_n4630));
  nor_5  g02282(.A(new_n4630), .B(new_n4621), .Y(new_n4631));
  and_5  g02283(.A(new_n4631), .B(new_n4619), .Y(new_n4632));
  or_5   g02284(.A(new_n4632), .B(new_n4618), .Y(new_n4633));
  and_5  g02285(.A(new_n4633), .B(new_n4616), .Y(new_n4634));
  or_5   g02286(.A(new_n4634), .B(new_n4615), .Y(new_n4635));
  xor_4  g02287(.A(new_n4635), .B(new_n4613), .Y(new_n4636));
  xnor_4 g02288(.A(n4119), .B(n1525), .Y(new_n4637));
  not_8  g02289(.A(n16988), .Y(new_n4638));
  nor_5  g02290(.A(new_n4638), .B(n14510), .Y(new_n4639));
  xnor_4 g02291(.A(n16988), .B(n14510), .Y(new_n4640));
  not_8  g02292(.A(n21779), .Y(new_n4641));
  nor_5  g02293(.A(new_n4641), .B(n13263), .Y(new_n4642));
  xnor_4 g02294(.A(n21779), .B(n13263), .Y(new_n4643));
  nor_5  g02295(.A(new_n3446), .B(n5376), .Y(new_n4644));
  not_8  g02296(.A(n5376), .Y(new_n4645));
  nor_5  g02297(.A(n20455), .B(new_n4645), .Y(new_n4646_1));
  nor_5  g02298(.A(n5128), .B(new_n3448), .Y(new_n4647));
  not_8  g02299(.A(n5128), .Y(new_n4648));
  nor_5  g02300(.A(new_n4648), .B(n1639), .Y(new_n4649));
  nor_5  g02301(.A(n23120), .B(new_n3451_1), .Y(new_n4650));
  not_8  g02302(.A(new_n4650), .Y(new_n4651));
  nor_5  g02303(.A(new_n4651), .B(new_n4649), .Y(new_n4652));
  nor_5  g02304(.A(new_n4652), .B(new_n4647), .Y(new_n4653));
  nor_5  g02305(.A(new_n4653), .B(new_n4646_1), .Y(new_n4654));
  nor_5  g02306(.A(new_n4654), .B(new_n4644), .Y(new_n4655));
  and_5  g02307(.A(new_n4655), .B(new_n4643), .Y(new_n4656));
  or_5   g02308(.A(new_n4656), .B(new_n4642), .Y(new_n4657));
  and_5  g02309(.A(new_n4657), .B(new_n4640), .Y(new_n4658));
  or_5   g02310(.A(new_n4658), .B(new_n4639), .Y(new_n4659));
  xor_4  g02311(.A(new_n4659), .B(new_n4637), .Y(new_n4660));
  xnor_4 g02312(.A(n12626), .B(n4272), .Y(new_n4661));
  not_8  g02313(.A(n24319), .Y(new_n4662));
  nor_5  g02314(.A(new_n4662), .B(n6971), .Y(new_n4663));
  xnor_4 g02315(.A(n24319), .B(n6971), .Y(new_n4664));
  not_8  g02316(.A(n7460), .Y(new_n4665_1));
  nor_5  g02317(.A(n22068), .B(new_n4665_1), .Y(new_n4666));
  xnor_4 g02318(.A(n22068), .B(n7460), .Y(new_n4667));
  not_8  g02319(.A(n196), .Y(new_n4668));
  and_5  g02320(.A(n9460), .B(new_n4668), .Y(new_n4669));
  nor_5  g02321(.A(n9460), .B(new_n4668), .Y(new_n4670));
  not_8  g02322(.A(n11749), .Y(new_n4671));
  and_5  g02323(.A(n14954), .B(new_n4671), .Y(new_n4672));
  nor_5  g02324(.A(n14954), .B(new_n4671), .Y(new_n4673));
  not_8  g02325(.A(n23831), .Y(new_n4674_1));
  nor_5  g02326(.A(new_n4674_1), .B(n13424), .Y(new_n4675));
  not_8  g02327(.A(new_n4675), .Y(new_n4676));
  nor_5  g02328(.A(new_n4676), .B(new_n4673), .Y(new_n4677));
  nor_5  g02329(.A(new_n4677), .B(new_n4672), .Y(new_n4678));
  nor_5  g02330(.A(new_n4678), .B(new_n4670), .Y(new_n4679));
  nor_5  g02331(.A(new_n4679), .B(new_n4669), .Y(new_n4680));
  and_5  g02332(.A(new_n4680), .B(new_n4667), .Y(new_n4681));
  or_5   g02333(.A(new_n4681), .B(new_n4666), .Y(new_n4682));
  and_5  g02334(.A(new_n4682), .B(new_n4664), .Y(new_n4683));
  or_5   g02335(.A(new_n4683), .B(new_n4663), .Y(new_n4684));
  xor_4  g02336(.A(new_n4684), .B(new_n4661), .Y(new_n4685));
  xnor_4 g02337(.A(new_n4685), .B(new_n4660), .Y(new_n4686));
  xor_4  g02338(.A(new_n4657), .B(new_n4640), .Y(new_n4687));
  xor_4  g02339(.A(new_n4682), .B(new_n4664), .Y(new_n4688));
  and_5  g02340(.A(new_n4688), .B(new_n4687), .Y(new_n4689));
  xor_4  g02341(.A(new_n4688), .B(new_n4687), .Y(new_n4690));
  xnor_4 g02342(.A(new_n4655), .B(new_n4643), .Y(new_n4691));
  not_8  g02343(.A(new_n4691), .Y(new_n4692));
  xnor_4 g02344(.A(new_n4680), .B(new_n4667), .Y(new_n4693_1));
  not_8  g02345(.A(new_n4693_1), .Y(new_n4694));
  nor_5  g02346(.A(new_n4694), .B(new_n4692), .Y(new_n4695));
  xnor_4 g02347(.A(new_n4694), .B(new_n4692), .Y(new_n4696));
  xnor_4 g02348(.A(n20455), .B(n5376), .Y(new_n4697));
  xnor_4 g02349(.A(new_n4697), .B(new_n4653), .Y(new_n4698));
  not_8  g02350(.A(new_n4698), .Y(new_n4699));
  xnor_4 g02351(.A(n9460), .B(n196), .Y(new_n4700));
  xnor_4 g02352(.A(new_n4700), .B(new_n4678), .Y(new_n4701));
  not_8  g02353(.A(new_n4701), .Y(new_n4702));
  nor_5  g02354(.A(new_n4702), .B(new_n4699), .Y(new_n4703));
  xnor_4 g02355(.A(new_n4701), .B(new_n4699), .Y(new_n4704));
  xnor_4 g02356(.A(n5128), .B(n1639), .Y(new_n4705));
  xnor_4 g02357(.A(new_n4705), .B(new_n4651), .Y(new_n4706));
  xnor_4 g02358(.A(n14954), .B(n11749), .Y(new_n4707));
  xnor_4 g02359(.A(new_n4707), .B(new_n4676), .Y(new_n4708));
  nor_5  g02360(.A(new_n4708), .B(new_n4706), .Y(new_n4709));
  xnor_4 g02361(.A(n23120), .B(n16968), .Y(new_n4710));
  xnor_4 g02362(.A(n23831), .B(n13424), .Y(new_n4711));
  nor_5  g02363(.A(new_n4711), .B(new_n4710), .Y(new_n4712));
  not_8  g02364(.A(new_n4706), .Y(new_n4713));
  xnor_4 g02365(.A(new_n4708), .B(new_n4713), .Y(new_n4714));
  and_5  g02366(.A(new_n4714), .B(new_n4712), .Y(new_n4715));
  nor_5  g02367(.A(new_n4715), .B(new_n4709), .Y(new_n4716));
  and_5  g02368(.A(new_n4716), .B(new_n4704), .Y(new_n4717));
  nor_5  g02369(.A(new_n4717), .B(new_n4703), .Y(new_n4718));
  nor_5  g02370(.A(new_n4718), .B(new_n4696), .Y(new_n4719));
  nor_5  g02371(.A(new_n4719), .B(new_n4695), .Y(new_n4720));
  and_5  g02372(.A(new_n4720), .B(new_n4690), .Y(new_n4721));
  nor_5  g02373(.A(new_n4721), .B(new_n4689), .Y(new_n4722_1));
  xnor_4 g02374(.A(new_n4722_1), .B(new_n4686), .Y(new_n4723));
  xnor_4 g02375(.A(new_n4723), .B(new_n4636), .Y(new_n4724));
  xor_4  g02376(.A(new_n4633), .B(new_n4616), .Y(new_n4725));
  xor_4  g02377(.A(new_n4720), .B(new_n4690), .Y(new_n4726));
  nor_5  g02378(.A(new_n4726), .B(new_n4725), .Y(new_n4727));
  xnor_4 g02379(.A(new_n4726), .B(new_n4725), .Y(new_n4728));
  xnor_4 g02380(.A(new_n4718), .B(new_n4696), .Y(new_n4729));
  not_8  g02381(.A(new_n4729), .Y(new_n4730));
  xnor_4 g02382(.A(new_n4631), .B(new_n4619), .Y(new_n4731_1));
  and_5  g02383(.A(new_n4731_1), .B(new_n4730), .Y(new_n4732));
  xnor_4 g02384(.A(new_n4716), .B(new_n4704), .Y(new_n4733));
  not_8  g02385(.A(new_n4733), .Y(new_n4734));
  xnor_4 g02386(.A(n18171), .B(n1738), .Y(new_n4735));
  xnor_4 g02387(.A(new_n4735), .B(new_n4629), .Y(new_n4736));
  and_5  g02388(.A(new_n4736), .B(new_n4734), .Y(new_n4737));
  xnor_4 g02389(.A(new_n4736), .B(new_n4734), .Y(new_n4738));
  xnor_4 g02390(.A(n22309), .B(n19107), .Y(new_n4739));
  xnor_4 g02391(.A(new_n4711), .B(new_n4710), .Y(new_n4740));
  nor_5  g02392(.A(new_n4740), .B(new_n4739), .Y(new_n4741));
  xnor_4 g02393(.A(n25073), .B(n12152), .Y(new_n4742));
  xnor_4 g02394(.A(new_n4742), .B(new_n4627), .Y(new_n4743));
  nor_5  g02395(.A(new_n4743), .B(new_n4741), .Y(new_n4744));
  xnor_4 g02396(.A(new_n4714), .B(new_n4712), .Y(new_n4745_1));
  not_8  g02397(.A(new_n4745_1), .Y(new_n4746));
  xnor_4 g02398(.A(new_n4743), .B(new_n4741), .Y(new_n4747_1));
  nor_5  g02399(.A(new_n4747_1), .B(new_n4746), .Y(new_n4748));
  nor_5  g02400(.A(new_n4748), .B(new_n4744), .Y(new_n4749));
  nor_5  g02401(.A(new_n4749), .B(new_n4738), .Y(new_n4750));
  nor_5  g02402(.A(new_n4750), .B(new_n4737), .Y(new_n4751));
  xnor_4 g02403(.A(new_n4731_1), .B(new_n4730), .Y(new_n4752));
  nor_5  g02404(.A(new_n4752), .B(new_n4751), .Y(new_n4753));
  nor_5  g02405(.A(new_n4753), .B(new_n4732), .Y(new_n4754));
  nor_5  g02406(.A(new_n4754), .B(new_n4728), .Y(new_n4755));
  nor_5  g02407(.A(new_n4755), .B(new_n4727), .Y(new_n4756));
  xor_4  g02408(.A(new_n4756), .B(new_n4724), .Y(n317));
  nor_5  g02409(.A(n9934), .B(n3506), .Y(new_n4758));
  xnor_4 g02410(.A(n9934), .B(n3506), .Y(new_n4759));
  nor_5  g02411(.A(n18496), .B(n14899), .Y(new_n4760));
  xnor_4 g02412(.A(n18496), .B(n14899), .Y(new_n4761));
  nor_5  g02413(.A(n26224), .B(n18444), .Y(new_n4762));
  xnor_4 g02414(.A(n26224), .B(n18444), .Y(new_n4763));
  nor_5  g02415(.A(n24638), .B(n19327), .Y(new_n4764));
  xnor_4 g02416(.A(n24638), .B(n19327), .Y(new_n4765));
  nor_5  g02417(.A(n22597), .B(n21674), .Y(new_n4766_1));
  xnor_4 g02418(.A(n22597), .B(n21674), .Y(new_n4767));
  nor_5  g02419(.A(n26107), .B(n17251), .Y(new_n4768));
  xnor_4 g02420(.A(n26107), .B(n17251), .Y(new_n4769));
  nor_5  g02421(.A(n14790), .B(n342), .Y(new_n4770_1));
  xnor_4 g02422(.A(n14790), .B(n342), .Y(new_n4771));
  nor_5  g02423(.A(n26553), .B(n10096), .Y(new_n4772));
  xnor_4 g02424(.A(n26553), .B(new_n3555_1), .Y(new_n4773));
  nor_5  g02425(.A(n16994), .B(n4964), .Y(new_n4774));
  nor_5  g02426(.A(new_n3562), .B(new_n3755_1), .Y(new_n4775));
  not_8  g02427(.A(n4964), .Y(new_n4776));
  xnor_4 g02428(.A(n16994), .B(new_n4776), .Y(new_n4777_1));
  not_8  g02429(.A(new_n4777_1), .Y(new_n4778));
  nor_5  g02430(.A(new_n4778), .B(new_n4775), .Y(new_n4779));
  or_5   g02431(.A(new_n4779), .B(new_n4774), .Y(new_n4780));
  and_5  g02432(.A(new_n4780), .B(new_n4773), .Y(new_n4781));
  nor_5  g02433(.A(new_n4781), .B(new_n4772), .Y(new_n4782));
  nor_5  g02434(.A(new_n4782), .B(new_n4771), .Y(new_n4783));
  nor_5  g02435(.A(new_n4783), .B(new_n4770_1), .Y(new_n4784));
  nor_5  g02436(.A(new_n4784), .B(new_n4769), .Y(new_n4785_1));
  nor_5  g02437(.A(new_n4785_1), .B(new_n4768), .Y(new_n4786));
  nor_5  g02438(.A(new_n4786), .B(new_n4767), .Y(new_n4787));
  nor_5  g02439(.A(new_n4787), .B(new_n4766_1), .Y(new_n4788));
  nor_5  g02440(.A(new_n4788), .B(new_n4765), .Y(new_n4789));
  nor_5  g02441(.A(new_n4789), .B(new_n4764), .Y(new_n4790));
  nor_5  g02442(.A(new_n4790), .B(new_n4763), .Y(new_n4791));
  nor_5  g02443(.A(new_n4791), .B(new_n4762), .Y(new_n4792));
  nor_5  g02444(.A(new_n4792), .B(new_n4761), .Y(new_n4793));
  nor_5  g02445(.A(new_n4793), .B(new_n4760), .Y(new_n4794));
  nor_5  g02446(.A(new_n4794), .B(new_n4759), .Y(new_n4795));
  nor_5  g02447(.A(new_n4795), .B(new_n4758), .Y(new_n4796));
  not_8  g02448(.A(n9259), .Y(new_n4797));
  not_8  g02449(.A(n2979), .Y(new_n4798));
  xnor_4 g02450(.A(n9554), .B(new_n4798), .Y(new_n4799));
  nor_5  g02451(.A(n26408), .B(n647), .Y(new_n4800));
  not_8  g02452(.A(n647), .Y(new_n4801));
  xnor_4 g02453(.A(n26408), .B(new_n4801), .Y(new_n4802));
  nor_5  g02454(.A(n20409), .B(n18227), .Y(new_n4803));
  not_8  g02455(.A(n18227), .Y(new_n4804_1));
  xnor_4 g02456(.A(n20409), .B(new_n4804_1), .Y(new_n4805));
  nor_5  g02457(.A(n25749), .B(n7377), .Y(new_n4806));
  not_8  g02458(.A(n7377), .Y(new_n4807));
  xnor_4 g02459(.A(n25749), .B(new_n4807), .Y(new_n4808));
  nor_5  g02460(.A(n11630), .B(n3161), .Y(new_n4809));
  xnor_4 g02461(.A(n11630), .B(new_n3774), .Y(new_n4810_1));
  nor_5  g02462(.A(n13453), .B(n9003), .Y(new_n4811));
  xnor_4 g02463(.A(n13453), .B(new_n3778), .Y(new_n4812_1));
  nor_5  g02464(.A(n7421), .B(n4957), .Y(new_n4813));
  xnor_4 g02465(.A(n7421), .B(new_n3784), .Y(new_n4814_1));
  nor_5  g02466(.A(n19680), .B(n7524), .Y(new_n4815));
  xnor_4 g02467(.A(n19680), .B(new_n3788), .Y(new_n4816));
  nor_5  g02468(.A(n15743), .B(n2809), .Y(new_n4817));
  not_8  g02469(.A(n15508), .Y(new_n4818));
  nor_5  g02470(.A(new_n3798), .B(new_n4818), .Y(new_n4819));
  xnor_4 g02471(.A(n15743), .B(n2809), .Y(new_n4820));
  nor_5  g02472(.A(new_n4820), .B(new_n4819), .Y(new_n4821));
  or_5   g02473(.A(new_n4821), .B(new_n4817), .Y(new_n4822));
  and_5  g02474(.A(new_n4822), .B(new_n4816), .Y(new_n4823));
  or_5   g02475(.A(new_n4823), .B(new_n4815), .Y(new_n4824));
  and_5  g02476(.A(new_n4824), .B(new_n4814_1), .Y(new_n4825));
  or_5   g02477(.A(new_n4825), .B(new_n4813), .Y(new_n4826));
  and_5  g02478(.A(new_n4826), .B(new_n4812_1), .Y(new_n4827));
  or_5   g02479(.A(new_n4827), .B(new_n4811), .Y(new_n4828));
  and_5  g02480(.A(new_n4828), .B(new_n4810_1), .Y(new_n4829));
  or_5   g02481(.A(new_n4829), .B(new_n4809), .Y(new_n4830));
  and_5  g02482(.A(new_n4830), .B(new_n4808), .Y(new_n4831));
  or_5   g02483(.A(new_n4831), .B(new_n4806), .Y(new_n4832));
  and_5  g02484(.A(new_n4832), .B(new_n4805), .Y(new_n4833));
  or_5   g02485(.A(new_n4833), .B(new_n4803), .Y(new_n4834));
  and_5  g02486(.A(new_n4834), .B(new_n4802), .Y(new_n4835));
  nor_5  g02487(.A(new_n4835), .B(new_n4800), .Y(new_n4836));
  xnor_4 g02488(.A(new_n4836), .B(new_n4799), .Y(new_n4837));
  nor_5  g02489(.A(new_n4837), .B(new_n4797), .Y(new_n4838));
  not_8  g02490(.A(new_n4837), .Y(new_n4839));
  xnor_4 g02491(.A(new_n4839), .B(new_n4797), .Y(new_n4840));
  xor_4  g02492(.A(new_n4834), .B(new_n4802), .Y(new_n4841));
  nor_5  g02493(.A(new_n4841), .B(new_n3583), .Y(new_n4842));
  xnor_4 g02494(.A(new_n4841), .B(new_n3583), .Y(new_n4843));
  not_8  g02495(.A(n20213), .Y(new_n4844));
  xor_4  g02496(.A(new_n4832), .B(new_n4805), .Y(new_n4845));
  nor_5  g02497(.A(new_n4845), .B(new_n4844), .Y(new_n4846));
  xnor_4 g02498(.A(new_n4845), .B(new_n4844), .Y(new_n4847));
  not_8  g02499(.A(n13912), .Y(new_n4848));
  nor_5  g02500(.A(new_n4829), .B(new_n4809), .Y(new_n4849));
  xnor_4 g02501(.A(new_n4849), .B(new_n4808), .Y(new_n4850_1));
  nor_5  g02502(.A(new_n4850_1), .B(new_n4848), .Y(new_n4851));
  xnor_4 g02503(.A(new_n4850_1), .B(new_n4848), .Y(new_n4852));
  not_8  g02504(.A(n7670), .Y(new_n4853));
  xor_4  g02505(.A(new_n4828), .B(new_n4810_1), .Y(new_n4854));
  nor_5  g02506(.A(new_n4854), .B(new_n4853), .Y(new_n4855));
  xnor_4 g02507(.A(new_n4854), .B(new_n4853), .Y(new_n4856));
  not_8  g02508(.A(n9598), .Y(new_n4857));
  nor_5  g02509(.A(new_n4825), .B(new_n4813), .Y(new_n4858_1));
  xnor_4 g02510(.A(new_n4858_1), .B(new_n4812_1), .Y(new_n4859));
  nor_5  g02511(.A(new_n4859), .B(new_n4857), .Y(new_n4860));
  not_8  g02512(.A(new_n4859), .Y(new_n4861));
  xnor_4 g02513(.A(new_n4861), .B(n9598), .Y(new_n4862));
  not_8  g02514(.A(n22290), .Y(new_n4863));
  xor_4  g02515(.A(new_n4824), .B(new_n4814_1), .Y(new_n4864));
  nor_5  g02516(.A(new_n4864), .B(new_n4863), .Y(new_n4865));
  xnor_4 g02517(.A(new_n4864), .B(new_n4863), .Y(new_n4866));
  not_8  g02518(.A(n11273), .Y(new_n4867));
  nor_5  g02519(.A(new_n4821), .B(new_n4817), .Y(new_n4868));
  xnor_4 g02520(.A(new_n4868), .B(new_n4816), .Y(new_n4869));
  nor_5  g02521(.A(new_n4869), .B(new_n4867), .Y(new_n4870));
  xor_4  g02522(.A(new_n4820), .B(new_n4819), .Y(new_n4871));
  not_8  g02523(.A(new_n4871), .Y(new_n4872));
  nor_5  g02524(.A(new_n4872), .B(n25565), .Y(new_n4873));
  xnor_4 g02525(.A(n20658), .B(n15508), .Y(new_n4874));
  nor_5  g02526(.A(new_n4874), .B(new_n3635), .Y(new_n4875));
  xnor_4 g02527(.A(new_n4872), .B(n25565), .Y(new_n4876));
  nor_5  g02528(.A(new_n4876), .B(new_n4875), .Y(new_n4877));
  nor_5  g02529(.A(new_n4877), .B(new_n4873), .Y(new_n4878));
  not_8  g02530(.A(new_n4878), .Y(new_n4879));
  not_8  g02531(.A(new_n4869), .Y(new_n4880));
  xnor_4 g02532(.A(new_n4880), .B(n11273), .Y(new_n4881));
  nor_5  g02533(.A(new_n4881), .B(new_n4879), .Y(new_n4882));
  nor_5  g02534(.A(new_n4882), .B(new_n4870), .Y(new_n4883));
  nor_5  g02535(.A(new_n4883), .B(new_n4866), .Y(new_n4884));
  nor_5  g02536(.A(new_n4884), .B(new_n4865), .Y(new_n4885));
  nor_5  g02537(.A(new_n4885), .B(new_n4862), .Y(new_n4886));
  nor_5  g02538(.A(new_n4886), .B(new_n4860), .Y(new_n4887));
  nor_5  g02539(.A(new_n4887), .B(new_n4856), .Y(new_n4888));
  nor_5  g02540(.A(new_n4888), .B(new_n4855), .Y(new_n4889));
  nor_5  g02541(.A(new_n4889), .B(new_n4852), .Y(new_n4890));
  nor_5  g02542(.A(new_n4890), .B(new_n4851), .Y(new_n4891_1));
  nor_5  g02543(.A(new_n4891_1), .B(new_n4847), .Y(new_n4892));
  nor_5  g02544(.A(new_n4892), .B(new_n4846), .Y(new_n4893));
  nor_5  g02545(.A(new_n4893), .B(new_n4843), .Y(new_n4894));
  or_5   g02546(.A(new_n4894), .B(new_n4842), .Y(new_n4895));
  and_5  g02547(.A(new_n4895), .B(new_n4840), .Y(new_n4896));
  nor_5  g02548(.A(new_n4896), .B(new_n4838), .Y(new_n4897));
  nor_5  g02549(.A(n9554), .B(n2979), .Y(new_n4898));
  or_5   g02550(.A(new_n4835), .B(new_n4800), .Y(new_n4899));
  and_5  g02551(.A(new_n4899), .B(new_n4799), .Y(new_n4900));
  nor_5  g02552(.A(new_n4900), .B(new_n4898), .Y(new_n4901));
  xnor_4 g02553(.A(new_n4901), .B(new_n4897), .Y(new_n4902));
  nor_5  g02554(.A(new_n4894), .B(new_n4842), .Y(new_n4903));
  xnor_4 g02555(.A(new_n4903), .B(new_n4840), .Y(new_n4904));
  not_8  g02556(.A(new_n4904), .Y(new_n4905));
  nor_5  g02557(.A(new_n4905), .B(n3740), .Y(new_n4906));
  not_8  g02558(.A(n3740), .Y(new_n4907));
  xnor_4 g02559(.A(new_n4905), .B(new_n4907), .Y(new_n4908));
  not_8  g02560(.A(n2858), .Y(new_n4909));
  xor_4  g02561(.A(new_n4893), .B(new_n4843), .Y(new_n4910));
  nor_5  g02562(.A(new_n4910), .B(new_n4909), .Y(new_n4911));
  xnor_4 g02563(.A(new_n4910), .B(new_n4909), .Y(new_n4912));
  not_8  g02564(.A(n2659), .Y(new_n4913_1));
  xor_4  g02565(.A(new_n4891_1), .B(new_n4847), .Y(new_n4914));
  nor_5  g02566(.A(new_n4914), .B(new_n4913_1), .Y(new_n4915));
  xnor_4 g02567(.A(new_n4914), .B(new_n4913_1), .Y(new_n4916));
  not_8  g02568(.A(n24327), .Y(new_n4917));
  xor_4  g02569(.A(new_n4889), .B(new_n4852), .Y(new_n4918));
  nor_5  g02570(.A(new_n4918), .B(new_n4917), .Y(new_n4919));
  not_8  g02571(.A(new_n4918), .Y(new_n4920));
  xnor_4 g02572(.A(new_n4920), .B(n24327), .Y(new_n4921));
  not_8  g02573(.A(n22198), .Y(new_n4922));
  xor_4  g02574(.A(new_n4887), .B(new_n4856), .Y(new_n4923));
  nor_5  g02575(.A(new_n4923), .B(new_n4922), .Y(new_n4924));
  not_8  g02576(.A(new_n4923), .Y(new_n4925_1));
  xnor_4 g02577(.A(new_n4925_1), .B(n22198), .Y(new_n4926));
  not_8  g02578(.A(n20826), .Y(new_n4927));
  xor_4  g02579(.A(new_n4885), .B(new_n4862), .Y(new_n4928));
  nor_5  g02580(.A(new_n4928), .B(new_n4927), .Y(new_n4929));
  not_8  g02581(.A(new_n4928), .Y(new_n4930));
  xnor_4 g02582(.A(new_n4930), .B(n20826), .Y(new_n4931));
  not_8  g02583(.A(n7305), .Y(new_n4932));
  xor_4  g02584(.A(new_n4883), .B(new_n4866), .Y(new_n4933));
  nor_5  g02585(.A(new_n4933), .B(new_n4932), .Y(new_n4934));
  xnor_4 g02586(.A(new_n4881), .B(new_n4878), .Y(new_n4935));
  not_8  g02587(.A(new_n4935), .Y(new_n4936));
  nor_5  g02588(.A(new_n4936), .B(n25872), .Y(new_n4937));
  xnor_4 g02589(.A(new_n4935), .B(n25872), .Y(new_n4938));
  not_8  g02590(.A(n20259), .Y(new_n4939_1));
  xnor_4 g02591(.A(new_n4876), .B(new_n4875), .Y(new_n4940));
  nor_5  g02592(.A(new_n4940), .B(new_n4939_1), .Y(new_n4941));
  xnor_4 g02593(.A(new_n4874), .B(n21993), .Y(new_n4942));
  not_8  g02594(.A(new_n4942), .Y(new_n4943));
  nor_5  g02595(.A(new_n4943), .B(n3925), .Y(new_n4944));
  xnor_4 g02596(.A(new_n4940), .B(new_n4939_1), .Y(new_n4945));
  nor_5  g02597(.A(new_n4945), .B(new_n4944), .Y(new_n4946));
  nor_5  g02598(.A(new_n4946), .B(new_n4941), .Y(new_n4947_1));
  and_5  g02599(.A(new_n4947_1), .B(new_n4938), .Y(new_n4948));
  nor_5  g02600(.A(new_n4948), .B(new_n4937), .Y(new_n4949));
  not_8  g02601(.A(new_n4933), .Y(new_n4950));
  xnor_4 g02602(.A(new_n4950), .B(new_n4932), .Y(new_n4951));
  and_5  g02603(.A(new_n4951), .B(new_n4949), .Y(new_n4952_1));
  nor_5  g02604(.A(new_n4952_1), .B(new_n4934), .Y(new_n4953));
  nor_5  g02605(.A(new_n4953), .B(new_n4931), .Y(new_n4954));
  nor_5  g02606(.A(new_n4954), .B(new_n4929), .Y(new_n4955));
  nor_5  g02607(.A(new_n4955), .B(new_n4926), .Y(new_n4956));
  nor_5  g02608(.A(new_n4956), .B(new_n4924), .Y(new_n4957_1));
  nor_5  g02609(.A(new_n4957_1), .B(new_n4921), .Y(new_n4958));
  nor_5  g02610(.A(new_n4958), .B(new_n4919), .Y(new_n4959));
  nor_5  g02611(.A(new_n4959), .B(new_n4916), .Y(new_n4960));
  nor_5  g02612(.A(new_n4960), .B(new_n4915), .Y(new_n4961));
  nor_5  g02613(.A(new_n4961), .B(new_n4912), .Y(new_n4962));
  nor_5  g02614(.A(new_n4962), .B(new_n4911), .Y(new_n4963));
  and_5  g02615(.A(new_n4963), .B(new_n4908), .Y(new_n4964_1));
  nor_5  g02616(.A(new_n4964_1), .B(new_n4906), .Y(new_n4965));
  xnor_4 g02617(.A(new_n4965), .B(new_n4902), .Y(new_n4966_1));
  xor_4  g02618(.A(new_n4966_1), .B(new_n4796), .Y(new_n4967_1));
  xnor_4 g02619(.A(new_n4794), .B(new_n4759), .Y(new_n4968));
  xnor_4 g02620(.A(new_n4963), .B(new_n4908), .Y(new_n4969));
  nor_5  g02621(.A(new_n4969), .B(new_n4968), .Y(new_n4970));
  xnor_4 g02622(.A(new_n4969), .B(new_n4968), .Y(new_n4971));
  xnor_4 g02623(.A(new_n4792), .B(new_n4761), .Y(new_n4972_1));
  xor_4  g02624(.A(new_n4961), .B(new_n4912), .Y(new_n4973));
  nor_5  g02625(.A(new_n4973), .B(new_n4972_1), .Y(new_n4974));
  xnor_4 g02626(.A(new_n4973), .B(new_n4972_1), .Y(new_n4975));
  xnor_4 g02627(.A(new_n4790), .B(new_n4763), .Y(new_n4976));
  xor_4  g02628(.A(new_n4959), .B(new_n4916), .Y(new_n4977));
  nor_5  g02629(.A(new_n4977), .B(new_n4976), .Y(new_n4978));
  xnor_4 g02630(.A(new_n4977), .B(new_n4976), .Y(new_n4979));
  xnor_4 g02631(.A(new_n4788), .B(new_n4765), .Y(new_n4980));
  xor_4  g02632(.A(new_n4957_1), .B(new_n4921), .Y(new_n4981));
  nor_5  g02633(.A(new_n4981), .B(new_n4980), .Y(new_n4982));
  xnor_4 g02634(.A(new_n4981), .B(new_n4980), .Y(new_n4983));
  xnor_4 g02635(.A(new_n4786), .B(new_n4767), .Y(new_n4984));
  xor_4  g02636(.A(new_n4955), .B(new_n4926), .Y(new_n4985));
  nor_5  g02637(.A(new_n4985), .B(new_n4984), .Y(new_n4986));
  xnor_4 g02638(.A(new_n4985), .B(new_n4984), .Y(new_n4987));
  xnor_4 g02639(.A(new_n4784), .B(new_n4769), .Y(new_n4988));
  xor_4  g02640(.A(new_n4953), .B(new_n4931), .Y(new_n4989));
  nor_5  g02641(.A(new_n4989), .B(new_n4988), .Y(new_n4990));
  xnor_4 g02642(.A(new_n4989), .B(new_n4988), .Y(new_n4991));
  xnor_4 g02643(.A(new_n4782), .B(new_n4771), .Y(new_n4992));
  xor_4  g02644(.A(new_n4951), .B(new_n4949), .Y(new_n4993));
  nor_5  g02645(.A(new_n4993), .B(new_n4992), .Y(new_n4994));
  xnor_4 g02646(.A(new_n4993), .B(new_n4992), .Y(new_n4995));
  xnor_4 g02647(.A(new_n4947_1), .B(new_n4938), .Y(new_n4996));
  nor_5  g02648(.A(new_n4779), .B(new_n4774), .Y(new_n4997));
  xnor_4 g02649(.A(new_n4997), .B(new_n4773), .Y(new_n4998));
  not_8  g02650(.A(new_n4998), .Y(new_n4999));
  nor_5  g02651(.A(new_n4999), .B(new_n4996), .Y(new_n5000));
  xnor_4 g02652(.A(new_n4998), .B(new_n4996), .Y(new_n5001));
  not_8  g02653(.A(n3925), .Y(new_n5002));
  xnor_4 g02654(.A(new_n4943), .B(new_n5002), .Y(new_n5003));
  xnor_4 g02655(.A(n9246), .B(n7876), .Y(new_n5004));
  nor_5  g02656(.A(new_n5004), .B(new_n5003), .Y(new_n5005));
  and_5  g02657(.A(new_n5005), .B(new_n4777_1), .Y(new_n5006));
  xor_4  g02658(.A(new_n4945), .B(new_n4944), .Y(new_n5007));
  xnor_4 g02659(.A(new_n4778), .B(new_n4775), .Y(new_n5008));
  nor_5  g02660(.A(new_n5008), .B(new_n5005), .Y(new_n5009));
  nor_5  g02661(.A(new_n5009), .B(new_n5006), .Y(new_n5010));
  and_5  g02662(.A(new_n5010), .B(new_n5007), .Y(new_n5011_1));
  nor_5  g02663(.A(new_n5011_1), .B(new_n5006), .Y(new_n5012));
  and_5  g02664(.A(new_n5012), .B(new_n5001), .Y(new_n5013));
  nor_5  g02665(.A(new_n5013), .B(new_n5000), .Y(new_n5014));
  nor_5  g02666(.A(new_n5014), .B(new_n4995), .Y(new_n5015));
  nor_5  g02667(.A(new_n5015), .B(new_n4994), .Y(new_n5016));
  nor_5  g02668(.A(new_n5016), .B(new_n4991), .Y(new_n5017));
  nor_5  g02669(.A(new_n5017), .B(new_n4990), .Y(new_n5018));
  nor_5  g02670(.A(new_n5018), .B(new_n4987), .Y(new_n5019));
  nor_5  g02671(.A(new_n5019), .B(new_n4986), .Y(new_n5020_1));
  nor_5  g02672(.A(new_n5020_1), .B(new_n4983), .Y(new_n5021));
  nor_5  g02673(.A(new_n5021), .B(new_n4982), .Y(new_n5022));
  nor_5  g02674(.A(new_n5022), .B(new_n4979), .Y(new_n5023));
  nor_5  g02675(.A(new_n5023), .B(new_n4978), .Y(new_n5024_1));
  nor_5  g02676(.A(new_n5024_1), .B(new_n4975), .Y(new_n5025_1));
  nor_5  g02677(.A(new_n5025_1), .B(new_n4974), .Y(new_n5026_1));
  nor_5  g02678(.A(new_n5026_1), .B(new_n4971), .Y(new_n5027));
  nor_5  g02679(.A(new_n5027), .B(new_n4970), .Y(new_n5028));
  xor_4  g02680(.A(new_n5028), .B(new_n4967_1), .Y(n332));
  xnor_4 g02681(.A(n18295), .B(new_n2361_1), .Y(new_n5030));
  nor_5  g02682(.A(n19494), .B(n6502), .Y(new_n5031_1));
  or_5   g02683(.A(new_n2907), .B(new_n3116), .Y(new_n5032));
  not_8  g02684(.A(n6502), .Y(new_n5033));
  xnor_4 g02685(.A(n19494), .B(new_n5033), .Y(new_n5034));
  and_5  g02686(.A(new_n5034), .B(new_n5032), .Y(new_n5035));
  nor_5  g02687(.A(new_n5035), .B(new_n5031_1), .Y(new_n5036));
  xnor_4 g02688(.A(new_n5036), .B(new_n5030), .Y(new_n5037));
  not_8  g02689(.A(new_n5037), .Y(new_n5038));
  xnor_4 g02690(.A(new_n5038), .B(n8381), .Y(new_n5039));
  not_8  g02691(.A(n20235), .Y(new_n5040));
  xnor_4 g02692(.A(n15780), .B(new_n3116), .Y(new_n5041));
  not_8  g02693(.A(new_n5041), .Y(new_n5042));
  nor_5  g02694(.A(new_n5042), .B(n12495), .Y(new_n5043));
  and_5  g02695(.A(new_n5043), .B(new_n5040), .Y(new_n5044));
  xnor_4 g02696(.A(new_n5043), .B(n20235), .Y(new_n5045));
  not_8  g02697(.A(new_n5045), .Y(new_n5046_1));
  nor_5  g02698(.A(new_n2907), .B(new_n3116), .Y(new_n5047));
  xnor_4 g02699(.A(new_n5034), .B(new_n5047), .Y(new_n5048));
  nor_5  g02700(.A(new_n5048), .B(new_n5046_1), .Y(new_n5049));
  nor_5  g02701(.A(new_n5049), .B(new_n5044), .Y(new_n5050));
  xnor_4 g02702(.A(new_n5050), .B(new_n5039), .Y(new_n5051));
  not_8  g02703(.A(new_n5051), .Y(new_n5052));
  not_8  g02704(.A(n23146), .Y(new_n5053));
  nor_5  g02705(.A(n21654), .B(new_n3304), .Y(new_n5054));
  xnor_4 g02706(.A(n25471), .B(n23842), .Y(new_n5055));
  xnor_4 g02707(.A(new_n5055), .B(new_n5054), .Y(new_n5056));
  not_8  g02708(.A(new_n5056), .Y(new_n5057));
  nor_5  g02709(.A(new_n5057), .B(new_n5053), .Y(new_n5058));
  xnor_4 g02710(.A(n21654), .B(new_n3304), .Y(new_n5059));
  and_5  g02711(.A(new_n5059), .B(n17968), .Y(new_n5060_1));
  xnor_4 g02712(.A(new_n5057), .B(n23146), .Y(new_n5061));
  and_5  g02713(.A(new_n5061), .B(new_n5060_1), .Y(new_n5062_1));
  nor_5  g02714(.A(new_n5062_1), .B(new_n5058), .Y(new_n5063));
  not_8  g02715(.A(n3828), .Y(new_n5064_1));
  xnor_4 g02716(.A(n15053), .B(new_n5064_1), .Y(new_n5065));
  not_8  g02717(.A(n25471), .Y(new_n5066));
  nor_5  g02718(.A(new_n5066), .B(n23842), .Y(new_n5067));
  and_5  g02719(.A(new_n5055), .B(new_n5054), .Y(new_n5068));
  nor_5  g02720(.A(new_n5068), .B(new_n5067), .Y(new_n5069));
  xor_4  g02721(.A(new_n5069), .B(new_n5065), .Y(new_n5070));
  xnor_4 g02722(.A(new_n5070), .B(n11184), .Y(new_n5071));
  xnor_4 g02723(.A(new_n5071), .B(new_n5063), .Y(new_n5072));
  xnor_4 g02724(.A(new_n5072), .B(new_n5052), .Y(new_n5073));
  not_8  g02725(.A(new_n5061), .Y(new_n5074));
  xnor_4 g02726(.A(new_n5074), .B(new_n5060_1), .Y(new_n5075));
  not_8  g02727(.A(new_n5048), .Y(new_n5076));
  xnor_4 g02728(.A(new_n5076), .B(new_n5046_1), .Y(new_n5077_1));
  not_8  g02729(.A(new_n5077_1), .Y(new_n5078));
  nor_5  g02730(.A(new_n5078), .B(new_n5075), .Y(new_n5079));
  not_8  g02731(.A(n12495), .Y(new_n5080));
  xnor_4 g02732(.A(new_n5042), .B(new_n5080), .Y(new_n5081));
  xnor_4 g02733(.A(n21654), .B(n16502), .Y(new_n5082_1));
  xnor_4 g02734(.A(new_n5082_1), .B(n17968), .Y(new_n5083));
  not_8  g02735(.A(new_n5083), .Y(new_n5084));
  nor_5  g02736(.A(new_n5084), .B(new_n5081), .Y(new_n5085));
  xnor_4 g02737(.A(new_n5078), .B(new_n5075), .Y(new_n5086));
  nor_5  g02738(.A(new_n5086), .B(new_n5085), .Y(new_n5087));
  nor_5  g02739(.A(new_n5087), .B(new_n5079), .Y(new_n5088));
  xnor_4 g02740(.A(new_n5088), .B(new_n5073), .Y(n357));
  xnor_4 g02741(.A(n22309), .B(new_n2367), .Y(new_n5090));
  nor_5  g02742(.A(new_n4626), .B(new_n2367), .Y(new_n5091));
  xnor_4 g02743(.A(n25073), .B(new_n2363_1), .Y(new_n5092));
  xnor_4 g02744(.A(new_n5092), .B(new_n5091), .Y(new_n5093));
  not_8  g02745(.A(new_n5093), .Y(new_n5094));
  nor_5  g02746(.A(new_n5094), .B(new_n5090), .Y(new_n5095));
  not_8  g02747(.A(new_n5095), .Y(new_n5096));
  xnor_4 g02748(.A(n18171), .B(new_n2359), .Y(new_n5097));
  nor_5  g02749(.A(n25073), .B(n20138), .Y(new_n5098_1));
  or_5   g02750(.A(new_n4626), .B(new_n2367), .Y(new_n5099));
  and_5  g02751(.A(new_n5092), .B(new_n5099), .Y(new_n5100));
  nor_5  g02752(.A(new_n5100), .B(new_n5098_1), .Y(new_n5101_1));
  xnor_4 g02753(.A(new_n5101_1), .B(new_n5097), .Y(new_n5102));
  not_8  g02754(.A(new_n5102), .Y(new_n5103));
  nor_5  g02755(.A(new_n5103), .B(new_n5096), .Y(new_n5104));
  not_8  g02756(.A(new_n5104), .Y(new_n5105));
  not_8  g02757(.A(n3136), .Y(new_n5106));
  xnor_4 g02758(.A(n5752), .B(new_n5106), .Y(new_n5107));
  nor_5  g02759(.A(n18171), .B(n6385), .Y(new_n5108));
  or_5   g02760(.A(new_n5100), .B(new_n5098_1), .Y(new_n5109));
  and_5  g02761(.A(new_n5109), .B(new_n5097), .Y(new_n5110));
  nor_5  g02762(.A(new_n5110), .B(new_n5108), .Y(new_n5111));
  xnor_4 g02763(.A(new_n5111), .B(new_n5107), .Y(new_n5112));
  not_8  g02764(.A(new_n5112), .Y(new_n5113));
  nor_5  g02765(.A(new_n5113), .B(new_n5105), .Y(new_n5114));
  not_8  g02766(.A(new_n5114), .Y(new_n5115_1));
  not_8  g02767(.A(n9557), .Y(new_n5116));
  xnor_4 g02768(.A(n16158), .B(new_n5116), .Y(new_n5117));
  nor_5  g02769(.A(n5752), .B(n3136), .Y(new_n5118));
  or_5   g02770(.A(new_n5110), .B(new_n5108), .Y(new_n5119));
  and_5  g02771(.A(new_n5119), .B(new_n5107), .Y(new_n5120_1));
  nor_5  g02772(.A(new_n5120_1), .B(new_n5118), .Y(new_n5121));
  xnor_4 g02773(.A(new_n5121), .B(new_n5117), .Y(new_n5122));
  not_8  g02774(.A(new_n5122), .Y(new_n5123));
  nor_5  g02775(.A(new_n5123), .B(new_n5115_1), .Y(new_n5124));
  not_8  g02776(.A(n20604), .Y(new_n5125));
  xnor_4 g02777(.A(n25643), .B(new_n5125), .Y(new_n5126));
  nor_5  g02778(.A(n16158), .B(n9557), .Y(new_n5127));
  or_5   g02779(.A(new_n5120_1), .B(new_n5118), .Y(new_n5128_1));
  and_5  g02780(.A(new_n5128_1), .B(new_n5117), .Y(new_n5129));
  nor_5  g02781(.A(new_n5129), .B(new_n5127), .Y(new_n5130));
  xnor_4 g02782(.A(new_n5130), .B(new_n5126), .Y(new_n5131_1));
  not_8  g02783(.A(new_n5131_1), .Y(new_n5132));
  xnor_4 g02784(.A(new_n5132), .B(new_n5124), .Y(new_n5133));
  xnor_4 g02785(.A(new_n5133), .B(new_n3153), .Y(new_n5134));
  xnor_4 g02786(.A(new_n5123), .B(new_n5114), .Y(new_n5135));
  nor_5  g02787(.A(new_n5135), .B(new_n3157), .Y(new_n5136));
  xnor_4 g02788(.A(new_n5135), .B(new_n3157), .Y(new_n5137));
  xnor_4 g02789(.A(new_n5113), .B(new_n5104), .Y(new_n5138));
  nor_5  g02790(.A(new_n5138), .B(new_n3163), .Y(new_n5139));
  xnor_4 g02791(.A(new_n5138), .B(new_n3160), .Y(new_n5140_1));
  xnor_4 g02792(.A(new_n5103), .B(new_n5095), .Y(new_n5141));
  and_5  g02793(.A(new_n5141), .B(new_n3165), .Y(new_n5142));
  not_8  g02794(.A(new_n5090), .Y(new_n5143));
  nor_5  g02795(.A(new_n5143), .B(new_n3170), .Y(new_n5144));
  nor_5  g02796(.A(new_n5144), .B(new_n3260_1), .Y(new_n5145));
  or_5   g02797(.A(n22309), .B(n9251), .Y(new_n5146));
  and_5  g02798(.A(new_n5100), .B(new_n5146), .Y(new_n5147));
  or_5   g02799(.A(new_n5147), .B(new_n5095), .Y(new_n5148));
  and_5  g02800(.A(new_n5144), .B(new_n3119), .Y(new_n5149));
  nor_5  g02801(.A(new_n5149), .B(new_n5145), .Y(new_n5150));
  and_5  g02802(.A(new_n5150), .B(new_n5148), .Y(new_n5151));
  nor_5  g02803(.A(new_n5151), .B(new_n5145), .Y(new_n5152));
  xnor_4 g02804(.A(new_n5141), .B(new_n3166), .Y(new_n5153));
  and_5  g02805(.A(new_n5153), .B(new_n5152), .Y(new_n5154));
  nor_5  g02806(.A(new_n5154), .B(new_n5142), .Y(new_n5155));
  and_5  g02807(.A(new_n5155), .B(new_n5140_1), .Y(new_n5156));
  nor_5  g02808(.A(new_n5156), .B(new_n5139), .Y(new_n5157));
  nor_5  g02809(.A(new_n5157), .B(new_n5137), .Y(new_n5158_1));
  nor_5  g02810(.A(new_n5158_1), .B(new_n5136), .Y(new_n5159));
  xnor_4 g02811(.A(new_n5159), .B(new_n5134), .Y(new_n5160));
  not_8  g02812(.A(new_n5160), .Y(new_n5161));
  xnor_4 g02813(.A(n5255), .B(n4119), .Y(new_n5162));
  not_8  g02814(.A(n21649), .Y(new_n5163));
  nor_5  g02815(.A(new_n5163), .B(n14510), .Y(new_n5164));
  xnor_4 g02816(.A(n21649), .B(n14510), .Y(new_n5165));
  not_8  g02817(.A(n18274), .Y(new_n5166));
  nor_5  g02818(.A(new_n5166), .B(n13263), .Y(new_n5167));
  xnor_4 g02819(.A(n18274), .B(n13263), .Y(new_n5168_1));
  nor_5  g02820(.A(new_n3446), .B(n3828), .Y(new_n5169));
  nor_5  g02821(.A(n20455), .B(new_n5064_1), .Y(new_n5170));
  nor_5  g02822(.A(n23842), .B(new_n3448), .Y(new_n5171));
  not_8  g02823(.A(n23842), .Y(new_n5172));
  nor_5  g02824(.A(new_n5172), .B(n1639), .Y(new_n5173));
  nor_5  g02825(.A(n21654), .B(new_n3451_1), .Y(new_n5174));
  not_8  g02826(.A(new_n5174), .Y(new_n5175));
  nor_5  g02827(.A(new_n5175), .B(new_n5173), .Y(new_n5176));
  nor_5  g02828(.A(new_n5176), .B(new_n5171), .Y(new_n5177));
  nor_5  g02829(.A(new_n5177), .B(new_n5170), .Y(new_n5178));
  nor_5  g02830(.A(new_n5178), .B(new_n5169), .Y(new_n5179));
  and_5  g02831(.A(new_n5179), .B(new_n5168_1), .Y(new_n5180));
  or_5   g02832(.A(new_n5180), .B(new_n5167), .Y(new_n5181));
  and_5  g02833(.A(new_n5181), .B(new_n5165), .Y(new_n5182));
  or_5   g02834(.A(new_n5182), .B(new_n5164), .Y(new_n5183));
  xor_4  g02835(.A(new_n5183), .B(new_n5162), .Y(new_n5184_1));
  xnor_4 g02836(.A(new_n5184_1), .B(new_n5161), .Y(new_n5185));
  xor_4  g02837(.A(new_n5181), .B(new_n5165), .Y(new_n5186));
  xnor_4 g02838(.A(new_n5157), .B(new_n5137), .Y(new_n5187));
  nor_5  g02839(.A(new_n5187), .B(new_n5186), .Y(new_n5188));
  xnor_4 g02840(.A(new_n5187), .B(new_n5186), .Y(new_n5189));
  xnor_4 g02841(.A(new_n5155), .B(new_n5140_1), .Y(new_n5190));
  not_8  g02842(.A(new_n5190), .Y(new_n5191));
  xnor_4 g02843(.A(new_n5179), .B(new_n5168_1), .Y(new_n5192));
  and_5  g02844(.A(new_n5192), .B(new_n5191), .Y(new_n5193));
  xnor_4 g02845(.A(new_n5192), .B(new_n5191), .Y(new_n5194));
  xnor_4 g02846(.A(new_n5153), .B(new_n5152), .Y(new_n5195));
  xnor_4 g02847(.A(n20455), .B(n3828), .Y(new_n5196));
  xnor_4 g02848(.A(new_n5196), .B(new_n5177), .Y(new_n5197));
  and_5  g02849(.A(new_n5197), .B(new_n5195), .Y(new_n5198));
  xnor_4 g02850(.A(new_n5197), .B(new_n5195), .Y(new_n5199));
  xnor_4 g02851(.A(n21654), .B(n16968), .Y(new_n5200));
  xnor_4 g02852(.A(new_n5090), .B(new_n3170), .Y(new_n5201));
  not_8  g02853(.A(new_n5201), .Y(new_n5202));
  or_5   g02854(.A(new_n5202), .B(new_n5200), .Y(new_n5203));
  xnor_4 g02855(.A(n23842), .B(n1639), .Y(new_n5204));
  xnor_4 g02856(.A(new_n5204), .B(new_n5175), .Y(new_n5205));
  and_5  g02857(.A(new_n5205), .B(new_n5203), .Y(new_n5206));
  xnor_4 g02858(.A(new_n5150), .B(new_n5148), .Y(new_n5207));
  not_8  g02859(.A(new_n5207), .Y(new_n5208));
  xor_4  g02860(.A(new_n5205), .B(new_n5203), .Y(new_n5209));
  and_5  g02861(.A(new_n5209), .B(new_n5208), .Y(new_n5210));
  nor_5  g02862(.A(new_n5210), .B(new_n5206), .Y(new_n5211_1));
  nor_5  g02863(.A(new_n5211_1), .B(new_n5199), .Y(new_n5212));
  nor_5  g02864(.A(new_n5212), .B(new_n5198), .Y(new_n5213_1));
  nor_5  g02865(.A(new_n5213_1), .B(new_n5194), .Y(new_n5214));
  nor_5  g02866(.A(new_n5214), .B(new_n5193), .Y(new_n5215));
  nor_5  g02867(.A(new_n5215), .B(new_n5189), .Y(new_n5216));
  nor_5  g02868(.A(new_n5216), .B(new_n5188), .Y(new_n5217));
  xor_4  g02869(.A(new_n5217), .B(new_n5185), .Y(n422));
  nor_5  g02870(.A(n23333), .B(n20794), .Y(new_n5219));
  not_8  g02871(.A(new_n5219), .Y(new_n5220));
  nor_5  g02872(.A(new_n5220), .B(n14603), .Y(new_n5221));
  not_8  g02873(.A(new_n5221), .Y(new_n5222));
  nor_5  g02874(.A(new_n5222), .B(n18737), .Y(new_n5223));
  not_8  g02875(.A(new_n5223), .Y(new_n5224));
  nor_5  g02876(.A(new_n5224), .B(n21471), .Y(new_n5225));
  not_8  g02877(.A(new_n5225), .Y(new_n5226_1));
  nor_5  g02878(.A(new_n5226_1), .B(n25738), .Y(new_n5227));
  not_8  g02879(.A(new_n5227), .Y(new_n5228_1));
  nor_5  g02880(.A(new_n5228_1), .B(n5302), .Y(new_n5229));
  not_8  g02881(.A(new_n5229), .Y(new_n5230));
  nor_5  g02882(.A(new_n5230), .B(n3228), .Y(new_n5231));
  xnor_4 g02883(.A(new_n5231), .B(n337), .Y(new_n5232));
  xnor_4 g02884(.A(new_n5232), .B(new_n3140), .Y(new_n5233));
  xnor_4 g02885(.A(new_n5229), .B(n3228), .Y(new_n5234));
  nor_5  g02886(.A(new_n5234), .B(n26036), .Y(new_n5235));
  xnor_4 g02887(.A(new_n5234), .B(n26036), .Y(new_n5236));
  xnor_4 g02888(.A(new_n5227), .B(n5302), .Y(new_n5237));
  nor_5  g02889(.A(new_n5237), .B(n19770), .Y(new_n5238));
  xnor_4 g02890(.A(new_n5237), .B(new_n3148), .Y(new_n5239));
  xnor_4 g02891(.A(new_n5225), .B(n25738), .Y(new_n5240));
  nor_5  g02892(.A(new_n5240), .B(n8782), .Y(new_n5241));
  xnor_4 g02893(.A(new_n5240), .B(new_n3152), .Y(new_n5242));
  xnor_4 g02894(.A(new_n5223), .B(n21471), .Y(new_n5243));
  nor_5  g02895(.A(new_n5243), .B(n8678), .Y(new_n5244));
  xnor_4 g02896(.A(new_n5243), .B(n8678), .Y(new_n5245));
  xnor_4 g02897(.A(new_n5221), .B(n18737), .Y(new_n5246));
  nor_5  g02898(.A(new_n5246), .B(n1432), .Y(new_n5247));
  xnor_4 g02899(.A(new_n5219), .B(n14603), .Y(new_n5248));
  nor_5  g02900(.A(new_n5248), .B(n21599), .Y(new_n5249));
  xor_4  g02901(.A(new_n5248), .B(n21599), .Y(new_n5250));
  xnor_4 g02902(.A(n23333), .B(new_n3307), .Y(new_n5251));
  nor_5  g02903(.A(new_n5251), .B(n25336), .Y(new_n5252));
  or_5   g02904(.A(new_n3305), .B(new_n3256), .Y(new_n5253));
  xnor_4 g02905(.A(new_n5251), .B(new_n3169), .Y(new_n5254));
  and_5  g02906(.A(new_n5254), .B(new_n5253), .Y(new_n5255_1));
  or_5   g02907(.A(new_n5255_1), .B(new_n5252), .Y(new_n5256_1));
  and_5  g02908(.A(new_n5256_1), .B(new_n5250), .Y(new_n5257));
  or_5   g02909(.A(new_n5257), .B(new_n5249), .Y(new_n5258));
  xnor_4 g02910(.A(new_n5246), .B(new_n3162), .Y(new_n5259));
  and_5  g02911(.A(new_n5259), .B(new_n5258), .Y(new_n5260));
  nor_5  g02912(.A(new_n5260), .B(new_n5247), .Y(new_n5261));
  nor_5  g02913(.A(new_n5261), .B(new_n5245), .Y(new_n5262));
  or_5   g02914(.A(new_n5262), .B(new_n5244), .Y(new_n5263));
  and_5  g02915(.A(new_n5263), .B(new_n5242), .Y(new_n5264));
  or_5   g02916(.A(new_n5264), .B(new_n5241), .Y(new_n5265_1));
  and_5  g02917(.A(new_n5265_1), .B(new_n5239), .Y(new_n5266));
  nor_5  g02918(.A(new_n5266), .B(new_n5238), .Y(new_n5267));
  nor_5  g02919(.A(new_n5267), .B(new_n5236), .Y(new_n5268));
  or_5   g02920(.A(new_n5268), .B(new_n5235), .Y(new_n5269));
  xor_4  g02921(.A(new_n5269), .B(new_n5233), .Y(new_n5270));
  xnor_4 g02922(.A(n22379), .B(n9967), .Y(new_n5271));
  nor_5  g02923(.A(n20946), .B(n1662), .Y(new_n5272));
  xnor_4 g02924(.A(n20946), .B(new_n2850), .Y(new_n5273_1));
  nor_5  g02925(.A(n12875), .B(n7751), .Y(new_n5274_1));
  not_8  g02926(.A(n7751), .Y(new_n5275));
  xnor_4 g02927(.A(n12875), .B(new_n5275), .Y(new_n5276));
  nor_5  g02928(.A(n26823), .B(n2035), .Y(new_n5277));
  xnor_4 g02929(.A(n26823), .B(new_n2856), .Y(new_n5278));
  nor_5  g02930(.A(n5213), .B(n4812), .Y(new_n5279));
  not_8  g02931(.A(n4812), .Y(new_n5280));
  xnor_4 g02932(.A(n5213), .B(new_n5280), .Y(new_n5281));
  nor_5  g02933(.A(n24278), .B(n4665), .Y(new_n5282));
  xnor_4 g02934(.A(n24278), .B(new_n2862), .Y(new_n5283));
  nor_5  g02935(.A(n24618), .B(n19005), .Y(new_n5284));
  xnor_4 g02936(.A(n24618), .B(new_n2866), .Y(new_n5285));
  nor_5  g02937(.A(n4326), .B(n3952), .Y(new_n5286));
  not_8  g02938(.A(n5438), .Y(new_n5287));
  or_5   g02939(.A(new_n2448), .B(new_n5287), .Y(new_n5288));
  xnor_4 g02940(.A(n4326), .B(new_n2443), .Y(new_n5289));
  and_5  g02941(.A(new_n5289), .B(new_n5288), .Y(new_n5290));
  or_5   g02942(.A(new_n5290), .B(new_n5286), .Y(new_n5291));
  and_5  g02943(.A(new_n5291), .B(new_n5285), .Y(new_n5292));
  or_5   g02944(.A(new_n5292), .B(new_n5284), .Y(new_n5293));
  and_5  g02945(.A(new_n5293), .B(new_n5283), .Y(new_n5294));
  or_5   g02946(.A(new_n5294), .B(new_n5282), .Y(new_n5295));
  and_5  g02947(.A(new_n5295), .B(new_n5281), .Y(new_n5296));
  or_5   g02948(.A(new_n5296), .B(new_n5279), .Y(new_n5297));
  and_5  g02949(.A(new_n5297), .B(new_n5278), .Y(new_n5298));
  or_5   g02950(.A(new_n5298), .B(new_n5277), .Y(new_n5299));
  and_5  g02951(.A(new_n5299), .B(new_n5276), .Y(new_n5300_1));
  or_5   g02952(.A(new_n5300_1), .B(new_n5274_1), .Y(new_n5301));
  and_5  g02953(.A(new_n5301), .B(new_n5273_1), .Y(new_n5302_1));
  nor_5  g02954(.A(new_n5302_1), .B(new_n5272), .Y(new_n5303));
  xnor_4 g02955(.A(new_n5303), .B(new_n5271), .Y(new_n5304));
  xnor_4 g02956(.A(n10763), .B(new_n3091), .Y(new_n5305));
  nor_5  g02957(.A(n13367), .B(n7437), .Y(new_n5306));
  xnor_4 g02958(.A(n13367), .B(new_n2890), .Y(new_n5307));
  nor_5  g02959(.A(n20700), .B(n932), .Y(new_n5308));
  xnor_4 g02960(.A(n20700), .B(n932), .Y(new_n5309));
  nor_5  g02961(.A(n7099), .B(n6691), .Y(new_n5310));
  xnor_4 g02962(.A(n7099), .B(n6691), .Y(new_n5311));
  nor_5  g02963(.A(n12811), .B(n3260), .Y(new_n5312));
  xnor_4 g02964(.A(n12811), .B(new_n3106), .Y(new_n5313));
  nor_5  g02965(.A(n20489), .B(n1118), .Y(new_n5314));
  xnor_4 g02966(.A(n20489), .B(n1118), .Y(new_n5315));
  nor_5  g02967(.A(n25974), .B(n2355), .Y(new_n5316));
  xnor_4 g02968(.A(n25974), .B(n2355), .Y(new_n5317));
  nor_5  g02969(.A(n11121), .B(n1630), .Y(new_n5318));
  nor_5  g02970(.A(new_n3117), .B(new_n2906), .Y(new_n5319));
  xnor_4 g02971(.A(n11121), .B(n1630), .Y(new_n5320));
  nor_5  g02972(.A(new_n5320), .B(new_n5319), .Y(new_n5321));
  nor_5  g02973(.A(new_n5321), .B(new_n5318), .Y(new_n5322));
  nor_5  g02974(.A(new_n5322), .B(new_n5317), .Y(new_n5323));
  nor_5  g02975(.A(new_n5323), .B(new_n5316), .Y(new_n5324));
  nor_5  g02976(.A(new_n5324), .B(new_n5315), .Y(new_n5325_1));
  or_5   g02977(.A(new_n5325_1), .B(new_n5314), .Y(new_n5326));
  and_5  g02978(.A(new_n5326), .B(new_n5313), .Y(new_n5327));
  nor_5  g02979(.A(new_n5327), .B(new_n5312), .Y(new_n5328));
  nor_5  g02980(.A(new_n5328), .B(new_n5311), .Y(new_n5329));
  nor_5  g02981(.A(new_n5329), .B(new_n5310), .Y(new_n5330_1));
  nor_5  g02982(.A(new_n5330_1), .B(new_n5309), .Y(new_n5331));
  or_5   g02983(.A(new_n5331), .B(new_n5308), .Y(new_n5332));
  and_5  g02984(.A(new_n5332), .B(new_n5307), .Y(new_n5333));
  or_5   g02985(.A(new_n5333), .B(new_n5306), .Y(new_n5334));
  xor_4  g02986(.A(new_n5334), .B(new_n5305), .Y(new_n5335));
  xnor_4 g02987(.A(new_n5335), .B(new_n5304), .Y(new_n5336));
  nor_5  g02988(.A(new_n5331), .B(new_n5308), .Y(new_n5337_1));
  xnor_4 g02989(.A(new_n5337_1), .B(new_n5307), .Y(new_n5338));
  nor_5  g02990(.A(new_n5300_1), .B(new_n5274_1), .Y(new_n5339));
  xnor_4 g02991(.A(new_n5339), .B(new_n5273_1), .Y(new_n5340));
  not_8  g02992(.A(new_n5340), .Y(new_n5341));
  nor_5  g02993(.A(new_n5341), .B(new_n5338), .Y(new_n5342));
  xnor_4 g02994(.A(new_n5340), .B(new_n5338), .Y(new_n5343));
  xnor_4 g02995(.A(new_n5330_1), .B(new_n5309), .Y(new_n5344));
  nor_5  g02996(.A(new_n5298), .B(new_n5277), .Y(new_n5345));
  xnor_4 g02997(.A(new_n5345), .B(new_n5276), .Y(new_n5346));
  nor_5  g02998(.A(new_n5346), .B(new_n5344), .Y(new_n5347));
  not_8  g02999(.A(new_n5346), .Y(new_n5348));
  xnor_4 g03000(.A(new_n5348), .B(new_n5344), .Y(new_n5349));
  xnor_4 g03001(.A(new_n5328), .B(new_n5311), .Y(new_n5350));
  nor_5  g03002(.A(new_n5296), .B(new_n5279), .Y(new_n5351_1));
  xnor_4 g03003(.A(new_n5351_1), .B(new_n5278), .Y(new_n5352));
  nor_5  g03004(.A(new_n5352), .B(new_n5350), .Y(new_n5353_1));
  xnor_4 g03005(.A(new_n5324), .B(new_n5315), .Y(new_n5354));
  nor_5  g03006(.A(new_n5292), .B(new_n5284), .Y(new_n5355));
  xnor_4 g03007(.A(new_n5355), .B(new_n5283), .Y(new_n5356));
  nor_5  g03008(.A(new_n5356), .B(new_n5354), .Y(new_n5357));
  not_8  g03009(.A(new_n5356), .Y(new_n5358));
  xnor_4 g03010(.A(new_n5358), .B(new_n5354), .Y(new_n5359));
  xnor_4 g03011(.A(new_n5322), .B(new_n5317), .Y(new_n5360));
  nor_5  g03012(.A(new_n5290), .B(new_n5286), .Y(new_n5361));
  xnor_4 g03013(.A(new_n5361), .B(new_n5285), .Y(new_n5362));
  nor_5  g03014(.A(new_n5362), .B(new_n5360), .Y(new_n5363));
  nor_5  g03015(.A(new_n2448), .B(new_n5287), .Y(new_n5364));
  xnor_4 g03016(.A(new_n5289), .B(new_n5364), .Y(new_n5365));
  xnor_4 g03017(.A(new_n5320), .B(new_n5319), .Y(new_n5366));
  nor_5  g03018(.A(new_n5366), .B(new_n5365), .Y(new_n5367));
  xnor_4 g03019(.A(n12315), .B(new_n5287), .Y(new_n5368));
  not_8  g03020(.A(new_n5368), .Y(new_n5369));
  xnor_4 g03021(.A(n16217), .B(new_n2906), .Y(new_n5370));
  nor_5  g03022(.A(new_n5370), .B(new_n5369), .Y(new_n5371));
  not_8  g03023(.A(new_n5365), .Y(new_n5372));
  xnor_4 g03024(.A(new_n5366), .B(new_n5372), .Y(new_n5373));
  and_5  g03025(.A(new_n5373), .B(new_n5371), .Y(new_n5374));
  or_5   g03026(.A(new_n5374), .B(new_n5367), .Y(new_n5375));
  not_8  g03027(.A(new_n5362), .Y(new_n5376_1));
  xnor_4 g03028(.A(new_n5376_1), .B(new_n5360), .Y(new_n5377));
  and_5  g03029(.A(new_n5377), .B(new_n5375), .Y(new_n5378));
  or_5   g03030(.A(new_n5378), .B(new_n5363), .Y(new_n5379));
  and_5  g03031(.A(new_n5379), .B(new_n5359), .Y(new_n5380));
  nor_5  g03032(.A(new_n5380), .B(new_n5357), .Y(new_n5381));
  xor_4  g03033(.A(new_n5326), .B(new_n5313), .Y(new_n5382));
  not_8  g03034(.A(new_n5382), .Y(new_n5383));
  and_5  g03035(.A(new_n5383), .B(new_n5381), .Y(new_n5384));
  xnor_4 g03036(.A(new_n5383), .B(new_n5381), .Y(new_n5385));
  nor_5  g03037(.A(new_n5294), .B(new_n5282), .Y(new_n5386_1));
  xnor_4 g03038(.A(new_n5386_1), .B(new_n5281), .Y(new_n5387));
  not_8  g03039(.A(new_n5387), .Y(new_n5388));
  nor_5  g03040(.A(new_n5388), .B(new_n5385), .Y(new_n5389));
  nor_5  g03041(.A(new_n5389), .B(new_n5384), .Y(new_n5390));
  not_8  g03042(.A(new_n5352), .Y(new_n5391));
  xnor_4 g03043(.A(new_n5391), .B(new_n5350), .Y(new_n5392));
  and_5  g03044(.A(new_n5392), .B(new_n5390), .Y(new_n5393));
  or_5   g03045(.A(new_n5393), .B(new_n5353_1), .Y(new_n5394));
  and_5  g03046(.A(new_n5394), .B(new_n5349), .Y(new_n5395));
  nor_5  g03047(.A(new_n5395), .B(new_n5347), .Y(new_n5396));
  and_5  g03048(.A(new_n5396), .B(new_n5343), .Y(new_n5397));
  nor_5  g03049(.A(new_n5397), .B(new_n5342), .Y(new_n5398));
  xnor_4 g03050(.A(new_n5398), .B(new_n5336), .Y(new_n5399_1));
  not_8  g03051(.A(new_n5399_1), .Y(new_n5400_1));
  xnor_4 g03052(.A(new_n5400_1), .B(new_n5270), .Y(new_n5401));
  xnor_4 g03053(.A(new_n5267), .B(new_n5236), .Y(new_n5402));
  xnor_4 g03054(.A(new_n5396), .B(new_n5343), .Y(new_n5403_1));
  not_8  g03055(.A(new_n5403_1), .Y(new_n5404));
  nor_5  g03056(.A(new_n5404), .B(new_n5402), .Y(new_n5405));
  xnor_4 g03057(.A(new_n5404), .B(new_n5402), .Y(new_n5406));
  xor_4  g03058(.A(new_n5265_1), .B(new_n5239), .Y(new_n5407));
  nor_5  g03059(.A(new_n5393), .B(new_n5353_1), .Y(new_n5408));
  xnor_4 g03060(.A(new_n5408), .B(new_n5349), .Y(new_n5409));
  and_5  g03061(.A(new_n5409), .B(new_n5407), .Y(new_n5410));
  xnor_4 g03062(.A(new_n5409), .B(new_n5407), .Y(new_n5411));
  xor_4  g03063(.A(new_n5263), .B(new_n5242), .Y(new_n5412));
  xnor_4 g03064(.A(new_n5392), .B(new_n5390), .Y(new_n5413));
  not_8  g03065(.A(new_n5413), .Y(new_n5414));
  and_5  g03066(.A(new_n5414), .B(new_n5412), .Y(new_n5415));
  xnor_4 g03067(.A(new_n5414), .B(new_n5412), .Y(new_n5416));
  xnor_4 g03068(.A(new_n5261), .B(new_n5245), .Y(new_n5417));
  xnor_4 g03069(.A(new_n5387), .B(new_n5385), .Y(new_n5418));
  nor_5  g03070(.A(new_n5418), .B(new_n5417), .Y(new_n5419));
  xnor_4 g03071(.A(new_n5418), .B(new_n5417), .Y(new_n5420));
  xor_4  g03072(.A(new_n5379), .B(new_n5359), .Y(new_n5421));
  xor_4  g03073(.A(new_n5259), .B(new_n5258), .Y(new_n5422));
  and_5  g03074(.A(new_n5422), .B(new_n5421), .Y(new_n5423));
  xnor_4 g03075(.A(new_n5422), .B(new_n5421), .Y(new_n5424));
  not_8  g03076(.A(new_n5424), .Y(new_n5425));
  xor_4  g03077(.A(new_n5256_1), .B(new_n5250), .Y(new_n5426));
  xor_4  g03078(.A(new_n5377), .B(new_n5375), .Y(new_n5427));
  nor_5  g03079(.A(new_n5427), .B(new_n5426), .Y(new_n5428));
  xor_4  g03080(.A(new_n5427), .B(new_n5426), .Y(new_n5429));
  xnor_4 g03081(.A(new_n5373), .B(new_n5371), .Y(new_n5430_1));
  nor_5  g03082(.A(new_n5430_1), .B(new_n5254), .Y(new_n5431));
  not_8  g03083(.A(new_n5430_1), .Y(new_n5432));
  xor_4  g03084(.A(new_n5254), .B(new_n5253), .Y(new_n5433));
  nor_5  g03085(.A(new_n5433), .B(new_n5432), .Y(new_n5434));
  xnor_4 g03086(.A(n23333), .B(n11424), .Y(new_n5435));
  xnor_4 g03087(.A(new_n5370), .B(new_n5368), .Y(new_n5436));
  nor_5  g03088(.A(new_n5436), .B(new_n5435), .Y(new_n5437));
  nor_5  g03089(.A(new_n5437), .B(new_n5434), .Y(new_n5438_1));
  nor_5  g03090(.A(new_n5438_1), .B(new_n5431), .Y(new_n5439_1));
  and_5  g03091(.A(new_n5439_1), .B(new_n5429), .Y(new_n5440));
  nor_5  g03092(.A(new_n5440), .B(new_n5428), .Y(new_n5441));
  and_5  g03093(.A(new_n5441), .B(new_n5425), .Y(new_n5442));
  nor_5  g03094(.A(new_n5442), .B(new_n5423), .Y(new_n5443_1));
  nor_5  g03095(.A(new_n5443_1), .B(new_n5420), .Y(new_n5444));
  nor_5  g03096(.A(new_n5444), .B(new_n5419), .Y(new_n5445));
  nor_5  g03097(.A(new_n5445), .B(new_n5416), .Y(new_n5446));
  nor_5  g03098(.A(new_n5446), .B(new_n5415), .Y(new_n5447));
  nor_5  g03099(.A(new_n5447), .B(new_n5411), .Y(new_n5448));
  nor_5  g03100(.A(new_n5448), .B(new_n5410), .Y(new_n5449));
  nor_5  g03101(.A(new_n5449), .B(new_n5406), .Y(new_n5450));
  nor_5  g03102(.A(new_n5450), .B(new_n5405), .Y(new_n5451_1));
  xor_4  g03103(.A(new_n5451_1), .B(new_n5401), .Y(n431));
  not_8  g03104(.A(n23895), .Y(new_n5453));
  nor_5  g03105(.A(new_n5453), .B(n8614), .Y(new_n5454));
  xnor_4 g03106(.A(n23895), .B(n8614), .Y(new_n5455));
  not_8  g03107(.A(n17351), .Y(new_n5456));
  nor_5  g03108(.A(new_n5456), .B(n15182), .Y(new_n5457));
  xnor_4 g03109(.A(n17351), .B(n15182), .Y(new_n5458));
  not_8  g03110(.A(n11736), .Y(new_n5459));
  nor_5  g03111(.A(n27037), .B(new_n5459), .Y(new_n5460));
  xnor_4 g03112(.A(n27037), .B(n11736), .Y(new_n5461));
  not_8  g03113(.A(n23200), .Y(new_n5462));
  nor_5  g03114(.A(new_n5462), .B(n8964), .Y(new_n5463));
  xnor_4 g03115(.A(n23200), .B(n8964), .Y(new_n5464));
  not_8  g03116(.A(n17959), .Y(new_n5465));
  nor_5  g03117(.A(n20151), .B(new_n5465), .Y(new_n5466));
  xnor_4 g03118(.A(n20151), .B(n17959), .Y(new_n5467));
  not_8  g03119(.A(n7566), .Y(new_n5468));
  nor_5  g03120(.A(n7693), .B(new_n5468), .Y(new_n5469));
  xnor_4 g03121(.A(n7693), .B(n7566), .Y(new_n5470));
  not_8  g03122(.A(n7731), .Y(new_n5471));
  nor_5  g03123(.A(n10405), .B(new_n5471), .Y(new_n5472_1));
  xnor_4 g03124(.A(n10405), .B(n7731), .Y(new_n5473));
  nor_5  g03125(.A(n12341), .B(new_n4106), .Y(new_n5474));
  not_8  g03126(.A(n12341), .Y(new_n5475));
  nor_5  g03127(.A(new_n5475), .B(n11302), .Y(new_n5476));
  nor_5  g03128(.A(n20986), .B(new_n4111), .Y(new_n5477));
  not_8  g03129(.A(n20986), .Y(new_n5478));
  or_5   g03130(.A(new_n5478), .B(n17090), .Y(new_n5479));
  nor_5  g03131(.A(n12384), .B(new_n4030), .Y(new_n5480));
  and_5  g03132(.A(new_n5480), .B(new_n5479), .Y(new_n5481));
  nor_5  g03133(.A(new_n5481), .B(new_n5477), .Y(new_n5482));
  nor_5  g03134(.A(new_n5482), .B(new_n5476), .Y(new_n5483));
  nor_5  g03135(.A(new_n5483), .B(new_n5474), .Y(new_n5484));
  and_5  g03136(.A(new_n5484), .B(new_n5473), .Y(new_n5485_1));
  or_5   g03137(.A(new_n5485_1), .B(new_n5472_1), .Y(new_n5486));
  and_5  g03138(.A(new_n5486), .B(new_n5470), .Y(new_n5487));
  or_5   g03139(.A(new_n5487), .B(new_n5469), .Y(new_n5488));
  and_5  g03140(.A(new_n5488), .B(new_n5467), .Y(new_n5489));
  or_5   g03141(.A(new_n5489), .B(new_n5466), .Y(new_n5490));
  and_5  g03142(.A(new_n5490), .B(new_n5464), .Y(new_n5491));
  or_5   g03143(.A(new_n5491), .B(new_n5463), .Y(new_n5492));
  and_5  g03144(.A(new_n5492), .B(new_n5461), .Y(new_n5493));
  or_5   g03145(.A(new_n5493), .B(new_n5460), .Y(new_n5494));
  and_5  g03146(.A(new_n5494), .B(new_n5458), .Y(new_n5495));
  or_5   g03147(.A(new_n5495), .B(new_n5457), .Y(new_n5496));
  and_5  g03148(.A(new_n5496), .B(new_n5455), .Y(new_n5497));
  nor_5  g03149(.A(new_n5497), .B(new_n5454), .Y(new_n5498));
  not_8  g03150(.A(new_n5498), .Y(new_n5499));
  not_8  g03151(.A(n13494), .Y(new_n5500));
  nor_5  g03152(.A(n18880), .B(new_n5500), .Y(new_n5501));
  xnor_4 g03153(.A(n18880), .B(n13494), .Y(new_n5502));
  not_8  g03154(.A(n25345), .Y(new_n5503));
  nor_5  g03155(.A(n25475), .B(new_n5503), .Y(new_n5504));
  xnor_4 g03156(.A(n25475), .B(n25345), .Y(new_n5505));
  not_8  g03157(.A(n9655), .Y(new_n5506));
  nor_5  g03158(.A(n23849), .B(new_n5506), .Y(new_n5507));
  xnor_4 g03159(.A(n23849), .B(n9655), .Y(new_n5508));
  and_5  g03160(.A(n13490), .B(new_n4442), .Y(new_n5509));
  xnor_4 g03161(.A(n13490), .B(n12446), .Y(new_n5510));
  not_8  g03162(.A(n22660), .Y(new_n5511));
  nor_5  g03163(.A(new_n5511), .B(n11011), .Y(new_n5512));
  xnor_4 g03164(.A(n22660), .B(n11011), .Y(new_n5513));
  not_8  g03165(.A(n1777), .Y(new_n5514));
  nor_5  g03166(.A(n16029), .B(new_n5514), .Y(new_n5515));
  xnor_4 g03167(.A(n16029), .B(n1777), .Y(new_n5516));
  not_8  g03168(.A(n8745), .Y(new_n5517_1));
  nor_5  g03169(.A(n16476), .B(new_n5517_1), .Y(new_n5518));
  xnor_4 g03170(.A(n16476), .B(n8745), .Y(new_n5519));
  nor_5  g03171(.A(n15636), .B(new_n3947), .Y(new_n5520));
  nor_5  g03172(.A(new_n2441), .B(n11615), .Y(new_n5521_1));
  nor_5  g03173(.A(new_n3949), .B(n20077), .Y(new_n5522));
  nor_5  g03174(.A(n22433), .B(new_n2444_1), .Y(new_n5523));
  or_5   g03175(.A(new_n3952_1), .B(n6794), .Y(new_n5524_1));
  nor_5  g03176(.A(new_n5524_1), .B(new_n5523), .Y(new_n5525));
  nor_5  g03177(.A(new_n5525), .B(new_n5522), .Y(new_n5526));
  nor_5  g03178(.A(new_n5526), .B(new_n5521_1), .Y(new_n5527));
  nor_5  g03179(.A(new_n5527), .B(new_n5520), .Y(new_n5528));
  and_5  g03180(.A(new_n5528), .B(new_n5519), .Y(new_n5529));
  or_5   g03181(.A(new_n5529), .B(new_n5518), .Y(new_n5530));
  and_5  g03182(.A(new_n5530), .B(new_n5516), .Y(new_n5531));
  or_5   g03183(.A(new_n5531), .B(new_n5515), .Y(new_n5532_1));
  and_5  g03184(.A(new_n5532_1), .B(new_n5513), .Y(new_n5533));
  or_5   g03185(.A(new_n5533), .B(new_n5512), .Y(new_n5534));
  and_5  g03186(.A(new_n5534), .B(new_n5510), .Y(new_n5535));
  or_5   g03187(.A(new_n5535), .B(new_n5509), .Y(new_n5536));
  and_5  g03188(.A(new_n5536), .B(new_n5508), .Y(new_n5537));
  or_5   g03189(.A(new_n5537), .B(new_n5507), .Y(new_n5538));
  and_5  g03190(.A(new_n5538), .B(new_n5505), .Y(new_n5539));
  or_5   g03191(.A(new_n5539), .B(new_n5504), .Y(new_n5540));
  and_5  g03192(.A(new_n5540), .B(new_n5502), .Y(new_n5541));
  nor_5  g03193(.A(new_n5541), .B(new_n5501), .Y(new_n5542));
  nor_5  g03194(.A(new_n5539), .B(new_n5504), .Y(new_n5543));
  xnor_4 g03195(.A(new_n5543), .B(new_n5502), .Y(new_n5544));
  nor_5  g03196(.A(n22173), .B(n583), .Y(new_n5545));
  not_8  g03197(.A(new_n5545), .Y(new_n5546));
  nor_5  g03198(.A(new_n5546), .B(n2146), .Y(new_n5547));
  not_8  g03199(.A(new_n5547), .Y(new_n5548));
  nor_5  g03200(.A(new_n5548), .B(n23974), .Y(new_n5549));
  not_8  g03201(.A(new_n5549), .Y(new_n5550));
  nor_5  g03202(.A(new_n5550), .B(n3909), .Y(new_n5551));
  not_8  g03203(.A(new_n5551), .Y(new_n5552));
  nor_5  g03204(.A(new_n5552), .B(n20429), .Y(new_n5553));
  not_8  g03205(.A(new_n5553), .Y(new_n5554));
  nor_5  g03206(.A(new_n5554), .B(n22554), .Y(new_n5555));
  not_8  g03207(.A(new_n5555), .Y(new_n5556));
  nor_5  g03208(.A(new_n5556), .B(n23913), .Y(new_n5557));
  xnor_4 g03209(.A(new_n5557), .B(n26797), .Y(new_n5558));
  nor_5  g03210(.A(new_n5558), .B(n10201), .Y(new_n5559));
  not_8  g03211(.A(n10201), .Y(new_n5560));
  xnor_4 g03212(.A(new_n5558), .B(new_n5560), .Y(new_n5561));
  xnor_4 g03213(.A(new_n5555), .B(n23913), .Y(new_n5562));
  nor_5  g03214(.A(new_n5562), .B(n10593), .Y(new_n5563));
  not_8  g03215(.A(n10593), .Y(new_n5564_1));
  xnor_4 g03216(.A(new_n5562), .B(new_n5564_1), .Y(new_n5565));
  xnor_4 g03217(.A(new_n5553), .B(n22554), .Y(new_n5566));
  nor_5  g03218(.A(new_n5566), .B(n18290), .Y(new_n5567));
  not_8  g03219(.A(n18290), .Y(new_n5568));
  xnor_4 g03220(.A(new_n5566), .B(new_n5568), .Y(new_n5569));
  xnor_4 g03221(.A(new_n5551), .B(n20429), .Y(new_n5570));
  nor_5  g03222(.A(new_n5570), .B(n11580), .Y(new_n5571));
  not_8  g03223(.A(n11580), .Y(new_n5572));
  xnor_4 g03224(.A(new_n5570), .B(new_n5572), .Y(new_n5573));
  xnor_4 g03225(.A(new_n5549), .B(n3909), .Y(new_n5574));
  nor_5  g03226(.A(new_n5574), .B(n15884), .Y(new_n5575));
  not_8  g03227(.A(n15884), .Y(new_n5576));
  xnor_4 g03228(.A(new_n5574), .B(new_n5576), .Y(new_n5577));
  xnor_4 g03229(.A(new_n5547), .B(n23974), .Y(new_n5578));
  nor_5  g03230(.A(new_n5578), .B(n6356), .Y(new_n5579_1));
  xnor_4 g03231(.A(new_n5545), .B(n2146), .Y(new_n5580));
  nor_5  g03232(.A(new_n5580), .B(n27104), .Y(new_n5581));
  not_8  g03233(.A(n27104), .Y(new_n5582));
  xnor_4 g03234(.A(new_n5580), .B(new_n5582), .Y(new_n5583));
  not_8  g03235(.A(n27188), .Y(new_n5584));
  xnor_4 g03236(.A(n22173), .B(n583), .Y(new_n5585));
  and_5  g03237(.A(new_n5585), .B(new_n5584), .Y(new_n5586));
  not_8  g03238(.A(n583), .Y(new_n5587));
  not_8  g03239(.A(n6611), .Y(new_n5588));
  or_5   g03240(.A(new_n5588), .B(new_n5587), .Y(new_n5589));
  xnor_4 g03241(.A(new_n5585), .B(n27188), .Y(new_n5590));
  and_5  g03242(.A(new_n5590), .B(new_n5589), .Y(new_n5591));
  or_5   g03243(.A(new_n5591), .B(new_n5586), .Y(new_n5592));
  and_5  g03244(.A(new_n5592), .B(new_n5583), .Y(new_n5593_1));
  or_5   g03245(.A(new_n5593_1), .B(new_n5581), .Y(new_n5594));
  not_8  g03246(.A(n6356), .Y(new_n5595));
  xnor_4 g03247(.A(new_n5578), .B(new_n5595), .Y(new_n5596));
  and_5  g03248(.A(new_n5596), .B(new_n5594), .Y(new_n5597));
  or_5   g03249(.A(new_n5597), .B(new_n5579_1), .Y(new_n5598));
  and_5  g03250(.A(new_n5598), .B(new_n5577), .Y(new_n5599));
  or_5   g03251(.A(new_n5599), .B(new_n5575), .Y(new_n5600));
  and_5  g03252(.A(new_n5600), .B(new_n5573), .Y(new_n5601));
  or_5   g03253(.A(new_n5601), .B(new_n5571), .Y(new_n5602));
  and_5  g03254(.A(new_n5602), .B(new_n5569), .Y(new_n5603_1));
  or_5   g03255(.A(new_n5603_1), .B(new_n5567), .Y(new_n5604));
  and_5  g03256(.A(new_n5604), .B(new_n5565), .Y(new_n5605_1));
  or_5   g03257(.A(new_n5605_1), .B(new_n5563), .Y(new_n5606));
  and_5  g03258(.A(new_n5606), .B(new_n5561), .Y(new_n5607));
  nor_5  g03259(.A(new_n5607), .B(new_n5559), .Y(new_n5608));
  not_8  g03260(.A(new_n5608), .Y(new_n5609_1));
  not_8  g03261(.A(n12650), .Y(new_n5610));
  not_8  g03262(.A(n26797), .Y(new_n5611));
  and_5  g03263(.A(new_n5557), .B(new_n5611), .Y(new_n5612));
  xnor_4 g03264(.A(new_n5612), .B(n12702), .Y(new_n5613));
  xnor_4 g03265(.A(new_n5613), .B(new_n5610), .Y(new_n5614));
  xnor_4 g03266(.A(new_n5614), .B(new_n5609_1), .Y(new_n5615));
  nor_5  g03267(.A(new_n5615), .B(new_n5544), .Y(new_n5616));
  xnor_4 g03268(.A(new_n5615), .B(new_n5544), .Y(new_n5617));
  nor_5  g03269(.A(new_n5537), .B(new_n5507), .Y(new_n5618));
  xnor_4 g03270(.A(new_n5618), .B(new_n5505), .Y(new_n5619));
  not_8  g03271(.A(new_n5619), .Y(new_n5620));
  xor_4  g03272(.A(new_n5606), .B(new_n5561), .Y(new_n5621));
  and_5  g03273(.A(new_n5621), .B(new_n5620), .Y(new_n5622));
  xnor_4 g03274(.A(new_n5621), .B(new_n5620), .Y(new_n5623));
  nor_5  g03275(.A(new_n5535), .B(new_n5509), .Y(new_n5624));
  xnor_4 g03276(.A(new_n5624), .B(new_n5508), .Y(new_n5625));
  not_8  g03277(.A(new_n5625), .Y(new_n5626));
  xor_4  g03278(.A(new_n5604), .B(new_n5565), .Y(new_n5627));
  and_5  g03279(.A(new_n5627), .B(new_n5626), .Y(new_n5628));
  xnor_4 g03280(.A(new_n5627), .B(new_n5626), .Y(new_n5629));
  nor_5  g03281(.A(new_n5533), .B(new_n5512), .Y(new_n5630));
  xnor_4 g03282(.A(new_n5630), .B(new_n5510), .Y(new_n5631));
  not_8  g03283(.A(new_n5631), .Y(new_n5632));
  xor_4  g03284(.A(new_n5602), .B(new_n5569), .Y(new_n5633));
  and_5  g03285(.A(new_n5633), .B(new_n5632), .Y(new_n5634_1));
  xnor_4 g03286(.A(new_n5633), .B(new_n5632), .Y(new_n5635));
  nor_5  g03287(.A(new_n5531), .B(new_n5515), .Y(new_n5636));
  xnor_4 g03288(.A(new_n5636), .B(new_n5513), .Y(new_n5637));
  not_8  g03289(.A(new_n5637), .Y(new_n5638));
  xor_4  g03290(.A(new_n5600), .B(new_n5573), .Y(new_n5639));
  and_5  g03291(.A(new_n5639), .B(new_n5638), .Y(new_n5640));
  xnor_4 g03292(.A(new_n5639), .B(new_n5638), .Y(new_n5641));
  nor_5  g03293(.A(new_n5529), .B(new_n5518), .Y(new_n5642));
  xnor_4 g03294(.A(new_n5642), .B(new_n5516), .Y(new_n5643_1));
  not_8  g03295(.A(new_n5643_1), .Y(new_n5644));
  xor_4  g03296(.A(new_n5598), .B(new_n5577), .Y(new_n5645));
  and_5  g03297(.A(new_n5645), .B(new_n5644), .Y(new_n5646));
  xnor_4 g03298(.A(new_n5645), .B(new_n5644), .Y(new_n5647));
  xor_4  g03299(.A(new_n5528), .B(new_n5519), .Y(new_n5648));
  not_8  g03300(.A(new_n5648), .Y(new_n5649));
  xor_4  g03301(.A(new_n5596), .B(new_n5594), .Y(new_n5650));
  and_5  g03302(.A(new_n5650), .B(new_n5649), .Y(new_n5651));
  xnor_4 g03303(.A(new_n5650), .B(new_n5648), .Y(new_n5652));
  xor_4  g03304(.A(new_n5592), .B(new_n5583), .Y(new_n5653));
  xnor_4 g03305(.A(n15636), .B(n11615), .Y(new_n5654));
  xnor_4 g03306(.A(new_n5654), .B(new_n5526), .Y(new_n5655));
  nor_5  g03307(.A(new_n5655), .B(new_n5653), .Y(new_n5656));
  xnor_4 g03308(.A(new_n5655), .B(new_n5653), .Y(new_n5657));
  nor_5  g03309(.A(new_n5588), .B(new_n5587), .Y(new_n5658));
  xnor_4 g03310(.A(new_n5590), .B(new_n5658), .Y(new_n5659));
  xnor_4 g03311(.A(n22433), .B(n20077), .Y(new_n5660));
  xnor_4 g03312(.A(new_n5660), .B(new_n5524_1), .Y(new_n5661));
  nor_5  g03313(.A(new_n5661), .B(new_n5659), .Y(new_n5662));
  xnor_4 g03314(.A(n14090), .B(n6794), .Y(new_n5663));
  xnor_4 g03315(.A(n6611), .B(n583), .Y(new_n5664));
  nor_5  g03316(.A(new_n5664), .B(new_n5663), .Y(new_n5665));
  not_8  g03317(.A(new_n5661), .Y(new_n5666));
  xnor_4 g03318(.A(new_n5666), .B(new_n5659), .Y(new_n5667));
  and_5  g03319(.A(new_n5667), .B(new_n5665), .Y(new_n5668));
  nor_5  g03320(.A(new_n5668), .B(new_n5662), .Y(new_n5669));
  nor_5  g03321(.A(new_n5669), .B(new_n5657), .Y(new_n5670));
  nor_5  g03322(.A(new_n5670), .B(new_n5656), .Y(new_n5671));
  and_5  g03323(.A(new_n5671), .B(new_n5652), .Y(new_n5672));
  nor_5  g03324(.A(new_n5672), .B(new_n5651), .Y(new_n5673));
  nor_5  g03325(.A(new_n5673), .B(new_n5647), .Y(new_n5674));
  nor_5  g03326(.A(new_n5674), .B(new_n5646), .Y(new_n5675));
  nor_5  g03327(.A(new_n5675), .B(new_n5641), .Y(new_n5676));
  nor_5  g03328(.A(new_n5676), .B(new_n5640), .Y(new_n5677));
  nor_5  g03329(.A(new_n5677), .B(new_n5635), .Y(new_n5678));
  nor_5  g03330(.A(new_n5678), .B(new_n5634_1), .Y(new_n5679));
  nor_5  g03331(.A(new_n5679), .B(new_n5629), .Y(new_n5680_1));
  nor_5  g03332(.A(new_n5680_1), .B(new_n5628), .Y(new_n5681));
  nor_5  g03333(.A(new_n5681), .B(new_n5623), .Y(new_n5682));
  nor_5  g03334(.A(new_n5682), .B(new_n5622), .Y(new_n5683));
  nor_5  g03335(.A(new_n5683), .B(new_n5617), .Y(new_n5684));
  nor_5  g03336(.A(new_n5684), .B(new_n5616), .Y(new_n5685));
  not_8  g03337(.A(n12702), .Y(new_n5686));
  and_5  g03338(.A(new_n5612), .B(new_n5686), .Y(new_n5687_1));
  and_5  g03339(.A(new_n5613), .B(n12650), .Y(new_n5688));
  nor_5  g03340(.A(new_n5613), .B(n12650), .Y(new_n5689));
  nor_5  g03341(.A(new_n5689), .B(new_n5609_1), .Y(new_n5690));
  or_5   g03342(.A(new_n5690), .B(new_n5688), .Y(new_n5691));
  nor_5  g03343(.A(new_n5691), .B(new_n5687_1), .Y(new_n5692));
  not_8  g03344(.A(new_n5692), .Y(new_n5693));
  and_5  g03345(.A(new_n5693), .B(new_n5685), .Y(new_n5694));
  and_5  g03346(.A(new_n5694), .B(new_n5542), .Y(new_n5695));
  or_5   g03347(.A(new_n5693), .B(new_n5685), .Y(new_n5696_1));
  nor_5  g03348(.A(new_n5696_1), .B(new_n5542), .Y(new_n5697));
  nor_5  g03349(.A(new_n5697), .B(new_n5695), .Y(new_n5698));
  not_8  g03350(.A(new_n5698), .Y(new_n5699));
  xnor_4 g03351(.A(new_n5699), .B(new_n5499), .Y(new_n5700_1));
  xnor_4 g03352(.A(new_n5692), .B(new_n5685), .Y(new_n5701));
  xnor_4 g03353(.A(new_n5701), .B(new_n5542), .Y(new_n5702));
  and_5  g03354(.A(new_n5702), .B(new_n5498), .Y(new_n5703));
  or_5   g03355(.A(new_n5702), .B(new_n5498), .Y(new_n5704_1));
  xor_4  g03356(.A(new_n5496), .B(new_n5455), .Y(new_n5705));
  xnor_4 g03357(.A(new_n5683), .B(new_n5617), .Y(new_n5706));
  nor_5  g03358(.A(new_n5706), .B(new_n5705), .Y(new_n5707));
  xnor_4 g03359(.A(new_n5706), .B(new_n5705), .Y(new_n5708));
  xor_4  g03360(.A(new_n5494), .B(new_n5458), .Y(new_n5709));
  xnor_4 g03361(.A(new_n5681), .B(new_n5623), .Y(new_n5710));
  nor_5  g03362(.A(new_n5710), .B(new_n5709), .Y(new_n5711));
  xnor_4 g03363(.A(new_n5710), .B(new_n5709), .Y(new_n5712));
  xor_4  g03364(.A(new_n5492), .B(new_n5461), .Y(new_n5713));
  xnor_4 g03365(.A(new_n5679), .B(new_n5629), .Y(new_n5714));
  nor_5  g03366(.A(new_n5714), .B(new_n5713), .Y(new_n5715));
  xnor_4 g03367(.A(new_n5714), .B(new_n5713), .Y(new_n5716));
  xor_4  g03368(.A(new_n5490), .B(new_n5464), .Y(new_n5717));
  xnor_4 g03369(.A(new_n5677), .B(new_n5635), .Y(new_n5718));
  nor_5  g03370(.A(new_n5718), .B(new_n5717), .Y(new_n5719));
  xnor_4 g03371(.A(new_n5718), .B(new_n5717), .Y(new_n5720));
  xor_4  g03372(.A(new_n5488), .B(new_n5467), .Y(new_n5721));
  xnor_4 g03373(.A(new_n5675), .B(new_n5641), .Y(new_n5722));
  nor_5  g03374(.A(new_n5722), .B(new_n5721), .Y(new_n5723));
  xnor_4 g03375(.A(new_n5722), .B(new_n5721), .Y(new_n5724));
  xor_4  g03376(.A(new_n5486), .B(new_n5470), .Y(new_n5725));
  xnor_4 g03377(.A(new_n5673), .B(new_n5647), .Y(new_n5726));
  nor_5  g03378(.A(new_n5726), .B(new_n5725), .Y(new_n5727));
  xnor_4 g03379(.A(new_n5726), .B(new_n5725), .Y(new_n5728));
  xnor_4 g03380(.A(new_n5671), .B(new_n5652), .Y(new_n5729));
  not_8  g03381(.A(new_n5729), .Y(new_n5730));
  xnor_4 g03382(.A(new_n5484), .B(new_n5473), .Y(new_n5731));
  and_5  g03383(.A(new_n5731), .B(new_n5730), .Y(new_n5732_1));
  xnor_4 g03384(.A(new_n5731), .B(new_n5730), .Y(new_n5733));
  xnor_4 g03385(.A(new_n5669), .B(new_n5657), .Y(new_n5734));
  xnor_4 g03386(.A(n12341), .B(n11302), .Y(new_n5735));
  xnor_4 g03387(.A(new_n5735), .B(new_n5482), .Y(new_n5736));
  and_5  g03388(.A(new_n5736), .B(new_n5734), .Y(new_n5737));
  xnor_4 g03389(.A(new_n5736), .B(new_n5734), .Y(new_n5738));
  xnor_4 g03390(.A(new_n5664), .B(new_n5663), .Y(new_n5739));
  xnor_4 g03391(.A(n12384), .B(n6773), .Y(new_n5740));
  nor_5  g03392(.A(new_n5740), .B(new_n5739), .Y(new_n5741));
  xnor_4 g03393(.A(n20986), .B(n17090), .Y(new_n5742_1));
  xnor_4 g03394(.A(new_n5742_1), .B(new_n5480), .Y(new_n5743));
  nor_5  g03395(.A(new_n5743), .B(new_n5741), .Y(new_n5744));
  xnor_4 g03396(.A(new_n5667), .B(new_n5665), .Y(new_n5745));
  not_8  g03397(.A(new_n5745), .Y(new_n5746));
  xnor_4 g03398(.A(new_n5743), .B(new_n5741), .Y(new_n5747));
  nor_5  g03399(.A(new_n5747), .B(new_n5746), .Y(new_n5748));
  nor_5  g03400(.A(new_n5748), .B(new_n5744), .Y(new_n5749));
  nor_5  g03401(.A(new_n5749), .B(new_n5738), .Y(new_n5750));
  nor_5  g03402(.A(new_n5750), .B(new_n5737), .Y(new_n5751));
  nor_5  g03403(.A(new_n5751), .B(new_n5733), .Y(new_n5752_1));
  nor_5  g03404(.A(new_n5752_1), .B(new_n5732_1), .Y(new_n5753));
  nor_5  g03405(.A(new_n5753), .B(new_n5728), .Y(new_n5754));
  nor_5  g03406(.A(new_n5754), .B(new_n5727), .Y(new_n5755));
  nor_5  g03407(.A(new_n5755), .B(new_n5724), .Y(new_n5756));
  nor_5  g03408(.A(new_n5756), .B(new_n5723), .Y(new_n5757));
  nor_5  g03409(.A(new_n5757), .B(new_n5720), .Y(new_n5758));
  nor_5  g03410(.A(new_n5758), .B(new_n5719), .Y(new_n5759));
  nor_5  g03411(.A(new_n5759), .B(new_n5716), .Y(new_n5760));
  nor_5  g03412(.A(new_n5760), .B(new_n5715), .Y(new_n5761));
  nor_5  g03413(.A(new_n5761), .B(new_n5712), .Y(new_n5762));
  nor_5  g03414(.A(new_n5762), .B(new_n5711), .Y(new_n5763));
  nor_5  g03415(.A(new_n5763), .B(new_n5708), .Y(new_n5764));
  nor_5  g03416(.A(new_n5764), .B(new_n5707), .Y(new_n5765_1));
  and_5  g03417(.A(new_n5765_1), .B(new_n5704_1), .Y(new_n5766));
  nor_5  g03418(.A(new_n5766), .B(new_n5703), .Y(new_n5767));
  xnor_4 g03419(.A(new_n5767), .B(new_n5700_1), .Y(n457));
  xnor_4 g03420(.A(n24323), .B(n1681), .Y(new_n5769));
  xnor_4 g03421(.A(n13781), .B(new_n2951), .Y(new_n5770));
  xnor_4 g03422(.A(new_n5770), .B(new_n5769), .Y(new_n5771));
  not_8  g03423(.A(new_n5771), .Y(new_n5772));
  nor_5  g03424(.A(new_n5772), .B(new_n5663), .Y(new_n5773));
  xnor_4 g03425(.A(new_n5773), .B(new_n5666), .Y(new_n5774));
  not_8  g03426(.A(new_n5770), .Y(new_n5775));
  nor_5  g03427(.A(new_n5775), .B(new_n5769), .Y(new_n5776_1));
  nor_5  g03428(.A(n24323), .B(new_n4394), .Y(new_n5777));
  xnor_4 g03429(.A(n26443), .B(n25877), .Y(new_n5778));
  xnor_4 g03430(.A(new_n5778), .B(new_n5777), .Y(new_n5779));
  xnor_4 g03431(.A(new_n5779), .B(new_n5776_1), .Y(new_n5780));
  xnor_4 g03432(.A(n9399), .B(new_n2951), .Y(new_n5781));
  nor_5  g03433(.A(new_n2383), .B(new_n2951), .Y(new_n5782_1));
  nor_5  g03434(.A(new_n5782_1), .B(n11486), .Y(new_n5783));
  not_8  g03435(.A(n11486), .Y(new_n5784));
  or_5   g03436(.A(new_n2383), .B(new_n5784), .Y(new_n5785));
  nor_5  g03437(.A(new_n5785), .B(new_n2951), .Y(new_n5786));
  nor_5  g03438(.A(new_n5786), .B(new_n5783), .Y(new_n5787));
  xnor_4 g03439(.A(new_n5787), .B(new_n5781), .Y(new_n5788));
  not_8  g03440(.A(new_n5788), .Y(new_n5789));
  xnor_4 g03441(.A(new_n5789), .B(new_n5780), .Y(new_n5790));
  xnor_4 g03442(.A(new_n5790), .B(new_n5774), .Y(n463));
  xnor_4 g03443(.A(n12121), .B(n6775), .Y(new_n5792));
  xnor_4 g03444(.A(new_n5792), .B(n8920), .Y(new_n5793));
  not_8  g03445(.A(new_n5793), .Y(new_n5794));
  xnor_4 g03446(.A(new_n3063), .B(n5438), .Y(new_n5795));
  xnor_4 g03447(.A(new_n5795), .B(new_n5794), .Y(n491));
  xnor_4 g03448(.A(new_n5751), .B(new_n5733), .Y(n496));
  not_8  g03449(.A(n12384), .Y(new_n5798));
  xnor_4 g03450(.A(n25926), .B(new_n5798), .Y(new_n5799));
  not_8  g03451(.A(new_n5799), .Y(new_n5800));
  xnor_4 g03452(.A(new_n5800), .B(new_n4030), .Y(new_n5801));
  xnor_4 g03453(.A(new_n5663), .B(n16167), .Y(new_n5802));
  not_8  g03454(.A(new_n5802), .Y(new_n5803));
  nor_5  g03455(.A(new_n5803), .B(new_n5801), .Y(new_n5804));
  not_8  g03456(.A(n16167), .Y(new_n5805));
  or_5   g03457(.A(new_n5663), .B(new_n5805), .Y(new_n5806));
  not_8  g03458(.A(n18745), .Y(new_n5807));
  xnor_4 g03459(.A(new_n5666), .B(new_n5807), .Y(new_n5808));
  xor_4  g03460(.A(new_n5808), .B(new_n5806), .Y(new_n5809));
  nor_5  g03461(.A(new_n3982), .B(new_n5798), .Y(new_n5810));
  xnor_4 g03462(.A(n25926), .B(n7657), .Y(new_n5811));
  xnor_4 g03463(.A(new_n5811), .B(n20986), .Y(new_n5812));
  xnor_4 g03464(.A(new_n5812), .B(new_n5810), .Y(new_n5813));
  not_8  g03465(.A(new_n5813), .Y(new_n5814));
  or_5   g03466(.A(new_n5800), .B(new_n4030), .Y(new_n5815));
  nor_5  g03467(.A(new_n5815), .B(n17090), .Y(new_n5816));
  nor_5  g03468(.A(n17090), .B(n6773), .Y(new_n5817));
  or_5   g03469(.A(new_n4111), .B(new_n4030), .Y(new_n5818));
  nor_5  g03470(.A(new_n5818), .B(new_n5799), .Y(new_n5819));
  or_5   g03471(.A(new_n5819), .B(new_n5817), .Y(new_n5820));
  nor_5  g03472(.A(new_n5820), .B(new_n5816), .Y(new_n5821));
  xnor_4 g03473(.A(new_n5821), .B(new_n5814), .Y(new_n5822_1));
  xnor_4 g03474(.A(new_n5822_1), .B(new_n5809), .Y(new_n5823));
  xnor_4 g03475(.A(new_n5823), .B(new_n5804), .Y(n498));
  xnor_4 g03476(.A(n25872), .B(new_n4237), .Y(new_n5825));
  nor_5  g03477(.A(n22043), .B(n20259), .Y(new_n5826));
  or_5   g03478(.A(new_n3875), .B(new_n5002), .Y(new_n5827));
  xnor_4 g03479(.A(n22043), .B(new_n4939_1), .Y(new_n5828));
  and_5  g03480(.A(new_n5828), .B(new_n5827), .Y(new_n5829));
  or_5   g03481(.A(new_n5829), .B(new_n5826), .Y(new_n5830));
  xor_4  g03482(.A(new_n5830), .B(new_n5825), .Y(new_n5831));
  xnor_4 g03483(.A(new_n5831), .B(new_n4880), .Y(new_n5832));
  nor_5  g03484(.A(new_n3875), .B(new_n5002), .Y(new_n5833_1));
  xnor_4 g03485(.A(new_n5828), .B(new_n5833_1), .Y(new_n5834_1));
  nor_5  g03486(.A(new_n5834_1), .B(new_n4872), .Y(new_n5835));
  xnor_4 g03487(.A(n12121), .B(new_n5002), .Y(new_n5836));
  or_5   g03488(.A(new_n5836), .B(new_n4874), .Y(new_n5837));
  not_8  g03489(.A(new_n5834_1), .Y(new_n5838));
  xnor_4 g03490(.A(new_n5838), .B(new_n4872), .Y(new_n5839));
  and_5  g03491(.A(new_n5839), .B(new_n5837), .Y(new_n5840_1));
  nor_5  g03492(.A(new_n5840_1), .B(new_n5835), .Y(new_n5841_1));
  xnor_4 g03493(.A(new_n5841_1), .B(new_n5832), .Y(new_n5842_1));
  xnor_4 g03494(.A(new_n5842_1), .B(new_n3792), .Y(new_n5843));
  xor_4  g03495(.A(new_n5839), .B(new_n5837), .Y(new_n5844));
  nor_5  g03496(.A(new_n5844), .B(new_n3759), .Y(new_n5845));
  not_8  g03497(.A(new_n3796), .Y(new_n5846));
  and_5  g03498(.A(new_n5844), .B(new_n5846), .Y(new_n5847));
  xnor_4 g03499(.A(new_n5836), .B(new_n4874), .Y(new_n5848));
  and_5  g03500(.A(new_n5848), .B(new_n3799), .Y(new_n5849));
  nor_5  g03501(.A(new_n5849), .B(new_n5847), .Y(new_n5850_1));
  nor_5  g03502(.A(new_n5850_1), .B(new_n5845), .Y(new_n5851));
  xor_4  g03503(.A(new_n5851), .B(new_n5843), .Y(n521));
  not_8  g03504(.A(new_n5739), .Y(new_n5853));
  xnor_4 g03505(.A(new_n5740), .B(new_n5853), .Y(n548));
  xor_4  g03506(.A(new_n4308), .B(new_n4289), .Y(n554));
  nor_5  g03507(.A(n20658), .B(n15743), .Y(new_n5856));
  not_8  g03508(.A(new_n5856), .Y(new_n5857));
  nor_5  g03509(.A(new_n5857), .B(n7524), .Y(new_n5858));
  not_8  g03510(.A(new_n5858), .Y(new_n5859));
  nor_5  g03511(.A(new_n5859), .B(n4957), .Y(new_n5860));
  not_8  g03512(.A(new_n5860), .Y(new_n5861));
  nor_5  g03513(.A(new_n5861), .B(n9003), .Y(new_n5862));
  not_8  g03514(.A(new_n5862), .Y(new_n5863));
  nor_5  g03515(.A(new_n5863), .B(n3161), .Y(new_n5864));
  not_8  g03516(.A(new_n5864), .Y(new_n5865));
  nor_5  g03517(.A(new_n5865), .B(n25749), .Y(new_n5866));
  not_8  g03518(.A(new_n5866), .Y(new_n5867));
  nor_5  g03519(.A(new_n5867), .B(n20409), .Y(new_n5868));
  not_8  g03520(.A(new_n5868), .Y(new_n5869));
  nor_5  g03521(.A(new_n5869), .B(n647), .Y(new_n5870));
  xnor_4 g03522(.A(new_n5870), .B(n2979), .Y(new_n5871));
  not_8  g03523(.A(n6456), .Y(new_n5872));
  xnor_4 g03524(.A(n9259), .B(new_n5872), .Y(new_n5873));
  nor_5  g03525(.A(n21489), .B(n4085), .Y(new_n5874));
  not_8  g03526(.A(n4085), .Y(new_n5875));
  xnor_4 g03527(.A(n21489), .B(new_n5875), .Y(new_n5876));
  nor_5  g03528(.A(n26725), .B(n20213), .Y(new_n5877));
  xnor_4 g03529(.A(n26725), .B(new_n4844), .Y(new_n5878));
  nor_5  g03530(.A(n13912), .B(n11980), .Y(new_n5879));
  not_8  g03531(.A(n11980), .Y(new_n5880));
  xnor_4 g03532(.A(n13912), .B(new_n5880), .Y(new_n5881));
  nor_5  g03533(.A(n7670), .B(n3253), .Y(new_n5882_1));
  not_8  g03534(.A(n3253), .Y(new_n5883));
  xnor_4 g03535(.A(n7670), .B(new_n5883), .Y(new_n5884));
  nor_5  g03536(.A(n9598), .B(n7759), .Y(new_n5885));
  not_8  g03537(.A(n7759), .Y(new_n5886));
  xnor_4 g03538(.A(n9598), .B(new_n5886), .Y(new_n5887));
  nor_5  g03539(.A(n22290), .B(n12562), .Y(new_n5888));
  not_8  g03540(.A(n12562), .Y(new_n5889));
  xnor_4 g03541(.A(n22290), .B(new_n5889), .Y(new_n5890));
  nor_5  g03542(.A(n11273), .B(n7949), .Y(new_n5891));
  not_8  g03543(.A(n7949), .Y(new_n5892));
  xnor_4 g03544(.A(n11273), .B(new_n5892), .Y(new_n5893));
  nor_5  g03545(.A(n25565), .B(n24374), .Y(new_n5894));
  not_8  g03546(.A(n14575), .Y(new_n5895));
  nor_5  g03547(.A(new_n3635), .B(new_n5895), .Y(new_n5896));
  xnor_4 g03548(.A(n25565), .B(n24374), .Y(new_n5897));
  nor_5  g03549(.A(new_n5897), .B(new_n5896), .Y(new_n5898));
  or_5   g03550(.A(new_n5898), .B(new_n5894), .Y(new_n5899));
  and_5  g03551(.A(new_n5899), .B(new_n5893), .Y(new_n5900));
  or_5   g03552(.A(new_n5900), .B(new_n5891), .Y(new_n5901));
  and_5  g03553(.A(new_n5901), .B(new_n5890), .Y(new_n5902));
  or_5   g03554(.A(new_n5902), .B(new_n5888), .Y(new_n5903_1));
  and_5  g03555(.A(new_n5903_1), .B(new_n5887), .Y(new_n5904_1));
  or_5   g03556(.A(new_n5904_1), .B(new_n5885), .Y(new_n5905));
  and_5  g03557(.A(new_n5905), .B(new_n5884), .Y(new_n5906));
  or_5   g03558(.A(new_n5906), .B(new_n5882_1), .Y(new_n5907));
  and_5  g03559(.A(new_n5907), .B(new_n5881), .Y(new_n5908));
  or_5   g03560(.A(new_n5908), .B(new_n5879), .Y(new_n5909));
  and_5  g03561(.A(new_n5909), .B(new_n5878), .Y(new_n5910));
  or_5   g03562(.A(new_n5910), .B(new_n5877), .Y(new_n5911_1));
  and_5  g03563(.A(new_n5911_1), .B(new_n5876), .Y(new_n5912));
  nor_5  g03564(.A(new_n5912), .B(new_n5874), .Y(new_n5913));
  xnor_4 g03565(.A(new_n5913), .B(new_n5873), .Y(new_n5914));
  not_8  g03566(.A(new_n5914), .Y(new_n5915));
  xnor_4 g03567(.A(new_n5915), .B(new_n5871), .Y(new_n5916));
  xnor_4 g03568(.A(new_n5868), .B(n647), .Y(new_n5917));
  nor_5  g03569(.A(new_n5910), .B(new_n5877), .Y(new_n5918));
  xnor_4 g03570(.A(new_n5918), .B(new_n5876), .Y(new_n5919));
  and_5  g03571(.A(new_n5919), .B(new_n5917), .Y(new_n5920));
  not_8  g03572(.A(new_n5919), .Y(new_n5921));
  xnor_4 g03573(.A(new_n5921), .B(new_n5917), .Y(new_n5922));
  xnor_4 g03574(.A(new_n5866), .B(n20409), .Y(new_n5923));
  nor_5  g03575(.A(new_n5908), .B(new_n5879), .Y(new_n5924));
  xnor_4 g03576(.A(new_n5924), .B(new_n5878), .Y(new_n5925));
  nor_5  g03577(.A(new_n5925), .B(new_n5923), .Y(new_n5926));
  xnor_4 g03578(.A(new_n5925), .B(new_n5923), .Y(new_n5927));
  xnor_4 g03579(.A(new_n5864), .B(n25749), .Y(new_n5928));
  nor_5  g03580(.A(new_n5906), .B(new_n5882_1), .Y(new_n5929));
  xnor_4 g03581(.A(new_n5929), .B(new_n5881), .Y(new_n5930));
  nor_5  g03582(.A(new_n5930), .B(new_n5928), .Y(new_n5931));
  xnor_4 g03583(.A(new_n5930), .B(new_n5928), .Y(new_n5932));
  xnor_4 g03584(.A(new_n5862), .B(n3161), .Y(new_n5933));
  nor_5  g03585(.A(new_n5904_1), .B(new_n5885), .Y(new_n5934));
  xnor_4 g03586(.A(new_n5934), .B(new_n5884), .Y(new_n5935));
  nor_5  g03587(.A(new_n5935), .B(new_n5933), .Y(new_n5936_1));
  xnor_4 g03588(.A(new_n5935), .B(new_n5933), .Y(new_n5937));
  xnor_4 g03589(.A(new_n5860), .B(n9003), .Y(new_n5938));
  nor_5  g03590(.A(new_n5902), .B(new_n5888), .Y(new_n5939));
  xnor_4 g03591(.A(new_n5939), .B(new_n5887), .Y(new_n5940));
  nor_5  g03592(.A(new_n5940), .B(new_n5938), .Y(new_n5941));
  xnor_4 g03593(.A(new_n5940), .B(new_n5938), .Y(new_n5942));
  xnor_4 g03594(.A(new_n5858), .B(n4957), .Y(new_n5943_1));
  nor_5  g03595(.A(new_n5900), .B(new_n5891), .Y(new_n5944));
  xnor_4 g03596(.A(new_n5944), .B(new_n5890), .Y(new_n5945));
  nor_5  g03597(.A(new_n5945), .B(new_n5943_1), .Y(new_n5946));
  not_8  g03598(.A(new_n5945), .Y(new_n5947));
  xnor_4 g03599(.A(new_n5947), .B(new_n5943_1), .Y(new_n5948));
  xnor_4 g03600(.A(new_n5856), .B(n7524), .Y(new_n5949));
  not_8  g03601(.A(new_n5949), .Y(new_n5950));
  nor_5  g03602(.A(new_n5898), .B(new_n5894), .Y(new_n5951));
  xnor_4 g03603(.A(new_n5951), .B(new_n5893), .Y(new_n5952));
  not_8  g03604(.A(new_n5952), .Y(new_n5953));
  nor_5  g03605(.A(new_n5953), .B(new_n5950), .Y(new_n5954));
  xnor_4 g03606(.A(new_n5953), .B(new_n5949), .Y(new_n5955));
  xnor_4 g03607(.A(n21993), .B(n14575), .Y(new_n5956));
  nor_5  g03608(.A(new_n5956), .B(n20658), .Y(new_n5957));
  and_5  g03609(.A(new_n5957), .B(new_n3794_1), .Y(new_n5958));
  xnor_4 g03610(.A(new_n5897), .B(new_n5896), .Y(new_n5959));
  xnor_4 g03611(.A(n20658), .B(new_n3794_1), .Y(new_n5960));
  not_8  g03612(.A(new_n5960), .Y(new_n5961));
  nor_5  g03613(.A(new_n5961), .B(new_n5957), .Y(new_n5962));
  nor_5  g03614(.A(new_n5962), .B(new_n5958), .Y(new_n5963));
  and_5  g03615(.A(new_n5963), .B(new_n5959), .Y(new_n5964_1));
  nor_5  g03616(.A(new_n5964_1), .B(new_n5958), .Y(new_n5965));
  and_5  g03617(.A(new_n5965), .B(new_n5955), .Y(new_n5966));
  nor_5  g03618(.A(new_n5966), .B(new_n5954), .Y(new_n5967));
  and_5  g03619(.A(new_n5967), .B(new_n5948), .Y(new_n5968));
  nor_5  g03620(.A(new_n5968), .B(new_n5946), .Y(new_n5969));
  nor_5  g03621(.A(new_n5969), .B(new_n5942), .Y(new_n5970));
  nor_5  g03622(.A(new_n5970), .B(new_n5941), .Y(new_n5971));
  nor_5  g03623(.A(new_n5971), .B(new_n5937), .Y(new_n5972));
  nor_5  g03624(.A(new_n5972), .B(new_n5936_1), .Y(new_n5973));
  nor_5  g03625(.A(new_n5973), .B(new_n5932), .Y(new_n5974));
  nor_5  g03626(.A(new_n5974), .B(new_n5931), .Y(new_n5975));
  nor_5  g03627(.A(new_n5975), .B(new_n5927), .Y(new_n5976));
  nor_5  g03628(.A(new_n5976), .B(new_n5926), .Y(new_n5977));
  and_5  g03629(.A(new_n5977), .B(new_n5922), .Y(new_n5978));
  or_5   g03630(.A(new_n5978), .B(new_n5920), .Y(new_n5979));
  xor_4  g03631(.A(new_n5979), .B(new_n5916), .Y(new_n5980_1));
  not_8  g03632(.A(n8526), .Y(new_n5981));
  not_8  g03633(.A(n3582), .Y(new_n5982));
  xnor_4 g03634(.A(n21784), .B(new_n5982), .Y(new_n5983));
  nor_5  g03635(.A(n5521), .B(n2145), .Y(new_n5984));
  not_8  g03636(.A(n2145), .Y(new_n5985));
  xnor_4 g03637(.A(n5521), .B(new_n5985), .Y(new_n5986));
  nor_5  g03638(.A(n11926), .B(n5031), .Y(new_n5987));
  not_8  g03639(.A(n5031), .Y(new_n5988));
  xnor_4 g03640(.A(n11926), .B(new_n5988), .Y(new_n5989));
  nor_5  g03641(.A(n11044), .B(n4325), .Y(new_n5990));
  not_8  g03642(.A(n4325), .Y(new_n5991));
  xnor_4 g03643(.A(n11044), .B(new_n5991), .Y(new_n5992));
  nor_5  g03644(.A(n5337), .B(n2421), .Y(new_n5993));
  not_8  g03645(.A(n2421), .Y(new_n5994));
  xnor_4 g03646(.A(n5337), .B(new_n5994), .Y(new_n5995));
  nor_5  g03647(.A(n987), .B(n626), .Y(new_n5996));
  xnor_4 g03648(.A(n987), .B(new_n4223), .Y(new_n5997));
  nor_5  g03649(.A(n20478), .B(n1204), .Y(new_n5998));
  xnor_4 g03650(.A(n20478), .B(new_n4233), .Y(new_n5999));
  nor_5  g03651(.A(n26882), .B(n19618), .Y(new_n6000));
  xnor_4 g03652(.A(n26882), .B(new_n4237), .Y(new_n6001));
  nor_5  g03653(.A(n22619), .B(n22043), .Y(new_n6002));
  not_8  g03654(.A(n6775), .Y(new_n6003));
  nor_5  g03655(.A(new_n3875), .B(new_n6003), .Y(new_n6004));
  xnor_4 g03656(.A(n22619), .B(n22043), .Y(new_n6005));
  nor_5  g03657(.A(new_n6005), .B(new_n6004), .Y(new_n6006));
  or_5   g03658(.A(new_n6006), .B(new_n6002), .Y(new_n6007));
  and_5  g03659(.A(new_n6007), .B(new_n6001), .Y(new_n6008));
  or_5   g03660(.A(new_n6008), .B(new_n6000), .Y(new_n6009));
  and_5  g03661(.A(new_n6009), .B(new_n5999), .Y(new_n6010));
  or_5   g03662(.A(new_n6010), .B(new_n5998), .Y(new_n6011));
  and_5  g03663(.A(new_n6011), .B(new_n5997), .Y(new_n6012_1));
  or_5   g03664(.A(new_n6012_1), .B(new_n5996), .Y(new_n6013));
  and_5  g03665(.A(new_n6013), .B(new_n5995), .Y(new_n6014));
  or_5   g03666(.A(new_n6014), .B(new_n5993), .Y(new_n6015));
  and_5  g03667(.A(new_n6015), .B(new_n5992), .Y(new_n6016));
  or_5   g03668(.A(new_n6016), .B(new_n5990), .Y(new_n6017));
  and_5  g03669(.A(new_n6017), .B(new_n5989), .Y(new_n6018));
  or_5   g03670(.A(new_n6018), .B(new_n5987), .Y(new_n6019));
  and_5  g03671(.A(new_n6019), .B(new_n5986), .Y(new_n6020));
  nor_5  g03672(.A(new_n6020), .B(new_n5984), .Y(new_n6021));
  xnor_4 g03673(.A(new_n6021), .B(new_n5983), .Y(new_n6022_1));
  not_8  g03674(.A(new_n6022_1), .Y(new_n6023));
  xnor_4 g03675(.A(new_n6023), .B(new_n5981), .Y(new_n6024));
  not_8  g03676(.A(n2816), .Y(new_n6025));
  nor_5  g03677(.A(new_n6018), .B(new_n5987), .Y(new_n6026));
  xnor_4 g03678(.A(new_n6026), .B(new_n5986), .Y(new_n6027));
  nor_5  g03679(.A(new_n6027), .B(new_n6025), .Y(new_n6028));
  not_8  g03680(.A(new_n6027), .Y(new_n6029));
  xnor_4 g03681(.A(new_n6029), .B(new_n6025), .Y(new_n6030));
  not_8  g03682(.A(n20359), .Y(new_n6031_1));
  nor_5  g03683(.A(new_n6016), .B(new_n5990), .Y(new_n6032));
  xnor_4 g03684(.A(new_n6032), .B(new_n5989), .Y(new_n6033));
  nor_5  g03685(.A(new_n6033), .B(new_n6031_1), .Y(new_n6034));
  not_8  g03686(.A(new_n6033), .Y(new_n6035));
  xnor_4 g03687(.A(new_n6035), .B(new_n6031_1), .Y(new_n6036));
  not_8  g03688(.A(n4409), .Y(new_n6037));
  nor_5  g03689(.A(new_n6014), .B(new_n5993), .Y(new_n6038));
  xnor_4 g03690(.A(new_n6038), .B(new_n5992), .Y(new_n6039));
  nor_5  g03691(.A(new_n6039), .B(new_n6037), .Y(new_n6040));
  not_8  g03692(.A(new_n6039), .Y(new_n6041));
  xnor_4 g03693(.A(new_n6041), .B(new_n6037), .Y(new_n6042));
  not_8  g03694(.A(n3570), .Y(new_n6043));
  nor_5  g03695(.A(new_n6012_1), .B(new_n5996), .Y(new_n6044_1));
  xnor_4 g03696(.A(new_n6044_1), .B(new_n5995), .Y(new_n6045));
  nor_5  g03697(.A(new_n6045), .B(new_n6043), .Y(new_n6046_1));
  not_8  g03698(.A(new_n6045), .Y(new_n6047));
  xnor_4 g03699(.A(new_n6047), .B(new_n6043), .Y(new_n6048));
  not_8  g03700(.A(n13668), .Y(new_n6049));
  nor_5  g03701(.A(new_n6010), .B(new_n5998), .Y(new_n6050));
  xnor_4 g03702(.A(new_n6050), .B(new_n5997), .Y(new_n6051));
  nor_5  g03703(.A(new_n6051), .B(new_n6049), .Y(new_n6052));
  not_8  g03704(.A(new_n6051), .Y(new_n6053));
  xnor_4 g03705(.A(new_n6053), .B(new_n6049), .Y(new_n6054));
  not_8  g03706(.A(n21276), .Y(new_n6055));
  nor_5  g03707(.A(new_n6008), .B(new_n6000), .Y(new_n6056));
  xnor_4 g03708(.A(new_n6056), .B(new_n5999), .Y(new_n6057));
  nor_5  g03709(.A(new_n6057), .B(new_n6055), .Y(new_n6058));
  not_8  g03710(.A(new_n6057), .Y(new_n6059));
  xnor_4 g03711(.A(new_n6059), .B(new_n6055), .Y(new_n6060));
  not_8  g03712(.A(n26748), .Y(new_n6061));
  nor_5  g03713(.A(new_n6006), .B(new_n6002), .Y(new_n6062));
  xnor_4 g03714(.A(new_n6062), .B(new_n6001), .Y(new_n6063));
  nor_5  g03715(.A(new_n6063), .B(new_n6061), .Y(new_n6064));
  xnor_4 g03716(.A(new_n6005), .B(new_n6004), .Y(new_n6065));
  nor_5  g03717(.A(new_n6065), .B(n10057), .Y(new_n6066));
  or_5   g03718(.A(new_n5792), .B(new_n4242), .Y(new_n6067));
  not_8  g03719(.A(n10057), .Y(new_n6068));
  xnor_4 g03720(.A(new_n6065), .B(new_n6068), .Y(new_n6069));
  and_5  g03721(.A(new_n6069), .B(new_n6067), .Y(new_n6070));
  nor_5  g03722(.A(new_n6070), .B(new_n6066), .Y(new_n6071));
  not_8  g03723(.A(new_n6063), .Y(new_n6072));
  xnor_4 g03724(.A(new_n6072), .B(new_n6061), .Y(new_n6073));
  and_5  g03725(.A(new_n6073), .B(new_n6071), .Y(new_n6074));
  or_5   g03726(.A(new_n6074), .B(new_n6064), .Y(new_n6075));
  and_5  g03727(.A(new_n6075), .B(new_n6060), .Y(new_n6076));
  or_5   g03728(.A(new_n6076), .B(new_n6058), .Y(new_n6077));
  and_5  g03729(.A(new_n6077), .B(new_n6054), .Y(new_n6078));
  or_5   g03730(.A(new_n6078), .B(new_n6052), .Y(new_n6079));
  and_5  g03731(.A(new_n6079), .B(new_n6048), .Y(new_n6080));
  or_5   g03732(.A(new_n6080), .B(new_n6046_1), .Y(new_n6081));
  and_5  g03733(.A(new_n6081), .B(new_n6042), .Y(new_n6082));
  or_5   g03734(.A(new_n6082), .B(new_n6040), .Y(new_n6083));
  and_5  g03735(.A(new_n6083), .B(new_n6036), .Y(new_n6084_1));
  or_5   g03736(.A(new_n6084_1), .B(new_n6034), .Y(new_n6085));
  and_5  g03737(.A(new_n6085), .B(new_n6030), .Y(new_n6086));
  nor_5  g03738(.A(new_n6086), .B(new_n6028), .Y(new_n6087));
  xnor_4 g03739(.A(new_n6087), .B(new_n6024), .Y(new_n6088));
  xnor_4 g03740(.A(new_n6088), .B(new_n5980_1), .Y(new_n6089));
  nor_5  g03741(.A(new_n6084_1), .B(new_n6034), .Y(new_n6090));
  xnor_4 g03742(.A(new_n6090), .B(new_n6030), .Y(new_n6091));
  xor_4  g03743(.A(new_n5977), .B(new_n5922), .Y(new_n6092));
  nor_5  g03744(.A(new_n6092), .B(new_n6091), .Y(new_n6093));
  xnor_4 g03745(.A(new_n6092), .B(new_n6091), .Y(new_n6094));
  xnor_4 g03746(.A(new_n5975), .B(new_n5927), .Y(new_n6095));
  nor_5  g03747(.A(new_n6082), .B(new_n6040), .Y(new_n6096));
  xnor_4 g03748(.A(new_n6096), .B(new_n6036), .Y(new_n6097));
  nor_5  g03749(.A(new_n6097), .B(new_n6095), .Y(new_n6098));
  xnor_4 g03750(.A(new_n6097), .B(new_n6095), .Y(new_n6099));
  xnor_4 g03751(.A(new_n5973), .B(new_n5932), .Y(new_n6100));
  nor_5  g03752(.A(new_n6080), .B(new_n6046_1), .Y(new_n6101));
  xnor_4 g03753(.A(new_n6101), .B(new_n6042), .Y(new_n6102));
  nor_5  g03754(.A(new_n6102), .B(new_n6100), .Y(new_n6103));
  xnor_4 g03755(.A(new_n6102), .B(new_n6100), .Y(new_n6104_1));
  xnor_4 g03756(.A(new_n5971), .B(new_n5937), .Y(new_n6105_1));
  nor_5  g03757(.A(new_n6078), .B(new_n6052), .Y(new_n6106));
  xnor_4 g03758(.A(new_n6106), .B(new_n6048), .Y(new_n6107));
  nor_5  g03759(.A(new_n6107), .B(new_n6105_1), .Y(new_n6108));
  xnor_4 g03760(.A(new_n6107), .B(new_n6105_1), .Y(new_n6109));
  xnor_4 g03761(.A(new_n5969), .B(new_n5942), .Y(new_n6110));
  nor_5  g03762(.A(new_n6076), .B(new_n6058), .Y(new_n6111));
  xnor_4 g03763(.A(new_n6111), .B(new_n6054), .Y(new_n6112));
  nor_5  g03764(.A(new_n6112), .B(new_n6110), .Y(new_n6113));
  xnor_4 g03765(.A(new_n6112), .B(new_n6110), .Y(new_n6114));
  xnor_4 g03766(.A(new_n5967), .B(new_n5948), .Y(new_n6115));
  xor_4  g03767(.A(new_n6075), .B(new_n6060), .Y(new_n6116));
  nor_5  g03768(.A(new_n6116), .B(new_n6115), .Y(new_n6117));
  xnor_4 g03769(.A(new_n6116), .B(new_n6115), .Y(new_n6118));
  xnor_4 g03770(.A(new_n5965), .B(new_n5955), .Y(new_n6119));
  not_8  g03771(.A(new_n6119), .Y(new_n6120));
  xnor_4 g03772(.A(new_n6073), .B(new_n6071), .Y(new_n6121));
  not_8  g03773(.A(new_n6121), .Y(new_n6122));
  nor_5  g03774(.A(new_n6122), .B(new_n6120), .Y(new_n6123));
  xnor_4 g03775(.A(new_n6121), .B(new_n6120), .Y(new_n6124));
  nor_5  g03776(.A(new_n5792), .B(new_n4242), .Y(new_n6125));
  xnor_4 g03777(.A(new_n6069), .B(new_n6125), .Y(new_n6126));
  not_8  g03778(.A(new_n5959), .Y(new_n6127));
  xnor_4 g03779(.A(new_n5963), .B(new_n6127), .Y(new_n6128));
  nor_5  g03780(.A(new_n6128), .B(new_n6126), .Y(new_n6129));
  xnor_4 g03781(.A(new_n5956), .B(new_n3798), .Y(new_n6130));
  nor_5  g03782(.A(new_n6130), .B(new_n5794), .Y(new_n6131));
  not_8  g03783(.A(new_n6126), .Y(new_n6132));
  xnor_4 g03784(.A(new_n6128), .B(new_n6132), .Y(new_n6133));
  and_5  g03785(.A(new_n6133), .B(new_n6131), .Y(new_n6134));
  nor_5  g03786(.A(new_n6134), .B(new_n6129), .Y(new_n6135));
  and_5  g03787(.A(new_n6135), .B(new_n6124), .Y(new_n6136));
  nor_5  g03788(.A(new_n6136), .B(new_n6123), .Y(new_n6137));
  nor_5  g03789(.A(new_n6137), .B(new_n6118), .Y(new_n6138));
  nor_5  g03790(.A(new_n6138), .B(new_n6117), .Y(new_n6139));
  nor_5  g03791(.A(new_n6139), .B(new_n6114), .Y(new_n6140));
  nor_5  g03792(.A(new_n6140), .B(new_n6113), .Y(new_n6141));
  nor_5  g03793(.A(new_n6141), .B(new_n6109), .Y(new_n6142));
  nor_5  g03794(.A(new_n6142), .B(new_n6108), .Y(new_n6143));
  nor_5  g03795(.A(new_n6143), .B(new_n6104_1), .Y(new_n6144));
  nor_5  g03796(.A(new_n6144), .B(new_n6103), .Y(new_n6145));
  nor_5  g03797(.A(new_n6145), .B(new_n6099), .Y(new_n6146));
  nor_5  g03798(.A(new_n6146), .B(new_n6098), .Y(new_n6147));
  nor_5  g03799(.A(new_n6147), .B(new_n6094), .Y(new_n6148));
  nor_5  g03800(.A(new_n6148), .B(new_n6093), .Y(new_n6149));
  xnor_4 g03801(.A(new_n6149), .B(new_n6089), .Y(n567));
  nor_5  g03802(.A(n10250), .B(n1831), .Y(new_n6151));
  not_8  g03803(.A(n1831), .Y(new_n6152));
  xnor_4 g03804(.A(n10250), .B(new_n6152), .Y(new_n6153));
  nor_5  g03805(.A(n13137), .B(n7674), .Y(new_n6154));
  not_8  g03806(.A(n7674), .Y(new_n6155));
  xnor_4 g03807(.A(n13137), .B(new_n6155), .Y(new_n6156));
  nor_5  g03808(.A(n18452), .B(n6397), .Y(new_n6157));
  not_8  g03809(.A(n6397), .Y(new_n6158));
  xnor_4 g03810(.A(n18452), .B(new_n6158), .Y(new_n6159));
  nor_5  g03811(.A(n21317), .B(n19196), .Y(new_n6160_1));
  not_8  g03812(.A(n19196), .Y(new_n6161));
  xnor_4 g03813(.A(n21317), .B(new_n6161), .Y(new_n6162));
  nor_5  g03814(.A(n23586), .B(n12398), .Y(new_n6163));
  not_8  g03815(.A(n12398), .Y(new_n6164));
  xnor_4 g03816(.A(n23586), .B(new_n6164), .Y(new_n6165));
  nor_5  g03817(.A(n21226), .B(n19789), .Y(new_n6166));
  not_8  g03818(.A(n19789), .Y(new_n6167));
  xnor_4 g03819(.A(n21226), .B(new_n6167), .Y(new_n6168));
  nor_5  g03820(.A(n20169), .B(n4426), .Y(new_n6169));
  not_8  g03821(.A(n4426), .Y(new_n6170));
  xnor_4 g03822(.A(n20169), .B(new_n6170), .Y(new_n6171_1));
  nor_5  g03823(.A(n20036), .B(n8285), .Y(new_n6172));
  not_8  g03824(.A(n8285), .Y(new_n6173));
  xnor_4 g03825(.A(n20036), .B(new_n6173), .Y(new_n6174));
  nor_5  g03826(.A(n11192), .B(n6729), .Y(new_n6175));
  not_8  g03827(.A(n9380), .Y(new_n6176));
  or_5   g03828(.A(new_n2548), .B(new_n6176), .Y(new_n6177));
  not_8  g03829(.A(n6729), .Y(new_n6178));
  xnor_4 g03830(.A(n11192), .B(new_n6178), .Y(new_n6179));
  and_5  g03831(.A(new_n6179), .B(new_n6177), .Y(new_n6180));
  or_5   g03832(.A(new_n6180), .B(new_n6175), .Y(new_n6181));
  and_5  g03833(.A(new_n6181), .B(new_n6174), .Y(new_n6182));
  or_5   g03834(.A(new_n6182), .B(new_n6172), .Y(new_n6183_1));
  and_5  g03835(.A(new_n6183_1), .B(new_n6171_1), .Y(new_n6184));
  or_5   g03836(.A(new_n6184), .B(new_n6169), .Y(new_n6185));
  and_5  g03837(.A(new_n6185), .B(new_n6168), .Y(new_n6186));
  or_5   g03838(.A(new_n6186), .B(new_n6166), .Y(new_n6187));
  and_5  g03839(.A(new_n6187), .B(new_n6165), .Y(new_n6188));
  or_5   g03840(.A(new_n6188), .B(new_n6163), .Y(new_n6189_1));
  and_5  g03841(.A(new_n6189_1), .B(new_n6162), .Y(new_n6190));
  or_5   g03842(.A(new_n6190), .B(new_n6160_1), .Y(new_n6191));
  and_5  g03843(.A(new_n6191), .B(new_n6159), .Y(new_n6192));
  or_5   g03844(.A(new_n6192), .B(new_n6157), .Y(new_n6193));
  and_5  g03845(.A(new_n6193), .B(new_n6156), .Y(new_n6194));
  or_5   g03846(.A(new_n6194), .B(new_n6154), .Y(new_n6195));
  and_5  g03847(.A(new_n6195), .B(new_n6153), .Y(new_n6196));
  nor_5  g03848(.A(new_n6196), .B(new_n6151), .Y(new_n6197));
  not_8  g03849(.A(n8614), .Y(new_n6198));
  not_8  g03850(.A(new_n4011), .Y(new_n6199));
  nor_5  g03851(.A(new_n6199), .B(n25694), .Y(new_n6200));
  not_8  g03852(.A(new_n6200), .Y(new_n6201));
  nor_5  g03853(.A(new_n6201), .B(n13110), .Y(new_n6202));
  not_8  g03854(.A(new_n6202), .Y(new_n6203));
  nor_5  g03855(.A(new_n6203), .B(n1752), .Y(new_n6204_1));
  not_8  g03856(.A(new_n6204_1), .Y(new_n6205));
  nor_5  g03857(.A(new_n6205), .B(n1288), .Y(new_n6206));
  xnor_4 g03858(.A(new_n6206), .B(n3320), .Y(new_n6207));
  not_8  g03859(.A(new_n6207), .Y(new_n6208));
  nor_5  g03860(.A(new_n6208), .B(new_n6198), .Y(new_n6209));
  not_8  g03861(.A(new_n6206), .Y(new_n6210));
  nor_5  g03862(.A(new_n6210), .B(n3320), .Y(new_n6211));
  or_5   g03863(.A(new_n6207), .B(n8614), .Y(new_n6212));
  xnor_4 g03864(.A(new_n6204_1), .B(n1288), .Y(new_n6213));
  nor_5  g03865(.A(new_n6213), .B(n15182), .Y(new_n6214));
  not_8  g03866(.A(n15182), .Y(new_n6215));
  not_8  g03867(.A(new_n6213), .Y(new_n6216));
  xnor_4 g03868(.A(new_n6216), .B(new_n6215), .Y(new_n6217));
  xnor_4 g03869(.A(new_n6202), .B(n1752), .Y(new_n6218_1));
  nor_5  g03870(.A(new_n6218_1), .B(n27037), .Y(new_n6219));
  not_8  g03871(.A(new_n6218_1), .Y(new_n6220));
  xnor_4 g03872(.A(new_n6220), .B(n27037), .Y(new_n6221));
  not_8  g03873(.A(n8964), .Y(new_n6222));
  xnor_4 g03874(.A(new_n6200), .B(n13110), .Y(new_n6223_1));
  not_8  g03875(.A(new_n6223_1), .Y(new_n6224));
  nor_5  g03876(.A(new_n6224), .B(new_n6222), .Y(new_n6225));
  xnor_4 g03877(.A(new_n6224), .B(n8964), .Y(new_n6226));
  not_8  g03878(.A(n20151), .Y(new_n6227));
  nor_5  g03879(.A(new_n4013), .B(new_n6227), .Y(new_n6228));
  or_5   g03880(.A(new_n4041), .B(new_n4018), .Y(new_n6229));
  and_5  g03881(.A(new_n6229), .B(new_n4014_1), .Y(new_n6230));
  or_5   g03882(.A(new_n6230), .B(new_n6228), .Y(new_n6231));
  and_5  g03883(.A(new_n6231), .B(new_n6226), .Y(new_n6232));
  nor_5  g03884(.A(new_n6232), .B(new_n6225), .Y(new_n6233_1));
  and_5  g03885(.A(new_n6233_1), .B(new_n6221), .Y(new_n6234));
  nor_5  g03886(.A(new_n6234), .B(new_n6219), .Y(new_n6235));
  nor_5  g03887(.A(new_n6235), .B(new_n6217), .Y(new_n6236));
  nor_5  g03888(.A(new_n6236), .B(new_n6214), .Y(new_n6237));
  and_5  g03889(.A(new_n6237), .B(new_n6212), .Y(new_n6238));
  or_5   g03890(.A(new_n6238), .B(new_n6211), .Y(new_n6239));
  nor_5  g03891(.A(new_n6239), .B(new_n6209), .Y(new_n6240));
  nor_5  g03892(.A(new_n6240), .B(new_n6197), .Y(new_n6241));
  not_8  g03893(.A(new_n6197), .Y(new_n6242));
  xnor_4 g03894(.A(new_n6240), .B(new_n6242), .Y(new_n6243));
  xor_4  g03895(.A(new_n6195), .B(new_n6153), .Y(new_n6244));
  xnor_4 g03896(.A(new_n6208), .B(n8614), .Y(new_n6245_1));
  xnor_4 g03897(.A(new_n6245_1), .B(new_n6237), .Y(new_n6246));
  nor_5  g03898(.A(new_n6246), .B(new_n6244), .Y(new_n6247));
  xnor_4 g03899(.A(new_n6235), .B(new_n6217), .Y(new_n6248_1));
  nor_5  g03900(.A(new_n6192), .B(new_n6157), .Y(new_n6249));
  xnor_4 g03901(.A(new_n6249), .B(new_n6156), .Y(new_n6250));
  not_8  g03902(.A(new_n6250), .Y(new_n6251));
  nor_5  g03903(.A(new_n6251), .B(new_n6248_1), .Y(new_n6252));
  xnor_4 g03904(.A(new_n6250), .B(new_n6248_1), .Y(new_n6253));
  xnor_4 g03905(.A(new_n6233_1), .B(new_n6221), .Y(new_n6254));
  nor_5  g03906(.A(new_n6190), .B(new_n6160_1), .Y(new_n6255));
  xnor_4 g03907(.A(new_n6255), .B(new_n6159), .Y(new_n6256_1));
  not_8  g03908(.A(new_n6256_1), .Y(new_n6257));
  nor_5  g03909(.A(new_n6257), .B(new_n6254), .Y(new_n6258));
  not_8  g03910(.A(new_n6254), .Y(new_n6259));
  xnor_4 g03911(.A(new_n6257), .B(new_n6259), .Y(new_n6260));
  nor_5  g03912(.A(new_n6188), .B(new_n6163), .Y(new_n6261));
  xnor_4 g03913(.A(new_n6261), .B(new_n6162), .Y(new_n6262));
  nor_5  g03914(.A(new_n6230), .B(new_n6228), .Y(new_n6263));
  xnor_4 g03915(.A(new_n6263), .B(new_n6226), .Y(new_n6264));
  not_8  g03916(.A(new_n6264), .Y(new_n6265));
  nor_5  g03917(.A(new_n6265), .B(new_n6262), .Y(new_n6266));
  nor_5  g03918(.A(new_n6186), .B(new_n6166), .Y(new_n6267));
  xnor_4 g03919(.A(new_n6267), .B(new_n6165), .Y(new_n6268));
  not_8  g03920(.A(new_n6268), .Y(new_n6269));
  nor_5  g03921(.A(new_n6269), .B(new_n4043), .Y(new_n6270));
  xnor_4 g03922(.A(new_n6269), .B(new_n4044), .Y(new_n6271_1));
  nor_5  g03923(.A(new_n6184), .B(new_n6169), .Y(new_n6272));
  xnor_4 g03924(.A(new_n6272), .B(new_n6168), .Y(new_n6273));
  not_8  g03925(.A(new_n6273), .Y(new_n6274));
  nor_5  g03926(.A(new_n6182), .B(new_n6172), .Y(new_n6275));
  xnor_4 g03927(.A(new_n6275), .B(new_n6171_1), .Y(new_n6276_1));
  not_8  g03928(.A(new_n6276_1), .Y(new_n6277));
  nor_5  g03929(.A(new_n6277), .B(new_n4052), .Y(new_n6278));
  nor_5  g03930(.A(new_n6180), .B(new_n6175), .Y(new_n6279));
  xnor_4 g03931(.A(new_n6279), .B(new_n6174), .Y(new_n6280));
  nor_5  g03932(.A(new_n6280), .B(new_n4057), .Y(new_n6281));
  not_8  g03933(.A(new_n6280), .Y(new_n6282));
  xnor_4 g03934(.A(new_n6282), .B(new_n4058), .Y(new_n6283));
  nor_5  g03935(.A(new_n2548), .B(new_n6176), .Y(new_n6284));
  xnor_4 g03936(.A(new_n6179), .B(new_n6284), .Y(new_n6285));
  nor_5  g03937(.A(new_n6285), .B(new_n4064), .Y(new_n6286));
  xnor_4 g03938(.A(n21687), .B(new_n6176), .Y(new_n6287));
  not_8  g03939(.A(new_n6287), .Y(new_n6288));
  nor_5  g03940(.A(new_n6288), .B(new_n2549), .Y(new_n6289));
  xnor_4 g03941(.A(new_n6285), .B(new_n4067), .Y(new_n6290));
  and_5  g03942(.A(new_n6290), .B(new_n6289), .Y(new_n6291));
  nor_5  g03943(.A(new_n6291), .B(new_n6286), .Y(new_n6292));
  nor_5  g03944(.A(new_n6292), .B(new_n6283), .Y(new_n6293));
  nor_5  g03945(.A(new_n6293), .B(new_n6281), .Y(new_n6294));
  xnor_4 g03946(.A(new_n6276_1), .B(new_n4052), .Y(new_n6295));
  and_5  g03947(.A(new_n6295), .B(new_n6294), .Y(new_n6296));
  nor_5  g03948(.A(new_n6296), .B(new_n6278), .Y(new_n6297));
  nor_5  g03949(.A(new_n6297), .B(new_n6274), .Y(new_n6298));
  xnor_4 g03950(.A(new_n6297), .B(new_n6273), .Y(new_n6299));
  and_5  g03951(.A(new_n6299), .B(new_n4049), .Y(new_n6300));
  or_5   g03952(.A(new_n6300), .B(new_n6298), .Y(new_n6301));
  and_5  g03953(.A(new_n6301), .B(new_n6271_1), .Y(new_n6302));
  nor_5  g03954(.A(new_n6302), .B(new_n6270), .Y(new_n6303));
  not_8  g03955(.A(new_n6262), .Y(new_n6304));
  xnor_4 g03956(.A(new_n6265), .B(new_n6304), .Y(new_n6305));
  and_5  g03957(.A(new_n6305), .B(new_n6303), .Y(new_n6306));
  nor_5  g03958(.A(new_n6306), .B(new_n6266), .Y(new_n6307));
  and_5  g03959(.A(new_n6307), .B(new_n6260), .Y(new_n6308_1));
  or_5   g03960(.A(new_n6308_1), .B(new_n6258), .Y(new_n6309));
  and_5  g03961(.A(new_n6309), .B(new_n6253), .Y(new_n6310));
  nor_5  g03962(.A(new_n6310), .B(new_n6252), .Y(new_n6311_1));
  not_8  g03963(.A(new_n6246), .Y(new_n6312));
  xnor_4 g03964(.A(new_n6312), .B(new_n6244), .Y(new_n6313));
  and_5  g03965(.A(new_n6313), .B(new_n6311_1), .Y(new_n6314));
  nor_5  g03966(.A(new_n6314), .B(new_n6247), .Y(new_n6315));
  and_5  g03967(.A(new_n6315), .B(new_n6243), .Y(new_n6316));
  nor_5  g03968(.A(new_n6316), .B(new_n6241), .Y(new_n6317));
  xnor_4 g03969(.A(new_n6315), .B(new_n6243), .Y(new_n6318));
  nor_5  g03970(.A(n15766), .B(n6105), .Y(new_n6319));
  not_8  g03971(.A(n15766), .Y(new_n6320));
  xnor_4 g03972(.A(new_n6320), .B(n6105), .Y(new_n6321));
  nor_5  g03973(.A(n25629), .B(n3795), .Y(new_n6322));
  not_8  g03974(.A(n3795), .Y(new_n6323_1));
  xnor_4 g03975(.A(n25629), .B(new_n6323_1), .Y(new_n6324));
  nor_5  g03976(.A(n25464), .B(n7692), .Y(new_n6325));
  not_8  g03977(.A(n7692), .Y(new_n6326));
  xnor_4 g03978(.A(n25464), .B(new_n6326), .Y(new_n6327));
  nor_5  g03979(.A(n23039), .B(n4590), .Y(new_n6328));
  not_8  g03980(.A(n23039), .Y(new_n6329));
  xnor_4 g03981(.A(new_n6329), .B(n4590), .Y(new_n6330_1));
  nor_5  g03982(.A(n26752), .B(n13677), .Y(new_n6331));
  xnor_4 g03983(.A(n26752), .B(n13677), .Y(new_n6332));
  nor_5  g03984(.A(n18926), .B(n6513), .Y(new_n6333));
  not_8  g03985(.A(n6513), .Y(new_n6334));
  xnor_4 g03986(.A(n18926), .B(new_n6334), .Y(new_n6335));
  not_8  g03987(.A(n3918), .Y(new_n6336));
  nor_5  g03988(.A(new_n3967), .B(new_n6336), .Y(new_n6337));
  or_5   g03989(.A(n5451), .B(n3918), .Y(new_n6338));
  nor_5  g03990(.A(n5330), .B(n919), .Y(new_n6339_1));
  or_5   g03991(.A(new_n4149), .B(new_n4145), .Y(new_n6340));
  and_5  g03992(.A(new_n6340), .B(new_n4144), .Y(new_n6341));
  nor_5  g03993(.A(new_n6341), .B(new_n6339_1), .Y(new_n6342));
  and_5  g03994(.A(new_n6342), .B(new_n6338), .Y(new_n6343));
  nor_5  g03995(.A(new_n6343), .B(new_n6337), .Y(new_n6344));
  and_5  g03996(.A(new_n6344), .B(new_n6335), .Y(new_n6345));
  nor_5  g03997(.A(new_n6345), .B(new_n6333), .Y(new_n6346));
  nor_5  g03998(.A(new_n6346), .B(new_n6332), .Y(new_n6347));
  or_5   g03999(.A(new_n6347), .B(new_n6331), .Y(new_n6348));
  and_5  g04000(.A(new_n6348), .B(new_n6330_1), .Y(new_n6349));
  or_5   g04001(.A(new_n6349), .B(new_n6328), .Y(new_n6350));
  and_5  g04002(.A(new_n6350), .B(new_n6327), .Y(new_n6351));
  or_5   g04003(.A(new_n6351), .B(new_n6325), .Y(new_n6352));
  and_5  g04004(.A(new_n6352), .B(new_n6324), .Y(new_n6353));
  or_5   g04005(.A(new_n6353), .B(new_n6322), .Y(new_n6354_1));
  and_5  g04006(.A(new_n6354_1), .B(new_n6321), .Y(new_n6355));
  nor_5  g04007(.A(new_n6355), .B(new_n6319), .Y(new_n6356_1));
  not_8  g04008(.A(new_n6356_1), .Y(new_n6357));
  nor_5  g04009(.A(new_n6357), .B(new_n6318), .Y(new_n6358));
  xnor_4 g04010(.A(new_n6357), .B(new_n6318), .Y(new_n6359));
  nor_5  g04011(.A(new_n6353), .B(new_n6322), .Y(new_n6360));
  xnor_4 g04012(.A(new_n6360), .B(new_n6321), .Y(new_n6361));
  not_8  g04013(.A(new_n6361), .Y(new_n6362));
  xnor_4 g04014(.A(new_n6313), .B(new_n6311_1), .Y(new_n6363));
  and_5  g04015(.A(new_n6363), .B(new_n6362), .Y(new_n6364));
  xnor_4 g04016(.A(new_n6363), .B(new_n6362), .Y(new_n6365));
  xor_4  g04017(.A(new_n6309), .B(new_n6253), .Y(new_n6366));
  xor_4  g04018(.A(new_n6352), .B(new_n6324), .Y(new_n6367));
  not_8  g04019(.A(new_n6367), .Y(new_n6368));
  and_5  g04020(.A(new_n6368), .B(new_n6366), .Y(new_n6369_1));
  xnor_4 g04021(.A(new_n6368), .B(new_n6366), .Y(new_n6370));
  xnor_4 g04022(.A(new_n6307), .B(new_n6260), .Y(new_n6371));
  nor_5  g04023(.A(new_n6349), .B(new_n6328), .Y(new_n6372));
  xnor_4 g04024(.A(new_n6372), .B(new_n6327), .Y(new_n6373));
  nor_5  g04025(.A(new_n6373), .B(new_n6371), .Y(new_n6374));
  xnor_4 g04026(.A(new_n6373), .B(new_n6371), .Y(new_n6375_1));
  xor_4  g04027(.A(new_n6348), .B(new_n6330_1), .Y(new_n6376));
  not_8  g04028(.A(new_n6376), .Y(new_n6377));
  xnor_4 g04029(.A(new_n6305), .B(new_n6303), .Y(new_n6378));
  and_5  g04030(.A(new_n6378), .B(new_n6377), .Y(new_n6379_1));
  xnor_4 g04031(.A(new_n6378), .B(new_n6377), .Y(new_n6380));
  xor_4  g04032(.A(new_n6301), .B(new_n6271_1), .Y(new_n6381_1));
  xnor_4 g04033(.A(new_n6346), .B(new_n6332), .Y(new_n6382));
  and_5  g04034(.A(new_n6382), .B(new_n6381_1), .Y(new_n6383_1));
  xnor_4 g04035(.A(new_n6382), .B(new_n6381_1), .Y(new_n6384));
  xnor_4 g04036(.A(new_n6299), .B(new_n4049), .Y(new_n6385_1));
  xor_4  g04037(.A(new_n6344), .B(new_n6335), .Y(new_n6386));
  nor_5  g04038(.A(new_n6386), .B(new_n6385_1), .Y(new_n6387));
  xnor_4 g04039(.A(new_n6386), .B(new_n6385_1), .Y(new_n6388));
  xnor_4 g04040(.A(new_n6295), .B(new_n6294), .Y(new_n6389));
  xnor_4 g04041(.A(n5451), .B(new_n6336), .Y(new_n6390));
  xnor_4 g04042(.A(new_n6390), .B(new_n6342), .Y(new_n6391));
  nor_5  g04043(.A(new_n6391), .B(new_n6389), .Y(new_n6392));
  xnor_4 g04044(.A(new_n6391), .B(new_n6389), .Y(new_n6393));
  not_8  g04045(.A(new_n4151_1), .Y(new_n6394));
  xnor_4 g04046(.A(new_n6292), .B(new_n6283), .Y(new_n6395));
  and_5  g04047(.A(new_n6395), .B(new_n6394), .Y(new_n6396));
  xnor_4 g04048(.A(new_n6395), .B(new_n6394), .Y(new_n6397_1));
  xnor_4 g04049(.A(new_n6290), .B(new_n6289), .Y(new_n6398));
  not_8  g04050(.A(new_n6398), .Y(new_n6399));
  nor_5  g04051(.A(new_n6399), .B(new_n4155), .Y(new_n6400));
  xnor_4 g04052(.A(new_n6287), .B(new_n2549), .Y(new_n6401));
  nor_5  g04053(.A(new_n6401), .B(new_n4157), .Y(new_n6402));
  xnor_4 g04054(.A(new_n6399), .B(new_n4160), .Y(new_n6403));
  and_5  g04055(.A(new_n6403), .B(new_n6402), .Y(new_n6404));
  nor_5  g04056(.A(new_n6404), .B(new_n6400), .Y(new_n6405));
  nor_5  g04057(.A(new_n6405), .B(new_n6397_1), .Y(new_n6406));
  nor_5  g04058(.A(new_n6406), .B(new_n6396), .Y(new_n6407_1));
  nor_5  g04059(.A(new_n6407_1), .B(new_n6393), .Y(new_n6408));
  nor_5  g04060(.A(new_n6408), .B(new_n6392), .Y(new_n6409));
  nor_5  g04061(.A(new_n6409), .B(new_n6388), .Y(new_n6410));
  nor_5  g04062(.A(new_n6410), .B(new_n6387), .Y(new_n6411));
  nor_5  g04063(.A(new_n6411), .B(new_n6384), .Y(new_n6412));
  nor_5  g04064(.A(new_n6412), .B(new_n6383_1), .Y(new_n6413));
  nor_5  g04065(.A(new_n6413), .B(new_n6380), .Y(new_n6414));
  nor_5  g04066(.A(new_n6414), .B(new_n6379_1), .Y(new_n6415));
  nor_5  g04067(.A(new_n6415), .B(new_n6375_1), .Y(new_n6416));
  nor_5  g04068(.A(new_n6416), .B(new_n6374), .Y(new_n6417));
  nor_5  g04069(.A(new_n6417), .B(new_n6370), .Y(new_n6418));
  nor_5  g04070(.A(new_n6418), .B(new_n6369_1), .Y(new_n6419));
  nor_5  g04071(.A(new_n6419), .B(new_n6365), .Y(new_n6420));
  nor_5  g04072(.A(new_n6420), .B(new_n6364), .Y(new_n6421));
  nor_5  g04073(.A(new_n6421), .B(new_n6359), .Y(new_n6422));
  nor_5  g04074(.A(new_n6422), .B(new_n6358), .Y(new_n6423));
  nor_5  g04075(.A(new_n6423), .B(new_n6317), .Y(n588));
  xnor_4 g04076(.A(n19803), .B(n18584), .Y(new_n6425));
  not_8  g04077(.A(n12626), .Y(new_n6426));
  nor_5  g04078(.A(new_n6426), .B(n4272), .Y(new_n6427_1));
  and_5  g04079(.A(new_n4684), .B(new_n4661), .Y(new_n6428));
  nor_5  g04080(.A(new_n6428), .B(new_n6427_1), .Y(new_n6429));
  xnor_4 g04081(.A(new_n6429), .B(new_n6425), .Y(new_n6430));
  not_8  g04082(.A(new_n6430), .Y(new_n6431_1));
  xnor_4 g04083(.A(n16911), .B(n7773), .Y(new_n6432));
  not_8  g04084(.A(n376), .Y(new_n6433));
  nor_5  g04085(.A(n7721), .B(new_n6433), .Y(new_n6434));
  xnor_4 g04086(.A(n7721), .B(n376), .Y(new_n6435));
  not_8  g04087(.A(n5517), .Y(new_n6436));
  nor_5  g04088(.A(n21981), .B(new_n6436), .Y(new_n6437_1));
  xnor_4 g04089(.A(n21981), .B(n5517), .Y(new_n6438));
  not_8  g04090(.A(n12113), .Y(new_n6439));
  nor_5  g04091(.A(n12917), .B(new_n6439), .Y(new_n6440));
  xnor_4 g04092(.A(n12917), .B(n12113), .Y(new_n6441));
  not_8  g04093(.A(n10614), .Y(new_n6442));
  and_5  g04094(.A(n21898), .B(new_n6442), .Y(new_n6443));
  nor_5  g04095(.A(n21898), .B(new_n6442), .Y(new_n6444));
  not_8  g04096(.A(n11266), .Y(new_n6445));
  and_5  g04097(.A(new_n6445), .B(n9926), .Y(new_n6446));
  nor_5  g04098(.A(new_n6445), .B(n9926), .Y(new_n6447));
  not_8  g04099(.A(n22072), .Y(new_n6448));
  nor_5  g04100(.A(new_n6448), .B(n2646), .Y(new_n6449));
  not_8  g04101(.A(new_n6449), .Y(new_n6450));
  nor_5  g04102(.A(new_n6450), .B(new_n6447), .Y(new_n6451));
  nor_5  g04103(.A(new_n6451), .B(new_n6446), .Y(new_n6452));
  nor_5  g04104(.A(new_n6452), .B(new_n6444), .Y(new_n6453));
  nor_5  g04105(.A(new_n6453), .B(new_n6443), .Y(new_n6454));
  and_5  g04106(.A(new_n6454), .B(new_n6441), .Y(new_n6455));
  or_5   g04107(.A(new_n6455), .B(new_n6440), .Y(new_n6456_1));
  and_5  g04108(.A(new_n6456_1), .B(new_n6438), .Y(new_n6457_1));
  or_5   g04109(.A(new_n6457_1), .B(new_n6437_1), .Y(new_n6458));
  and_5  g04110(.A(new_n6458), .B(new_n6435), .Y(new_n6459));
  or_5   g04111(.A(new_n6459), .B(new_n6434), .Y(new_n6460));
  xor_4  g04112(.A(new_n6460), .B(new_n6432), .Y(new_n6461));
  nor_5  g04113(.A(n15652), .B(n4939), .Y(new_n6462));
  not_8  g04114(.A(new_n6462), .Y(new_n6463));
  nor_5  g04115(.A(new_n6463), .B(n5605), .Y(new_n6464));
  not_8  g04116(.A(new_n6464), .Y(new_n6465_1));
  nor_5  g04117(.A(new_n6465_1), .B(n2985), .Y(new_n6466));
  not_8  g04118(.A(new_n6466), .Y(new_n6467));
  nor_5  g04119(.A(new_n6467), .B(n14576), .Y(new_n6468));
  not_8  g04120(.A(new_n6468), .Y(new_n6469));
  nor_5  g04121(.A(new_n6469), .B(n1269), .Y(new_n6470_1));
  xnor_4 g04122(.A(new_n6470_1), .B(n16818), .Y(new_n6471));
  not_8  g04123(.A(new_n6471), .Y(new_n6472));
  xnor_4 g04124(.A(new_n6472), .B(n1742), .Y(new_n6473));
  xnor_4 g04125(.A(new_n6468), .B(n1269), .Y(new_n6474));
  nor_5  g04126(.A(new_n6474), .B(n4858), .Y(new_n6475));
  not_8  g04127(.A(new_n6474), .Y(new_n6476_1));
  xnor_4 g04128(.A(new_n6476_1), .B(n4858), .Y(new_n6477));
  xnor_4 g04129(.A(new_n6466), .B(n14576), .Y(new_n6478));
  nor_5  g04130(.A(new_n6478), .B(n8244), .Y(new_n6479));
  not_8  g04131(.A(new_n6478), .Y(new_n6480));
  xnor_4 g04132(.A(new_n6480), .B(n8244), .Y(new_n6481));
  xnor_4 g04133(.A(new_n6464), .B(n2985), .Y(new_n6482));
  nor_5  g04134(.A(new_n6482), .B(n9493), .Y(new_n6483));
  xnor_4 g04135(.A(new_n6462), .B(n5605), .Y(new_n6484));
  nor_5  g04136(.A(new_n6484), .B(n15167), .Y(new_n6485_1));
  not_8  g04137(.A(new_n6484), .Y(new_n6486));
  xnor_4 g04138(.A(new_n6486), .B(n15167), .Y(new_n6487));
  xnor_4 g04139(.A(n15652), .B(n4939), .Y(new_n6488));
  not_8  g04140(.A(new_n6488), .Y(new_n6489));
  nor_5  g04141(.A(new_n6489), .B(n21095), .Y(new_n6490));
  not_8  g04142(.A(n4939), .Y(new_n6491));
  not_8  g04143(.A(n8656), .Y(new_n6492));
  or_5   g04144(.A(new_n6492), .B(new_n6491), .Y(new_n6493));
  xnor_4 g04145(.A(new_n6488), .B(n21095), .Y(new_n6494));
  and_5  g04146(.A(new_n6494), .B(new_n6493), .Y(new_n6495));
  or_5   g04147(.A(new_n6495), .B(new_n6490), .Y(new_n6496));
  and_5  g04148(.A(new_n6496), .B(new_n6487), .Y(new_n6497));
  or_5   g04149(.A(new_n6497), .B(new_n6485_1), .Y(new_n6498));
  not_8  g04150(.A(new_n6482), .Y(new_n6499));
  xnor_4 g04151(.A(new_n6499), .B(n9493), .Y(new_n6500));
  and_5  g04152(.A(new_n6500), .B(new_n6498), .Y(new_n6501));
  or_5   g04153(.A(new_n6501), .B(new_n6483), .Y(new_n6502_1));
  and_5  g04154(.A(new_n6502_1), .B(new_n6481), .Y(new_n6503));
  or_5   g04155(.A(new_n6503), .B(new_n6479), .Y(new_n6504));
  and_5  g04156(.A(new_n6504), .B(new_n6477), .Y(new_n6505));
  nor_5  g04157(.A(new_n6505), .B(new_n6475), .Y(new_n6506_1));
  xnor_4 g04158(.A(new_n6506_1), .B(new_n6473), .Y(new_n6507));
  not_8  g04159(.A(new_n6507), .Y(new_n6508));
  xnor_4 g04160(.A(new_n6508), .B(new_n6461), .Y(new_n6509));
  xor_4  g04161(.A(new_n6458), .B(new_n6435), .Y(new_n6510));
  not_8  g04162(.A(new_n6510), .Y(new_n6511));
  nor_5  g04163(.A(new_n6503), .B(new_n6479), .Y(new_n6512));
  xnor_4 g04164(.A(new_n6512), .B(new_n6477), .Y(new_n6513_1));
  nor_5  g04165(.A(new_n6513_1), .B(new_n6511), .Y(new_n6514_1));
  xnor_4 g04166(.A(new_n6513_1), .B(new_n6510), .Y(new_n6515));
  xnor_4 g04167(.A(new_n6456_1), .B(new_n6438), .Y(new_n6516));
  nor_5  g04168(.A(new_n6501), .B(new_n6483), .Y(new_n6517));
  xnor_4 g04169(.A(new_n6517), .B(new_n6481), .Y(new_n6518));
  and_5  g04170(.A(new_n6518), .B(new_n6516), .Y(new_n6519));
  xor_4  g04171(.A(new_n6456_1), .B(new_n6438), .Y(new_n6520));
  xnor_4 g04172(.A(new_n6518), .B(new_n6520), .Y(new_n6521));
  xnor_4 g04173(.A(new_n6454), .B(new_n6441), .Y(new_n6522));
  nor_5  g04174(.A(new_n6497), .B(new_n6485_1), .Y(new_n6523));
  xnor_4 g04175(.A(new_n6500), .B(new_n6523), .Y(new_n6524));
  nor_5  g04176(.A(new_n6524), .B(new_n6522), .Y(new_n6525));
  xor_4  g04177(.A(new_n6496), .B(new_n6487), .Y(new_n6526));
  xnor_4 g04178(.A(n21898), .B(n10614), .Y(new_n6527));
  xnor_4 g04179(.A(new_n6527), .B(new_n6452), .Y(new_n6528));
  and_5  g04180(.A(new_n6528), .B(new_n6526), .Y(new_n6529));
  xnor_4 g04181(.A(new_n6528), .B(new_n6526), .Y(new_n6530));
  xnor_4 g04182(.A(n8656), .B(n4939), .Y(new_n6531));
  xnor_4 g04183(.A(n22072), .B(n2646), .Y(new_n6532));
  nor_5  g04184(.A(new_n6532), .B(new_n6531), .Y(new_n6533));
  xnor_4 g04185(.A(n11266), .B(n9926), .Y(new_n6534));
  xnor_4 g04186(.A(new_n6534), .B(new_n6450), .Y(new_n6535));
  not_8  g04187(.A(new_n6535), .Y(new_n6536));
  nor_5  g04188(.A(new_n6536), .B(new_n6533), .Y(new_n6537));
  xor_4  g04189(.A(new_n6494), .B(new_n6493), .Y(new_n6538));
  xnor_4 g04190(.A(new_n6535), .B(new_n6533), .Y(new_n6539));
  and_5  g04191(.A(new_n6539), .B(new_n6538), .Y(new_n6540));
  nor_5  g04192(.A(new_n6540), .B(new_n6537), .Y(new_n6541));
  nor_5  g04193(.A(new_n6541), .B(new_n6530), .Y(new_n6542_1));
  nor_5  g04194(.A(new_n6542_1), .B(new_n6529), .Y(new_n6543));
  xor_4  g04195(.A(new_n6524), .B(new_n6522), .Y(new_n6544));
  and_5  g04196(.A(new_n6544), .B(new_n6543), .Y(new_n6545));
  nor_5  g04197(.A(new_n6545), .B(new_n6525), .Y(new_n6546));
  and_5  g04198(.A(new_n6546), .B(new_n6521), .Y(new_n6547));
  nor_5  g04199(.A(new_n6547), .B(new_n6519), .Y(new_n6548));
  and_5  g04200(.A(new_n6548), .B(new_n6515), .Y(new_n6549));
  nor_5  g04201(.A(new_n6549), .B(new_n6514_1), .Y(new_n6550));
  xnor_4 g04202(.A(new_n6550), .B(new_n6509), .Y(new_n6551));
  not_8  g04203(.A(new_n6551), .Y(new_n6552));
  xnor_4 g04204(.A(new_n6552), .B(new_n6431_1), .Y(new_n6553));
  xor_4  g04205(.A(new_n6548), .B(new_n6515), .Y(new_n6554));
  nor_5  g04206(.A(new_n6554), .B(new_n4685), .Y(new_n6555));
  xnor_4 g04207(.A(new_n6554), .B(new_n4685), .Y(new_n6556_1));
  xnor_4 g04208(.A(new_n6546), .B(new_n6521), .Y(new_n6557));
  nor_5  g04209(.A(new_n6557), .B(new_n4688), .Y(new_n6558_1));
  xnor_4 g04210(.A(new_n6557), .B(new_n4688), .Y(new_n6559));
  xnor_4 g04211(.A(new_n6544), .B(new_n6543), .Y(new_n6560_1));
  not_8  g04212(.A(new_n6560_1), .Y(new_n6561));
  nor_5  g04213(.A(new_n6561), .B(new_n4694), .Y(new_n6562));
  xnor_4 g04214(.A(new_n6561), .B(new_n4694), .Y(new_n6563));
  xnor_4 g04215(.A(new_n6541), .B(new_n6530), .Y(new_n6564));
  nor_5  g04216(.A(new_n6564), .B(new_n4702), .Y(new_n6565));
  not_8  g04217(.A(new_n6564), .Y(new_n6566));
  xnor_4 g04218(.A(new_n6566), .B(new_n4701), .Y(new_n6567_1));
  xnor_4 g04219(.A(new_n6532), .B(new_n6531), .Y(new_n6568));
  or_5   g04220(.A(new_n6568), .B(new_n4711), .Y(new_n6569));
  and_5  g04221(.A(new_n6569), .B(new_n4708), .Y(new_n6570));
  xnor_4 g04222(.A(new_n6539), .B(new_n6538), .Y(new_n6571));
  not_8  g04223(.A(new_n6571), .Y(new_n6572));
  xor_4  g04224(.A(new_n6569), .B(new_n4708), .Y(new_n6573));
  and_5  g04225(.A(new_n6573), .B(new_n6572), .Y(new_n6574));
  nor_5  g04226(.A(new_n6574), .B(new_n6570), .Y(new_n6575));
  nor_5  g04227(.A(new_n6575), .B(new_n6567_1), .Y(new_n6576_1));
  nor_5  g04228(.A(new_n6576_1), .B(new_n6565), .Y(new_n6577));
  nor_5  g04229(.A(new_n6577), .B(new_n6563), .Y(new_n6578));
  nor_5  g04230(.A(new_n6578), .B(new_n6562), .Y(new_n6579));
  nor_5  g04231(.A(new_n6579), .B(new_n6559), .Y(new_n6580));
  nor_5  g04232(.A(new_n6580), .B(new_n6558_1), .Y(new_n6581));
  nor_5  g04233(.A(new_n6581), .B(new_n6556_1), .Y(new_n6582));
  nor_5  g04234(.A(new_n6582), .B(new_n6555), .Y(new_n6583));
  xor_4  g04235(.A(new_n6583), .B(new_n6553), .Y(n597));
  not_8  g04236(.A(n9646), .Y(new_n6585));
  xnor_4 g04237(.A(n25926), .B(new_n6585), .Y(new_n6586));
  xnor_4 g04238(.A(new_n6586), .B(n14230), .Y(new_n6587_1));
  xnor_4 g04239(.A(new_n6587_1), .B(new_n5802), .Y(n637));
  not_8  g04240(.A(n7421), .Y(new_n6589));
  not_8  g04241(.A(n10611), .Y(new_n6590_1));
  xnor_4 g04242(.A(n25797), .B(new_n6590_1), .Y(new_n6591));
  nor_5  g04243(.A(n15967), .B(n2783), .Y(new_n6592));
  not_8  g04244(.A(n2783), .Y(new_n6593));
  xnor_4 g04245(.A(n15967), .B(new_n6593), .Y(new_n6594));
  nor_5  g04246(.A(n15490), .B(n13319), .Y(new_n6595));
  not_8  g04247(.A(n18), .Y(new_n6596_1));
  nor_5  g04248(.A(new_n3756), .B(new_n6596_1), .Y(new_n6597));
  xnor_4 g04249(.A(n15490), .B(n13319), .Y(new_n6598));
  nor_5  g04250(.A(new_n6598), .B(new_n6597), .Y(new_n6599));
  or_5   g04251(.A(new_n6599), .B(new_n6595), .Y(new_n6600));
  and_5  g04252(.A(new_n6600), .B(new_n6594), .Y(new_n6601));
  nor_5  g04253(.A(new_n6601), .B(new_n6592), .Y(new_n6602));
  xnor_4 g04254(.A(new_n6602), .B(new_n6591), .Y(new_n6603));
  not_8  g04255(.A(new_n6603), .Y(new_n6604));
  xnor_4 g04256(.A(new_n6604), .B(new_n6589), .Y(new_n6605));
  not_8  g04257(.A(n19680), .Y(new_n6606));
  nor_5  g04258(.A(new_n6599), .B(new_n6595), .Y(new_n6607));
  xnor_4 g04259(.A(new_n6607), .B(new_n6594), .Y(new_n6608));
  nor_5  g04260(.A(new_n6608), .B(new_n6606), .Y(new_n6609));
  not_8  g04261(.A(new_n6608), .Y(new_n6610));
  xnor_4 g04262(.A(new_n6610), .B(new_n6606), .Y(new_n6611_1));
  xnor_4 g04263(.A(new_n6598), .B(new_n6597), .Y(new_n6612_1));
  nor_5  g04264(.A(new_n6612_1), .B(n2809), .Y(new_n6613));
  xnor_4 g04265(.A(n25435), .B(n18), .Y(new_n6614));
  or_5   g04266(.A(new_n6614), .B(new_n4818), .Y(new_n6615));
  not_8  g04267(.A(n2809), .Y(new_n6616));
  xnor_4 g04268(.A(new_n6612_1), .B(new_n6616), .Y(new_n6617));
  and_5  g04269(.A(new_n6617), .B(new_n6615), .Y(new_n6618));
  nor_5  g04270(.A(new_n6618), .B(new_n6613), .Y(new_n6619));
  and_5  g04271(.A(new_n6619), .B(new_n6611_1), .Y(new_n6620));
  or_5   g04272(.A(new_n6620), .B(new_n6609), .Y(new_n6621));
  xor_4  g04273(.A(new_n6621), .B(new_n6605), .Y(new_n6622));
  not_8  g04274(.A(new_n6622), .Y(new_n6623));
  xnor_4 g04275(.A(n18157), .B(n11056), .Y(new_n6624));
  nor_5  g04276(.A(n15271), .B(n12161), .Y(new_n6625));
  xnor_4 g04277(.A(n15271), .B(n12161), .Y(new_n6626));
  nor_5  g04278(.A(n25877), .B(n5026), .Y(new_n6627));
  not_8  g04279(.A(n8581), .Y(new_n6628_1));
  not_8  g04280(.A(n24323), .Y(new_n6629));
  nor_5  g04281(.A(new_n6629), .B(new_n6628_1), .Y(new_n6630_1));
  xnor_4 g04282(.A(n25877), .B(n5026), .Y(new_n6631_1));
  nor_5  g04283(.A(new_n6631_1), .B(new_n6630_1), .Y(new_n6632));
  nor_5  g04284(.A(new_n6632), .B(new_n6627), .Y(new_n6633));
  nor_5  g04285(.A(new_n6633), .B(new_n6626), .Y(new_n6634_1));
  nor_5  g04286(.A(new_n6634_1), .B(new_n6625), .Y(new_n6635));
  xnor_4 g04287(.A(new_n6635), .B(new_n6624), .Y(new_n6636));
  xnor_4 g04288(.A(new_n6636), .B(n20250), .Y(new_n6637));
  xnor_4 g04289(.A(new_n6633), .B(new_n6626), .Y(new_n6638));
  nor_5  g04290(.A(new_n6638), .B(n5822), .Y(new_n6639));
  xnor_4 g04291(.A(new_n6631_1), .B(new_n6630_1), .Y(new_n6640));
  nor_5  g04292(.A(new_n6640), .B(n26443), .Y(new_n6641));
  xnor_4 g04293(.A(n24323), .B(n8581), .Y(new_n6642));
  or_5   g04294(.A(new_n6642), .B(new_n4394), .Y(new_n6643));
  not_8  g04295(.A(n26443), .Y(new_n6644));
  xnor_4 g04296(.A(new_n6640), .B(new_n6644), .Y(new_n6645));
  and_5  g04297(.A(new_n6645), .B(new_n6643), .Y(new_n6646));
  or_5   g04298(.A(new_n6646), .B(new_n6641), .Y(new_n6647));
  xnor_4 g04299(.A(new_n6638), .B(new_n4384), .Y(new_n6648));
  and_5  g04300(.A(new_n6648), .B(new_n6647), .Y(new_n6649));
  nor_5  g04301(.A(new_n6649), .B(new_n6639), .Y(new_n6650));
  xnor_4 g04302(.A(new_n6650), .B(new_n6637), .Y(new_n6651));
  not_8  g04303(.A(new_n6651), .Y(new_n6652_1));
  xnor_4 g04304(.A(new_n6652_1), .B(new_n6623), .Y(new_n6653));
  xnor_4 g04305(.A(new_n6619), .B(new_n6611_1), .Y(new_n6654));
  xnor_4 g04306(.A(new_n6648), .B(new_n6647), .Y(new_n6655_1));
  and_5  g04307(.A(new_n6655_1), .B(new_n6654), .Y(new_n6656));
  xor_4  g04308(.A(new_n6648), .B(new_n6647), .Y(new_n6657));
  xnor_4 g04309(.A(new_n6657), .B(new_n6654), .Y(new_n6658));
  nor_5  g04310(.A(new_n6614), .B(new_n4818), .Y(new_n6659_1));
  xnor_4 g04311(.A(new_n6617), .B(new_n6659_1), .Y(new_n6660));
  nor_5  g04312(.A(new_n6642), .B(new_n4394), .Y(new_n6661));
  xnor_4 g04313(.A(new_n6645), .B(new_n6661), .Y(new_n6662));
  not_8  g04314(.A(new_n6662), .Y(new_n6663));
  nor_5  g04315(.A(new_n6663), .B(new_n6660), .Y(new_n6664));
  xnor_4 g04316(.A(new_n6614), .B(new_n4818), .Y(new_n6665));
  xnor_4 g04317(.A(new_n6642), .B(n1681), .Y(new_n6666));
  nor_5  g04318(.A(new_n6666), .B(new_n6665), .Y(new_n6667));
  not_8  g04319(.A(new_n6660), .Y(new_n6668));
  xnor_4 g04320(.A(new_n6663), .B(new_n6668), .Y(new_n6669_1));
  and_5  g04321(.A(new_n6669_1), .B(new_n6667), .Y(new_n6670));
  nor_5  g04322(.A(new_n6670), .B(new_n6664), .Y(new_n6671_1));
  and_5  g04323(.A(new_n6671_1), .B(new_n6658), .Y(new_n6672));
  nor_5  g04324(.A(new_n6672), .B(new_n6656), .Y(new_n6673_1));
  xnor_4 g04325(.A(new_n6673_1), .B(new_n6653), .Y(n646));
  nor_5  g04326(.A(n19494), .B(n2387), .Y(new_n6675));
  not_8  g04327(.A(new_n6675), .Y(new_n6676));
  nor_5  g04328(.A(new_n6676), .B(n16223), .Y(new_n6677));
  not_8  g04329(.A(new_n6677), .Y(new_n6678));
  nor_5  g04330(.A(new_n6678), .B(n26913), .Y(new_n6679));
  xnor_4 g04331(.A(new_n6679), .B(n21832), .Y(new_n6680));
  xnor_4 g04332(.A(new_n2466), .B(new_n5468), .Y(new_n6681));
  nor_5  g04333(.A(new_n2470), .B(new_n5471), .Y(new_n6682));
  xnor_4 g04334(.A(new_n2470), .B(new_n5471), .Y(new_n6683));
  nor_5  g04335(.A(new_n2473), .B(new_n5475), .Y(new_n6684_1));
  xnor_4 g04336(.A(new_n2475), .B(n12341), .Y(new_n6685));
  nor_5  g04337(.A(new_n2478), .B(n12384), .Y(new_n6686));
  and_5  g04338(.A(new_n6686), .B(new_n5478), .Y(new_n6687));
  xor_4  g04339(.A(new_n2480), .B(new_n2449), .Y(new_n6688));
  xnor_4 g04340(.A(new_n6686), .B(new_n5478), .Y(new_n6689));
  nor_5  g04341(.A(new_n6689), .B(new_n6688), .Y(new_n6690));
  or_5   g04342(.A(new_n6690), .B(new_n6687), .Y(new_n6691_1));
  nor_5  g04343(.A(new_n6691_1), .B(new_n6685), .Y(new_n6692));
  nor_5  g04344(.A(new_n6692), .B(new_n6684_1), .Y(new_n6693));
  nor_5  g04345(.A(new_n6693), .B(new_n6683), .Y(new_n6694));
  nor_5  g04346(.A(new_n6694), .B(new_n6682), .Y(new_n6695));
  xor_4  g04347(.A(new_n6695), .B(new_n6681), .Y(new_n6696));
  xnor_4 g04348(.A(new_n6696), .B(new_n6680), .Y(new_n6697));
  xnor_4 g04349(.A(new_n6677), .B(n26913), .Y(new_n6698));
  xor_4  g04350(.A(new_n6693), .B(new_n6683), .Y(new_n6699));
  and_5  g04351(.A(new_n6699), .B(new_n6698), .Y(new_n6700));
  xnor_4 g04352(.A(new_n6699), .B(new_n6698), .Y(new_n6701));
  xnor_4 g04353(.A(new_n2478), .B(new_n5798), .Y(new_n6702));
  nor_5  g04354(.A(new_n6702), .B(new_n3116), .Y(new_n6703));
  and_5  g04355(.A(new_n6703), .B(new_n2365), .Y(new_n6704));
  xnor_4 g04356(.A(new_n6689), .B(new_n2481), .Y(new_n6705));
  xnor_4 g04357(.A(n19494), .B(new_n3116), .Y(new_n6706_1));
  nor_5  g04358(.A(new_n6706_1), .B(new_n6703), .Y(new_n6707_1));
  or_5   g04359(.A(new_n6707_1), .B(new_n6704), .Y(new_n6708));
  nor_5  g04360(.A(new_n6708), .B(new_n6705), .Y(new_n6709));
  nor_5  g04361(.A(new_n6709), .B(new_n6704), .Y(new_n6710));
  xnor_4 g04362(.A(new_n6675), .B(n16223), .Y(new_n6711));
  not_8  g04363(.A(new_n6711), .Y(new_n6712));
  nor_5  g04364(.A(new_n6712), .B(new_n6710), .Y(new_n6713));
  xnor_4 g04365(.A(new_n6691_1), .B(new_n6685), .Y(new_n6714));
  not_8  g04366(.A(new_n6714), .Y(new_n6715));
  xnor_4 g04367(.A(new_n6711), .B(new_n6710), .Y(new_n6716));
  and_5  g04368(.A(new_n6716), .B(new_n6715), .Y(new_n6717));
  nor_5  g04369(.A(new_n6717), .B(new_n6713), .Y(new_n6718));
  nor_5  g04370(.A(new_n6718), .B(new_n6701), .Y(new_n6719));
  nor_5  g04371(.A(new_n6719), .B(new_n6700), .Y(new_n6720));
  xor_4  g04372(.A(new_n6720), .B(new_n6697), .Y(new_n6721));
  xnor_4 g04373(.A(new_n6721), .B(new_n3354), .Y(new_n6722));
  xor_4  g04374(.A(new_n6718), .B(new_n6701), .Y(new_n6723));
  nor_5  g04375(.A(new_n6723), .B(new_n3358), .Y(new_n6724));
  xnor_4 g04376(.A(new_n6716), .B(new_n6714), .Y(new_n6725));
  and_5  g04377(.A(new_n6725), .B(new_n3364), .Y(new_n6726));
  xnor_4 g04378(.A(new_n6725), .B(new_n3363), .Y(new_n6727));
  xnor_4 g04379(.A(new_n6702), .B(n2387), .Y(new_n6728));
  and_5  g04380(.A(new_n6728), .B(new_n3367), .Y(new_n6729_1));
  nor_5  g04381(.A(new_n6729_1), .B(new_n3370), .Y(new_n6730));
  not_8  g04382(.A(new_n6705), .Y(new_n6731));
  xnor_4 g04383(.A(new_n6708), .B(new_n6731), .Y(new_n6732));
  not_8  g04384(.A(new_n6732), .Y(new_n6733));
  and_5  g04385(.A(new_n6729_1), .B(new_n3308), .Y(new_n6734));
  nor_5  g04386(.A(new_n6734), .B(new_n6730), .Y(new_n6735));
  and_5  g04387(.A(new_n6735), .B(new_n6733), .Y(new_n6736_1));
  nor_5  g04388(.A(new_n6736_1), .B(new_n6730), .Y(new_n6737));
  and_5  g04389(.A(new_n6737), .B(new_n6727), .Y(new_n6738));
  or_5   g04390(.A(new_n6738), .B(new_n6726), .Y(new_n6739));
  xnor_4 g04391(.A(new_n6723), .B(new_n3358), .Y(new_n6740));
  nor_5  g04392(.A(new_n6740), .B(new_n6739), .Y(new_n6741));
  nor_5  g04393(.A(new_n6741), .B(new_n6724), .Y(new_n6742));
  xnor_4 g04394(.A(new_n6742), .B(new_n6722), .Y(n696));
  not_8  g04395(.A(n23697), .Y(new_n6744));
  xnor_4 g04396(.A(n25475), .B(new_n6744), .Y(new_n6745));
  not_8  g04397(.A(new_n6745), .Y(new_n6746));
  nor_5  g04398(.A(n23849), .B(n2289), .Y(new_n6747));
  not_8  g04399(.A(n2289), .Y(new_n6748));
  xnor_4 g04400(.A(n23849), .B(new_n6748), .Y(new_n6749));
  not_8  g04401(.A(new_n6749), .Y(new_n6750));
  nor_5  g04402(.A(n12446), .B(n1112), .Y(new_n6751));
  not_8  g04403(.A(n1112), .Y(new_n6752));
  xnor_4 g04404(.A(n12446), .B(new_n6752), .Y(new_n6753));
  not_8  g04405(.A(new_n6753), .Y(new_n6754));
  nor_5  g04406(.A(n20179), .B(n11011), .Y(new_n6755));
  not_8  g04407(.A(n20179), .Y(new_n6756));
  xnor_4 g04408(.A(new_n6756), .B(n11011), .Y(new_n6757));
  not_8  g04409(.A(new_n6757), .Y(new_n6758));
  nor_5  g04410(.A(n19228), .B(n16029), .Y(new_n6759));
  xnor_4 g04411(.A(n19228), .B(new_n3939), .Y(new_n6760));
  not_8  g04412(.A(new_n6760), .Y(new_n6761));
  nor_5  g04413(.A(n16476), .B(n15539), .Y(new_n6762));
  not_8  g04414(.A(n15539), .Y(new_n6763));
  xnor_4 g04415(.A(n16476), .B(new_n6763), .Y(new_n6764));
  not_8  g04416(.A(new_n6764), .Y(new_n6765));
  nor_5  g04417(.A(n11615), .B(n8052), .Y(new_n6766));
  not_8  g04418(.A(n8052), .Y(new_n6767));
  xnor_4 g04419(.A(n11615), .B(new_n6767), .Y(new_n6768));
  not_8  g04420(.A(new_n6768), .Y(new_n6769));
  nor_5  g04421(.A(n22433), .B(n10158), .Y(new_n6770));
  not_8  g04422(.A(n18962), .Y(new_n6771));
  nor_5  g04423(.A(new_n6771), .B(new_n3952_1), .Y(new_n6772));
  xnor_4 g04424(.A(n22433), .B(n10158), .Y(new_n6773_1));
  nor_5  g04425(.A(new_n6773_1), .B(new_n6772), .Y(new_n6774));
  nor_5  g04426(.A(new_n6774), .B(new_n6770), .Y(new_n6775_1));
  nor_5  g04427(.A(new_n6775_1), .B(new_n6769), .Y(new_n6776));
  nor_5  g04428(.A(new_n6776), .B(new_n6766), .Y(new_n6777));
  nor_5  g04429(.A(new_n6777), .B(new_n6765), .Y(new_n6778));
  nor_5  g04430(.A(new_n6778), .B(new_n6762), .Y(new_n6779));
  nor_5  g04431(.A(new_n6779), .B(new_n6761), .Y(new_n6780));
  nor_5  g04432(.A(new_n6780), .B(new_n6759), .Y(new_n6781));
  nor_5  g04433(.A(new_n6781), .B(new_n6758), .Y(new_n6782));
  nor_5  g04434(.A(new_n6782), .B(new_n6755), .Y(new_n6783));
  nor_5  g04435(.A(new_n6783), .B(new_n6754), .Y(new_n6784));
  nor_5  g04436(.A(new_n6784), .B(new_n6751), .Y(new_n6785_1));
  nor_5  g04437(.A(new_n6785_1), .B(new_n6750), .Y(new_n6786));
  nor_5  g04438(.A(new_n6786), .B(new_n6747), .Y(new_n6787));
  xnor_4 g04439(.A(new_n6787), .B(new_n6746), .Y(new_n6788));
  not_8  g04440(.A(new_n6788), .Y(new_n6789));
  xnor_4 g04441(.A(new_n6789), .B(new_n5503), .Y(new_n6790_1));
  xnor_4 g04442(.A(new_n6785_1), .B(new_n6750), .Y(new_n6791_1));
  and_5  g04443(.A(new_n6791_1), .B(n9655), .Y(new_n6792));
  xnor_4 g04444(.A(new_n6791_1), .B(n9655), .Y(new_n6793));
  xnor_4 g04445(.A(new_n6783), .B(new_n6754), .Y(new_n6794_1));
  and_5  g04446(.A(new_n6794_1), .B(n13490), .Y(new_n6795));
  xnor_4 g04447(.A(new_n6794_1), .B(n13490), .Y(new_n6796));
  xnor_4 g04448(.A(new_n6781), .B(new_n6758), .Y(new_n6797));
  not_8  g04449(.A(new_n6797), .Y(new_n6798));
  nor_5  g04450(.A(new_n6798), .B(new_n5511), .Y(new_n6799));
  xnor_4 g04451(.A(new_n6779), .B(new_n6761), .Y(new_n6800));
  nor_5  g04452(.A(new_n6800), .B(n1777), .Y(new_n6801));
  not_8  g04453(.A(new_n6800), .Y(new_n6802_1));
  xnor_4 g04454(.A(new_n6802_1), .B(new_n5514), .Y(new_n6803));
  xnor_4 g04455(.A(new_n6777), .B(new_n6765), .Y(new_n6804));
  nor_5  g04456(.A(new_n6804), .B(n8745), .Y(new_n6805));
  not_8  g04457(.A(new_n6804), .Y(new_n6806));
  xnor_4 g04458(.A(new_n6806), .B(new_n5517_1), .Y(new_n6807));
  xnor_4 g04459(.A(new_n6775_1), .B(new_n6769), .Y(new_n6808));
  not_8  g04460(.A(new_n6808), .Y(new_n6809));
  nor_5  g04461(.A(new_n6809), .B(new_n2441), .Y(new_n6810));
  xnor_4 g04462(.A(new_n6809), .B(n15636), .Y(new_n6811));
  xnor_4 g04463(.A(n18962), .B(n14090), .Y(new_n6812));
  nor_5  g04464(.A(new_n6812), .B(new_n2447), .Y(new_n6813));
  nor_5  g04465(.A(new_n6813), .B(n20077), .Y(new_n6814_1));
  xor_4  g04466(.A(new_n6773_1), .B(new_n6772), .Y(new_n6815));
  xnor_4 g04467(.A(new_n6813), .B(new_n2444_1), .Y(new_n6816));
  and_5  g04468(.A(new_n6816), .B(new_n6815), .Y(new_n6817));
  nor_5  g04469(.A(new_n6817), .B(new_n6814_1), .Y(new_n6818));
  and_5  g04470(.A(new_n6818), .B(new_n6811), .Y(new_n6819));
  nor_5  g04471(.A(new_n6819), .B(new_n6810), .Y(new_n6820));
  not_8  g04472(.A(new_n6820), .Y(new_n6821));
  nor_5  g04473(.A(new_n6821), .B(new_n6807), .Y(new_n6822));
  nor_5  g04474(.A(new_n6822), .B(new_n6805), .Y(new_n6823));
  nor_5  g04475(.A(new_n6823), .B(new_n6803), .Y(new_n6824));
  or_5   g04476(.A(new_n6824), .B(new_n6801), .Y(new_n6825));
  xnor_4 g04477(.A(new_n6798), .B(new_n5511), .Y(new_n6826_1));
  nor_5  g04478(.A(new_n6826_1), .B(new_n6825), .Y(new_n6827));
  nor_5  g04479(.A(new_n6827), .B(new_n6799), .Y(new_n6828));
  nor_5  g04480(.A(new_n6828), .B(new_n6796), .Y(new_n6829));
  nor_5  g04481(.A(new_n6829), .B(new_n6795), .Y(new_n6830));
  nor_5  g04482(.A(new_n6830), .B(new_n6793), .Y(new_n6831));
  nor_5  g04483(.A(new_n6831), .B(new_n6792), .Y(new_n6832));
  xnor_4 g04484(.A(new_n6832), .B(new_n6790_1), .Y(new_n6833));
  xnor_4 g04485(.A(n21915), .B(new_n6215), .Y(new_n6834));
  nor_5  g04486(.A(n27037), .B(n13775), .Y(new_n6835_1));
  not_8  g04487(.A(n13775), .Y(new_n6836));
  xnor_4 g04488(.A(n27037), .B(new_n6836), .Y(new_n6837));
  nor_5  g04489(.A(n8964), .B(n1293), .Y(new_n6838));
  not_8  g04490(.A(n1293), .Y(new_n6839));
  xnor_4 g04491(.A(n8964), .B(new_n6839), .Y(new_n6840));
  nor_5  g04492(.A(n20151), .B(n19042), .Y(new_n6841));
  not_8  g04493(.A(n19042), .Y(new_n6842));
  xnor_4 g04494(.A(n20151), .B(new_n6842), .Y(new_n6843));
  nor_5  g04495(.A(n19472), .B(n7693), .Y(new_n6844));
  xnor_4 g04496(.A(n19472), .B(new_n4015), .Y(new_n6845));
  not_8  g04497(.A(n25370), .Y(new_n6846));
  nor_5  g04498(.A(new_n6846), .B(new_n4021), .Y(new_n6847));
  or_5   g04499(.A(n25370), .B(n10405), .Y(new_n6848));
  nor_5  g04500(.A(n24786), .B(n11302), .Y(new_n6849));
  or_5   g04501(.A(new_n4113), .B(new_n4108), .Y(new_n6850));
  and_5  g04502(.A(new_n6850), .B(new_n4107), .Y(new_n6851));
  nor_5  g04503(.A(new_n6851), .B(new_n6849), .Y(new_n6852));
  and_5  g04504(.A(new_n6852), .B(new_n6848), .Y(new_n6853_1));
  nor_5  g04505(.A(new_n6853_1), .B(new_n6847), .Y(new_n6854));
  and_5  g04506(.A(new_n6854), .B(new_n6845), .Y(new_n6855));
  or_5   g04507(.A(new_n6855), .B(new_n6844), .Y(new_n6856));
  and_5  g04508(.A(new_n6856), .B(new_n6843), .Y(new_n6857));
  or_5   g04509(.A(new_n6857), .B(new_n6841), .Y(new_n6858));
  and_5  g04510(.A(new_n6858), .B(new_n6840), .Y(new_n6859));
  or_5   g04511(.A(new_n6859), .B(new_n6838), .Y(new_n6860));
  and_5  g04512(.A(new_n6860), .B(new_n6837), .Y(new_n6861_1));
  nor_5  g04513(.A(new_n6861_1), .B(new_n6835_1), .Y(new_n6862_1));
  xnor_4 g04514(.A(new_n6862_1), .B(new_n6834), .Y(new_n6863_1));
  not_8  g04515(.A(new_n6863_1), .Y(new_n6864));
  xnor_4 g04516(.A(new_n6864), .B(new_n5456), .Y(new_n6865));
  nor_5  g04517(.A(new_n6859), .B(new_n6838), .Y(new_n6866));
  xnor_4 g04518(.A(new_n6866), .B(new_n6837), .Y(new_n6867_1));
  nor_5  g04519(.A(new_n6867_1), .B(new_n5459), .Y(new_n6868));
  not_8  g04520(.A(new_n6867_1), .Y(new_n6869));
  xnor_4 g04521(.A(new_n6869), .B(new_n5459), .Y(new_n6870));
  nor_5  g04522(.A(new_n6857), .B(new_n6841), .Y(new_n6871));
  xnor_4 g04523(.A(new_n6871), .B(new_n6840), .Y(new_n6872));
  nor_5  g04524(.A(new_n6872), .B(new_n5462), .Y(new_n6873));
  not_8  g04525(.A(new_n6872), .Y(new_n6874));
  xnor_4 g04526(.A(new_n6874), .B(new_n5462), .Y(new_n6875));
  nor_5  g04527(.A(new_n6855), .B(new_n6844), .Y(new_n6876));
  xnor_4 g04528(.A(new_n6876), .B(new_n6843), .Y(new_n6877));
  nor_5  g04529(.A(new_n6877), .B(new_n5465), .Y(new_n6878));
  not_8  g04530(.A(new_n6877), .Y(new_n6879));
  xnor_4 g04531(.A(new_n6879), .B(new_n5465), .Y(new_n6880));
  xnor_4 g04532(.A(new_n6854), .B(new_n6845), .Y(new_n6881));
  not_8  g04533(.A(new_n6881), .Y(new_n6882));
  nor_5  g04534(.A(new_n6882), .B(new_n5468), .Y(new_n6883));
  xnor_4 g04535(.A(new_n6882), .B(n7566), .Y(new_n6884));
  xnor_4 g04536(.A(n25370), .B(new_n4021), .Y(new_n6885));
  xnor_4 g04537(.A(new_n6885), .B(new_n6852), .Y(new_n6886));
  nor_5  g04538(.A(new_n6886), .B(new_n5471), .Y(new_n6887));
  not_8  g04539(.A(new_n6886), .Y(new_n6888));
  xnor_4 g04540(.A(new_n6888), .B(new_n5471), .Y(new_n6889));
  nor_5  g04541(.A(new_n4115), .B(new_n5475), .Y(new_n6890));
  nor_5  g04542(.A(new_n4138), .B(n20986), .Y(new_n6891));
  or_5   g04543(.A(new_n4135), .B(new_n5798), .Y(new_n6892));
  xnor_4 g04544(.A(new_n4138), .B(new_n5478), .Y(new_n6893));
  and_5  g04545(.A(new_n6893), .B(new_n6892), .Y(new_n6894));
  nor_5  g04546(.A(new_n6894), .B(new_n6891), .Y(new_n6895));
  xnor_4 g04547(.A(new_n4116), .B(new_n5475), .Y(new_n6896));
  and_5  g04548(.A(new_n6896), .B(new_n6895), .Y(new_n6897));
  or_5   g04549(.A(new_n6897), .B(new_n6890), .Y(new_n6898));
  and_5  g04550(.A(new_n6898), .B(new_n6889), .Y(new_n6899));
  or_5   g04551(.A(new_n6899), .B(new_n6887), .Y(new_n6900));
  and_5  g04552(.A(new_n6900), .B(new_n6884), .Y(new_n6901));
  or_5   g04553(.A(new_n6901), .B(new_n6883), .Y(new_n6902));
  and_5  g04554(.A(new_n6902), .B(new_n6880), .Y(new_n6903));
  or_5   g04555(.A(new_n6903), .B(new_n6878), .Y(new_n6904));
  and_5  g04556(.A(new_n6904), .B(new_n6875), .Y(new_n6905));
  or_5   g04557(.A(new_n6905), .B(new_n6873), .Y(new_n6906));
  and_5  g04558(.A(new_n6906), .B(new_n6870), .Y(new_n6907));
  or_5   g04559(.A(new_n6907), .B(new_n6868), .Y(new_n6908));
  xor_4  g04560(.A(new_n6908), .B(new_n6865), .Y(new_n6909));
  xnor_4 g04561(.A(new_n6909), .B(new_n6833), .Y(new_n6910));
  xor_4  g04562(.A(new_n6906), .B(new_n6870), .Y(new_n6911));
  not_8  g04563(.A(new_n6911), .Y(new_n6912));
  xor_4  g04564(.A(new_n6830), .B(new_n6793), .Y(new_n6913));
  and_5  g04565(.A(new_n6913), .B(new_n6912), .Y(new_n6914));
  xnor_4 g04566(.A(new_n6913), .B(new_n6912), .Y(new_n6915));
  xor_4  g04567(.A(new_n6904), .B(new_n6875), .Y(new_n6916));
  not_8  g04568(.A(new_n6916), .Y(new_n6917));
  xor_4  g04569(.A(new_n6828), .B(new_n6796), .Y(new_n6918));
  and_5  g04570(.A(new_n6918), .B(new_n6917), .Y(new_n6919));
  xnor_4 g04571(.A(new_n6918), .B(new_n6917), .Y(new_n6920));
  xor_4  g04572(.A(new_n6902), .B(new_n6880), .Y(new_n6921));
  not_8  g04573(.A(new_n6921), .Y(new_n6922));
  xor_4  g04574(.A(new_n6826_1), .B(new_n6825), .Y(new_n6923));
  and_5  g04575(.A(new_n6923), .B(new_n6922), .Y(new_n6924));
  xnor_4 g04576(.A(new_n6923), .B(new_n6922), .Y(new_n6925));
  xnor_4 g04577(.A(new_n6823), .B(new_n6803), .Y(new_n6926));
  not_8  g04578(.A(new_n6926), .Y(new_n6927));
  xor_4  g04579(.A(new_n6900), .B(new_n6884), .Y(new_n6928));
  nor_5  g04580(.A(new_n6928), .B(new_n6927), .Y(new_n6929));
  xnor_4 g04581(.A(new_n6928), .B(new_n6927), .Y(new_n6930));
  xnor_4 g04582(.A(new_n6820), .B(new_n6807), .Y(new_n6931));
  xor_4  g04583(.A(new_n6898), .B(new_n6889), .Y(new_n6932));
  nor_5  g04584(.A(new_n6932), .B(new_n6931), .Y(new_n6933));
  xnor_4 g04585(.A(new_n6932), .B(new_n6931), .Y(new_n6934));
  xnor_4 g04586(.A(new_n6896), .B(new_n6895), .Y(new_n6935));
  xnor_4 g04587(.A(new_n6818), .B(new_n6811), .Y(new_n6936));
  not_8  g04588(.A(new_n6936), .Y(new_n6937));
  and_5  g04589(.A(new_n6937), .B(new_n6935), .Y(new_n6938));
  xnor_4 g04590(.A(new_n6937), .B(new_n6935), .Y(new_n6939));
  nor_5  g04591(.A(new_n4135), .B(new_n5798), .Y(new_n6940));
  xnor_4 g04592(.A(new_n6893), .B(new_n6940), .Y(new_n6941));
  xnor_4 g04593(.A(new_n6773_1), .B(new_n6772), .Y(new_n6942));
  xnor_4 g04594(.A(new_n6816), .B(new_n6942), .Y(new_n6943));
  not_8  g04595(.A(new_n6943), .Y(new_n6944));
  and_5  g04596(.A(new_n6944), .B(new_n6941), .Y(new_n6945));
  xnor_4 g04597(.A(new_n6812), .B(n6794), .Y(new_n6946));
  not_8  g04598(.A(new_n6946), .Y(new_n6947));
  xnor_4 g04599(.A(new_n4135), .B(n12384), .Y(new_n6948));
  nor_5  g04600(.A(new_n6948), .B(new_n6947), .Y(new_n6949));
  xnor_4 g04601(.A(new_n6943), .B(new_n6941), .Y(new_n6950));
  and_5  g04602(.A(new_n6950), .B(new_n6949), .Y(new_n6951));
  nor_5  g04603(.A(new_n6951), .B(new_n6945), .Y(new_n6952));
  nor_5  g04604(.A(new_n6952), .B(new_n6939), .Y(new_n6953));
  nor_5  g04605(.A(new_n6953), .B(new_n6938), .Y(new_n6954));
  nor_5  g04606(.A(new_n6954), .B(new_n6934), .Y(new_n6955));
  nor_5  g04607(.A(new_n6955), .B(new_n6933), .Y(new_n6956));
  nor_5  g04608(.A(new_n6956), .B(new_n6930), .Y(new_n6957));
  nor_5  g04609(.A(new_n6957), .B(new_n6929), .Y(new_n6958));
  nor_5  g04610(.A(new_n6958), .B(new_n6925), .Y(new_n6959));
  nor_5  g04611(.A(new_n6959), .B(new_n6924), .Y(new_n6960));
  nor_5  g04612(.A(new_n6960), .B(new_n6920), .Y(new_n6961));
  nor_5  g04613(.A(new_n6961), .B(new_n6919), .Y(new_n6962));
  nor_5  g04614(.A(new_n6962), .B(new_n6915), .Y(new_n6963));
  nor_5  g04615(.A(new_n6963), .B(new_n6914), .Y(new_n6964));
  xnor_4 g04616(.A(new_n6964), .B(new_n6910), .Y(n723));
  xnor_4 g04617(.A(n26986), .B(n2272), .Y(new_n6966));
  not_8  g04618(.A(n25331), .Y(new_n6967_1));
  nor_5  g04619(.A(new_n6967_1), .B(n21287), .Y(new_n6968));
  xnor_4 g04620(.A(n25331), .B(n21287), .Y(new_n6969));
  not_8  g04621(.A(n18483), .Y(new_n6970));
  nor_5  g04622(.A(new_n6970), .B(n4256), .Y(new_n6971_1));
  xnor_4 g04623(.A(n18483), .B(n4256), .Y(new_n6972));
  not_8  g04624(.A(n21934), .Y(new_n6973));
  nor_5  g04625(.A(n22332), .B(new_n6973), .Y(new_n6974));
  xnor_4 g04626(.A(n22332), .B(n21934), .Y(new_n6975_1));
  not_8  g04627(.A(n18901), .Y(new_n6976));
  nor_5  g04628(.A(n18907), .B(new_n6976), .Y(new_n6977));
  xnor_4 g04629(.A(n18907), .B(n18901), .Y(new_n6978));
  not_8  g04630(.A(n4376), .Y(new_n6979));
  nor_5  g04631(.A(new_n6979), .B(n2731), .Y(new_n6980));
  xnor_4 g04632(.A(n4376), .B(n2731), .Y(new_n6981));
  not_8  g04633(.A(n14570), .Y(new_n6982));
  nor_5  g04634(.A(n19911), .B(new_n6982), .Y(new_n6983_1));
  xnor_4 g04635(.A(n19911), .B(n14570), .Y(new_n6984));
  nor_5  g04636(.A(n23775), .B(new_n2389), .Y(new_n6985_1));
  not_8  g04637(.A(n23775), .Y(new_n6986));
  nor_5  g04638(.A(new_n6986), .B(n13708), .Y(new_n6987));
  nor_5  g04639(.A(new_n3826), .B(n8259), .Y(new_n6988));
  not_8  g04640(.A(n8259), .Y(new_n6989));
  nor_5  g04641(.A(n18409), .B(new_n6989), .Y(new_n6990));
  nor_5  g04642(.A(n11479), .B(new_n2381), .Y(new_n6991));
  not_8  g04643(.A(new_n6991), .Y(new_n6992));
  nor_5  g04644(.A(new_n6992), .B(new_n6990), .Y(new_n6993));
  nor_5  g04645(.A(new_n6993), .B(new_n6988), .Y(new_n6994));
  nor_5  g04646(.A(new_n6994), .B(new_n6987), .Y(new_n6995));
  nor_5  g04647(.A(new_n6995), .B(new_n6985_1), .Y(new_n6996));
  and_5  g04648(.A(new_n6996), .B(new_n6984), .Y(new_n6997));
  or_5   g04649(.A(new_n6997), .B(new_n6983_1), .Y(new_n6998_1));
  and_5  g04650(.A(new_n6998_1), .B(new_n6981), .Y(new_n6999));
  or_5   g04651(.A(new_n6999), .B(new_n6980), .Y(new_n7000));
  and_5  g04652(.A(new_n7000), .B(new_n6978), .Y(new_n7001));
  or_5   g04653(.A(new_n7001), .B(new_n6977), .Y(new_n7002));
  and_5  g04654(.A(new_n7002), .B(new_n6975_1), .Y(new_n7003));
  or_5   g04655(.A(new_n7003), .B(new_n6974), .Y(new_n7004));
  and_5  g04656(.A(new_n7004), .B(new_n6972), .Y(new_n7005));
  or_5   g04657(.A(new_n7005), .B(new_n6971_1), .Y(new_n7006));
  and_5  g04658(.A(new_n7006), .B(new_n6969), .Y(new_n7007));
  or_5   g04659(.A(new_n7007), .B(new_n6968), .Y(new_n7008));
  xor_4  g04660(.A(new_n7008), .B(new_n6966), .Y(new_n7009));
  xnor_4 g04661(.A(n1255), .B(n468), .Y(new_n7010));
  nor_5  g04662(.A(n9512), .B(n5400), .Y(new_n7011));
  xnor_4 g04663(.A(n9512), .B(n5400), .Y(new_n7012));
  nor_5  g04664(.A(n23923), .B(n16608), .Y(new_n7013));
  xnor_4 g04665(.A(n23923), .B(n16608), .Y(new_n7014));
  nor_5  g04666(.A(n21735), .B(n329), .Y(new_n7015));
  xnor_4 g04667(.A(n21735), .B(n329), .Y(new_n7016));
  nor_5  g04668(.A(n24170), .B(n24085), .Y(new_n7017));
  xnor_4 g04669(.A(n24170), .B(n24085), .Y(new_n7018));
  nor_5  g04670(.A(n14071), .B(n2409), .Y(new_n7019));
  xnor_4 g04671(.A(n14071), .B(n2409), .Y(new_n7020));
  nor_5  g04672(.A(n8869), .B(n1738), .Y(new_n7021));
  xnor_4 g04673(.A(n8869), .B(n1738), .Y(new_n7022));
  nor_5  g04674(.A(n12152), .B(n10372), .Y(new_n7023));
  not_8  g04675(.A(n7428), .Y(new_n7024));
  not_8  g04676(.A(n19107), .Y(new_n7025));
  nor_5  g04677(.A(new_n7025), .B(new_n7024), .Y(new_n7026_1));
  xnor_4 g04678(.A(n12152), .B(n10372), .Y(new_n7027));
  nor_5  g04679(.A(new_n7027), .B(new_n7026_1), .Y(new_n7028));
  nor_5  g04680(.A(new_n7028), .B(new_n7023), .Y(new_n7029));
  nor_5  g04681(.A(new_n7029), .B(new_n7022), .Y(new_n7030));
  nor_5  g04682(.A(new_n7030), .B(new_n7021), .Y(new_n7031));
  nor_5  g04683(.A(new_n7031), .B(new_n7020), .Y(new_n7032_1));
  nor_5  g04684(.A(new_n7032_1), .B(new_n7019), .Y(new_n7033));
  nor_5  g04685(.A(new_n7033), .B(new_n7018), .Y(new_n7034));
  nor_5  g04686(.A(new_n7034), .B(new_n7017), .Y(new_n7035));
  nor_5  g04687(.A(new_n7035), .B(new_n7016), .Y(new_n7036));
  nor_5  g04688(.A(new_n7036), .B(new_n7015), .Y(new_n7037));
  nor_5  g04689(.A(new_n7037), .B(new_n7014), .Y(new_n7038_1));
  nor_5  g04690(.A(new_n7038_1), .B(new_n7013), .Y(new_n7039));
  nor_5  g04691(.A(new_n7039), .B(new_n7012), .Y(new_n7040));
  nor_5  g04692(.A(new_n7040), .B(new_n7011), .Y(new_n7041));
  xnor_4 g04693(.A(new_n7041), .B(new_n7010), .Y(new_n7042));
  not_8  g04694(.A(n12861), .Y(new_n7043));
  xnor_4 g04695(.A(n14130), .B(new_n7043), .Y(new_n7044));
  nor_5  g04696(.A(n16482), .B(n13333), .Y(new_n7045));
  not_8  g04697(.A(n13333), .Y(new_n7046));
  xnor_4 g04698(.A(n16482), .B(new_n7046), .Y(new_n7047));
  nor_5  g04699(.A(n9942), .B(n2210), .Y(new_n7048));
  not_8  g04700(.A(n2210), .Y(new_n7049));
  xnor_4 g04701(.A(n9942), .B(new_n7049), .Y(new_n7050));
  nor_5  g04702(.A(n25643), .B(n20604), .Y(new_n7051));
  or_5   g04703(.A(new_n5129), .B(new_n5127), .Y(new_n7052));
  and_5  g04704(.A(new_n7052), .B(new_n5126), .Y(new_n7053));
  or_5   g04705(.A(new_n7053), .B(new_n7051), .Y(new_n7054));
  and_5  g04706(.A(new_n7054), .B(new_n7050), .Y(new_n7055));
  or_5   g04707(.A(new_n7055), .B(new_n7048), .Y(new_n7056));
  and_5  g04708(.A(new_n7056), .B(new_n7047), .Y(new_n7057_1));
  nor_5  g04709(.A(new_n7057_1), .B(new_n7045), .Y(new_n7058));
  xnor_4 g04710(.A(new_n7058), .B(new_n7044), .Y(new_n7059));
  nor_5  g04711(.A(new_n7059), .B(new_n7042), .Y(new_n7060));
  xnor_4 g04712(.A(new_n7059), .B(new_n7042), .Y(new_n7061));
  xnor_4 g04713(.A(new_n7039), .B(new_n7012), .Y(new_n7062));
  nor_5  g04714(.A(new_n7055), .B(new_n7048), .Y(new_n7063));
  xnor_4 g04715(.A(new_n7063), .B(new_n7047), .Y(new_n7064));
  nor_5  g04716(.A(new_n7064), .B(new_n7062), .Y(new_n7065));
  xnor_4 g04717(.A(new_n7064), .B(new_n7062), .Y(new_n7066));
  nor_5  g04718(.A(new_n7053), .B(new_n7051), .Y(new_n7067));
  xnor_4 g04719(.A(new_n7067), .B(new_n7050), .Y(new_n7068));
  xnor_4 g04720(.A(new_n7037), .B(new_n7014), .Y(new_n7069));
  nor_5  g04721(.A(new_n7069), .B(new_n7068), .Y(new_n7070));
  xnor_4 g04722(.A(new_n7069), .B(new_n7068), .Y(new_n7071));
  xnor_4 g04723(.A(new_n7035), .B(new_n7016), .Y(new_n7072));
  nor_5  g04724(.A(new_n7072), .B(new_n5131_1), .Y(new_n7073));
  xnor_4 g04725(.A(new_n7072), .B(new_n5131_1), .Y(new_n7074));
  xnor_4 g04726(.A(new_n7033), .B(new_n7018), .Y(new_n7075));
  nor_5  g04727(.A(new_n7075), .B(new_n5122), .Y(new_n7076));
  xnor_4 g04728(.A(new_n7075), .B(new_n5122), .Y(new_n7077));
  xnor_4 g04729(.A(new_n7031), .B(new_n7020), .Y(new_n7078));
  nor_5  g04730(.A(new_n7078), .B(new_n5112), .Y(new_n7079_1));
  xnor_4 g04731(.A(new_n7078), .B(new_n5113), .Y(new_n7080));
  xnor_4 g04732(.A(new_n7029), .B(new_n7022), .Y(new_n7081));
  nor_5  g04733(.A(new_n7081), .B(new_n5102), .Y(new_n7082));
  xnor_4 g04734(.A(new_n7081), .B(new_n5102), .Y(new_n7083));
  xnor_4 g04735(.A(new_n7027), .B(new_n7026_1), .Y(new_n7084));
  nor_5  g04736(.A(new_n7084), .B(new_n5093), .Y(new_n7085));
  xnor_4 g04737(.A(n19107), .B(new_n7024), .Y(new_n7086));
  nor_5  g04738(.A(new_n7086), .B(new_n5143), .Y(new_n7087));
  xnor_4 g04739(.A(new_n7084), .B(new_n5094), .Y(new_n7088));
  and_5  g04740(.A(new_n7088), .B(new_n7087), .Y(new_n7089));
  nor_5  g04741(.A(new_n7089), .B(new_n7085), .Y(new_n7090));
  nor_5  g04742(.A(new_n7090), .B(new_n7083), .Y(new_n7091));
  or_5   g04743(.A(new_n7091), .B(new_n7082), .Y(new_n7092));
  and_5  g04744(.A(new_n7092), .B(new_n7080), .Y(new_n7093));
  nor_5  g04745(.A(new_n7093), .B(new_n7079_1), .Y(new_n7094));
  nor_5  g04746(.A(new_n7094), .B(new_n7077), .Y(new_n7095));
  nor_5  g04747(.A(new_n7095), .B(new_n7076), .Y(new_n7096));
  nor_5  g04748(.A(new_n7096), .B(new_n7074), .Y(new_n7097));
  nor_5  g04749(.A(new_n7097), .B(new_n7073), .Y(new_n7098));
  nor_5  g04750(.A(new_n7098), .B(new_n7071), .Y(new_n7099_1));
  nor_5  g04751(.A(new_n7099_1), .B(new_n7070), .Y(new_n7100));
  nor_5  g04752(.A(new_n7100), .B(new_n7066), .Y(new_n7101));
  nor_5  g04753(.A(new_n7101), .B(new_n7065), .Y(new_n7102));
  nor_5  g04754(.A(new_n7102), .B(new_n7061), .Y(new_n7103));
  nor_5  g04755(.A(new_n7103), .B(new_n7060), .Y(new_n7104));
  xnor_4 g04756(.A(n22442), .B(n22253), .Y(new_n7105));
  nor_5  g04757(.A(n1255), .B(n468), .Y(new_n7106));
  nor_5  g04758(.A(new_n7041), .B(new_n7010), .Y(new_n7107));
  nor_5  g04759(.A(new_n7107), .B(new_n7106), .Y(new_n7108));
  xnor_4 g04760(.A(new_n7108), .B(new_n7105), .Y(new_n7109));
  not_8  g04761(.A(n8305), .Y(new_n7110));
  xnor_4 g04762(.A(n8856), .B(new_n7110), .Y(new_n7111));
  nor_5  g04763(.A(n14130), .B(n12861), .Y(new_n7112));
  or_5   g04764(.A(new_n7057_1), .B(new_n7045), .Y(new_n7113));
  and_5  g04765(.A(new_n7113), .B(new_n7044), .Y(new_n7114));
  nor_5  g04766(.A(new_n7114), .B(new_n7112), .Y(new_n7115));
  xnor_4 g04767(.A(new_n7115), .B(new_n7111), .Y(new_n7116));
  xnor_4 g04768(.A(new_n7116), .B(new_n7109), .Y(new_n7117));
  xnor_4 g04769(.A(new_n7117), .B(new_n7104), .Y(new_n7118));
  nor_5  g04770(.A(new_n7118), .B(new_n7009), .Y(new_n7119));
  xnor_4 g04771(.A(new_n7118), .B(new_n7009), .Y(new_n7120));
  xor_4  g04772(.A(new_n7006), .B(new_n6969), .Y(new_n7121));
  xnor_4 g04773(.A(new_n7102), .B(new_n7061), .Y(new_n7122));
  nor_5  g04774(.A(new_n7122), .B(new_n7121), .Y(new_n7123));
  xnor_4 g04775(.A(new_n7122), .B(new_n7121), .Y(new_n7124));
  xor_4  g04776(.A(new_n7004), .B(new_n6972), .Y(new_n7125));
  xnor_4 g04777(.A(new_n7100), .B(new_n7066), .Y(new_n7126));
  nor_5  g04778(.A(new_n7126), .B(new_n7125), .Y(new_n7127));
  xnor_4 g04779(.A(new_n7126), .B(new_n7125), .Y(new_n7128));
  xor_4  g04780(.A(new_n7002), .B(new_n6975_1), .Y(new_n7129));
  xnor_4 g04781(.A(new_n7098), .B(new_n7071), .Y(new_n7130));
  nor_5  g04782(.A(new_n7130), .B(new_n7129), .Y(new_n7131));
  xnor_4 g04783(.A(new_n7130), .B(new_n7129), .Y(new_n7132));
  xor_4  g04784(.A(new_n7000), .B(new_n6978), .Y(new_n7133));
  xnor_4 g04785(.A(new_n7096), .B(new_n7074), .Y(new_n7134));
  nor_5  g04786(.A(new_n7134), .B(new_n7133), .Y(new_n7135));
  xnor_4 g04787(.A(new_n7134), .B(new_n7133), .Y(new_n7136));
  xor_4  g04788(.A(new_n6998_1), .B(new_n6981), .Y(new_n7137));
  xnor_4 g04789(.A(new_n7094), .B(new_n7077), .Y(new_n7138));
  nor_5  g04790(.A(new_n7138), .B(new_n7137), .Y(new_n7139_1));
  xnor_4 g04791(.A(new_n7138), .B(new_n7137), .Y(new_n7140));
  xor_4  g04792(.A(new_n7092), .B(new_n7080), .Y(new_n7141));
  xnor_4 g04793(.A(new_n6996), .B(new_n6984), .Y(new_n7142));
  and_5  g04794(.A(new_n7142), .B(new_n7141), .Y(new_n7143));
  xnor_4 g04795(.A(new_n7090), .B(new_n7083), .Y(new_n7144));
  not_8  g04796(.A(new_n7144), .Y(new_n7145));
  xnor_4 g04797(.A(n23775), .B(n13708), .Y(new_n7146));
  xnor_4 g04798(.A(new_n7146), .B(new_n6994), .Y(new_n7147));
  and_5  g04799(.A(new_n7147), .B(new_n7145), .Y(new_n7148));
  xnor_4 g04800(.A(new_n7147), .B(new_n7144), .Y(new_n7149_1));
  xnor_4 g04801(.A(new_n7086), .B(new_n5090), .Y(new_n7150));
  xnor_4 g04802(.A(n11479), .B(n5704), .Y(new_n7151));
  nor_5  g04803(.A(new_n7151), .B(new_n7150), .Y(new_n7152));
  xnor_4 g04804(.A(n18409), .B(n8259), .Y(new_n7153));
  xnor_4 g04805(.A(new_n7153), .B(new_n6992), .Y(new_n7154));
  not_8  g04806(.A(new_n7154), .Y(new_n7155));
  and_5  g04807(.A(new_n7155), .B(new_n7152), .Y(new_n7156));
  xnor_4 g04808(.A(new_n7088), .B(new_n7087), .Y(new_n7157));
  not_8  g04809(.A(new_n7157), .Y(new_n7158));
  xnor_4 g04810(.A(new_n7155), .B(new_n7152), .Y(new_n7159));
  nor_5  g04811(.A(new_n7159), .B(new_n7158), .Y(new_n7160));
  nor_5  g04812(.A(new_n7160), .B(new_n7156), .Y(new_n7161));
  and_5  g04813(.A(new_n7161), .B(new_n7149_1), .Y(new_n7162));
  nor_5  g04814(.A(new_n7162), .B(new_n7148), .Y(new_n7163));
  xnor_4 g04815(.A(new_n7142), .B(new_n7141), .Y(new_n7164));
  nor_5  g04816(.A(new_n7164), .B(new_n7163), .Y(new_n7165));
  nor_5  g04817(.A(new_n7165), .B(new_n7143), .Y(new_n7166));
  nor_5  g04818(.A(new_n7166), .B(new_n7140), .Y(new_n7167));
  nor_5  g04819(.A(new_n7167), .B(new_n7139_1), .Y(new_n7168));
  nor_5  g04820(.A(new_n7168), .B(new_n7136), .Y(new_n7169));
  nor_5  g04821(.A(new_n7169), .B(new_n7135), .Y(new_n7170));
  nor_5  g04822(.A(new_n7170), .B(new_n7132), .Y(new_n7171));
  nor_5  g04823(.A(new_n7171), .B(new_n7131), .Y(new_n7172));
  nor_5  g04824(.A(new_n7172), .B(new_n7128), .Y(new_n7173));
  nor_5  g04825(.A(new_n7173), .B(new_n7127), .Y(new_n7174));
  nor_5  g04826(.A(new_n7174), .B(new_n7124), .Y(new_n7175));
  nor_5  g04827(.A(new_n7175), .B(new_n7123), .Y(new_n7176));
  nor_5  g04828(.A(new_n7176), .B(new_n7120), .Y(new_n7177));
  nor_5  g04829(.A(new_n7177), .B(new_n7119), .Y(new_n7178));
  not_8  g04830(.A(n2272), .Y(new_n7179));
  nor_5  g04831(.A(n26986), .B(new_n7179), .Y(new_n7180));
  and_5  g04832(.A(new_n7008), .B(new_n6966), .Y(new_n7181));
  nor_5  g04833(.A(new_n7181), .B(new_n7180), .Y(new_n7182));
  nor_5  g04834(.A(n22442), .B(n22253), .Y(new_n7183));
  nor_5  g04835(.A(new_n7108), .B(new_n7105), .Y(new_n7184));
  nor_5  g04836(.A(new_n7184), .B(new_n7183), .Y(new_n7185));
  nor_5  g04837(.A(n8856), .B(n8305), .Y(new_n7186));
  or_5   g04838(.A(new_n7114), .B(new_n7112), .Y(new_n7187));
  and_5  g04839(.A(new_n7187), .B(new_n7111), .Y(new_n7188));
  nor_5  g04840(.A(new_n7188), .B(new_n7186), .Y(new_n7189));
  xnor_4 g04841(.A(new_n7189), .B(new_n7185), .Y(new_n7190_1));
  nor_5  g04842(.A(new_n7116), .B(new_n7109), .Y(new_n7191));
  nor_5  g04843(.A(new_n7117), .B(new_n7104), .Y(new_n7192));
  nor_5  g04844(.A(new_n7192), .B(new_n7191), .Y(new_n7193));
  xnor_4 g04845(.A(new_n7193), .B(new_n7190_1), .Y(new_n7194));
  not_8  g04846(.A(new_n7194), .Y(new_n7195));
  xnor_4 g04847(.A(new_n7195), .B(new_n7182), .Y(new_n7196));
  xnor_4 g04848(.A(new_n7196), .B(new_n7178), .Y(n735));
  xnor_4 g04849(.A(n21138), .B(n14230), .Y(new_n7198));
  xnor_4 g04850(.A(new_n6812), .B(n19234), .Y(new_n7199));
  not_8  g04851(.A(new_n7199), .Y(new_n7200));
  xnor_4 g04852(.A(new_n7200), .B(n26167), .Y(new_n7201));
  xnor_4 g04853(.A(new_n7201), .B(new_n7198), .Y(n779));
  nor_5  g04854(.A(n17458), .B(new_n5981), .Y(new_n7203));
  xnor_4 g04855(.A(n17458), .B(n8526), .Y(new_n7204));
  nor_5  g04856(.A(new_n6025), .B(n1222), .Y(new_n7205));
  xnor_4 g04857(.A(n2816), .B(n1222), .Y(new_n7206));
  nor_5  g04858(.A(n25240), .B(new_n6031_1), .Y(new_n7207));
  xnor_4 g04859(.A(n25240), .B(n20359), .Y(new_n7208));
  nor_5  g04860(.A(n10125), .B(new_n6037), .Y(new_n7209));
  xnor_4 g04861(.A(n10125), .B(n4409), .Y(new_n7210));
  nor_5  g04862(.A(n8067), .B(new_n6043), .Y(new_n7211));
  xnor_4 g04863(.A(n8067), .B(n3570), .Y(new_n7212));
  nor_5  g04864(.A(n20923), .B(new_n6049), .Y(new_n7213));
  xnor_4 g04865(.A(n20923), .B(n13668), .Y(new_n7214));
  nor_5  g04866(.A(new_n6055), .B(n18157), .Y(new_n7215));
  xnor_4 g04867(.A(n21276), .B(n18157), .Y(new_n7216));
  not_8  g04868(.A(n12161), .Y(new_n7217));
  nor_5  g04869(.A(n26748), .B(new_n7217), .Y(new_n7218));
  nor_5  g04870(.A(new_n6061), .B(n12161), .Y(new_n7219));
  not_8  g04871(.A(n5026), .Y(new_n7220));
  nor_5  g04872(.A(n10057), .B(new_n7220), .Y(new_n7221));
  nor_5  g04873(.A(new_n6068), .B(n5026), .Y(new_n7222));
  or_5   g04874(.A(n8920), .B(new_n6628_1), .Y(new_n7223));
  nor_5  g04875(.A(new_n7223), .B(new_n7222), .Y(new_n7224));
  nor_5  g04876(.A(new_n7224), .B(new_n7221), .Y(new_n7225));
  nor_5  g04877(.A(new_n7225), .B(new_n7219), .Y(new_n7226));
  nor_5  g04878(.A(new_n7226), .B(new_n7218), .Y(new_n7227));
  and_5  g04879(.A(new_n7227), .B(new_n7216), .Y(new_n7228));
  or_5   g04880(.A(new_n7228), .B(new_n7215), .Y(new_n7229_1));
  and_5  g04881(.A(new_n7229_1), .B(new_n7214), .Y(new_n7230_1));
  or_5   g04882(.A(new_n7230_1), .B(new_n7213), .Y(new_n7231));
  and_5  g04883(.A(new_n7231), .B(new_n7212), .Y(new_n7232));
  or_5   g04884(.A(new_n7232), .B(new_n7211), .Y(new_n7233_1));
  and_5  g04885(.A(new_n7233_1), .B(new_n7210), .Y(new_n7234));
  or_5   g04886(.A(new_n7234), .B(new_n7209), .Y(new_n7235));
  and_5  g04887(.A(new_n7235), .B(new_n7208), .Y(new_n7236_1));
  or_5   g04888(.A(new_n7236_1), .B(new_n7207), .Y(new_n7237));
  and_5  g04889(.A(new_n7237), .B(new_n7206), .Y(new_n7238));
  or_5   g04890(.A(new_n7238), .B(new_n7205), .Y(new_n7239));
  and_5  g04891(.A(new_n7239), .B(new_n7204), .Y(new_n7240));
  nor_5  g04892(.A(new_n7240), .B(new_n7203), .Y(new_n7241));
  not_8  g04893(.A(new_n7241), .Y(new_n7242));
  not_8  g04894(.A(n26986), .Y(new_n7243));
  nor_5  g04895(.A(new_n7243), .B(n19282), .Y(new_n7244));
  xnor_4 g04896(.A(n26986), .B(n19282), .Y(new_n7245));
  and_5  g04897(.A(n21287), .B(new_n2926), .Y(new_n7246));
  xnor_4 g04898(.A(n21287), .B(n12657), .Y(new_n7247));
  not_8  g04899(.A(n4256), .Y(new_n7248));
  nor_5  g04900(.A(n17077), .B(new_n7248), .Y(new_n7249));
  xnor_4 g04901(.A(n17077), .B(n4256), .Y(new_n7250));
  not_8  g04902(.A(n26510), .Y(new_n7251));
  and_5  g04903(.A(new_n7251), .B(n22332), .Y(new_n7252));
  and_5  g04904(.A(new_n3839), .B(new_n3814), .Y(new_n7253_1));
  or_5   g04905(.A(new_n7253_1), .B(new_n7252), .Y(new_n7254));
  and_5  g04906(.A(new_n7254), .B(new_n7250), .Y(new_n7255));
  or_5   g04907(.A(new_n7255), .B(new_n7249), .Y(new_n7256_1));
  and_5  g04908(.A(new_n7256_1), .B(new_n7247), .Y(new_n7257));
  or_5   g04909(.A(new_n7257), .B(new_n7246), .Y(new_n7258));
  and_5  g04910(.A(new_n7258), .B(new_n7245), .Y(new_n7259));
  nor_5  g04911(.A(new_n7259), .B(new_n7244), .Y(new_n7260));
  xnor_4 g04912(.A(new_n7260), .B(new_n7242), .Y(new_n7261));
  nor_5  g04913(.A(new_n7238), .B(new_n7205), .Y(new_n7262));
  xnor_4 g04914(.A(new_n7262), .B(new_n7204), .Y(new_n7263));
  xor_4  g04915(.A(new_n7258), .B(new_n7245), .Y(new_n7264));
  and_5  g04916(.A(new_n7264), .B(new_n7263), .Y(new_n7265));
  not_8  g04917(.A(new_n7263), .Y(new_n7266));
  xnor_4 g04918(.A(new_n7264), .B(new_n7266), .Y(new_n7267));
  nor_5  g04919(.A(new_n7236_1), .B(new_n7207), .Y(new_n7268_1));
  xnor_4 g04920(.A(new_n7268_1), .B(new_n7206), .Y(new_n7269));
  xor_4  g04921(.A(new_n7256_1), .B(new_n7247), .Y(new_n7270));
  nor_5  g04922(.A(new_n7270), .B(new_n7269), .Y(new_n7271));
  xnor_4 g04923(.A(new_n7270), .B(new_n7269), .Y(new_n7272));
  nor_5  g04924(.A(new_n7234), .B(new_n7209), .Y(new_n7273));
  xnor_4 g04925(.A(new_n7273), .B(new_n7208), .Y(new_n7274));
  xor_4  g04926(.A(new_n7254), .B(new_n7250), .Y(new_n7275));
  nor_5  g04927(.A(new_n7275), .B(new_n7274), .Y(new_n7276));
  xnor_4 g04928(.A(new_n7275), .B(new_n7274), .Y(new_n7277_1));
  xor_4  g04929(.A(new_n7233_1), .B(new_n7210), .Y(new_n7278));
  nor_5  g04930(.A(new_n7278), .B(new_n3840), .Y(new_n7279));
  xnor_4 g04931(.A(new_n7278), .B(new_n3840), .Y(new_n7280_1));
  nor_5  g04932(.A(new_n7230_1), .B(new_n7213), .Y(new_n7281));
  xnor_4 g04933(.A(new_n7281), .B(new_n7212), .Y(new_n7282));
  nor_5  g04934(.A(new_n7282), .B(new_n3852), .Y(new_n7283));
  xnor_4 g04935(.A(new_n7282), .B(new_n3852), .Y(new_n7284));
  xor_4  g04936(.A(new_n7229_1), .B(new_n7214), .Y(new_n7285));
  nor_5  g04937(.A(new_n7285), .B(new_n3856), .Y(new_n7286));
  xnor_4 g04938(.A(new_n7285), .B(new_n3856), .Y(new_n7287));
  xor_4  g04939(.A(new_n7227), .B(new_n7216), .Y(new_n7288));
  nor_5  g04940(.A(new_n7288), .B(new_n3862), .Y(new_n7289));
  not_8  g04941(.A(new_n7288), .Y(new_n7290));
  xnor_4 g04942(.A(new_n7290), .B(new_n3862), .Y(new_n7291));
  xnor_4 g04943(.A(n26748), .B(n12161), .Y(new_n7292));
  xor_4  g04944(.A(new_n7292), .B(new_n7225), .Y(new_n7293));
  nor_5  g04945(.A(new_n7293), .B(new_n3868), .Y(new_n7294));
  not_8  g04946(.A(new_n7293), .Y(new_n7295));
  xnor_4 g04947(.A(new_n7295), .B(new_n3868), .Y(new_n7296));
  xnor_4 g04948(.A(n10057), .B(n5026), .Y(new_n7297));
  xnor_4 g04949(.A(new_n7297), .B(new_n7223), .Y(new_n7298_1));
  nor_5  g04950(.A(new_n7298_1), .B(new_n3873), .Y(new_n7299));
  xnor_4 g04951(.A(n8920), .B(n8581), .Y(new_n7300));
  nor_5  g04952(.A(new_n7300), .B(new_n3876), .Y(new_n7301));
  not_8  g04953(.A(new_n7298_1), .Y(new_n7302));
  xnor_4 g04954(.A(new_n7302), .B(new_n3873), .Y(new_n7303));
  and_5  g04955(.A(new_n7303), .B(new_n7301), .Y(new_n7304));
  nor_5  g04956(.A(new_n7304), .B(new_n7299), .Y(new_n7305_1));
  and_5  g04957(.A(new_n7305_1), .B(new_n7296), .Y(new_n7306));
  or_5   g04958(.A(new_n7306), .B(new_n7294), .Y(new_n7307));
  and_5  g04959(.A(new_n7307), .B(new_n7291), .Y(new_n7308_1));
  nor_5  g04960(.A(new_n7308_1), .B(new_n7289), .Y(new_n7309));
  nor_5  g04961(.A(new_n7309), .B(new_n7287), .Y(new_n7310));
  nor_5  g04962(.A(new_n7310), .B(new_n7286), .Y(new_n7311));
  nor_5  g04963(.A(new_n7311), .B(new_n7284), .Y(new_n7312));
  nor_5  g04964(.A(new_n7312), .B(new_n7283), .Y(new_n7313_1));
  nor_5  g04965(.A(new_n7313_1), .B(new_n7280_1), .Y(new_n7314));
  nor_5  g04966(.A(new_n7314), .B(new_n7279), .Y(new_n7315));
  nor_5  g04967(.A(new_n7315), .B(new_n7277_1), .Y(new_n7316));
  nor_5  g04968(.A(new_n7316), .B(new_n7276), .Y(new_n7317));
  nor_5  g04969(.A(new_n7317), .B(new_n7272), .Y(new_n7318));
  nor_5  g04970(.A(new_n7318), .B(new_n7271), .Y(new_n7319));
  and_5  g04971(.A(new_n7319), .B(new_n7267), .Y(new_n7320));
  nor_5  g04972(.A(new_n7320), .B(new_n7265), .Y(new_n7321));
  xnor_4 g04973(.A(new_n7321), .B(new_n7261), .Y(new_n7322));
  not_8  g04974(.A(new_n7322), .Y(new_n7323));
  nor_5  g04975(.A(n11898), .B(new_n4798), .Y(new_n7324));
  xnor_4 g04976(.A(n11898), .B(n2979), .Y(new_n7325));
  nor_5  g04977(.A(n19941), .B(new_n4801), .Y(new_n7326));
  xnor_4 g04978(.A(n19941), .B(n647), .Y(new_n7327));
  not_8  g04979(.A(n20409), .Y(new_n7328));
  nor_5  g04980(.A(new_n7328), .B(n1099), .Y(new_n7329));
  xnor_4 g04981(.A(n20409), .B(n1099), .Y(new_n7330_1));
  nor_5  g04982(.A(new_n3725_1), .B(n2113), .Y(new_n7331));
  xnor_4 g04983(.A(n25749), .B(n2113), .Y(new_n7332));
  nor_5  g04984(.A(n21134), .B(new_n3774), .Y(new_n7333));
  xnor_4 g04985(.A(n21134), .B(n3161), .Y(new_n7334));
  nor_5  g04986(.A(new_n3778), .B(n6369), .Y(new_n7335_1));
  xnor_4 g04987(.A(n9003), .B(n6369), .Y(new_n7336));
  nor_5  g04988(.A(n25797), .B(new_n3784), .Y(new_n7337));
  xnor_4 g04989(.A(n25797), .B(n4957), .Y(new_n7338));
  nor_5  g04990(.A(new_n4178), .B(n7524), .Y(new_n7339_1));
  nor_5  g04991(.A(n15967), .B(new_n3788), .Y(new_n7340));
  nor_5  g04992(.A(n15743), .B(new_n3752), .Y(new_n7341));
  or_5   g04993(.A(new_n3794_1), .B(n13319), .Y(new_n7342));
  nor_5  g04994(.A(new_n3756), .B(n20658), .Y(new_n7343));
  and_5  g04995(.A(new_n7343), .B(new_n7342), .Y(new_n7344));
  nor_5  g04996(.A(new_n7344), .B(new_n7341), .Y(new_n7345));
  nor_5  g04997(.A(new_n7345), .B(new_n7340), .Y(new_n7346_1));
  nor_5  g04998(.A(new_n7346_1), .B(new_n7339_1), .Y(new_n7347));
  and_5  g04999(.A(new_n7347), .B(new_n7338), .Y(new_n7348));
  or_5   g05000(.A(new_n7348), .B(new_n7337), .Y(new_n7349_1));
  and_5  g05001(.A(new_n7349_1), .B(new_n7336), .Y(new_n7350));
  or_5   g05002(.A(new_n7350), .B(new_n7335_1), .Y(new_n7351));
  and_5  g05003(.A(new_n7351), .B(new_n7334), .Y(new_n7352));
  or_5   g05004(.A(new_n7352), .B(new_n7333), .Y(new_n7353));
  and_5  g05005(.A(new_n7353), .B(new_n7332), .Y(new_n7354));
  or_5   g05006(.A(new_n7354), .B(new_n7331), .Y(new_n7355));
  and_5  g05007(.A(new_n7355), .B(new_n7330_1), .Y(new_n7356));
  or_5   g05008(.A(new_n7356), .B(new_n7329), .Y(new_n7357));
  and_5  g05009(.A(new_n7357), .B(new_n7327), .Y(new_n7358));
  or_5   g05010(.A(new_n7358), .B(new_n7326), .Y(new_n7359));
  and_5  g05011(.A(new_n7359), .B(new_n7325), .Y(new_n7360));
  nor_5  g05012(.A(new_n7360), .B(new_n7324), .Y(new_n7361));
  not_8  g05013(.A(new_n7361), .Y(new_n7362));
  xnor_4 g05014(.A(new_n7362), .B(new_n7323), .Y(new_n7363_1));
  xor_4  g05015(.A(new_n7359), .B(new_n7325), .Y(new_n7364));
  xor_4  g05016(.A(new_n7319), .B(new_n7267), .Y(new_n7365));
  nor_5  g05017(.A(new_n7365), .B(new_n7364), .Y(new_n7366));
  xnor_4 g05018(.A(new_n7365), .B(new_n7364), .Y(new_n7367));
  xor_4  g05019(.A(new_n7357), .B(new_n7327), .Y(new_n7368));
  xnor_4 g05020(.A(new_n7317), .B(new_n7272), .Y(new_n7369));
  nor_5  g05021(.A(new_n7369), .B(new_n7368), .Y(new_n7370));
  xnor_4 g05022(.A(new_n7369), .B(new_n7368), .Y(new_n7371));
  xor_4  g05023(.A(new_n7355), .B(new_n7330_1), .Y(new_n7372));
  xnor_4 g05024(.A(new_n7315), .B(new_n7277_1), .Y(new_n7373));
  nor_5  g05025(.A(new_n7373), .B(new_n7372), .Y(new_n7374));
  xnor_4 g05026(.A(new_n7373), .B(new_n7372), .Y(new_n7375));
  xor_4  g05027(.A(new_n7353), .B(new_n7332), .Y(new_n7376));
  xnor_4 g05028(.A(new_n7313_1), .B(new_n7280_1), .Y(new_n7377_1));
  nor_5  g05029(.A(new_n7377_1), .B(new_n7376), .Y(new_n7378));
  xnor_4 g05030(.A(new_n7377_1), .B(new_n7376), .Y(new_n7379));
  xor_4  g05031(.A(new_n7351), .B(new_n7334), .Y(new_n7380));
  xnor_4 g05032(.A(new_n7311), .B(new_n7284), .Y(new_n7381));
  nor_5  g05033(.A(new_n7381), .B(new_n7380), .Y(new_n7382));
  xnor_4 g05034(.A(new_n7381), .B(new_n7380), .Y(new_n7383));
  xor_4  g05035(.A(new_n7349_1), .B(new_n7336), .Y(new_n7384));
  xnor_4 g05036(.A(new_n7309), .B(new_n7287), .Y(new_n7385));
  nor_5  g05037(.A(new_n7385), .B(new_n7384), .Y(new_n7386));
  xnor_4 g05038(.A(new_n7385), .B(new_n7384), .Y(new_n7387));
  nor_5  g05039(.A(new_n7306), .B(new_n7294), .Y(new_n7388));
  xnor_4 g05040(.A(new_n7388), .B(new_n7291), .Y(new_n7389));
  xnor_4 g05041(.A(new_n7347), .B(new_n7338), .Y(new_n7390_1));
  and_5  g05042(.A(new_n7390_1), .B(new_n7389), .Y(new_n7391));
  xnor_4 g05043(.A(new_n7305_1), .B(new_n7296), .Y(new_n7392));
  not_8  g05044(.A(new_n7392), .Y(new_n7393));
  xnor_4 g05045(.A(n15967), .B(n7524), .Y(new_n7394));
  xnor_4 g05046(.A(new_n7394), .B(new_n7345), .Y(new_n7395));
  and_5  g05047(.A(new_n7395), .B(new_n7393), .Y(new_n7396));
  xnor_4 g05048(.A(new_n7395), .B(new_n7393), .Y(new_n7397));
  xnor_4 g05049(.A(n25435), .B(n20658), .Y(new_n7398));
  not_8  g05050(.A(new_n7300), .Y(new_n7399));
  xnor_4 g05051(.A(new_n7399), .B(new_n3876), .Y(new_n7400));
  not_8  g05052(.A(new_n7400), .Y(new_n7401));
  nor_5  g05053(.A(new_n7401), .B(new_n7398), .Y(new_n7402));
  xnor_4 g05054(.A(n15743), .B(n13319), .Y(new_n7403_1));
  xnor_4 g05055(.A(new_n7403_1), .B(new_n7343), .Y(new_n7404));
  nor_5  g05056(.A(new_n7404), .B(new_n7402), .Y(new_n7405));
  xnor_4 g05057(.A(new_n7303), .B(new_n7301), .Y(new_n7406));
  not_8  g05058(.A(new_n7406), .Y(new_n7407));
  xnor_4 g05059(.A(new_n7404), .B(new_n7402), .Y(new_n7408_1));
  nor_5  g05060(.A(new_n7408_1), .B(new_n7407), .Y(new_n7409));
  nor_5  g05061(.A(new_n7409), .B(new_n7405), .Y(new_n7410));
  nor_5  g05062(.A(new_n7410), .B(new_n7397), .Y(new_n7411));
  nor_5  g05063(.A(new_n7411), .B(new_n7396), .Y(new_n7412));
  xnor_4 g05064(.A(new_n7390_1), .B(new_n7389), .Y(new_n7413));
  nor_5  g05065(.A(new_n7413), .B(new_n7412), .Y(new_n7414));
  nor_5  g05066(.A(new_n7414), .B(new_n7391), .Y(new_n7415));
  nor_5  g05067(.A(new_n7415), .B(new_n7387), .Y(new_n7416));
  nor_5  g05068(.A(new_n7416), .B(new_n7386), .Y(new_n7417));
  nor_5  g05069(.A(new_n7417), .B(new_n7383), .Y(new_n7418));
  nor_5  g05070(.A(new_n7418), .B(new_n7382), .Y(new_n7419));
  nor_5  g05071(.A(new_n7419), .B(new_n7379), .Y(new_n7420));
  nor_5  g05072(.A(new_n7420), .B(new_n7378), .Y(new_n7421_1));
  nor_5  g05073(.A(new_n7421_1), .B(new_n7375), .Y(new_n7422));
  nor_5  g05074(.A(new_n7422), .B(new_n7374), .Y(new_n7423));
  nor_5  g05075(.A(new_n7423), .B(new_n7371), .Y(new_n7424));
  nor_5  g05076(.A(new_n7424), .B(new_n7370), .Y(new_n7425));
  nor_5  g05077(.A(new_n7425), .B(new_n7367), .Y(new_n7426));
  nor_5  g05078(.A(new_n7426), .B(new_n7366), .Y(new_n7427));
  xnor_4 g05079(.A(new_n7427), .B(new_n7363_1), .Y(n809));
  not_8  g05080(.A(n2978), .Y(new_n7429));
  nor_5  g05081(.A(n19282), .B(new_n7429), .Y(new_n7430));
  xnor_4 g05082(.A(n19282), .B(n2978), .Y(new_n7431));
  nor_5  g05083(.A(new_n6744), .B(n12657), .Y(new_n7432_1));
  xnor_4 g05084(.A(n23697), .B(n12657), .Y(new_n7433));
  nor_5  g05085(.A(n17077), .B(new_n6748), .Y(new_n7434));
  xnor_4 g05086(.A(n17077), .B(n2289), .Y(new_n7435));
  nor_5  g05087(.A(n26510), .B(new_n6752), .Y(new_n7436));
  xnor_4 g05088(.A(n26510), .B(n1112), .Y(new_n7437_1));
  nor_5  g05089(.A(n23068), .B(new_n6756), .Y(new_n7438));
  xnor_4 g05090(.A(n23068), .B(n20179), .Y(new_n7439));
  not_8  g05091(.A(n19228), .Y(new_n7440));
  nor_5  g05092(.A(n19514), .B(new_n7440), .Y(new_n7441));
  xnor_4 g05093(.A(n19514), .B(n19228), .Y(new_n7442));
  nor_5  g05094(.A(new_n6763), .B(n10053), .Y(new_n7443));
  xnor_4 g05095(.A(n15539), .B(n10053), .Y(new_n7444));
  nor_5  g05096(.A(new_n2947), .B(n8052), .Y(new_n7445));
  nor_5  g05097(.A(n8399), .B(new_n6767), .Y(new_n7446));
  nor_5  g05098(.A(n10158), .B(new_n3824), .Y(new_n7447));
  not_8  g05099(.A(n10158), .Y(new_n7448));
  nor_5  g05100(.A(new_n7448), .B(n9507), .Y(new_n7449));
  nor_5  g05101(.A(new_n2952), .B(n18962), .Y(new_n7450));
  not_8  g05102(.A(new_n7450), .Y(new_n7451));
  nor_5  g05103(.A(new_n7451), .B(new_n7449), .Y(new_n7452));
  nor_5  g05104(.A(new_n7452), .B(new_n7447), .Y(new_n7453));
  nor_5  g05105(.A(new_n7453), .B(new_n7446), .Y(new_n7454));
  nor_5  g05106(.A(new_n7454), .B(new_n7445), .Y(new_n7455));
  and_5  g05107(.A(new_n7455), .B(new_n7444), .Y(new_n7456));
  or_5   g05108(.A(new_n7456), .B(new_n7443), .Y(new_n7457));
  and_5  g05109(.A(new_n7457), .B(new_n7442), .Y(new_n7458));
  or_5   g05110(.A(new_n7458), .B(new_n7441), .Y(new_n7459));
  and_5  g05111(.A(new_n7459), .B(new_n7439), .Y(new_n7460_1));
  or_5   g05112(.A(new_n7460_1), .B(new_n7438), .Y(new_n7461));
  and_5  g05113(.A(new_n7461), .B(new_n7437_1), .Y(new_n7462));
  or_5   g05114(.A(new_n7462), .B(new_n7436), .Y(new_n7463));
  and_5  g05115(.A(new_n7463), .B(new_n7435), .Y(new_n7464));
  or_5   g05116(.A(new_n7464), .B(new_n7434), .Y(new_n7465));
  and_5  g05117(.A(new_n7465), .B(new_n7433), .Y(new_n7466));
  or_5   g05118(.A(new_n7466), .B(new_n7432_1), .Y(new_n7467));
  and_5  g05119(.A(new_n7467), .B(new_n7431), .Y(new_n7468));
  nor_5  g05120(.A(new_n7468), .B(new_n7430), .Y(new_n7469));
  nor_5  g05121(.A(n26986), .B(n22626), .Y(new_n7470));
  not_8  g05122(.A(new_n2424), .Y(new_n7471));
  nor_5  g05123(.A(new_n2431), .B(new_n7471), .Y(new_n7472));
  not_8  g05124(.A(new_n7472), .Y(new_n7473));
  xnor_4 g05125(.A(n4256), .B(n1654), .Y(new_n7474));
  nor_5  g05126(.A(n22332), .B(n13783), .Y(new_n7475_1));
  or_5   g05127(.A(new_n2428), .B(new_n2427), .Y(new_n7476));
  and_5  g05128(.A(new_n7476), .B(new_n2426), .Y(new_n7477_1));
  nor_5  g05129(.A(new_n7477_1), .B(new_n7475_1), .Y(new_n7478));
  xnor_4 g05130(.A(new_n7478), .B(new_n7474), .Y(new_n7479));
  nor_5  g05131(.A(new_n7479), .B(new_n7473), .Y(new_n7480));
  not_8  g05132(.A(new_n7480), .Y(new_n7481));
  not_8  g05133(.A(n14440), .Y(new_n7482));
  xnor_4 g05134(.A(n21287), .B(new_n7482), .Y(new_n7483));
  nor_5  g05135(.A(n4256), .B(n1654), .Y(new_n7484));
  nor_5  g05136(.A(new_n7478), .B(new_n7474), .Y(new_n7485));
  nor_5  g05137(.A(new_n7485), .B(new_n7484), .Y(new_n7486));
  xnor_4 g05138(.A(new_n7486), .B(new_n7483), .Y(new_n7487));
  not_8  g05139(.A(new_n7487), .Y(new_n7488));
  nor_5  g05140(.A(new_n7488), .B(new_n7481), .Y(new_n7489));
  xnor_4 g05141(.A(n26986), .B(n22626), .Y(new_n7490));
  nor_5  g05142(.A(n21287), .B(n14440), .Y(new_n7491));
  or_5   g05143(.A(new_n7485), .B(new_n7484), .Y(new_n7492));
  and_5  g05144(.A(new_n7492), .B(new_n7483), .Y(new_n7493));
  nor_5  g05145(.A(new_n7493), .B(new_n7491), .Y(new_n7494));
  xor_4  g05146(.A(new_n7494), .B(new_n7490), .Y(new_n7495));
  and_5  g05147(.A(new_n7495), .B(new_n7489), .Y(new_n7496));
  and_5  g05148(.A(new_n7496), .B(new_n7470), .Y(new_n7497));
  nor_5  g05149(.A(new_n7494), .B(new_n7490), .Y(new_n7498));
  nor_5  g05150(.A(new_n7498), .B(new_n7470), .Y(new_n7499));
  not_8  g05151(.A(new_n7499), .Y(new_n7500));
  nor_5  g05152(.A(new_n7500), .B(new_n7496), .Y(new_n7501));
  nor_5  g05153(.A(new_n7501), .B(new_n7497), .Y(new_n7502));
  nor_5  g05154(.A(n13494), .B(n3425), .Y(new_n7503));
  xnor_4 g05155(.A(n13494), .B(new_n3217), .Y(new_n7504));
  not_8  g05156(.A(new_n7504), .Y(new_n7505));
  nor_5  g05157(.A(n25345), .B(n9967), .Y(new_n7506));
  xnor_4 g05158(.A(n25345), .B(new_n3198), .Y(new_n7507_1));
  not_8  g05159(.A(n20946), .Y(new_n7508));
  nor_5  g05160(.A(new_n7508), .B(new_n5506), .Y(new_n7509));
  or_5   g05161(.A(n20946), .B(n9655), .Y(new_n7510));
  nor_5  g05162(.A(n13490), .B(n7751), .Y(new_n7511));
  nor_5  g05163(.A(new_n2459), .B(new_n2433), .Y(new_n7512));
  nor_5  g05164(.A(new_n7512), .B(new_n7511), .Y(new_n7513));
  and_5  g05165(.A(new_n7513), .B(new_n7510), .Y(new_n7514_1));
  nor_5  g05166(.A(new_n7514_1), .B(new_n7509), .Y(new_n7515));
  and_5  g05167(.A(new_n7515), .B(new_n7507_1), .Y(new_n7516));
  nor_5  g05168(.A(new_n7516), .B(new_n7506), .Y(new_n7517));
  nor_5  g05169(.A(new_n7517), .B(new_n7505), .Y(new_n7518));
  nor_5  g05170(.A(new_n7518), .B(new_n7503), .Y(new_n7519));
  and_5  g05171(.A(new_n7519), .B(new_n7502), .Y(new_n7520));
  or_5   g05172(.A(new_n7519), .B(new_n7502), .Y(new_n7521));
  xnor_4 g05173(.A(new_n7494), .B(new_n7490), .Y(new_n7522));
  xnor_4 g05174(.A(new_n7522), .B(new_n7489), .Y(new_n7523));
  xnor_4 g05175(.A(new_n7517), .B(new_n7505), .Y(new_n7524_1));
  nor_5  g05176(.A(new_n7524_1), .B(new_n7523), .Y(new_n7525));
  xnor_4 g05177(.A(new_n7524_1), .B(new_n7523), .Y(new_n7526));
  xnor_4 g05178(.A(new_n7488), .B(new_n7480), .Y(new_n7527));
  xnor_4 g05179(.A(new_n7515), .B(new_n7507_1), .Y(new_n7528));
  nor_5  g05180(.A(new_n7528), .B(new_n7527), .Y(new_n7529));
  xnor_4 g05181(.A(new_n7528), .B(new_n7527), .Y(new_n7530));
  xnor_4 g05182(.A(new_n7479), .B(new_n7472), .Y(new_n7531));
  xnor_4 g05183(.A(n20946), .B(n9655), .Y(new_n7532));
  xnor_4 g05184(.A(new_n7532), .B(new_n7513), .Y(new_n7533));
  nor_5  g05185(.A(new_n7533), .B(new_n7531), .Y(new_n7534));
  xnor_4 g05186(.A(new_n7533), .B(new_n7531), .Y(new_n7535));
  nor_5  g05187(.A(new_n2460), .B(new_n2432), .Y(new_n7536));
  nor_5  g05188(.A(new_n2500), .B(new_n2461), .Y(new_n7537));
  nor_5  g05189(.A(new_n7537), .B(new_n7536), .Y(new_n7538));
  nor_5  g05190(.A(new_n7538), .B(new_n7535), .Y(new_n7539));
  nor_5  g05191(.A(new_n7539), .B(new_n7534), .Y(new_n7540));
  nor_5  g05192(.A(new_n7540), .B(new_n7530), .Y(new_n7541));
  nor_5  g05193(.A(new_n7541), .B(new_n7529), .Y(new_n7542));
  nor_5  g05194(.A(new_n7542), .B(new_n7526), .Y(new_n7543));
  nor_5  g05195(.A(new_n7543), .B(new_n7525), .Y(new_n7544));
  and_5  g05196(.A(new_n7544), .B(new_n7521), .Y(new_n7545));
  or_5   g05197(.A(new_n7545), .B(new_n7497), .Y(new_n7546));
  nor_5  g05198(.A(new_n7546), .B(new_n7520), .Y(new_n7547));
  xnor_4 g05199(.A(new_n7547), .B(new_n7469), .Y(new_n7548));
  xnor_4 g05200(.A(new_n7519), .B(new_n7502), .Y(new_n7549));
  xnor_4 g05201(.A(new_n7549), .B(new_n7544), .Y(new_n7550));
  nor_5  g05202(.A(new_n7550), .B(new_n7469), .Y(new_n7551));
  xnor_4 g05203(.A(new_n7550), .B(new_n7469), .Y(new_n7552));
  xor_4  g05204(.A(new_n7467), .B(new_n7431), .Y(new_n7553));
  xnor_4 g05205(.A(new_n7542), .B(new_n7526), .Y(new_n7554));
  nor_5  g05206(.A(new_n7554), .B(new_n7553), .Y(new_n7555));
  xnor_4 g05207(.A(new_n7554), .B(new_n7553), .Y(new_n7556));
  xor_4  g05208(.A(new_n7465), .B(new_n7433), .Y(new_n7557));
  xnor_4 g05209(.A(new_n7540), .B(new_n7530), .Y(new_n7558_1));
  nor_5  g05210(.A(new_n7558_1), .B(new_n7557), .Y(new_n7559));
  xnor_4 g05211(.A(new_n7558_1), .B(new_n7557), .Y(new_n7560));
  xor_4  g05212(.A(new_n7463), .B(new_n7435), .Y(new_n7561));
  xnor_4 g05213(.A(new_n7538), .B(new_n7535), .Y(new_n7562));
  nor_5  g05214(.A(new_n7562), .B(new_n7561), .Y(new_n7563));
  xnor_4 g05215(.A(new_n7562), .B(new_n7561), .Y(new_n7564));
  xor_4  g05216(.A(new_n7461), .B(new_n7437_1), .Y(new_n7565));
  nor_5  g05217(.A(new_n7565), .B(new_n2501), .Y(new_n7566_1));
  xnor_4 g05218(.A(new_n7565), .B(new_n2501), .Y(new_n7567));
  xor_4  g05219(.A(new_n7459), .B(new_n7439), .Y(new_n7568));
  nor_5  g05220(.A(new_n7568), .B(new_n2504), .Y(new_n7569_1));
  xnor_4 g05221(.A(new_n7568), .B(new_n2504), .Y(new_n7570));
  xor_4  g05222(.A(new_n7457), .B(new_n7442), .Y(new_n7571));
  nor_5  g05223(.A(new_n7571), .B(new_n2508), .Y(new_n7572_1));
  xnor_4 g05224(.A(new_n7571), .B(new_n2508), .Y(new_n7573));
  xnor_4 g05225(.A(new_n7455), .B(new_n7444), .Y(new_n7574));
  and_5  g05226(.A(new_n7574), .B(new_n2513_1), .Y(new_n7575_1));
  xnor_4 g05227(.A(new_n7574), .B(new_n2513_1), .Y(new_n7576));
  xnor_4 g05228(.A(n8399), .B(n8052), .Y(new_n7577));
  xnor_4 g05229(.A(new_n7577), .B(new_n7453), .Y(new_n7578));
  and_5  g05230(.A(new_n7578), .B(new_n2516), .Y(new_n7579));
  xnor_4 g05231(.A(new_n7578), .B(new_n2516), .Y(new_n7580));
  xnor_4 g05232(.A(n26979), .B(n18962), .Y(new_n7581));
  or_5   g05233(.A(new_n7581), .B(new_n2523), .Y(new_n7582));
  xnor_4 g05234(.A(n10158), .B(n9507), .Y(new_n7583));
  xnor_4 g05235(.A(new_n7583), .B(new_n7451), .Y(new_n7584));
  and_5  g05236(.A(new_n7584), .B(new_n7582), .Y(new_n7585_1));
  xor_4  g05237(.A(new_n7584), .B(new_n7582), .Y(new_n7586));
  and_5  g05238(.A(new_n7586), .B(new_n2529), .Y(new_n7587));
  nor_5  g05239(.A(new_n7587), .B(new_n7585_1), .Y(new_n7588_1));
  nor_5  g05240(.A(new_n7588_1), .B(new_n7580), .Y(new_n7589));
  nor_5  g05241(.A(new_n7589), .B(new_n7579), .Y(new_n7590));
  nor_5  g05242(.A(new_n7590), .B(new_n7576), .Y(new_n7591));
  nor_5  g05243(.A(new_n7591), .B(new_n7575_1), .Y(new_n7592));
  nor_5  g05244(.A(new_n7592), .B(new_n7573), .Y(new_n7593_1));
  nor_5  g05245(.A(new_n7593_1), .B(new_n7572_1), .Y(new_n7594));
  nor_5  g05246(.A(new_n7594), .B(new_n7570), .Y(new_n7595));
  nor_5  g05247(.A(new_n7595), .B(new_n7569_1), .Y(new_n7596));
  nor_5  g05248(.A(new_n7596), .B(new_n7567), .Y(new_n7597));
  nor_5  g05249(.A(new_n7597), .B(new_n7566_1), .Y(new_n7598_1));
  nor_5  g05250(.A(new_n7598_1), .B(new_n7564), .Y(new_n7599));
  nor_5  g05251(.A(new_n7599), .B(new_n7563), .Y(new_n7600));
  nor_5  g05252(.A(new_n7600), .B(new_n7560), .Y(new_n7601));
  nor_5  g05253(.A(new_n7601), .B(new_n7559), .Y(new_n7602));
  nor_5  g05254(.A(new_n7602), .B(new_n7556), .Y(new_n7603));
  nor_5  g05255(.A(new_n7603), .B(new_n7555), .Y(new_n7604));
  nor_5  g05256(.A(new_n7604), .B(new_n7552), .Y(new_n7605));
  nor_5  g05257(.A(new_n7605), .B(new_n7551), .Y(new_n7606));
  xnor_4 g05258(.A(new_n7606), .B(new_n7548), .Y(n819));
  not_8  g05259(.A(n8856), .Y(new_n7608));
  nor_5  g05260(.A(n22626), .B(new_n7608), .Y(new_n7609));
  xnor_4 g05261(.A(n22626), .B(n8856), .Y(new_n7610_1));
  nor_5  g05262(.A(n14440), .B(new_n3405), .Y(new_n7611));
  xnor_4 g05263(.A(n14440), .B(n14130), .Y(new_n7612));
  not_8  g05264(.A(n1654), .Y(new_n7613));
  and_5  g05265(.A(n16482), .B(new_n7613), .Y(new_n7614));
  xnor_4 g05266(.A(n16482), .B(n1654), .Y(new_n7615));
  and_5  g05267(.A(new_n2425), .B(n9942), .Y(new_n7616_1));
  xnor_4 g05268(.A(n13783), .B(n9942), .Y(new_n7617));
  not_8  g05269(.A(n26660), .Y(new_n7618));
  and_5  g05270(.A(new_n7618), .B(n25643), .Y(new_n7619));
  xnor_4 g05271(.A(n26660), .B(n25643), .Y(new_n7620));
  nor_5  g05272(.A(new_n5116), .B(n3018), .Y(new_n7621));
  xnor_4 g05273(.A(n9557), .B(n3018), .Y(new_n7622));
  nor_5  g05274(.A(n3480), .B(new_n5106), .Y(new_n7623));
  xnor_4 g05275(.A(n3480), .B(n3136), .Y(new_n7624));
  not_8  g05276(.A(n16722), .Y(new_n7625));
  nor_5  g05277(.A(new_n7625), .B(n6385), .Y(new_n7626));
  nor_5  g05278(.A(n16722), .B(new_n2359), .Y(new_n7627));
  nor_5  g05279(.A(n20138), .B(new_n5784), .Y(new_n7628));
  nor_5  g05280(.A(new_n2363_1), .B(n11486), .Y(new_n7629));
  nor_5  g05281(.A(new_n2383), .B(n9251), .Y(new_n7630_1));
  not_8  g05282(.A(new_n7630_1), .Y(new_n7631));
  nor_5  g05283(.A(new_n7631), .B(new_n7629), .Y(new_n7632));
  nor_5  g05284(.A(new_n7632), .B(new_n7628), .Y(new_n7633));
  nor_5  g05285(.A(new_n7633), .B(new_n7627), .Y(new_n7634));
  nor_5  g05286(.A(new_n7634), .B(new_n7626), .Y(new_n7635));
  and_5  g05287(.A(new_n7635), .B(new_n7624), .Y(new_n7636));
  or_5   g05288(.A(new_n7636), .B(new_n7623), .Y(new_n7637));
  and_5  g05289(.A(new_n7637), .B(new_n7622), .Y(new_n7638));
  or_5   g05290(.A(new_n7638), .B(new_n7621), .Y(new_n7639));
  and_5  g05291(.A(new_n7639), .B(new_n7620), .Y(new_n7640));
  or_5   g05292(.A(new_n7640), .B(new_n7619), .Y(new_n7641));
  and_5  g05293(.A(new_n7641), .B(new_n7617), .Y(new_n7642));
  or_5   g05294(.A(new_n7642), .B(new_n7616_1), .Y(new_n7643_1));
  and_5  g05295(.A(new_n7643_1), .B(new_n7615), .Y(new_n7644));
  or_5   g05296(.A(new_n7644), .B(new_n7614), .Y(new_n7645));
  and_5  g05297(.A(new_n7645), .B(new_n7612), .Y(new_n7646));
  or_5   g05298(.A(new_n7646), .B(new_n7611), .Y(new_n7647_1));
  and_5  g05299(.A(new_n7647_1), .B(new_n7610_1), .Y(new_n7648));
  nor_5  g05300(.A(new_n7648), .B(new_n7609), .Y(new_n7649));
  not_8  g05301(.A(new_n7649), .Y(new_n7650));
  nor_5  g05302(.A(n25120), .B(new_n5982), .Y(new_n7651));
  xnor_4 g05303(.A(n25120), .B(n3582), .Y(new_n7652));
  nor_5  g05304(.A(n8363), .B(new_n5985), .Y(new_n7653));
  xnor_4 g05305(.A(n8363), .B(n2145), .Y(new_n7654));
  nor_5  g05306(.A(n14680), .B(new_n5988), .Y(new_n7655));
  xnor_4 g05307(.A(n14680), .B(n5031), .Y(new_n7656));
  not_8  g05308(.A(n11044), .Y(new_n7657_1));
  nor_5  g05309(.A(n17250), .B(new_n7657_1), .Y(new_n7658));
  xnor_4 g05310(.A(n17250), .B(n11044), .Y(new_n7659));
  nor_5  g05311(.A(n23160), .B(new_n5994), .Y(new_n7660));
  xnor_4 g05312(.A(n23160), .B(n2421), .Y(new_n7661));
  not_8  g05313(.A(n987), .Y(new_n7662));
  nor_5  g05314(.A(n16524), .B(new_n7662), .Y(new_n7663));
  xnor_4 g05315(.A(n16524), .B(n987), .Y(new_n7664));
  not_8  g05316(.A(n20478), .Y(new_n7665));
  nor_5  g05317(.A(new_n7665), .B(n11056), .Y(new_n7666));
  xnor_4 g05318(.A(n20478), .B(n11056), .Y(new_n7667));
  not_8  g05319(.A(n15271), .Y(new_n7668));
  nor_5  g05320(.A(n26882), .B(new_n7668), .Y(new_n7669));
  not_8  g05321(.A(n26882), .Y(new_n7670_1));
  nor_5  g05322(.A(new_n7670_1), .B(n15271), .Y(new_n7671));
  not_8  g05323(.A(n22619), .Y(new_n7672));
  and_5  g05324(.A(n25877), .B(new_n7672), .Y(new_n7673));
  nor_5  g05325(.A(n25877), .B(new_n7672), .Y(new_n7674_1));
  nor_5  g05326(.A(new_n6629), .B(n6775), .Y(new_n7675));
  not_8  g05327(.A(new_n7675), .Y(new_n7676));
  nor_5  g05328(.A(new_n7676), .B(new_n7674_1), .Y(new_n7677));
  nor_5  g05329(.A(new_n7677), .B(new_n7673), .Y(new_n7678_1));
  nor_5  g05330(.A(new_n7678_1), .B(new_n7671), .Y(new_n7679_1));
  nor_5  g05331(.A(new_n7679_1), .B(new_n7669), .Y(new_n7680));
  and_5  g05332(.A(new_n7680), .B(new_n7667), .Y(new_n7681));
  or_5   g05333(.A(new_n7681), .B(new_n7666), .Y(new_n7682));
  and_5  g05334(.A(new_n7682), .B(new_n7664), .Y(new_n7683));
  or_5   g05335(.A(new_n7683), .B(new_n7663), .Y(new_n7684));
  and_5  g05336(.A(new_n7684), .B(new_n7661), .Y(new_n7685));
  or_5   g05337(.A(new_n7685), .B(new_n7660), .Y(new_n7686_1));
  and_5  g05338(.A(new_n7686_1), .B(new_n7659), .Y(new_n7687));
  or_5   g05339(.A(new_n7687), .B(new_n7658), .Y(new_n7688));
  and_5  g05340(.A(new_n7688), .B(new_n7656), .Y(new_n7689));
  or_5   g05341(.A(new_n7689), .B(new_n7655), .Y(new_n7690));
  and_5  g05342(.A(new_n7690), .B(new_n7654), .Y(new_n7691));
  or_5   g05343(.A(new_n7691), .B(new_n7653), .Y(new_n7692_1));
  and_5  g05344(.A(new_n7692_1), .B(new_n7652), .Y(new_n7693_1));
  nor_5  g05345(.A(new_n7693_1), .B(new_n7651), .Y(new_n7694));
  not_8  g05346(.A(new_n7694), .Y(new_n7695));
  xnor_4 g05347(.A(new_n7695), .B(new_n7650), .Y(new_n7696));
  nor_5  g05348(.A(new_n7691), .B(new_n7653), .Y(new_n7697));
  xnor_4 g05349(.A(new_n7697), .B(new_n7652), .Y(new_n7698_1));
  nor_5  g05350(.A(new_n7646), .B(new_n7611), .Y(new_n7699));
  xnor_4 g05351(.A(new_n7699), .B(new_n7610_1), .Y(new_n7700));
  nor_5  g05352(.A(new_n7700), .B(new_n7698_1), .Y(new_n7701));
  not_8  g05353(.A(new_n7698_1), .Y(new_n7702));
  not_8  g05354(.A(new_n7700), .Y(new_n7703));
  xnor_4 g05355(.A(new_n7703), .B(new_n7702), .Y(new_n7704));
  xor_4  g05356(.A(new_n7690), .B(new_n7654), .Y(new_n7705));
  xor_4  g05357(.A(new_n7645), .B(new_n7612), .Y(new_n7706));
  nor_5  g05358(.A(new_n7706), .B(new_n7705), .Y(new_n7707));
  xnor_4 g05359(.A(new_n7706), .B(new_n7705), .Y(new_n7708_1));
  nor_5  g05360(.A(new_n7687), .B(new_n7658), .Y(new_n7709));
  xnor_4 g05361(.A(new_n7709), .B(new_n7656), .Y(new_n7710));
  nor_5  g05362(.A(new_n7642), .B(new_n7616_1), .Y(new_n7711));
  xnor_4 g05363(.A(new_n7711), .B(new_n7615), .Y(new_n7712));
  nor_5  g05364(.A(new_n7712), .B(new_n7710), .Y(new_n7713));
  not_8  g05365(.A(new_n7710), .Y(new_n7714));
  not_8  g05366(.A(new_n7712), .Y(new_n7715));
  xnor_4 g05367(.A(new_n7715), .B(new_n7714), .Y(new_n7716));
  xor_4  g05368(.A(new_n7686_1), .B(new_n7659), .Y(new_n7717));
  xor_4  g05369(.A(new_n7641), .B(new_n7617), .Y(new_n7718));
  nor_5  g05370(.A(new_n7718), .B(new_n7717), .Y(new_n7719));
  xnor_4 g05371(.A(new_n7718), .B(new_n7717), .Y(new_n7720));
  xor_4  g05372(.A(new_n7684), .B(new_n7661), .Y(new_n7721_1));
  xor_4  g05373(.A(new_n7639), .B(new_n7620), .Y(new_n7722));
  nor_5  g05374(.A(new_n7722), .B(new_n7721_1), .Y(new_n7723));
  xnor_4 g05375(.A(new_n7722), .B(new_n7721_1), .Y(new_n7724));
  xor_4  g05376(.A(new_n7682), .B(new_n7664), .Y(new_n7725));
  xor_4  g05377(.A(new_n7637), .B(new_n7622), .Y(new_n7726));
  nor_5  g05378(.A(new_n7726), .B(new_n7725), .Y(new_n7727));
  xnor_4 g05379(.A(new_n7726), .B(new_n7725), .Y(new_n7728));
  xnor_4 g05380(.A(new_n7680), .B(new_n7667), .Y(new_n7729));
  not_8  g05381(.A(new_n7729), .Y(new_n7730));
  xor_4  g05382(.A(new_n7635), .B(new_n7624), .Y(new_n7731_1));
  nor_5  g05383(.A(new_n7731_1), .B(new_n7730), .Y(new_n7732));
  xnor_4 g05384(.A(new_n7731_1), .B(new_n7730), .Y(new_n7733));
  xnor_4 g05385(.A(n26882), .B(n15271), .Y(new_n7734));
  xnor_4 g05386(.A(new_n7734), .B(new_n7678_1), .Y(new_n7735));
  xnor_4 g05387(.A(n16722), .B(n6385), .Y(new_n7736));
  xnor_4 g05388(.A(new_n7736), .B(new_n7633), .Y(new_n7737));
  and_5  g05389(.A(new_n7737), .B(new_n7735), .Y(new_n7738));
  not_8  g05390(.A(new_n7735), .Y(new_n7739));
  xnor_4 g05391(.A(new_n7737), .B(new_n7739), .Y(new_n7740));
  xnor_4 g05392(.A(n25877), .B(n22619), .Y(new_n7741));
  xnor_4 g05393(.A(new_n7741), .B(new_n7676), .Y(new_n7742));
  not_8  g05394(.A(new_n7742), .Y(new_n7743));
  xnor_4 g05395(.A(n20138), .B(n11486), .Y(new_n7744));
  xnor_4 g05396(.A(new_n7744), .B(new_n7631), .Y(new_n7745));
  not_8  g05397(.A(new_n7745), .Y(new_n7746));
  nor_5  g05398(.A(new_n7746), .B(new_n7743), .Y(new_n7747));
  xnor_4 g05399(.A(n24323), .B(n6775), .Y(new_n7748));
  xnor_4 g05400(.A(n13781), .B(n9251), .Y(new_n7749));
  or_5   g05401(.A(new_n7749), .B(new_n7748), .Y(new_n7750));
  xnor_4 g05402(.A(new_n7745), .B(new_n7743), .Y(new_n7751_1));
  and_5  g05403(.A(new_n7751_1), .B(new_n7750), .Y(new_n7752));
  or_5   g05404(.A(new_n7752), .B(new_n7747), .Y(new_n7753));
  and_5  g05405(.A(new_n7753), .B(new_n7740), .Y(new_n7754));
  nor_5  g05406(.A(new_n7754), .B(new_n7738), .Y(new_n7755));
  nor_5  g05407(.A(new_n7755), .B(new_n7733), .Y(new_n7756));
  nor_5  g05408(.A(new_n7756), .B(new_n7732), .Y(new_n7757));
  nor_5  g05409(.A(new_n7757), .B(new_n7728), .Y(new_n7758));
  nor_5  g05410(.A(new_n7758), .B(new_n7727), .Y(new_n7759_1));
  nor_5  g05411(.A(new_n7759_1), .B(new_n7724), .Y(new_n7760));
  nor_5  g05412(.A(new_n7760), .B(new_n7723), .Y(new_n7761));
  nor_5  g05413(.A(new_n7761), .B(new_n7720), .Y(new_n7762));
  nor_5  g05414(.A(new_n7762), .B(new_n7719), .Y(new_n7763));
  nor_5  g05415(.A(new_n7763), .B(new_n7716), .Y(new_n7764));
  nor_5  g05416(.A(new_n7764), .B(new_n7713), .Y(new_n7765));
  nor_5  g05417(.A(new_n7765), .B(new_n7708_1), .Y(new_n7766));
  nor_5  g05418(.A(new_n7766), .B(new_n7707), .Y(new_n7767));
  nor_5  g05419(.A(new_n7767), .B(new_n7704), .Y(new_n7768));
  nor_5  g05420(.A(new_n7768), .B(new_n7701), .Y(new_n7769_1));
  xnor_4 g05421(.A(new_n7769_1), .B(new_n7696), .Y(new_n7770));
  not_8  g05422(.A(new_n7770), .Y(new_n7771));
  not_8  g05423(.A(n9554), .Y(new_n7772));
  not_8  g05424(.A(n26408), .Y(new_n7773_1));
  nor_5  g05425(.A(n15508), .B(n2809), .Y(new_n7774));
  not_8  g05426(.A(new_n7774), .Y(new_n7775));
  nor_5  g05427(.A(new_n7775), .B(n19680), .Y(new_n7776));
  not_8  g05428(.A(new_n7776), .Y(new_n7777));
  nor_5  g05429(.A(new_n7777), .B(n7421), .Y(new_n7778));
  not_8  g05430(.A(new_n7778), .Y(new_n7779));
  nor_5  g05431(.A(new_n7779), .B(n13453), .Y(new_n7780_1));
  not_8  g05432(.A(new_n7780_1), .Y(new_n7781));
  nor_5  g05433(.A(new_n7781), .B(n11630), .Y(new_n7782));
  not_8  g05434(.A(new_n7782), .Y(new_n7783));
  nor_5  g05435(.A(new_n7783), .B(n7377), .Y(new_n7784));
  not_8  g05436(.A(new_n7784), .Y(new_n7785));
  nor_5  g05437(.A(new_n7785), .B(n18227), .Y(new_n7786));
  and_5  g05438(.A(new_n7786), .B(new_n7773_1), .Y(new_n7787));
  and_5  g05439(.A(new_n7787), .B(new_n7772), .Y(new_n7788_1));
  xnor_4 g05440(.A(new_n7787), .B(n9554), .Y(new_n7789));
  nor_5  g05441(.A(new_n7789), .B(n9259), .Y(new_n7790));
  xnor_4 g05442(.A(new_n7786), .B(n26408), .Y(new_n7791));
  nor_5  g05443(.A(new_n7791), .B(n21489), .Y(new_n7792));
  xnor_4 g05444(.A(new_n7791), .B(new_n3583), .Y(new_n7793));
  xnor_4 g05445(.A(new_n7784), .B(n18227), .Y(new_n7794_1));
  nor_5  g05446(.A(new_n7794_1), .B(n20213), .Y(new_n7795));
  xnor_4 g05447(.A(new_n7794_1), .B(new_n4844), .Y(new_n7796));
  xnor_4 g05448(.A(new_n7782), .B(n7377), .Y(new_n7797));
  nor_5  g05449(.A(new_n7797), .B(n13912), .Y(new_n7798));
  xnor_4 g05450(.A(new_n7797), .B(new_n4848), .Y(new_n7799));
  xnor_4 g05451(.A(new_n7780_1), .B(n11630), .Y(new_n7800));
  nor_5  g05452(.A(new_n7800), .B(n7670), .Y(new_n7801));
  xnor_4 g05453(.A(new_n7800), .B(new_n4853), .Y(new_n7802));
  xnor_4 g05454(.A(new_n7778), .B(n13453), .Y(new_n7803));
  nor_5  g05455(.A(new_n7803), .B(n9598), .Y(new_n7804));
  xnor_4 g05456(.A(new_n7803), .B(new_n4857), .Y(new_n7805));
  xnor_4 g05457(.A(new_n7776), .B(n7421), .Y(new_n7806));
  nor_5  g05458(.A(new_n7806), .B(n22290), .Y(new_n7807));
  xnor_4 g05459(.A(new_n7774), .B(n19680), .Y(new_n7808));
  nor_5  g05460(.A(new_n7808), .B(n11273), .Y(new_n7809));
  xnor_4 g05461(.A(new_n7808), .B(new_n4867), .Y(new_n7810));
  xnor_4 g05462(.A(n15508), .B(new_n6616), .Y(new_n7811_1));
  nor_5  g05463(.A(new_n7811_1), .B(n25565), .Y(new_n7812));
  nor_5  g05464(.A(new_n3635), .B(new_n4818), .Y(new_n7813));
  xnor_4 g05465(.A(new_n7811_1), .B(n25565), .Y(new_n7814));
  nor_5  g05466(.A(new_n7814), .B(new_n7813), .Y(new_n7815));
  or_5   g05467(.A(new_n7815), .B(new_n7812), .Y(new_n7816));
  and_5  g05468(.A(new_n7816), .B(new_n7810), .Y(new_n7817));
  or_5   g05469(.A(new_n7817), .B(new_n7809), .Y(new_n7818));
  xnor_4 g05470(.A(new_n7806), .B(new_n4863), .Y(new_n7819));
  and_5  g05471(.A(new_n7819), .B(new_n7818), .Y(new_n7820));
  or_5   g05472(.A(new_n7820), .B(new_n7807), .Y(new_n7821));
  and_5  g05473(.A(new_n7821), .B(new_n7805), .Y(new_n7822));
  or_5   g05474(.A(new_n7822), .B(new_n7804), .Y(new_n7823));
  and_5  g05475(.A(new_n7823), .B(new_n7802), .Y(new_n7824));
  or_5   g05476(.A(new_n7824), .B(new_n7801), .Y(new_n7825));
  and_5  g05477(.A(new_n7825), .B(new_n7799), .Y(new_n7826));
  or_5   g05478(.A(new_n7826), .B(new_n7798), .Y(new_n7827));
  and_5  g05479(.A(new_n7827), .B(new_n7796), .Y(new_n7828));
  or_5   g05480(.A(new_n7828), .B(new_n7795), .Y(new_n7829));
  and_5  g05481(.A(new_n7829), .B(new_n7793), .Y(new_n7830_1));
  nor_5  g05482(.A(new_n7830_1), .B(new_n7792), .Y(new_n7831));
  and_5  g05483(.A(new_n7789), .B(n9259), .Y(new_n7832));
  nor_5  g05484(.A(new_n7832), .B(new_n7831), .Y(new_n7833));
  nor_5  g05485(.A(new_n7833), .B(new_n7790), .Y(new_n7834_1));
  nor_5  g05486(.A(new_n7834_1), .B(new_n7788_1), .Y(new_n7835));
  xnor_4 g05487(.A(new_n7835), .B(new_n7771), .Y(new_n7836));
  xnor_4 g05488(.A(new_n7767), .B(new_n7704), .Y(new_n7837));
  xnor_4 g05489(.A(new_n7789), .B(new_n4797), .Y(new_n7838));
  xnor_4 g05490(.A(new_n7838), .B(new_n7831), .Y(new_n7839));
  not_8  g05491(.A(new_n7839), .Y(new_n7840));
  nor_5  g05492(.A(new_n7840), .B(new_n7837), .Y(new_n7841_1));
  not_8  g05493(.A(new_n7837), .Y(new_n7842));
  xnor_4 g05494(.A(new_n7840), .B(new_n7842), .Y(new_n7843));
  xnor_4 g05495(.A(new_n7765), .B(new_n7708_1), .Y(new_n7844));
  not_8  g05496(.A(new_n7844), .Y(new_n7845));
  nor_5  g05497(.A(new_n7828), .B(new_n7795), .Y(new_n7846));
  xnor_4 g05498(.A(new_n7846), .B(new_n7793), .Y(new_n7847));
  nor_5  g05499(.A(new_n7847), .B(new_n7845), .Y(new_n7848));
  not_8  g05500(.A(new_n7847), .Y(new_n7849));
  xnor_4 g05501(.A(new_n7849), .B(new_n7845), .Y(new_n7850));
  xnor_4 g05502(.A(new_n7763), .B(new_n7716), .Y(new_n7851));
  not_8  g05503(.A(new_n7851), .Y(new_n7852));
  nor_5  g05504(.A(new_n7826), .B(new_n7798), .Y(new_n7853));
  xnor_4 g05505(.A(new_n7853), .B(new_n7796), .Y(new_n7854));
  nor_5  g05506(.A(new_n7854), .B(new_n7852), .Y(new_n7855));
  not_8  g05507(.A(new_n7854), .Y(new_n7856));
  xnor_4 g05508(.A(new_n7856), .B(new_n7852), .Y(new_n7857));
  xnor_4 g05509(.A(new_n7761), .B(new_n7720), .Y(new_n7858));
  nor_5  g05510(.A(new_n7824), .B(new_n7801), .Y(new_n7859));
  xnor_4 g05511(.A(new_n7859), .B(new_n7799), .Y(new_n7860));
  not_8  g05512(.A(new_n7860), .Y(new_n7861));
  nor_5  g05513(.A(new_n7861), .B(new_n7858), .Y(new_n7862));
  and_5  g05514(.A(new_n7861), .B(new_n7858), .Y(new_n7863));
  xnor_4 g05515(.A(new_n7759_1), .B(new_n7724), .Y(new_n7864));
  not_8  g05516(.A(new_n7864), .Y(new_n7865));
  xor_4  g05517(.A(new_n7823), .B(new_n7802), .Y(new_n7866));
  and_5  g05518(.A(new_n7866), .B(new_n7865), .Y(new_n7867));
  xnor_4 g05519(.A(new_n7866), .B(new_n7865), .Y(new_n7868));
  xor_4  g05520(.A(new_n7821), .B(new_n7805), .Y(new_n7869));
  not_8  g05521(.A(new_n7869), .Y(new_n7870));
  xnor_4 g05522(.A(new_n7757), .B(new_n7728), .Y(new_n7871));
  nor_5  g05523(.A(new_n7871), .B(new_n7870), .Y(new_n7872));
  xnor_4 g05524(.A(new_n7871), .B(new_n7870), .Y(new_n7873));
  xnor_4 g05525(.A(new_n7755), .B(new_n7733), .Y(new_n7874));
  nor_5  g05526(.A(new_n7817), .B(new_n7809), .Y(new_n7875));
  xnor_4 g05527(.A(new_n7819), .B(new_n7875), .Y(new_n7876_1));
  not_8  g05528(.A(new_n7876_1), .Y(new_n7877));
  nor_5  g05529(.A(new_n7877), .B(new_n7874), .Y(new_n7878));
  not_8  g05530(.A(new_n7874), .Y(new_n7879));
  or_5   g05531(.A(new_n7876_1), .B(new_n7879), .Y(new_n7880));
  nor_5  g05532(.A(new_n7752), .B(new_n7747), .Y(new_n7881));
  xnor_4 g05533(.A(new_n7881), .B(new_n7740), .Y(new_n7882));
  xor_4  g05534(.A(new_n7751_1), .B(new_n7750), .Y(new_n7883));
  not_8  g05535(.A(new_n7883), .Y(new_n7884_1));
  xnor_4 g05536(.A(new_n7814), .B(new_n7813), .Y(new_n7885));
  nor_5  g05537(.A(new_n7885), .B(new_n7884_1), .Y(new_n7886));
  xnor_4 g05538(.A(n21993), .B(n15508), .Y(new_n7887));
  not_8  g05539(.A(new_n7748), .Y(new_n7888));
  xnor_4 g05540(.A(new_n7749), .B(new_n7888), .Y(new_n7889));
  not_8  g05541(.A(new_n7889), .Y(new_n7890));
  nor_5  g05542(.A(new_n7890), .B(new_n7887), .Y(new_n7891));
  xnor_4 g05543(.A(new_n7885), .B(new_n7884_1), .Y(new_n7892));
  nor_5  g05544(.A(new_n7892), .B(new_n7891), .Y(new_n7893));
  nor_5  g05545(.A(new_n7893), .B(new_n7886), .Y(new_n7894));
  not_8  g05546(.A(new_n7894), .Y(new_n7895));
  nor_5  g05547(.A(new_n7895), .B(new_n7882), .Y(new_n7896));
  nor_5  g05548(.A(new_n7815), .B(new_n7812), .Y(new_n7897));
  xnor_4 g05549(.A(new_n7897), .B(new_n7810), .Y(new_n7898));
  not_8  g05550(.A(new_n7898), .Y(new_n7899));
  xnor_4 g05551(.A(new_n7894), .B(new_n7882), .Y(new_n7900));
  and_5  g05552(.A(new_n7900), .B(new_n7899), .Y(new_n7901));
  nor_5  g05553(.A(new_n7901), .B(new_n7896), .Y(new_n7902));
  and_5  g05554(.A(new_n7902), .B(new_n7880), .Y(new_n7903));
  nor_5  g05555(.A(new_n7903), .B(new_n7878), .Y(new_n7904));
  nor_5  g05556(.A(new_n7904), .B(new_n7873), .Y(new_n7905));
  nor_5  g05557(.A(new_n7905), .B(new_n7872), .Y(new_n7906));
  nor_5  g05558(.A(new_n7906), .B(new_n7868), .Y(new_n7907));
  nor_5  g05559(.A(new_n7907), .B(new_n7867), .Y(new_n7908));
  nor_5  g05560(.A(new_n7908), .B(new_n7863), .Y(new_n7909));
  nor_5  g05561(.A(new_n7909), .B(new_n7862), .Y(new_n7910));
  and_5  g05562(.A(new_n7910), .B(new_n7857), .Y(new_n7911));
  or_5   g05563(.A(new_n7911), .B(new_n7855), .Y(new_n7912));
  and_5  g05564(.A(new_n7912), .B(new_n7850), .Y(new_n7913));
  nor_5  g05565(.A(new_n7913), .B(new_n7848), .Y(new_n7914));
  and_5  g05566(.A(new_n7914), .B(new_n7843), .Y(new_n7915));
  nor_5  g05567(.A(new_n7915), .B(new_n7841_1), .Y(new_n7916));
  xor_4  g05568(.A(new_n7916), .B(new_n7836), .Y(n829));
  not_8  g05569(.A(n14826), .Y(new_n7918));
  xnor_4 g05570(.A(n23272), .B(new_n7918), .Y(new_n7919));
  nor_5  g05571(.A(n23493), .B(n11481), .Y(new_n7920));
  xnor_4 g05572(.A(n23493), .B(new_n4361), .Y(new_n7921));
  nor_5  g05573(.A(n16439), .B(n10275), .Y(new_n7922));
  not_8  g05574(.A(n10275), .Y(new_n7923));
  xnor_4 g05575(.A(n16439), .B(new_n7923), .Y(new_n7924));
  nor_5  g05576(.A(n15241), .B(n15146), .Y(new_n7925));
  not_8  g05577(.A(n15146), .Y(new_n7926));
  xnor_4 g05578(.A(n15241), .B(new_n7926), .Y(new_n7927));
  nor_5  g05579(.A(n11579), .B(n7678), .Y(new_n7928));
  xnor_4 g05580(.A(n11579), .B(new_n4373), .Y(new_n7929));
  nor_5  g05581(.A(n3785), .B(n21), .Y(new_n7930));
  not_8  g05582(.A(n21), .Y(new_n7931));
  xnor_4 g05583(.A(n3785), .B(new_n7931), .Y(new_n7932));
  nor_5  g05584(.A(n20250), .B(n1682), .Y(new_n7933));
  not_8  g05585(.A(n1682), .Y(new_n7934));
  xnor_4 g05586(.A(n20250), .B(new_n7934), .Y(new_n7935));
  nor_5  g05587(.A(n7963), .B(n5822), .Y(new_n7936));
  xnor_4 g05588(.A(n7963), .B(new_n4384), .Y(new_n7937_1));
  nor_5  g05589(.A(n26443), .B(n10017), .Y(new_n7938));
  not_8  g05590(.A(n3618), .Y(new_n7939));
  or_5   g05591(.A(new_n7939), .B(new_n4394), .Y(new_n7940));
  not_8  g05592(.A(n10017), .Y(new_n7941));
  xnor_4 g05593(.A(n26443), .B(new_n7941), .Y(new_n7942));
  and_5  g05594(.A(new_n7942), .B(new_n7940), .Y(new_n7943_1));
  or_5   g05595(.A(new_n7943_1), .B(new_n7938), .Y(new_n7944));
  and_5  g05596(.A(new_n7944), .B(new_n7937_1), .Y(new_n7945));
  or_5   g05597(.A(new_n7945), .B(new_n7936), .Y(new_n7946));
  and_5  g05598(.A(new_n7946), .B(new_n7935), .Y(new_n7947));
  or_5   g05599(.A(new_n7947), .B(new_n7933), .Y(new_n7948));
  and_5  g05600(.A(new_n7948), .B(new_n7932), .Y(new_n7949_1));
  or_5   g05601(.A(new_n7949_1), .B(new_n7930), .Y(new_n7950_1));
  and_5  g05602(.A(new_n7950_1), .B(new_n7929), .Y(new_n7951));
  or_5   g05603(.A(new_n7951), .B(new_n7928), .Y(new_n7952));
  and_5  g05604(.A(new_n7952), .B(new_n7927), .Y(new_n7953));
  or_5   g05605(.A(new_n7953), .B(new_n7925), .Y(new_n7954));
  and_5  g05606(.A(new_n7954), .B(new_n7924), .Y(new_n7955));
  or_5   g05607(.A(new_n7955), .B(new_n7922), .Y(new_n7956));
  and_5  g05608(.A(new_n7956), .B(new_n7921), .Y(new_n7957));
  nor_5  g05609(.A(new_n7957), .B(new_n7920), .Y(new_n7958));
  xnor_4 g05610(.A(new_n7958), .B(new_n7919), .Y(new_n7959_1));
  nor_5  g05611(.A(new_n7959_1), .B(n22764), .Y(new_n7960));
  not_8  g05612(.A(new_n7959_1), .Y(new_n7961));
  xnor_4 g05613(.A(new_n7961), .B(n22764), .Y(new_n7962));
  nor_5  g05614(.A(new_n7955), .B(new_n7922), .Y(new_n7963_1));
  xnor_4 g05615(.A(new_n7963_1), .B(new_n7921), .Y(new_n7964));
  nor_5  g05616(.A(new_n7964), .B(n26264), .Y(new_n7965));
  not_8  g05617(.A(new_n7964), .Y(new_n7966));
  xnor_4 g05618(.A(new_n7966), .B(n26264), .Y(new_n7967));
  nor_5  g05619(.A(new_n7953), .B(new_n7925), .Y(new_n7968_1));
  xnor_4 g05620(.A(new_n7968_1), .B(new_n7924), .Y(new_n7969));
  nor_5  g05621(.A(new_n7969), .B(n7841), .Y(new_n7970));
  not_8  g05622(.A(new_n7969), .Y(new_n7971));
  xnor_4 g05623(.A(new_n7971), .B(n7841), .Y(new_n7972));
  nor_5  g05624(.A(new_n7951), .B(new_n7928), .Y(new_n7973));
  xnor_4 g05625(.A(new_n7973), .B(new_n7927), .Y(new_n7974));
  nor_5  g05626(.A(new_n7974), .B(n16812), .Y(new_n7975));
  not_8  g05627(.A(new_n7974), .Y(new_n7976));
  xnor_4 g05628(.A(new_n7976), .B(n16812), .Y(new_n7977));
  nor_5  g05629(.A(new_n7949_1), .B(new_n7930), .Y(new_n7978));
  xnor_4 g05630(.A(new_n7978), .B(new_n7929), .Y(new_n7979));
  nor_5  g05631(.A(new_n7979), .B(n25068), .Y(new_n7980));
  not_8  g05632(.A(new_n7979), .Y(new_n7981));
  xnor_4 g05633(.A(new_n7981), .B(n25068), .Y(new_n7982));
  nor_5  g05634(.A(new_n7947), .B(new_n7933), .Y(new_n7983));
  xnor_4 g05635(.A(new_n7983), .B(new_n7932), .Y(new_n7984));
  nor_5  g05636(.A(new_n7984), .B(n2331), .Y(new_n7985));
  not_8  g05637(.A(new_n7984), .Y(new_n7986));
  xnor_4 g05638(.A(new_n7986), .B(n2331), .Y(new_n7987));
  nor_5  g05639(.A(new_n7945), .B(new_n7936), .Y(new_n7988));
  xnor_4 g05640(.A(new_n7988), .B(new_n7935), .Y(new_n7989));
  nor_5  g05641(.A(new_n7989), .B(n22631), .Y(new_n7990));
  not_8  g05642(.A(new_n7989), .Y(new_n7991));
  xnor_4 g05643(.A(new_n7991), .B(n22631), .Y(new_n7992_1));
  not_8  g05644(.A(n16743), .Y(new_n7993));
  xor_4  g05645(.A(new_n7944), .B(new_n7937_1), .Y(new_n7994));
  not_8  g05646(.A(new_n7994), .Y(new_n7995));
  nor_5  g05647(.A(new_n7995), .B(new_n7993), .Y(new_n7996));
  xnor_4 g05648(.A(new_n7995), .B(n16743), .Y(new_n7997));
  not_8  g05649(.A(n15258), .Y(new_n7998));
  nor_5  g05650(.A(new_n2543), .B(n4588), .Y(new_n7999_1));
  and_5  g05651(.A(new_n7999_1), .B(new_n7998), .Y(new_n8000));
  nor_5  g05652(.A(new_n7939), .B(new_n4394), .Y(new_n8001));
  xnor_4 g05653(.A(new_n7942), .B(new_n8001), .Y(new_n8002));
  not_8  g05654(.A(new_n8002), .Y(new_n8003));
  xnor_4 g05655(.A(new_n7999_1), .B(n15258), .Y(new_n8004));
  and_5  g05656(.A(new_n8004), .B(new_n8003), .Y(new_n8005));
  nor_5  g05657(.A(new_n8005), .B(new_n8000), .Y(new_n8006_1));
  and_5  g05658(.A(new_n8006_1), .B(new_n7997), .Y(new_n8007));
  nor_5  g05659(.A(new_n8007), .B(new_n7996), .Y(new_n8008));
  and_5  g05660(.A(new_n8008), .B(new_n7992_1), .Y(new_n8009));
  or_5   g05661(.A(new_n8009), .B(new_n7990), .Y(new_n8010));
  and_5  g05662(.A(new_n8010), .B(new_n7987), .Y(new_n8011));
  or_5   g05663(.A(new_n8011), .B(new_n7985), .Y(new_n8012));
  and_5  g05664(.A(new_n8012), .B(new_n7982), .Y(new_n8013));
  or_5   g05665(.A(new_n8013), .B(new_n7980), .Y(new_n8014));
  and_5  g05666(.A(new_n8014), .B(new_n7977), .Y(new_n8015));
  or_5   g05667(.A(new_n8015), .B(new_n7975), .Y(new_n8016));
  and_5  g05668(.A(new_n8016), .B(new_n7972), .Y(new_n8017));
  or_5   g05669(.A(new_n8017), .B(new_n7970), .Y(new_n8018));
  and_5  g05670(.A(new_n8018), .B(new_n7967), .Y(new_n8019));
  or_5   g05671(.A(new_n8019), .B(new_n7965), .Y(new_n8020));
  and_5  g05672(.A(new_n8020), .B(new_n7962), .Y(new_n8021));
  nor_5  g05673(.A(new_n8021), .B(new_n7960), .Y(new_n8022));
  nor_5  g05674(.A(n23272), .B(n14826), .Y(new_n8023));
  or_5   g05675(.A(new_n7957), .B(new_n7920), .Y(new_n8024));
  and_5  g05676(.A(new_n8024), .B(new_n7919), .Y(new_n8025));
  nor_5  g05677(.A(new_n8025), .B(new_n8023), .Y(new_n8026));
  not_8  g05678(.A(new_n8026), .Y(new_n8027_1));
  and_5  g05679(.A(new_n8027_1), .B(new_n8022), .Y(new_n8028));
  nor_5  g05680(.A(n18105), .B(new_n5686), .Y(new_n8029));
  xnor_4 g05681(.A(n18105), .B(n12702), .Y(new_n8030));
  nor_5  g05682(.A(new_n5611), .B(n24196), .Y(new_n8031_1));
  xnor_4 g05683(.A(n26797), .B(n24196), .Y(new_n8032));
  not_8  g05684(.A(n23913), .Y(new_n8033));
  nor_5  g05685(.A(new_n8033), .B(n16376), .Y(new_n8034));
  xnor_4 g05686(.A(n23913), .B(n16376), .Y(new_n8035));
  not_8  g05687(.A(n22554), .Y(new_n8036));
  nor_5  g05688(.A(n25381), .B(new_n8036), .Y(new_n8037));
  xnor_4 g05689(.A(n25381), .B(n22554), .Y(new_n8038));
  not_8  g05690(.A(n20429), .Y(new_n8039));
  nor_5  g05691(.A(new_n8039), .B(n12587), .Y(new_n8040));
  xnor_4 g05692(.A(n20429), .B(n12587), .Y(new_n8041));
  not_8  g05693(.A(n3909), .Y(new_n8042_1));
  nor_5  g05694(.A(new_n8042_1), .B(n268), .Y(new_n8043));
  xnor_4 g05695(.A(n3909), .B(n268), .Y(new_n8044));
  not_8  g05696(.A(n23974), .Y(new_n8045));
  nor_5  g05697(.A(n24879), .B(new_n8045), .Y(new_n8046));
  xnor_4 g05698(.A(n24879), .B(n23974), .Y(new_n8047));
  not_8  g05699(.A(n6785), .Y(new_n8048));
  nor_5  g05700(.A(new_n8048), .B(n2146), .Y(new_n8049));
  not_8  g05701(.A(n2146), .Y(new_n8050));
  nor_5  g05702(.A(n6785), .B(new_n8050), .Y(new_n8051));
  not_8  g05703(.A(n24032), .Y(new_n8052_1));
  nor_5  g05704(.A(new_n8052_1), .B(n22173), .Y(new_n8053));
  nor_5  g05705(.A(new_n4507), .B(n583), .Y(new_n8054));
  not_8  g05706(.A(n22173), .Y(new_n8055));
  or_5   g05707(.A(n24032), .B(new_n8055), .Y(new_n8056));
  and_5  g05708(.A(new_n8056), .B(new_n8054), .Y(new_n8057));
  nor_5  g05709(.A(new_n8057), .B(new_n8053), .Y(new_n8058));
  nor_5  g05710(.A(new_n8058), .B(new_n8051), .Y(new_n8059));
  nor_5  g05711(.A(new_n8059), .B(new_n8049), .Y(new_n8060));
  and_5  g05712(.A(new_n8060), .B(new_n8047), .Y(new_n8061));
  or_5   g05713(.A(new_n8061), .B(new_n8046), .Y(new_n8062));
  and_5  g05714(.A(new_n8062), .B(new_n8044), .Y(new_n8063));
  or_5   g05715(.A(new_n8063), .B(new_n8043), .Y(new_n8064));
  and_5  g05716(.A(new_n8064), .B(new_n8041), .Y(new_n8065));
  or_5   g05717(.A(new_n8065), .B(new_n8040), .Y(new_n8066));
  and_5  g05718(.A(new_n8066), .B(new_n8038), .Y(new_n8067_1));
  or_5   g05719(.A(new_n8067_1), .B(new_n8037), .Y(new_n8068));
  and_5  g05720(.A(new_n8068), .B(new_n8035), .Y(new_n8069));
  or_5   g05721(.A(new_n8069), .B(new_n8034), .Y(new_n8070));
  and_5  g05722(.A(new_n8070), .B(new_n8032), .Y(new_n8071));
  or_5   g05723(.A(new_n8071), .B(new_n8031_1), .Y(new_n8072));
  and_5  g05724(.A(new_n8072), .B(new_n8030), .Y(new_n8073));
  nor_5  g05725(.A(new_n8073), .B(new_n8029), .Y(new_n8074));
  not_8  g05726(.A(new_n8074), .Y(new_n8075));
  nor_5  g05727(.A(new_n8071), .B(new_n8031_1), .Y(new_n8076));
  xnor_4 g05728(.A(new_n8076), .B(new_n8030), .Y(new_n8077));
  nor_5  g05729(.A(new_n8077), .B(n1536), .Y(new_n8078));
  not_8  g05730(.A(new_n8077), .Y(new_n8079));
  xnor_4 g05731(.A(new_n8079), .B(n1536), .Y(new_n8080));
  xor_4  g05732(.A(new_n8070), .B(new_n8032), .Y(new_n8081));
  nor_5  g05733(.A(new_n8081), .B(n19454), .Y(new_n8082));
  xnor_4 g05734(.A(new_n8081), .B(n19454), .Y(new_n8083));
  xor_4  g05735(.A(new_n8068), .B(new_n8035), .Y(new_n8084));
  nor_5  g05736(.A(new_n8084), .B(n9445), .Y(new_n8085));
  xnor_4 g05737(.A(new_n8084), .B(n9445), .Y(new_n8086));
  xor_4  g05738(.A(new_n8066), .B(new_n8038), .Y(new_n8087));
  nor_5  g05739(.A(new_n8087), .B(n1279), .Y(new_n8088));
  xnor_4 g05740(.A(new_n8087), .B(n1279), .Y(new_n8089));
  nor_5  g05741(.A(new_n8063), .B(new_n8043), .Y(new_n8090));
  xnor_4 g05742(.A(new_n8090), .B(new_n8041), .Y(new_n8091));
  nor_5  g05743(.A(new_n8091), .B(n8324), .Y(new_n8092));
  not_8  g05744(.A(new_n8091), .Y(new_n8093));
  xnor_4 g05745(.A(new_n8093), .B(n8324), .Y(new_n8094));
  xor_4  g05746(.A(new_n8062), .B(new_n8044), .Y(new_n8095_1));
  nor_5  g05747(.A(new_n8095_1), .B(n12546), .Y(new_n8096));
  xnor_4 g05748(.A(new_n8095_1), .B(n12546), .Y(new_n8097));
  xnor_4 g05749(.A(new_n8060), .B(new_n8047), .Y(new_n8098));
  not_8  g05750(.A(new_n8098), .Y(new_n8099));
  nor_5  g05751(.A(new_n8099), .B(n21078), .Y(new_n8100));
  xnor_4 g05752(.A(new_n8098), .B(n21078), .Y(new_n8101));
  xnor_4 g05753(.A(n6785), .B(n2146), .Y(new_n8102));
  xnor_4 g05754(.A(new_n8102), .B(new_n8058), .Y(new_n8103_1));
  not_8  g05755(.A(new_n8103_1), .Y(new_n8104));
  and_5  g05756(.A(new_n8104), .B(n24485), .Y(new_n8105));
  or_5   g05757(.A(new_n8104), .B(n24485), .Y(new_n8106));
  xnor_4 g05758(.A(n24032), .B(n22173), .Y(new_n8107));
  xnor_4 g05759(.A(new_n8107), .B(new_n8054), .Y(new_n8108));
  nor_5  g05760(.A(new_n8108), .B(n2420), .Y(new_n8109_1));
  not_8  g05761(.A(n22201), .Y(new_n8110));
  or_5   g05762(.A(new_n2545), .B(new_n8110), .Y(new_n8111));
  not_8  g05763(.A(n2420), .Y(new_n8112));
  xnor_4 g05764(.A(new_n8108), .B(new_n8112), .Y(new_n8113));
  and_5  g05765(.A(new_n8113), .B(new_n8111), .Y(new_n8114));
  nor_5  g05766(.A(new_n8114), .B(new_n8109_1), .Y(new_n8115));
  and_5  g05767(.A(new_n8115), .B(new_n8106), .Y(new_n8116));
  nor_5  g05768(.A(new_n8116), .B(new_n8105), .Y(new_n8117));
  and_5  g05769(.A(new_n8117), .B(new_n8101), .Y(new_n8118));
  nor_5  g05770(.A(new_n8118), .B(new_n8100), .Y(new_n8119));
  nor_5  g05771(.A(new_n8119), .B(new_n8097), .Y(new_n8120));
  or_5   g05772(.A(new_n8120), .B(new_n8096), .Y(new_n8121));
  and_5  g05773(.A(new_n8121), .B(new_n8094), .Y(new_n8122));
  nor_5  g05774(.A(new_n8122), .B(new_n8092), .Y(new_n8123));
  nor_5  g05775(.A(new_n8123), .B(new_n8089), .Y(new_n8124));
  nor_5  g05776(.A(new_n8124), .B(new_n8088), .Y(new_n8125));
  nor_5  g05777(.A(new_n8125), .B(new_n8086), .Y(new_n8126));
  nor_5  g05778(.A(new_n8126), .B(new_n8085), .Y(new_n8127_1));
  nor_5  g05779(.A(new_n8127_1), .B(new_n8083), .Y(new_n8128));
  or_5   g05780(.A(new_n8128), .B(new_n8082), .Y(new_n8129));
  and_5  g05781(.A(new_n8129), .B(new_n8080), .Y(new_n8130_1));
  nor_5  g05782(.A(new_n8130_1), .B(new_n8078), .Y(new_n8131));
  not_8  g05783(.A(new_n8131), .Y(new_n8132));
  nor_5  g05784(.A(new_n8132), .B(new_n8075), .Y(new_n8133));
  xnor_4 g05785(.A(new_n8026), .B(new_n8022), .Y(new_n8134));
  xnor_4 g05786(.A(new_n8132), .B(new_n8074), .Y(new_n8135_1));
  nor_5  g05787(.A(new_n8135_1), .B(new_n8134), .Y(new_n8136));
  xnor_4 g05788(.A(new_n8135_1), .B(new_n8134), .Y(new_n8137));
  nor_5  g05789(.A(new_n8019), .B(new_n7965), .Y(new_n8138));
  xnor_4 g05790(.A(new_n8138), .B(new_n7962), .Y(new_n8139_1));
  xor_4  g05791(.A(new_n8129), .B(new_n8080), .Y(new_n8140));
  and_5  g05792(.A(new_n8140), .B(new_n8139_1), .Y(new_n8141));
  xnor_4 g05793(.A(new_n8140), .B(new_n8139_1), .Y(new_n8142));
  xor_4  g05794(.A(new_n8018), .B(new_n7967), .Y(new_n8143));
  not_8  g05795(.A(new_n8143), .Y(new_n8144));
  xnor_4 g05796(.A(new_n8127_1), .B(new_n8083), .Y(new_n8145));
  nor_5  g05797(.A(new_n8145), .B(new_n8144), .Y(new_n8146));
  xnor_4 g05798(.A(new_n8145), .B(new_n8144), .Y(new_n8147));
  xor_4  g05799(.A(new_n8016), .B(new_n7972), .Y(new_n8148_1));
  not_8  g05800(.A(new_n8148_1), .Y(new_n8149_1));
  xnor_4 g05801(.A(new_n8125), .B(new_n8086), .Y(new_n8150));
  nor_5  g05802(.A(new_n8150), .B(new_n8149_1), .Y(new_n8151));
  xnor_4 g05803(.A(new_n8150), .B(new_n8149_1), .Y(new_n8152));
  xor_4  g05804(.A(new_n8014), .B(new_n7977), .Y(new_n8153));
  not_8  g05805(.A(new_n8153), .Y(new_n8154));
  xnor_4 g05806(.A(new_n8123), .B(new_n8089), .Y(new_n8155));
  nor_5  g05807(.A(new_n8155), .B(new_n8154), .Y(new_n8156));
  xnor_4 g05808(.A(new_n8155), .B(new_n8154), .Y(new_n8157));
  nor_5  g05809(.A(new_n8011), .B(new_n7985), .Y(new_n8158));
  xnor_4 g05810(.A(new_n8158), .B(new_n7982), .Y(new_n8159_1));
  xor_4  g05811(.A(new_n8121), .B(new_n8094), .Y(new_n8160));
  and_5  g05812(.A(new_n8160), .B(new_n8159_1), .Y(new_n8161));
  xnor_4 g05813(.A(new_n8160), .B(new_n8159_1), .Y(new_n8162));
  xor_4  g05814(.A(new_n8010), .B(new_n7987), .Y(new_n8163));
  not_8  g05815(.A(new_n8163), .Y(new_n8164));
  xnor_4 g05816(.A(new_n8119), .B(new_n8097), .Y(new_n8165));
  nor_5  g05817(.A(new_n8165), .B(new_n8164), .Y(new_n8166));
  xnor_4 g05818(.A(new_n8165), .B(new_n8164), .Y(new_n8167));
  xnor_4 g05819(.A(new_n8008), .B(new_n7992_1), .Y(new_n8168));
  xnor_4 g05820(.A(new_n8117), .B(new_n8101), .Y(new_n8169));
  nor_5  g05821(.A(new_n8169), .B(new_n8168), .Y(new_n8170));
  xnor_4 g05822(.A(new_n8169), .B(new_n8168), .Y(new_n8171));
  xnor_4 g05823(.A(new_n8006_1), .B(new_n7997), .Y(new_n8172));
  not_8  g05824(.A(new_n8172), .Y(new_n8173));
  xnor_4 g05825(.A(new_n8104), .B(n24485), .Y(new_n8174));
  xnor_4 g05826(.A(new_n8174), .B(new_n8115), .Y(new_n8175));
  nor_5  g05827(.A(new_n8175), .B(new_n8173), .Y(new_n8176));
  xnor_4 g05828(.A(new_n8175), .B(new_n8172), .Y(new_n8177));
  xor_4  g05829(.A(new_n8113), .B(new_n8111), .Y(new_n8178));
  xnor_4 g05830(.A(new_n8004), .B(new_n8002), .Y(new_n8179_1));
  nor_5  g05831(.A(new_n8179_1), .B(new_n8178), .Y(new_n8180));
  not_8  g05832(.A(new_n2544), .Y(new_n8181));
  and_5  g05833(.A(new_n2546), .B(new_n8181), .Y(new_n8182));
  not_8  g05834(.A(new_n8179_1), .Y(new_n8183));
  xnor_4 g05835(.A(new_n8183), .B(new_n8178), .Y(new_n8184));
  and_5  g05836(.A(new_n8184), .B(new_n8182), .Y(new_n8185));
  nor_5  g05837(.A(new_n8185), .B(new_n8180), .Y(new_n8186));
  and_5  g05838(.A(new_n8186), .B(new_n8177), .Y(new_n8187));
  nor_5  g05839(.A(new_n8187), .B(new_n8176), .Y(new_n8188));
  nor_5  g05840(.A(new_n8188), .B(new_n8171), .Y(new_n8189));
  nor_5  g05841(.A(new_n8189), .B(new_n8170), .Y(new_n8190));
  nor_5  g05842(.A(new_n8190), .B(new_n8167), .Y(new_n8191));
  nor_5  g05843(.A(new_n8191), .B(new_n8166), .Y(new_n8192));
  nor_5  g05844(.A(new_n8192), .B(new_n8162), .Y(new_n8193));
  nor_5  g05845(.A(new_n8193), .B(new_n8161), .Y(new_n8194_1));
  nor_5  g05846(.A(new_n8194_1), .B(new_n8157), .Y(new_n8195));
  nor_5  g05847(.A(new_n8195), .B(new_n8156), .Y(new_n8196));
  nor_5  g05848(.A(new_n8196), .B(new_n8152), .Y(new_n8197));
  nor_5  g05849(.A(new_n8197), .B(new_n8151), .Y(new_n8198));
  nor_5  g05850(.A(new_n8198), .B(new_n8147), .Y(new_n8199));
  nor_5  g05851(.A(new_n8199), .B(new_n8146), .Y(new_n8200));
  nor_5  g05852(.A(new_n8200), .B(new_n8142), .Y(new_n8201));
  nor_5  g05853(.A(new_n8201), .B(new_n8141), .Y(new_n8202));
  nor_5  g05854(.A(new_n8202), .B(new_n8137), .Y(new_n8203));
  nor_5  g05855(.A(new_n8203), .B(new_n8136), .Y(new_n8204));
  xor_4  g05856(.A(new_n8204), .B(new_n8133), .Y(new_n8205));
  xnor_4 g05857(.A(new_n8205), .B(new_n8028), .Y(n849));
  xnor_4 g05858(.A(new_n2530), .B(new_n2529), .Y(n858));
  nor_5  g05859(.A(n16994), .B(n9246), .Y(new_n8208));
  not_8  g05860(.A(new_n8208), .Y(new_n8209));
  nor_5  g05861(.A(new_n8209), .B(n10096), .Y(new_n8210));
  not_8  g05862(.A(new_n8210), .Y(new_n8211));
  nor_5  g05863(.A(new_n8211), .B(n14790), .Y(new_n8212));
  not_8  g05864(.A(new_n8212), .Y(new_n8213));
  nor_5  g05865(.A(new_n8213), .B(n17251), .Y(new_n8214));
  not_8  g05866(.A(new_n8214), .Y(new_n8215_1));
  nor_5  g05867(.A(new_n8215_1), .B(n21674), .Y(new_n8216));
  not_8  g05868(.A(new_n8216), .Y(new_n8217));
  nor_5  g05869(.A(new_n8217), .B(n24638), .Y(new_n8218));
  not_8  g05870(.A(new_n8218), .Y(new_n8219));
  nor_5  g05871(.A(new_n8219), .B(n18444), .Y(new_n8220));
  not_8  g05872(.A(new_n8220), .Y(new_n8221));
  nor_5  g05873(.A(new_n8221), .B(n14899), .Y(new_n8222));
  xnor_4 g05874(.A(new_n8222), .B(n3506), .Y(new_n8223));
  xnor_4 g05875(.A(new_n8223), .B(n1314), .Y(new_n8224));
  xnor_4 g05876(.A(new_n8220), .B(n14899), .Y(new_n8225));
  and_5  g05877(.A(new_n8225), .B(n3306), .Y(new_n8226));
  or_5   g05878(.A(new_n8225), .B(n3306), .Y(new_n8227));
  xnor_4 g05879(.A(new_n8218), .B(n18444), .Y(new_n8228));
  nor_5  g05880(.A(new_n8228), .B(n22335), .Y(new_n8229));
  not_8  g05881(.A(n22335), .Y(new_n8230));
  xnor_4 g05882(.A(new_n8228), .B(new_n8230), .Y(new_n8231));
  xnor_4 g05883(.A(new_n8216), .B(n24638), .Y(new_n8232));
  nor_5  g05884(.A(new_n8232), .B(n24048), .Y(new_n8233));
  not_8  g05885(.A(n24048), .Y(new_n8234));
  xnor_4 g05886(.A(new_n8232), .B(new_n8234), .Y(new_n8235));
  xnor_4 g05887(.A(new_n8214), .B(n21674), .Y(new_n8236));
  nor_5  g05888(.A(new_n8236), .B(n1525), .Y(new_n8237));
  not_8  g05889(.A(n1525), .Y(new_n8238));
  xnor_4 g05890(.A(new_n8236), .B(new_n8238), .Y(new_n8239));
  xnor_4 g05891(.A(new_n8212), .B(n17251), .Y(new_n8240));
  nor_5  g05892(.A(new_n8240), .B(n16988), .Y(new_n8241));
  xnor_4 g05893(.A(new_n8240), .B(new_n4638), .Y(new_n8242));
  xnor_4 g05894(.A(new_n8210), .B(n14790), .Y(new_n8243));
  nor_5  g05895(.A(new_n8243), .B(n21779), .Y(new_n8244_1));
  xnor_4 g05896(.A(new_n8208), .B(n10096), .Y(new_n8245));
  nor_5  g05897(.A(new_n8245), .B(n5376), .Y(new_n8246));
  xnor_4 g05898(.A(new_n8245), .B(new_n4645), .Y(new_n8247));
  xnor_4 g05899(.A(n16994), .B(n9246), .Y(new_n8248));
  and_5  g05900(.A(new_n8248), .B(new_n4648), .Y(new_n8249));
  and_5  g05901(.A(n23120), .B(n9246), .Y(new_n8250));
  xnor_4 g05902(.A(new_n8248), .B(new_n4648), .Y(new_n8251));
  nor_5  g05903(.A(new_n8251), .B(new_n8250), .Y(new_n8252));
  or_5   g05904(.A(new_n8252), .B(new_n8249), .Y(new_n8253));
  and_5  g05905(.A(new_n8253), .B(new_n8247), .Y(new_n8254));
  or_5   g05906(.A(new_n8254), .B(new_n8246), .Y(new_n8255_1));
  xnor_4 g05907(.A(new_n8243), .B(new_n4641), .Y(new_n8256_1));
  and_5  g05908(.A(new_n8256_1), .B(new_n8255_1), .Y(new_n8257));
  or_5   g05909(.A(new_n8257), .B(new_n8244_1), .Y(new_n8258));
  and_5  g05910(.A(new_n8258), .B(new_n8242), .Y(new_n8259_1));
  or_5   g05911(.A(new_n8259_1), .B(new_n8241), .Y(new_n8260));
  and_5  g05912(.A(new_n8260), .B(new_n8239), .Y(new_n8261));
  or_5   g05913(.A(new_n8261), .B(new_n8237), .Y(new_n8262));
  and_5  g05914(.A(new_n8262), .B(new_n8235), .Y(new_n8263));
  or_5   g05915(.A(new_n8263), .B(new_n8233), .Y(new_n8264));
  and_5  g05916(.A(new_n8264), .B(new_n8231), .Y(new_n8265));
  nor_5  g05917(.A(new_n8265), .B(new_n8229), .Y(new_n8266));
  and_5  g05918(.A(new_n8266), .B(new_n8227), .Y(new_n8267_1));
  nor_5  g05919(.A(new_n8267_1), .B(new_n8226), .Y(new_n8268));
  xnor_4 g05920(.A(new_n8268), .B(new_n8224), .Y(new_n8269));
  nor_5  g05921(.A(new_n8269), .B(n22442), .Y(new_n8270));
  not_8  g05922(.A(n22442), .Y(new_n8271));
  xnor_4 g05923(.A(new_n8269), .B(new_n8271), .Y(new_n8272));
  not_8  g05924(.A(n468), .Y(new_n8273));
  xnor_4 g05925(.A(new_n8225), .B(n3306), .Y(new_n8274));
  xnor_4 g05926(.A(new_n8274), .B(new_n8266), .Y(new_n8275));
  nor_5  g05927(.A(new_n8275), .B(new_n8273), .Y(new_n8276_1));
  xnor_4 g05928(.A(new_n8275), .B(n468), .Y(new_n8277));
  xor_4  g05929(.A(new_n8264), .B(new_n8231), .Y(new_n8278));
  nor_5  g05930(.A(new_n8278), .B(n5400), .Y(new_n8279));
  not_8  g05931(.A(n5400), .Y(new_n8280));
  xnor_4 g05932(.A(new_n8278), .B(new_n8280), .Y(new_n8281));
  xor_4  g05933(.A(new_n8262), .B(new_n8235), .Y(new_n8282));
  nor_5  g05934(.A(new_n8282), .B(n23923), .Y(new_n8283));
  not_8  g05935(.A(n23923), .Y(new_n8284));
  xnor_4 g05936(.A(new_n8282), .B(new_n8284), .Y(new_n8285_1));
  xor_4  g05937(.A(new_n8260), .B(new_n8239), .Y(new_n8286));
  and_5  g05938(.A(new_n8286), .B(n329), .Y(new_n8287));
  or_5   g05939(.A(new_n8286), .B(n329), .Y(new_n8288_1));
  xor_4  g05940(.A(new_n8256_1), .B(new_n8255_1), .Y(new_n8289));
  nor_5  g05941(.A(new_n8289), .B(n2409), .Y(new_n8290));
  xnor_4 g05942(.A(new_n8289), .B(n2409), .Y(new_n8291));
  xor_4  g05943(.A(new_n8253), .B(new_n8247), .Y(new_n8292));
  nor_5  g05944(.A(new_n8292), .B(n8869), .Y(new_n8293));
  xor_4  g05945(.A(new_n8251), .B(new_n8250), .Y(new_n8294));
  nor_5  g05946(.A(new_n8294), .B(n10372), .Y(new_n8295));
  xnor_4 g05947(.A(n23120), .B(new_n3562), .Y(new_n8296));
  nor_5  g05948(.A(new_n8296), .B(new_n7024), .Y(new_n8297));
  xnor_4 g05949(.A(new_n8294), .B(n10372), .Y(new_n8298));
  nor_5  g05950(.A(new_n8298), .B(new_n8297), .Y(new_n8299));
  nor_5  g05951(.A(new_n8299), .B(new_n8295), .Y(new_n8300));
  xnor_4 g05952(.A(new_n8292), .B(n8869), .Y(new_n8301));
  nor_5  g05953(.A(new_n8301), .B(new_n8300), .Y(new_n8302));
  nor_5  g05954(.A(new_n8302), .B(new_n8293), .Y(new_n8303));
  nor_5  g05955(.A(new_n8303), .B(new_n8291), .Y(new_n8304));
  nor_5  g05956(.A(new_n8304), .B(new_n8290), .Y(new_n8305_1));
  nor_5  g05957(.A(new_n8305_1), .B(n24170), .Y(new_n8306_1));
  xor_4  g05958(.A(new_n8258), .B(new_n8242), .Y(new_n8307));
  xnor_4 g05959(.A(new_n8305_1), .B(n24170), .Y(new_n8308));
  nor_5  g05960(.A(new_n8308), .B(new_n8307), .Y(new_n8309_1));
  nor_5  g05961(.A(new_n8309_1), .B(new_n8306_1), .Y(new_n8310));
  and_5  g05962(.A(new_n8310), .B(new_n8288_1), .Y(new_n8311));
  nor_5  g05963(.A(new_n8311), .B(new_n8287), .Y(new_n8312));
  and_5  g05964(.A(new_n8312), .B(new_n8285_1), .Y(new_n8313));
  or_5   g05965(.A(new_n8313), .B(new_n8283), .Y(new_n8314));
  and_5  g05966(.A(new_n8314), .B(new_n8281), .Y(new_n8315));
  nor_5  g05967(.A(new_n8315), .B(new_n8279), .Y(new_n8316));
  and_5  g05968(.A(new_n8316), .B(new_n8277), .Y(new_n8317));
  nor_5  g05969(.A(new_n8317), .B(new_n8276_1), .Y(new_n8318));
  and_5  g05970(.A(new_n8318), .B(new_n8272), .Y(new_n8319));
  nor_5  g05971(.A(new_n8319), .B(new_n8270), .Y(new_n8320_1));
  nor_5  g05972(.A(new_n8223), .B(n1314), .Y(new_n8321_1));
  nor_5  g05973(.A(new_n8268), .B(new_n8321_1), .Y(new_n8322));
  not_8  g05974(.A(n3506), .Y(new_n8323));
  and_5  g05975(.A(new_n8222), .B(new_n8323), .Y(new_n8324_1));
  and_5  g05976(.A(new_n8223), .B(n1314), .Y(new_n8325));
  or_5   g05977(.A(new_n8325), .B(new_n8324_1), .Y(new_n8326));
  nor_5  g05978(.A(new_n8326), .B(new_n8322), .Y(new_n8327));
  xor_4  g05979(.A(new_n8327), .B(new_n8320_1), .Y(new_n8328));
  not_8  g05980(.A(new_n8328), .Y(new_n8329));
  nor_5  g05981(.A(new_n3472), .B(n26180), .Y(new_n8330));
  nor_5  g05982(.A(new_n3534), .B(new_n3473), .Y(new_n8331));
  nor_5  g05983(.A(new_n8331), .B(new_n8330), .Y(new_n8332));
  not_8  g05984(.A(new_n8332), .Y(new_n8333));
  and_5  g05985(.A(new_n3419), .B(new_n7608), .Y(new_n8334));
  nor_5  g05986(.A(new_n3420), .B(n25494), .Y(new_n8335));
  and_5  g05987(.A(new_n3420), .B(n25494), .Y(new_n8336));
  nor_5  g05988(.A(new_n3471), .B(new_n8336), .Y(new_n8337));
  nor_5  g05989(.A(new_n8337), .B(new_n8335), .Y(new_n8338));
  nor_5  g05990(.A(new_n8338), .B(new_n8334), .Y(new_n8339_1));
  xnor_4 g05991(.A(new_n8339_1), .B(new_n8333), .Y(new_n8340));
  xnor_4 g05992(.A(new_n8340), .B(new_n8329), .Y(new_n8341));
  xor_4  g05993(.A(new_n8318), .B(new_n8272), .Y(new_n8342));
  nor_5  g05994(.A(new_n8342), .B(new_n3535), .Y(new_n8343));
  xnor_4 g05995(.A(new_n8342), .B(new_n3535), .Y(new_n8344));
  xor_4  g05996(.A(new_n8316), .B(new_n8277), .Y(new_n8345));
  and_5  g05997(.A(new_n8345), .B(new_n3665_1), .Y(new_n8346));
  xnor_4 g05998(.A(new_n8345), .B(new_n3665_1), .Y(new_n8347));
  xor_4  g05999(.A(new_n8314), .B(new_n8281), .Y(new_n8348));
  nor_5  g06000(.A(new_n8348), .B(new_n3671), .Y(new_n8349));
  xnor_4 g06001(.A(new_n8348), .B(new_n3671), .Y(new_n8350));
  xor_4  g06002(.A(new_n8312), .B(new_n8285_1), .Y(new_n8351));
  nor_5  g06003(.A(new_n8351), .B(new_n3676), .Y(new_n8352));
  not_8  g06004(.A(n329), .Y(new_n8353));
  xnor_4 g06005(.A(new_n8286), .B(new_n8353), .Y(new_n8354));
  xnor_4 g06006(.A(new_n8354), .B(new_n8310), .Y(new_n8355));
  nor_5  g06007(.A(new_n8355), .B(new_n3681), .Y(new_n8356));
  xnor_4 g06008(.A(new_n8355), .B(new_n3681), .Y(new_n8357));
  xor_4  g06009(.A(new_n8308), .B(new_n8307), .Y(new_n8358));
  nor_5  g06010(.A(new_n8358), .B(new_n3686), .Y(new_n8359));
  xor_4  g06011(.A(new_n8303), .B(new_n8291), .Y(new_n8360));
  nor_5  g06012(.A(new_n8360), .B(new_n3690), .Y(new_n8361));
  xnor_4 g06013(.A(new_n8360), .B(new_n3690), .Y(new_n8362));
  xor_4  g06014(.A(new_n8301), .B(new_n8300), .Y(new_n8363_1));
  nor_5  g06015(.A(new_n8363_1), .B(new_n3696), .Y(new_n8364));
  xor_4  g06016(.A(new_n8298), .B(new_n8297), .Y(new_n8365));
  nor_5  g06017(.A(new_n8365), .B(new_n3702), .Y(new_n8366));
  not_8  g06018(.A(new_n3704), .Y(new_n8367));
  xnor_4 g06019(.A(new_n8296), .B(n7428), .Y(new_n8368));
  nor_5  g06020(.A(new_n8368), .B(new_n8367), .Y(new_n8369));
  xnor_4 g06021(.A(new_n8365), .B(new_n3702), .Y(new_n8370));
  nor_5  g06022(.A(new_n8370), .B(new_n8369), .Y(new_n8371));
  nor_5  g06023(.A(new_n8371), .B(new_n8366), .Y(new_n8372));
  xnor_4 g06024(.A(new_n8363_1), .B(new_n3696), .Y(new_n8373));
  nor_5  g06025(.A(new_n8373), .B(new_n8372), .Y(new_n8374));
  nor_5  g06026(.A(new_n8374), .B(new_n8364), .Y(new_n8375));
  nor_5  g06027(.A(new_n8375), .B(new_n8362), .Y(new_n8376_1));
  nor_5  g06028(.A(new_n8376_1), .B(new_n8361), .Y(new_n8377));
  xnor_4 g06029(.A(new_n8358), .B(new_n3686), .Y(new_n8378));
  nor_5  g06030(.A(new_n8378), .B(new_n8377), .Y(new_n8379));
  nor_5  g06031(.A(new_n8379), .B(new_n8359), .Y(new_n8380));
  nor_5  g06032(.A(new_n8380), .B(new_n8357), .Y(new_n8381_1));
  nor_5  g06033(.A(new_n8381_1), .B(new_n8356), .Y(new_n8382));
  xnor_4 g06034(.A(new_n8351), .B(new_n3676), .Y(new_n8383));
  nor_5  g06035(.A(new_n8383), .B(new_n8382), .Y(new_n8384));
  nor_5  g06036(.A(new_n8384), .B(new_n8352), .Y(new_n8385));
  nor_5  g06037(.A(new_n8385), .B(new_n8350), .Y(new_n8386));
  nor_5  g06038(.A(new_n8386), .B(new_n8349), .Y(new_n8387));
  nor_5  g06039(.A(new_n8387), .B(new_n8347), .Y(new_n8388));
  nor_5  g06040(.A(new_n8388), .B(new_n8346), .Y(new_n8389));
  nor_5  g06041(.A(new_n8389), .B(new_n8344), .Y(new_n8390));
  or_5   g06042(.A(new_n8390), .B(new_n8343), .Y(new_n8391));
  xnor_4 g06043(.A(new_n8391), .B(new_n8341), .Y(n873));
  xnor_4 g06044(.A(n4812), .B(n2731), .Y(new_n8393));
  not_8  g06045(.A(n24278), .Y(new_n8394));
  nor_5  g06046(.A(new_n8394), .B(n19911), .Y(new_n8395));
  xnor_4 g06047(.A(n24278), .B(n19911), .Y(new_n8396));
  nor_5  g06048(.A(n24618), .B(new_n2389), .Y(new_n8397));
  not_8  g06049(.A(n24618), .Y(new_n8398));
  nor_5  g06050(.A(new_n8398), .B(n13708), .Y(new_n8399_1));
  nor_5  g06051(.A(new_n3826), .B(n3952), .Y(new_n8400));
  nor_5  g06052(.A(n18409), .B(new_n2443), .Y(new_n8401));
  nor_5  g06053(.A(n12315), .B(new_n2381), .Y(new_n8402));
  not_8  g06054(.A(new_n8402), .Y(new_n8403));
  nor_5  g06055(.A(new_n8403), .B(new_n8401), .Y(new_n8404));
  nor_5  g06056(.A(new_n8404), .B(new_n8400), .Y(new_n8405_1));
  nor_5  g06057(.A(new_n8405_1), .B(new_n8399_1), .Y(new_n8406));
  nor_5  g06058(.A(new_n8406), .B(new_n8397), .Y(new_n8407));
  and_5  g06059(.A(new_n8407), .B(new_n8396), .Y(new_n8408_1));
  or_5   g06060(.A(new_n8408_1), .B(new_n8395), .Y(new_n8409));
  xor_4  g06061(.A(new_n8409), .B(new_n8393), .Y(new_n8410));
  xor_4  g06062(.A(new_n8410), .B(new_n5187), .Y(new_n8411));
  xnor_4 g06063(.A(new_n8407), .B(new_n8396), .Y(new_n8412));
  and_5  g06064(.A(new_n8412), .B(new_n5191), .Y(new_n8413));
  xnor_4 g06065(.A(n24618), .B(n13708), .Y(new_n8414));
  xnor_4 g06066(.A(new_n8414), .B(new_n8405_1), .Y(new_n8415));
  nor_5  g06067(.A(new_n8415), .B(new_n5195), .Y(new_n8416));
  xnor_4 g06068(.A(new_n8415), .B(new_n5195), .Y(new_n8417_1));
  xnor_4 g06069(.A(n12315), .B(n5704), .Y(new_n8418));
  nor_5  g06070(.A(new_n8418), .B(new_n5202), .Y(new_n8419));
  and_5  g06071(.A(new_n8419), .B(new_n5207), .Y(new_n8420));
  xnor_4 g06072(.A(new_n8419), .B(new_n5207), .Y(new_n8421));
  xnor_4 g06073(.A(n18409), .B(n3952), .Y(new_n8422));
  xnor_4 g06074(.A(new_n8422), .B(new_n8403), .Y(new_n8423));
  nor_5  g06075(.A(new_n8423), .B(new_n8421), .Y(new_n8424));
  nor_5  g06076(.A(new_n8424), .B(new_n8420), .Y(new_n8425));
  nor_5  g06077(.A(new_n8425), .B(new_n8417_1), .Y(new_n8426));
  nor_5  g06078(.A(new_n8426), .B(new_n8416), .Y(new_n8427));
  xnor_4 g06079(.A(new_n8412), .B(new_n5190), .Y(new_n8428));
  and_5  g06080(.A(new_n8428), .B(new_n8427), .Y(new_n8429));
  nor_5  g06081(.A(new_n8429), .B(new_n8413), .Y(new_n8430));
  xor_4  g06082(.A(new_n8430), .B(new_n8411), .Y(n879));
  not_8  g06083(.A(n18157), .Y(new_n8432_1));
  xnor_4 g06084(.A(new_n7991), .B(new_n8432_1), .Y(new_n8433));
  nor_5  g06085(.A(new_n7995), .B(n12161), .Y(new_n8434));
  nor_5  g06086(.A(new_n8002), .B(new_n7220), .Y(new_n8435));
  nor_5  g06087(.A(new_n2543), .B(new_n6628_1), .Y(new_n8436));
  xnor_4 g06088(.A(new_n8003), .B(new_n7220), .Y(new_n8437));
  and_5  g06089(.A(new_n8437), .B(new_n8436), .Y(new_n8438));
  nor_5  g06090(.A(new_n8438), .B(new_n8435), .Y(new_n8439_1));
  xnor_4 g06091(.A(new_n7995), .B(new_n7217), .Y(new_n8440));
  and_5  g06092(.A(new_n8440), .B(new_n8439_1), .Y(new_n8441));
  nor_5  g06093(.A(new_n8441), .B(new_n8434), .Y(new_n8442));
  xnor_4 g06094(.A(new_n8442), .B(new_n8433), .Y(new_n8443));
  xnor_4 g06095(.A(new_n8440), .B(new_n8439_1), .Y(new_n8444));
  not_8  g06096(.A(n14684), .Y(new_n8445));
  xnor_4 g06097(.A(new_n6610), .B(new_n8445), .Y(new_n8446));
  nor_5  g06098(.A(new_n6612_1), .B(n6631), .Y(new_n8447));
  or_5   g06099(.A(new_n6614), .B(new_n4183), .Y(new_n8448));
  xnor_4 g06100(.A(new_n6612_1), .B(new_n4180), .Y(new_n8449));
  and_5  g06101(.A(new_n8449), .B(new_n8448), .Y(new_n8450));
  or_5   g06102(.A(new_n8450), .B(new_n8447), .Y(new_n8451));
  xor_4  g06103(.A(new_n8451), .B(new_n8446), .Y(new_n8452));
  nor_5  g06104(.A(new_n8452), .B(new_n8444), .Y(new_n8453_1));
  xnor_4 g06105(.A(new_n8452), .B(new_n8444), .Y(new_n8454));
  xor_4  g06106(.A(new_n8449), .B(new_n8448), .Y(new_n8455));
  xor_4  g06107(.A(new_n8437), .B(new_n8436), .Y(new_n8456));
  nor_5  g06108(.A(new_n8456), .B(new_n8455), .Y(new_n8457));
  xnor_4 g06109(.A(new_n6614), .B(n24732), .Y(new_n8458));
  not_8  g06110(.A(new_n8458), .Y(new_n8459));
  xnor_4 g06111(.A(new_n2543), .B(n8581), .Y(new_n8460));
  nor_5  g06112(.A(new_n8460), .B(new_n8459), .Y(new_n8461));
  xnor_4 g06113(.A(new_n8456), .B(new_n8455), .Y(new_n8462));
  not_8  g06114(.A(new_n8462), .Y(new_n8463));
  and_5  g06115(.A(new_n8463), .B(new_n8461), .Y(new_n8464));
  nor_5  g06116(.A(new_n8464), .B(new_n8457), .Y(new_n8465));
  nor_5  g06117(.A(new_n8465), .B(new_n8454), .Y(new_n8466));
  nor_5  g06118(.A(new_n8466), .B(new_n8453_1), .Y(new_n8467));
  xnor_4 g06119(.A(new_n8467), .B(new_n8443), .Y(new_n8468));
  not_8  g06120(.A(n17035), .Y(new_n8469));
  xnor_4 g06121(.A(new_n6604), .B(new_n8469), .Y(new_n8470));
  nor_5  g06122(.A(new_n6610), .B(n14684), .Y(new_n8471));
  and_5  g06123(.A(new_n8451), .B(new_n8446), .Y(new_n8472));
  nor_5  g06124(.A(new_n8472), .B(new_n8471), .Y(new_n8473));
  xnor_4 g06125(.A(new_n8473), .B(new_n8470), .Y(new_n8474));
  xor_4  g06126(.A(new_n8474), .B(new_n8468), .Y(n887));
  xnor_4 g06127(.A(new_n6041), .B(new_n4917), .Y(new_n8476));
  nor_5  g06128(.A(new_n6045), .B(new_n4922), .Y(new_n8477));
  xnor_4 g06129(.A(new_n6047), .B(new_n4922), .Y(new_n8478));
  nor_5  g06130(.A(new_n6051), .B(new_n4927), .Y(new_n8479));
  xnor_4 g06131(.A(new_n6053), .B(new_n4927), .Y(new_n8480_1));
  nor_5  g06132(.A(new_n6057), .B(new_n4932), .Y(new_n8481));
  xnor_4 g06133(.A(new_n6059), .B(new_n4932), .Y(new_n8482));
  not_8  g06134(.A(n25872), .Y(new_n8483));
  nor_5  g06135(.A(new_n6063), .B(new_n8483), .Y(new_n8484));
  nor_5  g06136(.A(new_n6065), .B(n20259), .Y(new_n8485));
  or_5   g06137(.A(new_n5792), .B(new_n5002), .Y(new_n8486));
  xnor_4 g06138(.A(new_n6065), .B(new_n4939_1), .Y(new_n8487));
  and_5  g06139(.A(new_n8487), .B(new_n8486), .Y(new_n8488));
  nor_5  g06140(.A(new_n8488), .B(new_n8485), .Y(new_n8489_1));
  xnor_4 g06141(.A(new_n6072), .B(new_n8483), .Y(new_n8490));
  and_5  g06142(.A(new_n8490), .B(new_n8489_1), .Y(new_n8491));
  or_5   g06143(.A(new_n8491), .B(new_n8484), .Y(new_n8492));
  and_5  g06144(.A(new_n8492), .B(new_n8482), .Y(new_n8493));
  or_5   g06145(.A(new_n8493), .B(new_n8481), .Y(new_n8494));
  and_5  g06146(.A(new_n8494), .B(new_n8480_1), .Y(new_n8495));
  or_5   g06147(.A(new_n8495), .B(new_n8479), .Y(new_n8496));
  and_5  g06148(.A(new_n8496), .B(new_n8478), .Y(new_n8497));
  nor_5  g06149(.A(new_n8497), .B(new_n8477), .Y(new_n8498));
  xnor_4 g06150(.A(new_n8498), .B(new_n8476), .Y(new_n8499));
  not_8  g06151(.A(new_n8499), .Y(new_n8500));
  not_8  g06152(.A(n25119), .Y(new_n8501));
  xnor_4 g06153(.A(new_n2980), .B(new_n8501), .Y(new_n8502));
  not_8  g06154(.A(n1163), .Y(new_n8503));
  nor_5  g06155(.A(new_n2985_1), .B(new_n8503), .Y(new_n8504));
  nor_5  g06156(.A(new_n2990), .B(n18537), .Y(new_n8505_1));
  not_8  g06157(.A(n18537), .Y(new_n8506));
  xnor_4 g06158(.A(new_n2990), .B(new_n8506), .Y(new_n8507));
  nor_5  g06159(.A(new_n2996), .B(n7057), .Y(new_n8508));
  xor_4  g06160(.A(new_n2996), .B(n7057), .Y(new_n8509));
  not_8  g06161(.A(n8381), .Y(new_n8510_1));
  nor_5  g06162(.A(new_n3002), .B(new_n8510_1), .Y(new_n8511));
  xnor_4 g06163(.A(new_n3002), .B(n8381), .Y(new_n8512));
  nor_5  g06164(.A(new_n3063), .B(new_n5080), .Y(new_n8513));
  nor_5  g06165(.A(new_n8513), .B(n20235), .Y(new_n8514));
  xnor_4 g06166(.A(new_n8513), .B(new_n5040), .Y(new_n8515));
  and_5  g06167(.A(new_n8515), .B(new_n3008), .Y(new_n8516));
  nor_5  g06168(.A(new_n8516), .B(new_n8514), .Y(new_n8517));
  and_5  g06169(.A(new_n8517), .B(new_n8512), .Y(new_n8518));
  nor_5  g06170(.A(new_n8518), .B(new_n8511), .Y(new_n8519_1));
  and_5  g06171(.A(new_n8519_1), .B(new_n8509), .Y(new_n8520));
  or_5   g06172(.A(new_n8520), .B(new_n8508), .Y(new_n8521));
  and_5  g06173(.A(new_n8521), .B(new_n8507), .Y(new_n8522));
  nor_5  g06174(.A(new_n8522), .B(new_n8505_1), .Y(new_n8523));
  xnor_4 g06175(.A(new_n2986), .B(new_n8503), .Y(new_n8524));
  and_5  g06176(.A(new_n8524), .B(new_n8523), .Y(new_n8525));
  nor_5  g06177(.A(new_n8525), .B(new_n8504), .Y(new_n8526_1));
  xnor_4 g06178(.A(new_n8526_1), .B(new_n8502), .Y(new_n8527));
  xnor_4 g06179(.A(new_n8527), .B(new_n8500), .Y(new_n8528));
  nor_5  g06180(.A(new_n8495), .B(new_n8479), .Y(new_n8529));
  xnor_4 g06181(.A(new_n8529), .B(new_n8478), .Y(new_n8530));
  not_8  g06182(.A(new_n8530), .Y(new_n8531));
  xor_4  g06183(.A(new_n8524), .B(new_n8523), .Y(new_n8532));
  nor_5  g06184(.A(new_n8532), .B(new_n8531), .Y(new_n8533));
  xnor_4 g06185(.A(new_n8532), .B(new_n8531), .Y(new_n8534));
  xor_4  g06186(.A(new_n8521), .B(new_n8507), .Y(new_n8535_1));
  nor_5  g06187(.A(new_n8493), .B(new_n8481), .Y(new_n8536));
  xnor_4 g06188(.A(new_n8536), .B(new_n8480_1), .Y(new_n8537));
  and_5  g06189(.A(new_n8537), .B(new_n8535_1), .Y(new_n8538));
  xnor_4 g06190(.A(new_n8537), .B(new_n8535_1), .Y(new_n8539));
  xnor_4 g06191(.A(new_n8519_1), .B(new_n8509), .Y(new_n8540));
  nor_5  g06192(.A(new_n8491), .B(new_n8484), .Y(new_n8541));
  xnor_4 g06193(.A(new_n8541), .B(new_n8482), .Y(new_n8542));
  not_8  g06194(.A(new_n8542), .Y(new_n8543));
  nor_5  g06195(.A(new_n8543), .B(new_n8540), .Y(new_n8544));
  xnor_4 g06196(.A(new_n8543), .B(new_n8540), .Y(new_n8545));
  xnor_4 g06197(.A(new_n8517), .B(new_n8512), .Y(new_n8546));
  xnor_4 g06198(.A(new_n8490), .B(new_n8489_1), .Y(new_n8547));
  not_8  g06199(.A(new_n8547), .Y(new_n8548));
  and_5  g06200(.A(new_n8548), .B(new_n8546), .Y(new_n8549));
  xnor_4 g06201(.A(new_n8548), .B(new_n8546), .Y(new_n8550_1));
  nor_5  g06202(.A(new_n5792), .B(new_n5002), .Y(new_n8551));
  xnor_4 g06203(.A(new_n8487), .B(new_n8551), .Y(new_n8552));
  not_8  g06204(.A(new_n8552), .Y(new_n8553));
  xnor_4 g06205(.A(new_n8515), .B(new_n3009), .Y(new_n8554));
  and_5  g06206(.A(new_n8554), .B(new_n8553), .Y(new_n8555));
  xnor_4 g06207(.A(new_n5792), .B(n3925), .Y(new_n8556));
  not_8  g06208(.A(new_n8556), .Y(new_n8557));
  xnor_4 g06209(.A(new_n3063), .B(n12495), .Y(new_n8558));
  nor_5  g06210(.A(new_n8558), .B(new_n8557), .Y(new_n8559));
  xnor_4 g06211(.A(new_n8554), .B(new_n8552), .Y(new_n8560));
  and_5  g06212(.A(new_n8560), .B(new_n8559), .Y(new_n8561));
  nor_5  g06213(.A(new_n8561), .B(new_n8555), .Y(new_n8562));
  nor_5  g06214(.A(new_n8562), .B(new_n8550_1), .Y(new_n8563_1));
  nor_5  g06215(.A(new_n8563_1), .B(new_n8549), .Y(new_n8564));
  nor_5  g06216(.A(new_n8564), .B(new_n8545), .Y(new_n8565));
  nor_5  g06217(.A(new_n8565), .B(new_n8544), .Y(new_n8566));
  nor_5  g06218(.A(new_n8566), .B(new_n8539), .Y(new_n8567));
  nor_5  g06219(.A(new_n8567), .B(new_n8538), .Y(new_n8568));
  nor_5  g06220(.A(new_n8568), .B(new_n8534), .Y(new_n8569));
  nor_5  g06221(.A(new_n8569), .B(new_n8533), .Y(new_n8570));
  xnor_4 g06222(.A(new_n8570), .B(new_n8528), .Y(n904));
  not_8  g06223(.A(n19472), .Y(new_n8572));
  nor_5  g06224(.A(n18962), .B(n10158), .Y(new_n8573));
  not_8  g06225(.A(new_n8573), .Y(new_n8574));
  nor_5  g06226(.A(new_n8574), .B(n8052), .Y(new_n8575));
  not_8  g06227(.A(new_n8575), .Y(new_n8576));
  nor_5  g06228(.A(new_n8576), .B(n15539), .Y(new_n8577));
  xnor_4 g06229(.A(new_n8577), .B(n19228), .Y(new_n8578));
  xnor_4 g06230(.A(new_n8578), .B(n21471), .Y(new_n8579));
  xnor_4 g06231(.A(new_n8575), .B(n15539), .Y(new_n8580));
  and_5  g06232(.A(new_n8580), .B(n18737), .Y(new_n8581_1));
  xnor_4 g06233(.A(new_n8580), .B(n18737), .Y(new_n8582));
  xnor_4 g06234(.A(new_n8573), .B(n8052), .Y(new_n8583));
  not_8  g06235(.A(new_n8583), .Y(new_n8584));
  nor_5  g06236(.A(new_n8584), .B(new_n3301_1), .Y(new_n8585));
  xnor_4 g06237(.A(new_n8584), .B(n14603), .Y(new_n8586));
  xnor_4 g06238(.A(n18962), .B(n10158), .Y(new_n8587));
  not_8  g06239(.A(new_n8587), .Y(new_n8588));
  nor_5  g06240(.A(new_n8588), .B(n20794), .Y(new_n8589));
  nor_5  g06241(.A(new_n3305), .B(new_n6771), .Y(new_n8590));
  xnor_4 g06242(.A(new_n8587), .B(n20794), .Y(new_n8591));
  not_8  g06243(.A(new_n8591), .Y(new_n8592));
  nor_5  g06244(.A(new_n8592), .B(new_n8590), .Y(new_n8593));
  nor_5  g06245(.A(new_n8593), .B(new_n8589), .Y(new_n8594_1));
  and_5  g06246(.A(new_n8594_1), .B(new_n8586), .Y(new_n8595));
  nor_5  g06247(.A(new_n8595), .B(new_n8585), .Y(new_n8596));
  nor_5  g06248(.A(new_n8596), .B(new_n8582), .Y(new_n8597));
  nor_5  g06249(.A(new_n8597), .B(new_n8581_1), .Y(new_n8598));
  xnor_4 g06250(.A(new_n8598), .B(new_n8579), .Y(new_n8599));
  not_8  g06251(.A(new_n8599), .Y(new_n8600));
  xnor_4 g06252(.A(new_n8600), .B(new_n8572), .Y(new_n8601));
  xnor_4 g06253(.A(new_n8596), .B(new_n8582), .Y(new_n8602));
  not_8  g06254(.A(new_n8602), .Y(new_n8603));
  nor_5  g06255(.A(new_n8603), .B(n25370), .Y(new_n8604));
  not_8  g06256(.A(n24786), .Y(new_n8605));
  xnor_4 g06257(.A(new_n8594_1), .B(new_n8586), .Y(new_n8606));
  nor_5  g06258(.A(new_n8606), .B(new_n8605), .Y(new_n8607));
  not_8  g06259(.A(new_n8606), .Y(new_n8608_1));
  xnor_4 g06260(.A(new_n8608_1), .B(new_n8605), .Y(new_n8609));
  xnor_4 g06261(.A(n23333), .B(n18962), .Y(new_n8610));
  nor_5  g06262(.A(new_n8610), .B(new_n4109), .Y(new_n8611));
  and_5  g06263(.A(new_n8611), .B(new_n8591), .Y(new_n8612));
  xnor_4 g06264(.A(new_n8592), .B(new_n8590), .Y(new_n8613));
  nor_5  g06265(.A(new_n8613), .B(new_n8611), .Y(new_n8614_1));
  nor_5  g06266(.A(new_n8614_1), .B(new_n8612), .Y(new_n8615));
  and_5  g06267(.A(new_n8615), .B(n27120), .Y(new_n8616));
  or_5   g06268(.A(new_n8616), .B(new_n8612), .Y(new_n8617));
  and_5  g06269(.A(new_n8617), .B(new_n8609), .Y(new_n8618));
  nor_5  g06270(.A(new_n8618), .B(new_n8607), .Y(new_n8619));
  xnor_4 g06271(.A(new_n8603), .B(new_n6846), .Y(new_n8620_1));
  and_5  g06272(.A(new_n8620_1), .B(new_n8619), .Y(new_n8621));
  nor_5  g06273(.A(new_n8621), .B(new_n8604), .Y(new_n8622));
  xor_4  g06274(.A(new_n8622), .B(new_n8601), .Y(new_n8623));
  xnor_4 g06275(.A(new_n8623), .B(new_n6696), .Y(new_n8624));
  xnor_4 g06276(.A(new_n8620_1), .B(new_n8619), .Y(new_n8625));
  nor_5  g06277(.A(new_n8625), .B(new_n6699), .Y(new_n8626));
  xnor_4 g06278(.A(new_n8625), .B(new_n6699), .Y(new_n8627));
  not_8  g06279(.A(n27120), .Y(new_n8628));
  xnor_4 g06280(.A(new_n8615), .B(new_n8628), .Y(new_n8629));
  nor_5  g06281(.A(new_n8629), .B(new_n6731), .Y(new_n8630));
  xnor_4 g06282(.A(new_n8610), .B(n23065), .Y(new_n8631));
  not_8  g06283(.A(new_n8631), .Y(new_n8632));
  nor_5  g06284(.A(new_n8632), .B(new_n6702), .Y(new_n8633));
  xnor_4 g06285(.A(new_n8629), .B(new_n6731), .Y(new_n8634));
  nor_5  g06286(.A(new_n8634), .B(new_n8633), .Y(new_n8635));
  nor_5  g06287(.A(new_n8635), .B(new_n8630), .Y(new_n8636));
  nor_5  g06288(.A(new_n8636), .B(new_n6715), .Y(new_n8637_1));
  xor_4  g06289(.A(new_n8617), .B(new_n8609), .Y(new_n8638_1));
  xnor_4 g06290(.A(new_n8636), .B(new_n6715), .Y(new_n8639));
  nor_5  g06291(.A(new_n8639), .B(new_n8638_1), .Y(new_n8640));
  nor_5  g06292(.A(new_n8640), .B(new_n8637_1), .Y(new_n8641));
  nor_5  g06293(.A(new_n8641), .B(new_n8627), .Y(new_n8642));
  nor_5  g06294(.A(new_n8642), .B(new_n8626), .Y(new_n8643));
  xnor_4 g06295(.A(new_n8643), .B(new_n8624), .Y(n948));
  xnor_4 g06296(.A(n25972), .B(n10250), .Y(new_n8645));
  not_8  g06297(.A(n21915), .Y(new_n8646));
  nor_5  g06298(.A(new_n8646), .B(n7674), .Y(new_n8647));
  xnor_4 g06299(.A(n21915), .B(n7674), .Y(new_n8648));
  nor_5  g06300(.A(new_n6836), .B(n6397), .Y(new_n8649));
  xnor_4 g06301(.A(n13775), .B(n6397), .Y(new_n8650));
  nor_5  g06302(.A(n19196), .B(new_n6839), .Y(new_n8651));
  xnor_4 g06303(.A(n19196), .B(n1293), .Y(new_n8652));
  nor_5  g06304(.A(n23586), .B(new_n6842), .Y(new_n8653));
  xnor_4 g06305(.A(n23586), .B(n19042), .Y(new_n8654));
  nor_5  g06306(.A(n21226), .B(new_n8572), .Y(new_n8655));
  xnor_4 g06307(.A(n21226), .B(n19472), .Y(new_n8656_1));
  nor_5  g06308(.A(new_n6846), .B(n4426), .Y(new_n8657));
  xnor_4 g06309(.A(n25370), .B(n4426), .Y(new_n8658));
  not_8  g06310(.A(n20036), .Y(new_n8659));
  nor_5  g06311(.A(n24786), .B(new_n8659), .Y(new_n8660));
  nor_5  g06312(.A(new_n8605), .B(n20036), .Y(new_n8661));
  nor_5  g06313(.A(n27120), .B(new_n4120), .Y(new_n8662_1));
  or_5   g06314(.A(new_n8628), .B(n11192), .Y(new_n8663));
  nor_5  g06315(.A(n23065), .B(new_n6176), .Y(new_n8664));
  and_5  g06316(.A(new_n8664), .B(new_n8663), .Y(new_n8665));
  nor_5  g06317(.A(new_n8665), .B(new_n8662_1), .Y(new_n8666));
  nor_5  g06318(.A(new_n8666), .B(new_n8661), .Y(new_n8667));
  nor_5  g06319(.A(new_n8667), .B(new_n8660), .Y(new_n8668));
  and_5  g06320(.A(new_n8668), .B(new_n8658), .Y(new_n8669));
  or_5   g06321(.A(new_n8669), .B(new_n8657), .Y(new_n8670));
  and_5  g06322(.A(new_n8670), .B(new_n8656_1), .Y(new_n8671));
  or_5   g06323(.A(new_n8671), .B(new_n8655), .Y(new_n8672));
  and_5  g06324(.A(new_n8672), .B(new_n8654), .Y(new_n8673));
  or_5   g06325(.A(new_n8673), .B(new_n8653), .Y(new_n8674));
  and_5  g06326(.A(new_n8674), .B(new_n8652), .Y(new_n8675));
  or_5   g06327(.A(new_n8675), .B(new_n8651), .Y(new_n8676));
  and_5  g06328(.A(new_n8676), .B(new_n8650), .Y(new_n8677));
  or_5   g06329(.A(new_n8677), .B(new_n8649), .Y(new_n8678_1));
  and_5  g06330(.A(new_n8678_1), .B(new_n8648), .Y(new_n8679));
  or_5   g06331(.A(new_n8679), .B(new_n8647), .Y(new_n8680));
  xor_4  g06332(.A(new_n8680), .B(new_n8645), .Y(new_n8681));
  xnor_4 g06333(.A(n20040), .B(n2978), .Y(new_n8682));
  nor_5  g06334(.A(new_n6744), .B(n19531), .Y(new_n8683));
  xnor_4 g06335(.A(n23697), .B(n19531), .Y(new_n8684));
  nor_5  g06336(.A(n18345), .B(new_n6748), .Y(new_n8685));
  xnor_4 g06337(.A(n18345), .B(n2289), .Y(new_n8686));
  nor_5  g06338(.A(n13190), .B(new_n6752), .Y(new_n8687_1));
  xnor_4 g06339(.A(n13190), .B(n1112), .Y(new_n8688));
  nor_5  g06340(.A(new_n6756), .B(n3460), .Y(new_n8689));
  xnor_4 g06341(.A(n20179), .B(n3460), .Y(new_n8690));
  nor_5  g06342(.A(new_n7440), .B(n5226), .Y(new_n8691));
  xnor_4 g06343(.A(n19228), .B(n5226), .Y(new_n8692));
  nor_5  g06344(.A(n17664), .B(new_n6763), .Y(new_n8693));
  xnor_4 g06345(.A(n17664), .B(n15539), .Y(new_n8694_1));
  nor_5  g06346(.A(new_n2578_1), .B(n8052), .Y(new_n8695));
  nor_5  g06347(.A(n23369), .B(new_n6767), .Y(new_n8696));
  not_8  g06348(.A(n1136), .Y(new_n8697));
  nor_5  g06349(.A(n10158), .B(new_n8697), .Y(new_n8698));
  nor_5  g06350(.A(new_n7448), .B(n1136), .Y(new_n8699));
  nor_5  g06351(.A(new_n2582_1), .B(n18962), .Y(new_n8700));
  not_8  g06352(.A(new_n8700), .Y(new_n8701));
  nor_5  g06353(.A(new_n8701), .B(new_n8699), .Y(new_n8702));
  nor_5  g06354(.A(new_n8702), .B(new_n8698), .Y(new_n8703));
  nor_5  g06355(.A(new_n8703), .B(new_n8696), .Y(new_n8704));
  nor_5  g06356(.A(new_n8704), .B(new_n8695), .Y(new_n8705));
  and_5  g06357(.A(new_n8705), .B(new_n8694_1), .Y(new_n8706));
  or_5   g06358(.A(new_n8706), .B(new_n8693), .Y(new_n8707));
  and_5  g06359(.A(new_n8707), .B(new_n8692), .Y(new_n8708));
  or_5   g06360(.A(new_n8708), .B(new_n8691), .Y(new_n8709));
  and_5  g06361(.A(new_n8709), .B(new_n8690), .Y(new_n8710));
  or_5   g06362(.A(new_n8710), .B(new_n8689), .Y(new_n8711));
  and_5  g06363(.A(new_n8711), .B(new_n8688), .Y(new_n8712));
  or_5   g06364(.A(new_n8712), .B(new_n8687_1), .Y(new_n8713));
  and_5  g06365(.A(new_n8713), .B(new_n8686), .Y(new_n8714));
  or_5   g06366(.A(new_n8714), .B(new_n8685), .Y(new_n8715));
  and_5  g06367(.A(new_n8715), .B(new_n8684), .Y(new_n8716_1));
  nor_5  g06368(.A(new_n8716_1), .B(new_n8683), .Y(new_n8717));
  xnor_4 g06369(.A(new_n8717), .B(new_n8682), .Y(new_n8718));
  not_8  g06370(.A(n12507), .Y(new_n8719));
  nor_5  g06371(.A(n15258), .B(n4588), .Y(new_n8720));
  not_8  g06372(.A(new_n8720), .Y(new_n8721_1));
  nor_5  g06373(.A(new_n8721_1), .B(n16743), .Y(new_n8722));
  not_8  g06374(.A(new_n8722), .Y(new_n8723));
  nor_5  g06375(.A(new_n8723), .B(n22631), .Y(new_n8724));
  not_8  g06376(.A(new_n8724), .Y(new_n8725));
  nor_5  g06377(.A(new_n8725), .B(n2331), .Y(new_n8726));
  not_8  g06378(.A(new_n8726), .Y(new_n8727));
  nor_5  g06379(.A(new_n8727), .B(n25068), .Y(new_n8728));
  not_8  g06380(.A(new_n8728), .Y(new_n8729));
  nor_5  g06381(.A(new_n8729), .B(n16812), .Y(new_n8730));
  not_8  g06382(.A(new_n8730), .Y(new_n8731));
  nor_5  g06383(.A(new_n8731), .B(n7841), .Y(new_n8732));
  not_8  g06384(.A(new_n8732), .Y(new_n8733));
  nor_5  g06385(.A(new_n8733), .B(n26264), .Y(new_n8734));
  xnor_4 g06386(.A(new_n8734), .B(n22764), .Y(new_n8735));
  xnor_4 g06387(.A(new_n8735), .B(new_n8719), .Y(new_n8736));
  xnor_4 g06388(.A(new_n8732), .B(n26264), .Y(new_n8737));
  and_5  g06389(.A(new_n8737), .B(n15077), .Y(new_n8738));
  nor_5  g06390(.A(new_n8737), .B(n15077), .Y(new_n8739));
  xnor_4 g06391(.A(new_n8730), .B(n7841), .Y(new_n8740));
  and_5  g06392(.A(new_n8740), .B(n3710), .Y(new_n8741));
  or_5   g06393(.A(new_n8740), .B(n3710), .Y(new_n8742));
  xnor_4 g06394(.A(new_n8728), .B(n16812), .Y(new_n8743));
  nor_5  g06395(.A(new_n8743), .B(n26318), .Y(new_n8744_1));
  not_8  g06396(.A(n26318), .Y(new_n8745_1));
  xnor_4 g06397(.A(new_n8743), .B(new_n8745_1), .Y(new_n8746));
  xnor_4 g06398(.A(new_n8726), .B(n25068), .Y(new_n8747));
  nor_5  g06399(.A(new_n8747), .B(n26054), .Y(new_n8748));
  not_8  g06400(.A(n26054), .Y(new_n8749));
  xnor_4 g06401(.A(new_n8747), .B(new_n8749), .Y(new_n8750));
  xnor_4 g06402(.A(new_n8724), .B(n2331), .Y(new_n8751));
  nor_5  g06403(.A(new_n8751), .B(n19081), .Y(new_n8752));
  not_8  g06404(.A(n19081), .Y(new_n8753));
  xnor_4 g06405(.A(new_n8751), .B(new_n8753), .Y(new_n8754));
  xnor_4 g06406(.A(new_n8722), .B(n22631), .Y(new_n8755));
  nor_5  g06407(.A(new_n8755), .B(n8309), .Y(new_n8756));
  xnor_4 g06408(.A(new_n8720), .B(n16743), .Y(new_n8757));
  nor_5  g06409(.A(new_n8757), .B(n19144), .Y(new_n8758));
  not_8  g06410(.A(n19144), .Y(new_n8759));
  xnor_4 g06411(.A(new_n8757), .B(new_n8759), .Y(new_n8760));
  xnor_4 g06412(.A(n15258), .B(new_n2542), .Y(new_n8761));
  nor_5  g06413(.A(new_n8761), .B(n12593), .Y(new_n8762));
  not_8  g06414(.A(n13714), .Y(new_n8763));
  or_5   g06415(.A(new_n8763), .B(new_n2542), .Y(new_n8764));
  not_8  g06416(.A(new_n8761), .Y(new_n8765));
  xnor_4 g06417(.A(new_n8765), .B(n12593), .Y(new_n8766));
  and_5  g06418(.A(new_n8766), .B(new_n8764), .Y(new_n8767));
  or_5   g06419(.A(new_n8767), .B(new_n8762), .Y(new_n8768));
  and_5  g06420(.A(new_n8768), .B(new_n8760), .Y(new_n8769));
  or_5   g06421(.A(new_n8769), .B(new_n8758), .Y(new_n8770));
  not_8  g06422(.A(n8309), .Y(new_n8771));
  xnor_4 g06423(.A(new_n8755), .B(new_n8771), .Y(new_n8772));
  and_5  g06424(.A(new_n8772), .B(new_n8770), .Y(new_n8773));
  or_5   g06425(.A(new_n8773), .B(new_n8756), .Y(new_n8774));
  and_5  g06426(.A(new_n8774), .B(new_n8754), .Y(new_n8775));
  or_5   g06427(.A(new_n8775), .B(new_n8752), .Y(new_n8776));
  and_5  g06428(.A(new_n8776), .B(new_n8750), .Y(new_n8777));
  or_5   g06429(.A(new_n8777), .B(new_n8748), .Y(new_n8778));
  and_5  g06430(.A(new_n8778), .B(new_n8746), .Y(new_n8779));
  nor_5  g06431(.A(new_n8779), .B(new_n8744_1), .Y(new_n8780));
  and_5  g06432(.A(new_n8780), .B(new_n8742), .Y(new_n8781));
  nor_5  g06433(.A(new_n8781), .B(new_n8741), .Y(new_n8782_1));
  nor_5  g06434(.A(new_n8782_1), .B(new_n8739), .Y(new_n8783));
  nor_5  g06435(.A(new_n8783), .B(new_n8738), .Y(new_n8784));
  xnor_4 g06436(.A(new_n8784), .B(new_n8736), .Y(new_n8785));
  xnor_4 g06437(.A(new_n8785), .B(new_n8718), .Y(new_n8786));
  nor_5  g06438(.A(new_n8714), .B(new_n8685), .Y(new_n8787));
  xnor_4 g06439(.A(new_n8787), .B(new_n8684), .Y(new_n8788));
  not_8  g06440(.A(n15077), .Y(new_n8789));
  xnor_4 g06441(.A(new_n8737), .B(new_n8789), .Y(new_n8790));
  xnor_4 g06442(.A(new_n8790), .B(new_n8782_1), .Y(new_n8791));
  and_5  g06443(.A(new_n8791), .B(new_n8788), .Y(new_n8792));
  not_8  g06444(.A(new_n8788), .Y(new_n8793));
  xnor_4 g06445(.A(new_n8791), .B(new_n8793), .Y(new_n8794));
  xor_4  g06446(.A(new_n8713), .B(new_n8686), .Y(new_n8795));
  xnor_4 g06447(.A(new_n8740), .B(n3710), .Y(new_n8796));
  xnor_4 g06448(.A(new_n8796), .B(new_n8780), .Y(new_n8797));
  nor_5  g06449(.A(new_n8797), .B(new_n8795), .Y(new_n8798));
  xnor_4 g06450(.A(new_n8797), .B(new_n8795), .Y(new_n8799));
  nor_5  g06451(.A(new_n8710), .B(new_n8689), .Y(new_n8800));
  xnor_4 g06452(.A(new_n8800), .B(new_n8688), .Y(new_n8801));
  not_8  g06453(.A(new_n8801), .Y(new_n8802));
  xor_4  g06454(.A(new_n8778), .B(new_n8746), .Y(new_n8803_1));
  and_5  g06455(.A(new_n8803_1), .B(new_n8802), .Y(new_n8804));
  xnor_4 g06456(.A(new_n8803_1), .B(new_n8802), .Y(new_n8805));
  nor_5  g06457(.A(new_n8708), .B(new_n8691), .Y(new_n8806_1));
  xnor_4 g06458(.A(new_n8806_1), .B(new_n8690), .Y(new_n8807));
  not_8  g06459(.A(new_n8807), .Y(new_n8808));
  xor_4  g06460(.A(new_n8776), .B(new_n8750), .Y(new_n8809_1));
  and_5  g06461(.A(new_n8809_1), .B(new_n8808), .Y(new_n8810));
  xnor_4 g06462(.A(new_n8809_1), .B(new_n8808), .Y(new_n8811));
  nor_5  g06463(.A(new_n8706), .B(new_n8693), .Y(new_n8812));
  xnor_4 g06464(.A(new_n8812), .B(new_n8692), .Y(new_n8813));
  not_8  g06465(.A(new_n8813), .Y(new_n8814));
  xor_4  g06466(.A(new_n8774), .B(new_n8754), .Y(new_n8815));
  and_5  g06467(.A(new_n8815), .B(new_n8814), .Y(new_n8816));
  xnor_4 g06468(.A(new_n8815), .B(new_n8814), .Y(new_n8817));
  xnor_4 g06469(.A(new_n8705), .B(new_n8694_1), .Y(new_n8818));
  xor_4  g06470(.A(new_n8772), .B(new_n8770), .Y(new_n8819));
  and_5  g06471(.A(new_n8819), .B(new_n8818), .Y(new_n8820));
  not_8  g06472(.A(new_n8818), .Y(new_n8821_1));
  xnor_4 g06473(.A(new_n8819), .B(new_n8821_1), .Y(new_n8822));
  xor_4  g06474(.A(new_n8768), .B(new_n8760), .Y(new_n8823));
  xnor_4 g06475(.A(n23369), .B(n8052), .Y(new_n8824_1));
  xnor_4 g06476(.A(new_n8824_1), .B(new_n8703), .Y(new_n8825));
  nor_5  g06477(.A(new_n8825), .B(new_n8823), .Y(new_n8826));
  xnor_4 g06478(.A(new_n8825), .B(new_n8823), .Y(new_n8827_1));
  xor_4  g06479(.A(new_n8766), .B(new_n8764), .Y(new_n8828));
  xnor_4 g06480(.A(n10158), .B(n1136), .Y(new_n8829));
  xnor_4 g06481(.A(new_n8829), .B(new_n8701), .Y(new_n8830));
  nor_5  g06482(.A(new_n8830), .B(new_n8828), .Y(new_n8831));
  xnor_4 g06483(.A(n19234), .B(n18962), .Y(new_n8832));
  xnor_4 g06484(.A(n13714), .B(n4588), .Y(new_n8833));
  nor_5  g06485(.A(new_n8833), .B(new_n8832), .Y(new_n8834));
  not_8  g06486(.A(new_n8830), .Y(new_n8835));
  xnor_4 g06487(.A(new_n8835), .B(new_n8828), .Y(new_n8836));
  and_5  g06488(.A(new_n8836), .B(new_n8834), .Y(new_n8837));
  nor_5  g06489(.A(new_n8837), .B(new_n8831), .Y(new_n8838));
  nor_5  g06490(.A(new_n8838), .B(new_n8827_1), .Y(new_n8839));
  nor_5  g06491(.A(new_n8839), .B(new_n8826), .Y(new_n8840));
  and_5  g06492(.A(new_n8840), .B(new_n8822), .Y(new_n8841));
  nor_5  g06493(.A(new_n8841), .B(new_n8820), .Y(new_n8842));
  nor_5  g06494(.A(new_n8842), .B(new_n8817), .Y(new_n8843));
  nor_5  g06495(.A(new_n8843), .B(new_n8816), .Y(new_n8844));
  nor_5  g06496(.A(new_n8844), .B(new_n8811), .Y(new_n8845));
  nor_5  g06497(.A(new_n8845), .B(new_n8810), .Y(new_n8846));
  nor_5  g06498(.A(new_n8846), .B(new_n8805), .Y(new_n8847));
  nor_5  g06499(.A(new_n8847), .B(new_n8804), .Y(new_n8848));
  nor_5  g06500(.A(new_n8848), .B(new_n8799), .Y(new_n8849_1));
  nor_5  g06501(.A(new_n8849_1), .B(new_n8798), .Y(new_n8850));
  and_5  g06502(.A(new_n8850), .B(new_n8794), .Y(new_n8851));
  nor_5  g06503(.A(new_n8851), .B(new_n8792), .Y(new_n8852));
  xnor_4 g06504(.A(new_n8852), .B(new_n8786), .Y(new_n8853));
  xnor_4 g06505(.A(new_n8853), .B(new_n8681), .Y(new_n8854));
  xor_4  g06506(.A(new_n8678_1), .B(new_n8648), .Y(new_n8855));
  xor_4  g06507(.A(new_n8850), .B(new_n8794), .Y(new_n8856_1));
  nor_5  g06508(.A(new_n8856_1), .B(new_n8855), .Y(new_n8857));
  xnor_4 g06509(.A(new_n8856_1), .B(new_n8855), .Y(new_n8858));
  xor_4  g06510(.A(new_n8676), .B(new_n8650), .Y(new_n8859));
  xnor_4 g06511(.A(new_n8848), .B(new_n8799), .Y(new_n8860));
  nor_5  g06512(.A(new_n8860), .B(new_n8859), .Y(new_n8861_1));
  xnor_4 g06513(.A(new_n8860), .B(new_n8859), .Y(new_n8862_1));
  xor_4  g06514(.A(new_n8674), .B(new_n8652), .Y(new_n8863));
  xnor_4 g06515(.A(new_n8846), .B(new_n8805), .Y(new_n8864));
  nor_5  g06516(.A(new_n8864), .B(new_n8863), .Y(new_n8865));
  xnor_4 g06517(.A(new_n8864), .B(new_n8863), .Y(new_n8866));
  xor_4  g06518(.A(new_n8672), .B(new_n8654), .Y(new_n8867));
  xnor_4 g06519(.A(new_n8844), .B(new_n8811), .Y(new_n8868));
  nor_5  g06520(.A(new_n8868), .B(new_n8867), .Y(new_n8869_1));
  xnor_4 g06521(.A(new_n8868), .B(new_n8867), .Y(new_n8870));
  xor_4  g06522(.A(new_n8670), .B(new_n8656_1), .Y(new_n8871));
  xnor_4 g06523(.A(new_n8842), .B(new_n8817), .Y(new_n8872));
  nor_5  g06524(.A(new_n8872), .B(new_n8871), .Y(new_n8873));
  xnor_4 g06525(.A(new_n8872), .B(new_n8871), .Y(new_n8874));
  xnor_4 g06526(.A(new_n8840), .B(new_n8822), .Y(new_n8875));
  not_8  g06527(.A(new_n8875), .Y(new_n8876));
  xnor_4 g06528(.A(new_n8668), .B(new_n8658), .Y(new_n8877));
  and_5  g06529(.A(new_n8877), .B(new_n8876), .Y(new_n8878));
  xnor_4 g06530(.A(new_n8877), .B(new_n8876), .Y(new_n8879));
  xnor_4 g06531(.A(new_n8838), .B(new_n8827_1), .Y(new_n8880));
  xnor_4 g06532(.A(n24786), .B(n20036), .Y(new_n8881));
  xnor_4 g06533(.A(new_n8881), .B(new_n8666), .Y(new_n8882));
  and_5  g06534(.A(new_n8882), .B(new_n8880), .Y(new_n8883));
  xnor_4 g06535(.A(new_n8882), .B(new_n8880), .Y(new_n8884_1));
  xnor_4 g06536(.A(n23065), .B(n9380), .Y(new_n8885));
  xnor_4 g06537(.A(new_n8833), .B(new_n8832), .Y(new_n8886));
  nor_5  g06538(.A(new_n8886), .B(new_n8885), .Y(new_n8887));
  xnor_4 g06539(.A(n27120), .B(n11192), .Y(new_n8888));
  xnor_4 g06540(.A(new_n8888), .B(new_n8664), .Y(new_n8889));
  nor_5  g06541(.A(new_n8889), .B(new_n8887), .Y(new_n8890));
  xnor_4 g06542(.A(new_n8836), .B(new_n8834), .Y(new_n8891));
  not_8  g06543(.A(new_n8891), .Y(new_n8892));
  xnor_4 g06544(.A(new_n8889), .B(new_n8887), .Y(new_n8893));
  nor_5  g06545(.A(new_n8893), .B(new_n8892), .Y(new_n8894));
  nor_5  g06546(.A(new_n8894), .B(new_n8890), .Y(new_n8895));
  nor_5  g06547(.A(new_n8895), .B(new_n8884_1), .Y(new_n8896));
  nor_5  g06548(.A(new_n8896), .B(new_n8883), .Y(new_n8897));
  nor_5  g06549(.A(new_n8897), .B(new_n8879), .Y(new_n8898));
  nor_5  g06550(.A(new_n8898), .B(new_n8878), .Y(new_n8899));
  nor_5  g06551(.A(new_n8899), .B(new_n8874), .Y(new_n8900));
  nor_5  g06552(.A(new_n8900), .B(new_n8873), .Y(new_n8901));
  nor_5  g06553(.A(new_n8901), .B(new_n8870), .Y(new_n8902));
  nor_5  g06554(.A(new_n8902), .B(new_n8869_1), .Y(new_n8903));
  nor_5  g06555(.A(new_n8903), .B(new_n8866), .Y(new_n8904));
  nor_5  g06556(.A(new_n8904), .B(new_n8865), .Y(new_n8905));
  nor_5  g06557(.A(new_n8905), .B(new_n8862_1), .Y(new_n8906));
  nor_5  g06558(.A(new_n8906), .B(new_n8861_1), .Y(new_n8907));
  nor_5  g06559(.A(new_n8907), .B(new_n8858), .Y(new_n8908));
  nor_5  g06560(.A(new_n8908), .B(new_n8857), .Y(new_n8909_1));
  xor_4  g06561(.A(new_n8909_1), .B(new_n8854), .Y(n957));
  xnor_4 g06562(.A(new_n8832), .B(n20385), .Y(new_n8911_1));
  xnor_4 g06563(.A(n26167), .B(new_n4122), .Y(new_n8912));
  xnor_4 g06564(.A(new_n8912), .B(n21138), .Y(new_n8913));
  xnor_4 g06565(.A(new_n8913), .B(new_n8911_1), .Y(n980));
  nor_5  g06566(.A(new_n7702), .B(new_n4357), .Y(new_n8915));
  xnor_4 g06567(.A(new_n7698_1), .B(new_n4357), .Y(new_n8916));
  nor_5  g06568(.A(new_n7705), .B(new_n4359), .Y(new_n8917));
  xnor_4 g06569(.A(new_n7705), .B(new_n4359), .Y(new_n8918));
  nor_5  g06570(.A(new_n7710), .B(new_n4363), .Y(new_n8919));
  xnor_4 g06571(.A(new_n7710), .B(new_n4363), .Y(new_n8920_1));
  nor_5  g06572(.A(new_n7717), .B(new_n4367), .Y(new_n8921));
  xnor_4 g06573(.A(new_n7717), .B(new_n4367), .Y(new_n8922));
  nor_5  g06574(.A(new_n7721_1), .B(new_n4371), .Y(new_n8923));
  xnor_4 g06575(.A(new_n7721_1), .B(new_n4371), .Y(new_n8924));
  nor_5  g06576(.A(new_n7725), .B(new_n4375), .Y(new_n8925));
  xnor_4 g06577(.A(new_n7725), .B(new_n4375), .Y(new_n8926));
  nor_5  g06578(.A(new_n7730), .B(new_n4380), .Y(new_n8927));
  xnor_4 g06579(.A(new_n7730), .B(new_n4380), .Y(new_n8928));
  nor_5  g06580(.A(new_n7739), .B(new_n4388), .Y(new_n8929));
  xnor_4 g06581(.A(new_n7735), .B(new_n4388), .Y(new_n8930));
  nor_5  g06582(.A(new_n7742), .B(new_n4391), .Y(new_n8931));
  nor_5  g06583(.A(new_n7748), .B(new_n4395), .Y(new_n8932));
  xnor_4 g06584(.A(new_n7742), .B(new_n4392), .Y(new_n8933));
  and_5  g06585(.A(new_n8933), .B(new_n8932), .Y(new_n8934));
  nor_5  g06586(.A(new_n8934), .B(new_n8931), .Y(new_n8935));
  and_5  g06587(.A(new_n8935), .B(new_n8930), .Y(new_n8936));
  nor_5  g06588(.A(new_n8936), .B(new_n8929), .Y(new_n8937));
  nor_5  g06589(.A(new_n8937), .B(new_n8928), .Y(new_n8938));
  nor_5  g06590(.A(new_n8938), .B(new_n8927), .Y(new_n8939));
  nor_5  g06591(.A(new_n8939), .B(new_n8926), .Y(new_n8940));
  nor_5  g06592(.A(new_n8940), .B(new_n8925), .Y(new_n8941));
  nor_5  g06593(.A(new_n8941), .B(new_n8924), .Y(new_n8942));
  nor_5  g06594(.A(new_n8942), .B(new_n8923), .Y(new_n8943_1));
  nor_5  g06595(.A(new_n8943_1), .B(new_n8922), .Y(new_n8944));
  nor_5  g06596(.A(new_n8944), .B(new_n8921), .Y(new_n8945));
  nor_5  g06597(.A(new_n8945), .B(new_n8920_1), .Y(new_n8946));
  nor_5  g06598(.A(new_n8946), .B(new_n8919), .Y(new_n8947));
  nor_5  g06599(.A(new_n8947), .B(new_n8918), .Y(new_n8948));
  nor_5  g06600(.A(new_n8948), .B(new_n8917), .Y(new_n8949));
  and_5  g06601(.A(new_n8949), .B(new_n8916), .Y(new_n8950));
  or_5   g06602(.A(new_n8950), .B(new_n8915), .Y(new_n8951));
  xnor_4 g06603(.A(new_n7695), .B(new_n4353), .Y(new_n8952));
  xor_4  g06604(.A(new_n8952), .B(new_n8951), .Y(new_n8953));
  not_8  g06605(.A(n16544), .Y(new_n8954));
  nor_5  g06606(.A(new_n8954), .B(n12650), .Y(new_n8955));
  xnor_4 g06607(.A(n16544), .B(n12650), .Y(new_n8956));
  nor_5  g06608(.A(n10201), .B(new_n2887_1), .Y(new_n8957));
  xnor_4 g06609(.A(n10201), .B(n6814), .Y(new_n8958));
  not_8  g06610(.A(n19701), .Y(new_n8959));
  nor_5  g06611(.A(new_n8959), .B(n10593), .Y(new_n8960));
  xnor_4 g06612(.A(n19701), .B(n10593), .Y(new_n8961));
  not_8  g06613(.A(n23529), .Y(new_n8962));
  nor_5  g06614(.A(new_n8962), .B(n18290), .Y(new_n8963));
  xnor_4 g06615(.A(n23529), .B(n18290), .Y(new_n8964_1));
  not_8  g06616(.A(n24620), .Y(new_n8965));
  nor_5  g06617(.A(new_n8965), .B(n11580), .Y(new_n8966));
  xnor_4 g06618(.A(n24620), .B(n11580), .Y(new_n8967));
  not_8  g06619(.A(n5211), .Y(new_n8968));
  nor_5  g06620(.A(n15884), .B(new_n8968), .Y(new_n8969));
  xnor_4 g06621(.A(n15884), .B(n5211), .Y(new_n8970));
  not_8  g06622(.A(n12956), .Y(new_n8971_1));
  nor_5  g06623(.A(new_n8971_1), .B(n6356), .Y(new_n8972));
  xnor_4 g06624(.A(n12956), .B(n6356), .Y(new_n8973));
  nor_5  g06625(.A(new_n5582), .B(n18295), .Y(new_n8974));
  nor_5  g06626(.A(n27104), .B(new_n2903), .Y(new_n8975));
  nor_5  g06627(.A(new_n5584), .B(n6502), .Y(new_n8976));
  or_5   g06628(.A(n27188), .B(new_n5033), .Y(new_n8977));
  nor_5  g06629(.A(n15780), .B(new_n5588), .Y(new_n8978));
  and_5  g06630(.A(new_n8978), .B(new_n8977), .Y(new_n8979));
  nor_5  g06631(.A(new_n8979), .B(new_n8976), .Y(new_n8980));
  nor_5  g06632(.A(new_n8980), .B(new_n8975), .Y(new_n8981));
  nor_5  g06633(.A(new_n8981), .B(new_n8974), .Y(new_n8982_1));
  and_5  g06634(.A(new_n8982_1), .B(new_n8973), .Y(new_n8983));
  or_5   g06635(.A(new_n8983), .B(new_n8972), .Y(new_n8984));
  and_5  g06636(.A(new_n8984), .B(new_n8970), .Y(new_n8985));
  or_5   g06637(.A(new_n8985), .B(new_n8969), .Y(new_n8986));
  and_5  g06638(.A(new_n8986), .B(new_n8967), .Y(new_n8987));
  or_5   g06639(.A(new_n8987), .B(new_n8966), .Y(new_n8988));
  and_5  g06640(.A(new_n8988), .B(new_n8964_1), .Y(new_n8989));
  or_5   g06641(.A(new_n8989), .B(new_n8963), .Y(new_n8990));
  and_5  g06642(.A(new_n8990), .B(new_n8961), .Y(new_n8991));
  or_5   g06643(.A(new_n8991), .B(new_n8960), .Y(new_n8992));
  and_5  g06644(.A(new_n8992), .B(new_n8958), .Y(new_n8993_1));
  or_5   g06645(.A(new_n8993_1), .B(new_n8957), .Y(new_n8994));
  and_5  g06646(.A(new_n8994), .B(new_n8956), .Y(new_n8995));
  nor_5  g06647(.A(new_n8995), .B(new_n8955), .Y(new_n8996));
  xnor_4 g06648(.A(new_n8996), .B(new_n8953), .Y(new_n8997));
  xor_4  g06649(.A(new_n8994), .B(new_n8956), .Y(new_n8998));
  xor_4  g06650(.A(new_n8949), .B(new_n8916), .Y(new_n8999));
  nor_5  g06651(.A(new_n8999), .B(new_n8998), .Y(new_n9000));
  xnor_4 g06652(.A(new_n8999), .B(new_n8998), .Y(new_n9001));
  xor_4  g06653(.A(new_n8992), .B(new_n8958), .Y(new_n9002));
  xnor_4 g06654(.A(new_n8947), .B(new_n8918), .Y(new_n9003_1));
  nor_5  g06655(.A(new_n9003_1), .B(new_n9002), .Y(new_n9004));
  xnor_4 g06656(.A(new_n9003_1), .B(new_n9002), .Y(new_n9005));
  xor_4  g06657(.A(new_n8990), .B(new_n8961), .Y(new_n9006));
  xnor_4 g06658(.A(new_n8945), .B(new_n8920_1), .Y(new_n9007));
  nor_5  g06659(.A(new_n9007), .B(new_n9006), .Y(new_n9008));
  xnor_4 g06660(.A(new_n9007), .B(new_n9006), .Y(new_n9009));
  xor_4  g06661(.A(new_n8988), .B(new_n8964_1), .Y(new_n9010));
  xnor_4 g06662(.A(new_n8943_1), .B(new_n8922), .Y(new_n9011));
  nor_5  g06663(.A(new_n9011), .B(new_n9010), .Y(new_n9012_1));
  xnor_4 g06664(.A(new_n9011), .B(new_n9010), .Y(new_n9013));
  xor_4  g06665(.A(new_n8986), .B(new_n8967), .Y(new_n9014));
  xnor_4 g06666(.A(new_n8941), .B(new_n8924), .Y(new_n9015));
  nor_5  g06667(.A(new_n9015), .B(new_n9014), .Y(new_n9016));
  xnor_4 g06668(.A(new_n9015), .B(new_n9014), .Y(new_n9017));
  xor_4  g06669(.A(new_n8984), .B(new_n8970), .Y(new_n9018));
  xnor_4 g06670(.A(new_n8939), .B(new_n8926), .Y(new_n9019));
  nor_5  g06671(.A(new_n9019), .B(new_n9018), .Y(new_n9020));
  xnor_4 g06672(.A(new_n9019), .B(new_n9018), .Y(new_n9021));
  xnor_4 g06673(.A(new_n8937), .B(new_n8928), .Y(new_n9022));
  not_8  g06674(.A(new_n9022), .Y(new_n9023));
  xnor_4 g06675(.A(new_n8982_1), .B(new_n8973), .Y(new_n9024));
  and_5  g06676(.A(new_n9024), .B(new_n9023), .Y(new_n9025));
  xnor_4 g06677(.A(new_n8935), .B(new_n8930), .Y(new_n9026));
  not_8  g06678(.A(new_n9026), .Y(new_n9027));
  xnor_4 g06679(.A(n27104), .B(n18295), .Y(new_n9028));
  xnor_4 g06680(.A(new_n9028), .B(new_n8980), .Y(new_n9029));
  and_5  g06681(.A(new_n9029), .B(new_n9027), .Y(new_n9030));
  xnor_4 g06682(.A(new_n9029), .B(new_n9027), .Y(new_n9031));
  xnor_4 g06683(.A(n15780), .B(n6611), .Y(new_n9032_1));
  xnor_4 g06684(.A(new_n7888), .B(new_n4395), .Y(new_n9033));
  not_8  g06685(.A(new_n9033), .Y(new_n9034));
  nor_5  g06686(.A(new_n9034), .B(new_n9032_1), .Y(new_n9035));
  xnor_4 g06687(.A(n27188), .B(n6502), .Y(new_n9036));
  xnor_4 g06688(.A(new_n9036), .B(new_n8978), .Y(new_n9037));
  nor_5  g06689(.A(new_n9037), .B(new_n9035), .Y(new_n9038));
  xor_4  g06690(.A(new_n8933), .B(new_n8932), .Y(new_n9039));
  xnor_4 g06691(.A(new_n9037), .B(new_n9035), .Y(new_n9040));
  nor_5  g06692(.A(new_n9040), .B(new_n9039), .Y(new_n9041));
  nor_5  g06693(.A(new_n9041), .B(new_n9038), .Y(new_n9042_1));
  nor_5  g06694(.A(new_n9042_1), .B(new_n9031), .Y(new_n9043));
  nor_5  g06695(.A(new_n9043), .B(new_n9030), .Y(new_n9044));
  xnor_4 g06696(.A(new_n9024), .B(new_n9023), .Y(new_n9045));
  nor_5  g06697(.A(new_n9045), .B(new_n9044), .Y(new_n9046_1));
  nor_5  g06698(.A(new_n9046_1), .B(new_n9025), .Y(new_n9047_1));
  nor_5  g06699(.A(new_n9047_1), .B(new_n9021), .Y(new_n9048));
  nor_5  g06700(.A(new_n9048), .B(new_n9020), .Y(new_n9049));
  nor_5  g06701(.A(new_n9049), .B(new_n9017), .Y(new_n9050));
  nor_5  g06702(.A(new_n9050), .B(new_n9016), .Y(new_n9051));
  nor_5  g06703(.A(new_n9051), .B(new_n9013), .Y(new_n9052));
  nor_5  g06704(.A(new_n9052), .B(new_n9012_1), .Y(new_n9053));
  nor_5  g06705(.A(new_n9053), .B(new_n9009), .Y(new_n9054));
  nor_5  g06706(.A(new_n9054), .B(new_n9008), .Y(new_n9055));
  nor_5  g06707(.A(new_n9055), .B(new_n9005), .Y(new_n9056));
  nor_5  g06708(.A(new_n9056), .B(new_n9004), .Y(new_n9057));
  nor_5  g06709(.A(new_n9057), .B(new_n9001), .Y(new_n9058));
  nor_5  g06710(.A(new_n9058), .B(new_n9000), .Y(new_n9059));
  xnor_4 g06711(.A(new_n9059), .B(new_n8997), .Y(n982));
  not_8  g06712(.A(new_n4544), .Y(new_n9061));
  not_8  g06713(.A(n3279), .Y(new_n9062));
  nor_5  g06714(.A(n26808), .B(n7339), .Y(new_n9063));
  not_8  g06715(.A(new_n9063), .Y(new_n9064));
  nor_5  g06716(.A(new_n9064), .B(n1667), .Y(new_n9065));
  not_8  g06717(.A(new_n9065), .Y(new_n9066));
  nor_5  g06718(.A(new_n9066), .B(n2680), .Y(new_n9067));
  not_8  g06719(.A(new_n9067), .Y(new_n9068));
  nor_5  g06720(.A(new_n9068), .B(n2547), .Y(new_n9069));
  not_8  g06721(.A(new_n9069), .Y(new_n9070));
  nor_5  g06722(.A(new_n9070), .B(n2999), .Y(new_n9071));
  not_8  g06723(.A(new_n9071), .Y(new_n9072));
  nor_5  g06724(.A(new_n9072), .B(n14702), .Y(new_n9073));
  not_8  g06725(.A(new_n9073), .Y(new_n9074));
  nor_5  g06726(.A(new_n9074), .B(n13914), .Y(new_n9075));
  and_5  g06727(.A(new_n9075), .B(new_n9062), .Y(new_n9076));
  xnor_4 g06728(.A(new_n9076), .B(n4306), .Y(new_n9077));
  xnor_4 g06729(.A(n23166), .B(n18105), .Y(new_n9078));
  not_8  g06730(.A(n10577), .Y(new_n9079));
  nor_5  g06731(.A(n24196), .B(new_n9079), .Y(new_n9080));
  xnor_4 g06732(.A(n24196), .B(n10577), .Y(new_n9081));
  not_8  g06733(.A(n6381), .Y(new_n9082));
  nor_5  g06734(.A(n16376), .B(new_n9082), .Y(new_n9083));
  xnor_4 g06735(.A(n16376), .B(n6381), .Y(new_n9084));
  not_8  g06736(.A(n14345), .Y(new_n9085));
  nor_5  g06737(.A(n25381), .B(new_n9085), .Y(new_n9086));
  xnor_4 g06738(.A(n25381), .B(n14345), .Y(new_n9087));
  not_8  g06739(.A(n11356), .Y(new_n9088));
  nor_5  g06740(.A(n12587), .B(new_n9088), .Y(new_n9089));
  xnor_4 g06741(.A(n12587), .B(n11356), .Y(new_n9090_1));
  not_8  g06742(.A(n3164), .Y(new_n9091));
  nor_5  g06743(.A(new_n9091), .B(n268), .Y(new_n9092));
  xnor_4 g06744(.A(n3164), .B(n268), .Y(new_n9093));
  nor_5  g06745(.A(n24879), .B(new_n6590_1), .Y(new_n9094));
  xnor_4 g06746(.A(n24879), .B(n10611), .Y(new_n9095));
  nor_5  g06747(.A(new_n8048), .B(n2783), .Y(new_n9096));
  nor_5  g06748(.A(n6785), .B(new_n6593), .Y(new_n9097));
  nor_5  g06749(.A(new_n8052_1), .B(n15490), .Y(new_n9098));
  not_8  g06750(.A(n15490), .Y(new_n9099));
  nor_5  g06751(.A(n24032), .B(new_n9099), .Y(new_n9100));
  nor_5  g06752(.A(new_n4507), .B(n18), .Y(new_n9101));
  not_8  g06753(.A(new_n9101), .Y(new_n9102));
  nor_5  g06754(.A(new_n9102), .B(new_n9100), .Y(new_n9103));
  nor_5  g06755(.A(new_n9103), .B(new_n9098), .Y(new_n9104_1));
  nor_5  g06756(.A(new_n9104_1), .B(new_n9097), .Y(new_n9105));
  nor_5  g06757(.A(new_n9105), .B(new_n9096), .Y(new_n9106));
  and_5  g06758(.A(new_n9106), .B(new_n9095), .Y(new_n9107));
  or_5   g06759(.A(new_n9107), .B(new_n9094), .Y(new_n9108));
  and_5  g06760(.A(new_n9108), .B(new_n9093), .Y(new_n9109));
  or_5   g06761(.A(new_n9109), .B(new_n9092), .Y(new_n9110));
  and_5  g06762(.A(new_n9110), .B(new_n9090_1), .Y(new_n9111));
  or_5   g06763(.A(new_n9111), .B(new_n9089), .Y(new_n9112));
  and_5  g06764(.A(new_n9112), .B(new_n9087), .Y(new_n9113));
  or_5   g06765(.A(new_n9113), .B(new_n9086), .Y(new_n9114));
  and_5  g06766(.A(new_n9114), .B(new_n9084), .Y(new_n9115));
  or_5   g06767(.A(new_n9115), .B(new_n9083), .Y(new_n9116));
  and_5  g06768(.A(new_n9116), .B(new_n9081), .Y(new_n9117));
  nor_5  g06769(.A(new_n9117), .B(new_n9080), .Y(new_n9118));
  xnor_4 g06770(.A(new_n9118), .B(new_n9078), .Y(new_n9119));
  xor_4  g06771(.A(new_n9119), .B(new_n9077), .Y(new_n9120));
  xnor_4 g06772(.A(new_n9075), .B(n3279), .Y(new_n9121));
  nor_5  g06773(.A(new_n9115), .B(new_n9083), .Y(new_n9122));
  xnor_4 g06774(.A(new_n9122), .B(new_n9081), .Y(new_n9123));
  and_5  g06775(.A(new_n9123), .B(new_n9121), .Y(new_n9124));
  xor_4  g06776(.A(new_n9123), .B(new_n9121), .Y(new_n9125));
  xnor_4 g06777(.A(new_n9073), .B(n13914), .Y(new_n9126));
  xor_4  g06778(.A(new_n9114), .B(new_n9084), .Y(new_n9127));
  nor_5  g06779(.A(new_n9127), .B(new_n9126), .Y(new_n9128));
  xnor_4 g06780(.A(new_n9127), .B(new_n9126), .Y(new_n9129_1));
  xnor_4 g06781(.A(new_n9071), .B(n14702), .Y(new_n9130));
  xor_4  g06782(.A(new_n9112), .B(new_n9087), .Y(new_n9131));
  nor_5  g06783(.A(new_n9131), .B(new_n9130), .Y(new_n9132));
  xnor_4 g06784(.A(new_n9131), .B(new_n9130), .Y(new_n9133));
  xnor_4 g06785(.A(new_n9069), .B(n2999), .Y(new_n9134));
  xor_4  g06786(.A(new_n9110), .B(new_n9090_1), .Y(new_n9135));
  nor_5  g06787(.A(new_n9135), .B(new_n9134), .Y(new_n9136));
  xnor_4 g06788(.A(new_n9067), .B(n2547), .Y(new_n9137));
  xor_4  g06789(.A(new_n9108), .B(new_n9093), .Y(new_n9138));
  nor_5  g06790(.A(new_n9138), .B(new_n9137), .Y(new_n9139));
  xnor_4 g06791(.A(new_n9138), .B(new_n9137), .Y(new_n9140));
  xnor_4 g06792(.A(new_n9065), .B(n2680), .Y(new_n9141));
  xnor_4 g06793(.A(new_n9106), .B(new_n9095), .Y(new_n9142));
  not_8  g06794(.A(new_n9142), .Y(new_n9143));
  nor_5  g06795(.A(new_n9143), .B(new_n9141), .Y(new_n9144));
  xnor_4 g06796(.A(new_n9063), .B(n1667), .Y(new_n9145));
  xnor_4 g06797(.A(n6785), .B(n2783), .Y(new_n9146_1));
  xnor_4 g06798(.A(new_n9146_1), .B(new_n9104_1), .Y(new_n9147));
  not_8  g06799(.A(new_n9147), .Y(new_n9148));
  nor_5  g06800(.A(new_n9148), .B(new_n9145), .Y(new_n9149));
  xnor_4 g06801(.A(new_n9147), .B(new_n9145), .Y(new_n9150));
  xnor_4 g06802(.A(n26808), .B(n7339), .Y(new_n9151));
  xnor_4 g06803(.A(n24032), .B(n15490), .Y(new_n9152));
  xnor_4 g06804(.A(new_n9152), .B(new_n9102), .Y(new_n9153));
  nor_5  g06805(.A(new_n9153), .B(new_n9151), .Y(new_n9154));
  not_8  g06806(.A(n26808), .Y(new_n9155));
  xnor_4 g06807(.A(n22843), .B(n18), .Y(new_n9156));
  nor_5  g06808(.A(new_n9156), .B(new_n9155), .Y(new_n9157));
  not_8  g06809(.A(new_n9153), .Y(new_n9158));
  xnor_4 g06810(.A(new_n9158), .B(new_n9151), .Y(new_n9159));
  and_5  g06811(.A(new_n9159), .B(new_n9157), .Y(new_n9160));
  nor_5  g06812(.A(new_n9160), .B(new_n9154), .Y(new_n9161));
  and_5  g06813(.A(new_n9161), .B(new_n9150), .Y(new_n9162));
  or_5   g06814(.A(new_n9162), .B(new_n9149), .Y(new_n9163));
  xnor_4 g06815(.A(new_n9142), .B(new_n9141), .Y(new_n9164_1));
  and_5  g06816(.A(new_n9164_1), .B(new_n9163), .Y(new_n9165));
  nor_5  g06817(.A(new_n9165), .B(new_n9144), .Y(new_n9166_1));
  nor_5  g06818(.A(new_n9166_1), .B(new_n9140), .Y(new_n9167));
  nor_5  g06819(.A(new_n9167), .B(new_n9139), .Y(new_n9168));
  xnor_4 g06820(.A(new_n9135), .B(new_n9134), .Y(new_n9169));
  nor_5  g06821(.A(new_n9169), .B(new_n9168), .Y(new_n9170));
  nor_5  g06822(.A(new_n9170), .B(new_n9136), .Y(new_n9171));
  nor_5  g06823(.A(new_n9171), .B(new_n9133), .Y(new_n9172_1));
  nor_5  g06824(.A(new_n9172_1), .B(new_n9132), .Y(new_n9173));
  nor_5  g06825(.A(new_n9173), .B(new_n9129_1), .Y(new_n9174));
  nor_5  g06826(.A(new_n9174), .B(new_n9128), .Y(new_n9175));
  and_5  g06827(.A(new_n9175), .B(new_n9125), .Y(new_n9176));
  or_5   g06828(.A(new_n9176), .B(new_n9124), .Y(new_n9177));
  xor_4  g06829(.A(new_n9177), .B(new_n9120), .Y(new_n9178));
  xnor_4 g06830(.A(new_n9178), .B(new_n9061), .Y(new_n9179));
  xor_4  g06831(.A(new_n9175), .B(new_n9125), .Y(new_n9180));
  nor_5  g06832(.A(new_n9180), .B(new_n4549), .Y(new_n9181));
  xnor_4 g06833(.A(new_n9180), .B(new_n4549), .Y(new_n9182_1));
  xnor_4 g06834(.A(new_n9173), .B(new_n9129_1), .Y(new_n9183));
  nor_5  g06835(.A(new_n9183), .B(new_n4554), .Y(new_n9184));
  xnor_4 g06836(.A(new_n9183), .B(new_n4554), .Y(new_n9185));
  xnor_4 g06837(.A(new_n9171), .B(new_n9133), .Y(new_n9186));
  nor_5  g06838(.A(new_n9186), .B(new_n4559), .Y(new_n9187));
  xnor_4 g06839(.A(new_n9186), .B(new_n4559), .Y(new_n9188));
  xnor_4 g06840(.A(new_n9169), .B(new_n9168), .Y(new_n9189));
  nor_5  g06841(.A(new_n9189), .B(new_n4564), .Y(new_n9190));
  xnor_4 g06842(.A(new_n9189), .B(new_n4564), .Y(new_n9191_1));
  xnor_4 g06843(.A(new_n9166_1), .B(new_n9140), .Y(new_n9192));
  nor_5  g06844(.A(new_n9192), .B(new_n4568), .Y(new_n9193));
  xnor_4 g06845(.A(new_n9192), .B(new_n4568), .Y(new_n9194));
  xor_4  g06846(.A(new_n9164_1), .B(new_n9163), .Y(new_n9195));
  and_5  g06847(.A(new_n9195), .B(new_n4575), .Y(new_n9196));
  xnor_4 g06848(.A(new_n9195), .B(new_n4573), .Y(new_n9197));
  xor_4  g06849(.A(new_n9161), .B(new_n9150), .Y(new_n9198));
  nor_5  g06850(.A(new_n9198), .B(new_n4579), .Y(new_n9199));
  xnor_4 g06851(.A(new_n9198), .B(new_n4591), .Y(new_n9200));
  xnor_4 g06852(.A(new_n9159), .B(new_n9157), .Y(new_n9201));
  nor_5  g06853(.A(new_n9201), .B(new_n4581), .Y(new_n9202));
  xnor_4 g06854(.A(new_n9156), .B(n26808), .Y(new_n9203));
  and_5  g06855(.A(new_n9203), .B(new_n4585), .Y(new_n9204));
  xor_4  g06856(.A(new_n9201), .B(new_n4581), .Y(new_n9205));
  and_5  g06857(.A(new_n9205), .B(new_n9204), .Y(new_n9206));
  or_5   g06858(.A(new_n9206), .B(new_n9202), .Y(new_n9207));
  and_5  g06859(.A(new_n9207), .B(new_n9200), .Y(new_n9208));
  nor_5  g06860(.A(new_n9208), .B(new_n9199), .Y(new_n9209));
  and_5  g06861(.A(new_n9209), .B(new_n9197), .Y(new_n9210));
  nor_5  g06862(.A(new_n9210), .B(new_n9196), .Y(new_n9211));
  nor_5  g06863(.A(new_n9211), .B(new_n9194), .Y(new_n9212));
  nor_5  g06864(.A(new_n9212), .B(new_n9193), .Y(new_n9213));
  nor_5  g06865(.A(new_n9213), .B(new_n9191_1), .Y(new_n9214));
  nor_5  g06866(.A(new_n9214), .B(new_n9190), .Y(new_n9215));
  nor_5  g06867(.A(new_n9215), .B(new_n9188), .Y(new_n9216));
  nor_5  g06868(.A(new_n9216), .B(new_n9187), .Y(new_n9217_1));
  nor_5  g06869(.A(new_n9217_1), .B(new_n9185), .Y(new_n9218));
  nor_5  g06870(.A(new_n9218), .B(new_n9184), .Y(new_n9219));
  nor_5  g06871(.A(new_n9219), .B(new_n9182_1), .Y(new_n9220_1));
  nor_5  g06872(.A(new_n9220_1), .B(new_n9181), .Y(new_n9221));
  xnor_4 g06873(.A(new_n9221), .B(new_n9179), .Y(n984));
  xnor_4 g06874(.A(new_n9215), .B(new_n9188), .Y(n1005));
  xnor_4 g06875(.A(new_n3387), .B(new_n3344), .Y(n1016));
  xnor_4 g06876(.A(new_n4100_1), .B(new_n4086), .Y(n1020));
  xnor_4 g06877(.A(n18290), .B(new_n2853_1), .Y(new_n9226));
  nor_5  g06878(.A(n11580), .B(n2035), .Y(new_n9227));
  xnor_4 g06879(.A(n11580), .B(n2035), .Y(new_n9228));
  nor_5  g06880(.A(n15884), .B(n5213), .Y(new_n9229));
  xnor_4 g06881(.A(n15884), .B(new_n2859), .Y(new_n9230));
  nor_5  g06882(.A(n6356), .B(n4665), .Y(new_n9231));
  xnor_4 g06883(.A(n6356), .B(new_n2862), .Y(new_n9232));
  nor_5  g06884(.A(n27104), .B(n19005), .Y(new_n9233));
  xnor_4 g06885(.A(n27104), .B(new_n2866), .Y(new_n9234));
  nor_5  g06886(.A(n27188), .B(n4326), .Y(new_n9235));
  or_5   g06887(.A(new_n5588), .B(new_n5287), .Y(new_n9236));
  xnor_4 g06888(.A(n27188), .B(new_n2869), .Y(new_n9237));
  and_5  g06889(.A(new_n9237), .B(new_n9236), .Y(new_n9238));
  or_5   g06890(.A(new_n9238), .B(new_n9235), .Y(new_n9239));
  and_5  g06891(.A(new_n9239), .B(new_n9234), .Y(new_n9240));
  or_5   g06892(.A(new_n9240), .B(new_n9233), .Y(new_n9241));
  and_5  g06893(.A(new_n9241), .B(new_n9232), .Y(new_n9242));
  or_5   g06894(.A(new_n9242), .B(new_n9231), .Y(new_n9243));
  and_5  g06895(.A(new_n9243), .B(new_n9230), .Y(new_n9244));
  nor_5  g06896(.A(new_n9244), .B(new_n9229), .Y(new_n9245));
  nor_5  g06897(.A(new_n9245), .B(new_n9228), .Y(new_n9246_1));
  or_5   g06898(.A(new_n9246_1), .B(new_n9227), .Y(new_n9247));
  xor_4  g06899(.A(new_n9247), .B(new_n9226), .Y(new_n9248));
  not_8  g06900(.A(new_n9248), .Y(new_n9249));
  xnor_4 g06901(.A(new_n9249), .B(new_n8962), .Y(new_n9250));
  xnor_4 g06902(.A(new_n9245), .B(new_n9228), .Y(new_n9251_1));
  nor_5  g06903(.A(new_n9251_1), .B(n24620), .Y(new_n9252));
  xnor_4 g06904(.A(new_n9251_1), .B(new_n8965), .Y(new_n9253));
  nor_5  g06905(.A(new_n9242), .B(new_n9231), .Y(new_n9254));
  xnor_4 g06906(.A(new_n9254), .B(new_n9230), .Y(new_n9255));
  not_8  g06907(.A(new_n9255), .Y(new_n9256));
  nor_5  g06908(.A(new_n9256), .B(n5211), .Y(new_n9257));
  xnor_4 g06909(.A(new_n9256), .B(new_n8968), .Y(new_n9258));
  nor_5  g06910(.A(new_n9240), .B(new_n9233), .Y(new_n9259_1));
  xnor_4 g06911(.A(new_n9259_1), .B(new_n9232), .Y(new_n9260));
  not_8  g06912(.A(new_n9260), .Y(new_n9261_1));
  nor_5  g06913(.A(new_n9261_1), .B(n12956), .Y(new_n9262));
  xnor_4 g06914(.A(new_n9261_1), .B(new_n8971_1), .Y(new_n9263));
  nor_5  g06915(.A(new_n9238), .B(new_n9235), .Y(new_n9264));
  xnor_4 g06916(.A(new_n9264), .B(new_n9234), .Y(new_n9265));
  not_8  g06917(.A(new_n9265), .Y(new_n9266));
  nor_5  g06918(.A(new_n9266), .B(n18295), .Y(new_n9267));
  nor_5  g06919(.A(new_n5588), .B(new_n5287), .Y(new_n9268));
  xnor_4 g06920(.A(new_n9237), .B(new_n9268), .Y(new_n9269));
  nor_5  g06921(.A(new_n9269), .B(new_n5033), .Y(new_n9270));
  xnor_4 g06922(.A(n6611), .B(new_n5287), .Y(new_n9271));
  not_8  g06923(.A(new_n9271), .Y(new_n9272));
  nor_5  g06924(.A(new_n9272), .B(new_n2907), .Y(new_n9273));
  not_8  g06925(.A(new_n9269), .Y(new_n9274));
  xnor_4 g06926(.A(new_n9274), .B(new_n5033), .Y(new_n9275));
  and_5  g06927(.A(new_n9275), .B(new_n9273), .Y(new_n9276));
  nor_5  g06928(.A(new_n9276), .B(new_n9270), .Y(new_n9277));
  xnor_4 g06929(.A(new_n9266), .B(new_n2903), .Y(new_n9278));
  and_5  g06930(.A(new_n9278), .B(new_n9277), .Y(new_n9279));
  or_5   g06931(.A(new_n9279), .B(new_n9267), .Y(new_n9280));
  and_5  g06932(.A(new_n9280), .B(new_n9263), .Y(new_n9281));
  or_5   g06933(.A(new_n9281), .B(new_n9262), .Y(new_n9282));
  and_5  g06934(.A(new_n9282), .B(new_n9258), .Y(new_n9283));
  or_5   g06935(.A(new_n9283), .B(new_n9257), .Y(new_n9284));
  and_5  g06936(.A(new_n9284), .B(new_n9253), .Y(new_n9285));
  or_5   g06937(.A(new_n9285), .B(new_n9252), .Y(new_n9286));
  xor_4  g06938(.A(new_n9286), .B(new_n9250), .Y(new_n9287_1));
  xnor_4 g06939(.A(n17250), .B(new_n6037), .Y(new_n9288));
  nor_5  g06940(.A(n23160), .B(n3570), .Y(new_n9289));
  xnor_4 g06941(.A(n23160), .B(new_n6043), .Y(new_n9290));
  nor_5  g06942(.A(n16524), .B(n13668), .Y(new_n9291));
  xnor_4 g06943(.A(n16524), .B(new_n6049), .Y(new_n9292));
  nor_5  g06944(.A(n21276), .B(n11056), .Y(new_n9293));
  not_8  g06945(.A(n11056), .Y(new_n9294));
  xnor_4 g06946(.A(n21276), .B(new_n9294), .Y(new_n9295));
  nor_5  g06947(.A(n26748), .B(n15271), .Y(new_n9296));
  xnor_4 g06948(.A(n26748), .B(new_n7668), .Y(new_n9297));
  nor_5  g06949(.A(n25877), .B(n10057), .Y(new_n9298));
  nor_5  g06950(.A(new_n6629), .B(new_n4242), .Y(new_n9299));
  xnor_4 g06951(.A(n25877), .B(n10057), .Y(new_n9300));
  nor_5  g06952(.A(new_n9300), .B(new_n9299), .Y(new_n9301));
  or_5   g06953(.A(new_n9301), .B(new_n9298), .Y(new_n9302));
  and_5  g06954(.A(new_n9302), .B(new_n9297), .Y(new_n9303));
  or_5   g06955(.A(new_n9303), .B(new_n9296), .Y(new_n9304));
  and_5  g06956(.A(new_n9304), .B(new_n9295), .Y(new_n9305));
  or_5   g06957(.A(new_n9305), .B(new_n9293), .Y(new_n9306));
  and_5  g06958(.A(new_n9306), .B(new_n9292), .Y(new_n9307));
  or_5   g06959(.A(new_n9307), .B(new_n9291), .Y(new_n9308_1));
  and_5  g06960(.A(new_n9308_1), .B(new_n9290), .Y(new_n9309));
  nor_5  g06961(.A(new_n9309), .B(new_n9289), .Y(new_n9310));
  xnor_4 g06962(.A(new_n9310), .B(new_n9288), .Y(new_n9311));
  not_8  g06963(.A(new_n9311), .Y(new_n9312));
  xnor_4 g06964(.A(new_n9312), .B(n11044), .Y(new_n9313));
  nor_5  g06965(.A(new_n9307), .B(new_n9291), .Y(new_n9314));
  xnor_4 g06966(.A(new_n9314), .B(new_n9290), .Y(new_n9315));
  nor_5  g06967(.A(new_n9315), .B(new_n5994), .Y(new_n9316));
  not_8  g06968(.A(new_n9315), .Y(new_n9317));
  xnor_4 g06969(.A(new_n9317), .B(n2421), .Y(new_n9318_1));
  nor_5  g06970(.A(new_n9305), .B(new_n9293), .Y(new_n9319));
  xnor_4 g06971(.A(new_n9319), .B(new_n9292), .Y(new_n9320));
  nor_5  g06972(.A(new_n9320), .B(new_n7662), .Y(new_n9321));
  not_8  g06973(.A(new_n9320), .Y(new_n9322));
  xnor_4 g06974(.A(new_n9322), .B(n987), .Y(new_n9323_1));
  nor_5  g06975(.A(new_n9303), .B(new_n9296), .Y(new_n9324));
  xnor_4 g06976(.A(new_n9324), .B(new_n9295), .Y(new_n9325));
  nor_5  g06977(.A(new_n9325), .B(new_n7665), .Y(new_n9326));
  not_8  g06978(.A(new_n9325), .Y(new_n9327));
  xnor_4 g06979(.A(new_n9327), .B(n20478), .Y(new_n9328));
  nor_5  g06980(.A(new_n9301), .B(new_n9298), .Y(new_n9329));
  xnor_4 g06981(.A(new_n9329), .B(new_n9297), .Y(new_n9330));
  nor_5  g06982(.A(new_n9330), .B(new_n7670_1), .Y(new_n9331));
  xnor_4 g06983(.A(new_n9300), .B(new_n9299), .Y(new_n9332));
  nor_5  g06984(.A(new_n9332), .B(n22619), .Y(new_n9333));
  xnor_4 g06985(.A(n24323), .B(new_n4242), .Y(new_n9334));
  not_8  g06986(.A(new_n9334), .Y(new_n9335));
  nor_5  g06987(.A(new_n9335), .B(new_n6003), .Y(new_n9336));
  xnor_4 g06988(.A(new_n9332), .B(n22619), .Y(new_n9337));
  nor_5  g06989(.A(new_n9337), .B(new_n9336), .Y(new_n9338));
  or_5   g06990(.A(new_n9338), .B(new_n9333), .Y(new_n9339));
  not_8  g06991(.A(new_n9330), .Y(new_n9340));
  xnor_4 g06992(.A(new_n9340), .B(n26882), .Y(new_n9341));
  nor_5  g06993(.A(new_n9341), .B(new_n9339), .Y(new_n9342));
  nor_5  g06994(.A(new_n9342), .B(new_n9331), .Y(new_n9343));
  nor_5  g06995(.A(new_n9343), .B(new_n9328), .Y(new_n9344_1));
  nor_5  g06996(.A(new_n9344_1), .B(new_n9326), .Y(new_n9345));
  nor_5  g06997(.A(new_n9345), .B(new_n9323_1), .Y(new_n9346));
  nor_5  g06998(.A(new_n9346), .B(new_n9321), .Y(new_n9347));
  nor_5  g06999(.A(new_n9347), .B(new_n9318_1), .Y(new_n9348));
  nor_5  g07000(.A(new_n9348), .B(new_n9316), .Y(new_n9349));
  xnor_4 g07001(.A(new_n9349), .B(new_n9313), .Y(new_n9350));
  not_8  g07002(.A(new_n9350), .Y(new_n9351));
  xnor_4 g07003(.A(new_n9351), .B(new_n9287_1), .Y(new_n9352));
  xor_4  g07004(.A(new_n9284), .B(new_n9253), .Y(new_n9353));
  xnor_4 g07005(.A(new_n9347), .B(new_n9318_1), .Y(new_n9354));
  not_8  g07006(.A(new_n9354), .Y(new_n9355));
  and_5  g07007(.A(new_n9355), .B(new_n9353), .Y(new_n9356));
  xnor_4 g07008(.A(new_n9355), .B(new_n9353), .Y(new_n9357));
  xor_4  g07009(.A(new_n9282), .B(new_n9258), .Y(new_n9358));
  xnor_4 g07010(.A(new_n9345), .B(new_n9323_1), .Y(new_n9359));
  not_8  g07011(.A(new_n9359), .Y(new_n9360));
  and_5  g07012(.A(new_n9360), .B(new_n9358), .Y(new_n9361));
  xnor_4 g07013(.A(new_n9360), .B(new_n9358), .Y(new_n9362));
  xor_4  g07014(.A(new_n9280), .B(new_n9263), .Y(new_n9363));
  xnor_4 g07015(.A(new_n9343), .B(new_n9328), .Y(new_n9364_1));
  not_8  g07016(.A(new_n9364_1), .Y(new_n9365));
  and_5  g07017(.A(new_n9365), .B(new_n9363), .Y(new_n9366));
  xnor_4 g07018(.A(new_n9365), .B(new_n9363), .Y(new_n9367));
  xnor_4 g07019(.A(new_n9278), .B(new_n9277), .Y(new_n9368));
  not_8  g07020(.A(new_n9368), .Y(new_n9369));
  xor_4  g07021(.A(new_n9341), .B(new_n9339), .Y(new_n9370));
  and_5  g07022(.A(new_n9370), .B(new_n9369), .Y(new_n9371_1));
  xnor_4 g07023(.A(new_n9370), .B(new_n9369), .Y(new_n9372_1));
  xor_4  g07024(.A(new_n9337), .B(new_n9336), .Y(new_n9373));
  xor_4  g07025(.A(new_n9275), .B(new_n9273), .Y(new_n9374));
  nor_5  g07026(.A(new_n9374), .B(new_n9373), .Y(new_n9375));
  xnor_4 g07027(.A(new_n9335), .B(n6775), .Y(new_n9376));
  not_8  g07028(.A(new_n9376), .Y(new_n9377));
  xnor_4 g07029(.A(new_n9272), .B(n15780), .Y(new_n9378));
  nor_5  g07030(.A(new_n9378), .B(new_n9377), .Y(new_n9379));
  not_8  g07031(.A(new_n9373), .Y(new_n9380_1));
  xnor_4 g07032(.A(new_n9374), .B(new_n9380_1), .Y(new_n9381));
  and_5  g07033(.A(new_n9381), .B(new_n9379), .Y(new_n9382_1));
  nor_5  g07034(.A(new_n9382_1), .B(new_n9375), .Y(new_n9383));
  nor_5  g07035(.A(new_n9383), .B(new_n9372_1), .Y(new_n9384));
  nor_5  g07036(.A(new_n9384), .B(new_n9371_1), .Y(new_n9385));
  nor_5  g07037(.A(new_n9385), .B(new_n9367), .Y(new_n9386));
  nor_5  g07038(.A(new_n9386), .B(new_n9366), .Y(new_n9387));
  nor_5  g07039(.A(new_n9387), .B(new_n9362), .Y(new_n9388));
  nor_5  g07040(.A(new_n9388), .B(new_n9361), .Y(new_n9389));
  nor_5  g07041(.A(new_n9389), .B(new_n9357), .Y(new_n9390));
  nor_5  g07042(.A(new_n9390), .B(new_n9356), .Y(new_n9391));
  xnor_4 g07043(.A(new_n9391), .B(new_n9352), .Y(n1044));
  nor_5  g07044(.A(n22619), .B(n6775), .Y(new_n9393));
  not_8  g07045(.A(new_n9393), .Y(new_n9394));
  nor_5  g07046(.A(new_n9394), .B(n26882), .Y(new_n9395));
  xnor_4 g07047(.A(new_n9395), .B(n20478), .Y(new_n9396_1));
  xnor_4 g07048(.A(new_n9396_1), .B(new_n4932), .Y(new_n9397));
  xnor_4 g07049(.A(new_n9393), .B(n26882), .Y(new_n9398));
  and_5  g07050(.A(new_n9398), .B(n25872), .Y(new_n9399_1));
  xnor_4 g07051(.A(new_n9398), .B(new_n8483), .Y(new_n9400));
  xnor_4 g07052(.A(n22619), .B(n6775), .Y(new_n9401));
  nor_5  g07053(.A(new_n9401), .B(new_n4939_1), .Y(new_n9402));
  nor_5  g07054(.A(new_n6003), .B(new_n5002), .Y(new_n9403_1));
  xnor_4 g07055(.A(new_n9401), .B(n20259), .Y(new_n9404));
  and_5  g07056(.A(new_n9404), .B(new_n9403_1), .Y(new_n9405));
  or_5   g07057(.A(new_n9405), .B(new_n9402), .Y(new_n9406));
  and_5  g07058(.A(new_n9406), .B(new_n9400), .Y(new_n9407));
  nor_5  g07059(.A(new_n9407), .B(new_n9399_1), .Y(new_n9408));
  xnor_4 g07060(.A(new_n9408), .B(new_n9397), .Y(new_n9409));
  nor_5  g07061(.A(n9399), .B(n2088), .Y(new_n9410));
  not_8  g07062(.A(new_n9410), .Y(new_n9411));
  nor_5  g07063(.A(new_n9411), .B(n16396), .Y(new_n9412));
  xnor_4 g07064(.A(new_n9412), .B(n25074), .Y(new_n9413));
  xnor_4 g07065(.A(new_n9413), .B(new_n2398), .Y(new_n9414));
  xnor_4 g07066(.A(new_n9410), .B(n16396), .Y(new_n9415));
  and_5  g07067(.A(new_n9415), .B(n16722), .Y(new_n9416));
  xnor_4 g07068(.A(new_n9415), .B(new_n7625), .Y(new_n9417));
  not_8  g07069(.A(new_n5781), .Y(new_n9418));
  and_5  g07070(.A(new_n5787), .B(new_n9418), .Y(new_n9419_1));
  nor_5  g07071(.A(new_n9419_1), .B(new_n5783), .Y(new_n9420));
  and_5  g07072(.A(new_n9420), .B(new_n9417), .Y(new_n9421));
  nor_5  g07073(.A(new_n9421), .B(new_n9416), .Y(new_n9422));
  xnor_4 g07074(.A(new_n9422), .B(new_n9414), .Y(new_n9423_1));
  xnor_4 g07075(.A(new_n9423_1), .B(new_n9409), .Y(new_n9424));
  xnor_4 g07076(.A(new_n9420), .B(new_n9417), .Y(new_n9425));
  nor_5  g07077(.A(new_n9405), .B(new_n9402), .Y(new_n9426));
  xnor_4 g07078(.A(new_n9426), .B(new_n9400), .Y(new_n9427));
  not_8  g07079(.A(new_n9427), .Y(new_n9428));
  nor_5  g07080(.A(new_n9428), .B(new_n9425), .Y(new_n9429));
  xnor_4 g07081(.A(new_n9428), .B(new_n9425), .Y(new_n9430_1));
  xnor_4 g07082(.A(new_n9404), .B(new_n9403_1), .Y(new_n9431));
  nor_5  g07083(.A(new_n9431), .B(new_n5788), .Y(new_n9432));
  xnor_4 g07084(.A(n6775), .B(new_n5002), .Y(new_n9433));
  not_8  g07085(.A(new_n9433), .Y(new_n9434));
  nor_5  g07086(.A(new_n9434), .B(new_n5775), .Y(new_n9435_1));
  xnor_4 g07087(.A(new_n9431), .B(new_n5789), .Y(new_n9436));
  and_5  g07088(.A(new_n9436), .B(new_n9435_1), .Y(new_n9437));
  nor_5  g07089(.A(new_n9437), .B(new_n9432), .Y(new_n9438));
  nor_5  g07090(.A(new_n9438), .B(new_n9430_1), .Y(new_n9439));
  nor_5  g07091(.A(new_n9439), .B(new_n9429), .Y(new_n9440));
  xor_4  g07092(.A(new_n9440), .B(new_n9424), .Y(new_n9441));
  xnor_4 g07093(.A(n12956), .B(n7057), .Y(new_n9442));
  nor_5  g07094(.A(new_n2903), .B(n8381), .Y(new_n9443));
  nor_5  g07095(.A(n18295), .B(new_n8510_1), .Y(new_n9444));
  nor_5  g07096(.A(n20235), .B(new_n5033), .Y(new_n9445_1));
  or_5   g07097(.A(new_n5040), .B(n6502), .Y(new_n9446));
  nor_5  g07098(.A(new_n2907), .B(n12495), .Y(new_n9447));
  and_5  g07099(.A(new_n9447), .B(new_n9446), .Y(new_n9448));
  nor_5  g07100(.A(new_n9448), .B(new_n9445_1), .Y(new_n9449));
  nor_5  g07101(.A(new_n9449), .B(new_n9444), .Y(new_n9450));
  or_5   g07102(.A(new_n9450), .B(new_n9443), .Y(new_n9451_1));
  xnor_4 g07103(.A(new_n9451_1), .B(new_n9442), .Y(new_n9452));
  xor_4  g07104(.A(new_n9452), .B(new_n9441), .Y(new_n9453));
  xor_4  g07105(.A(new_n9438), .B(new_n9430_1), .Y(new_n9454));
  not_8  g07106(.A(new_n9454), .Y(new_n9455));
  xnor_4 g07107(.A(n18295), .B(n8381), .Y(new_n9456));
  xnor_4 g07108(.A(new_n9456), .B(new_n9449), .Y(new_n9457));
  and_5  g07109(.A(new_n9457), .B(new_n9455), .Y(new_n9458_1));
  xnor_4 g07110(.A(new_n9457), .B(new_n9455), .Y(new_n9459_1));
  xnor_4 g07111(.A(n15780), .B(n12495), .Y(new_n9460_1));
  xnor_4 g07112(.A(new_n9433), .B(new_n5775), .Y(new_n9461));
  not_8  g07113(.A(new_n9461), .Y(new_n9462));
  nor_5  g07114(.A(new_n9462), .B(new_n9460_1), .Y(new_n9463));
  xnor_4 g07115(.A(n20235), .B(n6502), .Y(new_n9464));
  xnor_4 g07116(.A(new_n9464), .B(new_n9447), .Y(new_n9465));
  nor_5  g07117(.A(new_n9465), .B(new_n9463), .Y(new_n9466));
  xnor_4 g07118(.A(new_n9436), .B(new_n9435_1), .Y(new_n9467));
  not_8  g07119(.A(new_n9467), .Y(new_n9468));
  xnor_4 g07120(.A(new_n9465), .B(new_n9463), .Y(new_n9469));
  nor_5  g07121(.A(new_n9469), .B(new_n9468), .Y(new_n9470));
  nor_5  g07122(.A(new_n9470), .B(new_n9466), .Y(new_n9471));
  nor_5  g07123(.A(new_n9471), .B(new_n9459_1), .Y(new_n9472));
  nor_5  g07124(.A(new_n9472), .B(new_n9458_1), .Y(new_n9473));
  xor_4  g07125(.A(new_n9473), .B(new_n9453), .Y(n1060));
  xnor_4 g07126(.A(new_n3385), .B(new_n3348), .Y(n1069));
  not_8  g07127(.A(n3959), .Y(new_n9476));
  xnor_4 g07128(.A(n9832), .B(new_n9476), .Y(new_n9477));
  nor_5  g07129(.A(n11566), .B(n1558), .Y(new_n9478));
  not_8  g07130(.A(n1558), .Y(new_n9479));
  xnor_4 g07131(.A(n11566), .B(new_n9479), .Y(new_n9480));
  nor_5  g07132(.A(n26744), .B(n21749), .Y(new_n9481));
  xnor_4 g07133(.A(n26744), .B(n21749), .Y(new_n9482));
  nor_5  g07134(.A(n26625), .B(n7769), .Y(new_n9483));
  not_8  g07135(.A(n14230), .Y(new_n9484));
  not_8  g07136(.A(n21138), .Y(new_n9485));
  or_5   g07137(.A(new_n9485), .B(new_n9484), .Y(new_n9486));
  not_8  g07138(.A(n7769), .Y(new_n9487));
  xnor_4 g07139(.A(n26625), .B(new_n9487), .Y(new_n9488));
  and_5  g07140(.A(new_n9488), .B(new_n9486), .Y(new_n9489));
  nor_5  g07141(.A(new_n9489), .B(new_n9483), .Y(new_n9490));
  nor_5  g07142(.A(new_n9490), .B(new_n9482), .Y(new_n9491));
  or_5   g07143(.A(new_n9491), .B(new_n9481), .Y(new_n9492));
  and_5  g07144(.A(new_n9492), .B(new_n9480), .Y(new_n9493_1));
  nor_5  g07145(.A(new_n9493_1), .B(new_n9478), .Y(new_n9494));
  xnor_4 g07146(.A(new_n9494), .B(new_n9477), .Y(new_n9495));
  nor_5  g07147(.A(n26167), .B(n22591), .Y(new_n9496));
  not_8  g07148(.A(new_n9496), .Y(new_n9497));
  nor_5  g07149(.A(new_n9497), .B(n17095), .Y(new_n9498));
  not_8  g07150(.A(new_n9498), .Y(new_n9499));
  nor_5  g07151(.A(new_n9499), .B(n15378), .Y(new_n9500));
  xnor_4 g07152(.A(new_n9500), .B(n19575), .Y(new_n9501));
  not_8  g07153(.A(n5226), .Y(new_n9502));
  xnor_4 g07154(.A(new_n6802_1), .B(new_n9502), .Y(new_n9503));
  nor_5  g07155(.A(new_n6806), .B(new_n2574), .Y(new_n9504));
  xnor_4 g07156(.A(new_n6806), .B(new_n2574), .Y(new_n9505));
  nor_5  g07157(.A(new_n6809), .B(new_n2578_1), .Y(new_n9506));
  xnor_4 g07158(.A(new_n6809), .B(new_n2578_1), .Y(new_n9507_1));
  nor_5  g07159(.A(new_n6942), .B(n1136), .Y(new_n9508_1));
  nor_5  g07160(.A(new_n6812), .B(new_n2582_1), .Y(new_n9509));
  xnor_4 g07161(.A(new_n6942), .B(n1136), .Y(new_n9510));
  nor_5  g07162(.A(new_n9510), .B(new_n9509), .Y(new_n9511));
  or_5   g07163(.A(new_n9511), .B(new_n9508_1), .Y(new_n9512_1));
  nor_5  g07164(.A(new_n9512_1), .B(new_n9507_1), .Y(new_n9513));
  nor_5  g07165(.A(new_n9513), .B(new_n9506), .Y(new_n9514));
  nor_5  g07166(.A(new_n9514), .B(new_n9505), .Y(new_n9515));
  nor_5  g07167(.A(new_n9515), .B(new_n9504), .Y(new_n9516));
  xor_4  g07168(.A(new_n9516), .B(new_n9503), .Y(new_n9517));
  not_8  g07169(.A(new_n9517), .Y(new_n9518));
  xnor_4 g07170(.A(new_n9518), .B(new_n9501), .Y(new_n9519));
  xor_4  g07171(.A(new_n9514), .B(new_n9505), .Y(new_n9520));
  xnor_4 g07172(.A(new_n9498), .B(n15378), .Y(new_n9521));
  nor_5  g07173(.A(new_n9521), .B(new_n9520), .Y(new_n9522));
  xnor_4 g07174(.A(new_n9521), .B(new_n9520), .Y(new_n9523));
  nor_5  g07175(.A(new_n9511), .B(new_n9508_1), .Y(new_n9524));
  xnor_4 g07176(.A(new_n9524), .B(new_n9507_1), .Y(new_n9525));
  xnor_4 g07177(.A(new_n9496), .B(n17095), .Y(new_n9526));
  nor_5  g07178(.A(new_n9526), .B(new_n9525), .Y(new_n9527));
  not_8  g07179(.A(new_n9525), .Y(new_n9528));
  xnor_4 g07180(.A(new_n9526), .B(new_n9528), .Y(new_n9529));
  xnor_4 g07181(.A(new_n9510), .B(new_n9509), .Y(new_n9530));
  not_8  g07182(.A(n22591), .Y(new_n9531));
  not_8  g07183(.A(n26167), .Y(new_n9532));
  nor_5  g07184(.A(new_n7199), .B(new_n9532), .Y(new_n9533));
  xnor_4 g07185(.A(new_n9533), .B(new_n9531), .Y(new_n9534));
  and_5  g07186(.A(new_n9534), .B(new_n9530), .Y(new_n9535));
  or_5   g07187(.A(new_n7200), .B(new_n9532), .Y(new_n9536));
  nor_5  g07188(.A(new_n9536), .B(n22591), .Y(new_n9537));
  nor_5  g07189(.A(new_n9537), .B(new_n9535), .Y(new_n9538));
  and_5  g07190(.A(new_n9538), .B(new_n9529), .Y(new_n9539));
  nor_5  g07191(.A(new_n9539), .B(new_n9527), .Y(new_n9540));
  nor_5  g07192(.A(new_n9540), .B(new_n9523), .Y(new_n9541));
  or_5   g07193(.A(new_n9541), .B(new_n9522), .Y(new_n9542));
  xor_4  g07194(.A(new_n9542), .B(new_n9519), .Y(new_n9543));
  xnor_4 g07195(.A(new_n9543), .B(new_n9495), .Y(new_n9544));
  xnor_4 g07196(.A(new_n9540), .B(new_n9523), .Y(new_n9545));
  xor_4  g07197(.A(new_n9492), .B(new_n9480), .Y(new_n9546));
  nor_5  g07198(.A(new_n9546), .B(new_n9545), .Y(new_n9547));
  xnor_4 g07199(.A(new_n9546), .B(new_n9545), .Y(new_n9548));
  not_8  g07200(.A(new_n9548), .Y(new_n9549));
  xor_4  g07201(.A(new_n9538), .B(new_n9529), .Y(new_n9550));
  xnor_4 g07202(.A(new_n9490), .B(new_n9482), .Y(new_n9551));
  nor_5  g07203(.A(new_n9551), .B(new_n9550), .Y(new_n9552_1));
  xor_4  g07204(.A(new_n9551), .B(new_n9550), .Y(new_n9553));
  not_8  g07205(.A(new_n9530), .Y(new_n9554_1));
  xnor_4 g07206(.A(new_n9534), .B(new_n9554_1), .Y(new_n9555));
  nor_5  g07207(.A(new_n9485), .B(new_n9484), .Y(new_n9556_1));
  xnor_4 g07208(.A(new_n9488), .B(new_n9556_1), .Y(new_n9557_1));
  nor_5  g07209(.A(new_n9557_1), .B(new_n9555), .Y(new_n9558_1));
  nor_5  g07210(.A(new_n7201), .B(new_n7198), .Y(new_n9559));
  not_8  g07211(.A(new_n9557_1), .Y(new_n9560));
  xnor_4 g07212(.A(new_n9560), .B(new_n9555), .Y(new_n9561));
  and_5  g07213(.A(new_n9561), .B(new_n9559), .Y(new_n9562));
  nor_5  g07214(.A(new_n9562), .B(new_n9558_1), .Y(new_n9563));
  and_5  g07215(.A(new_n9563), .B(new_n9553), .Y(new_n9564));
  nor_5  g07216(.A(new_n9564), .B(new_n9552_1), .Y(new_n9565));
  and_5  g07217(.A(new_n9565), .B(new_n9549), .Y(new_n9566));
  nor_5  g07218(.A(new_n9566), .B(new_n9547), .Y(new_n9567));
  xor_4  g07219(.A(new_n9567), .B(new_n9544), .Y(n1111));
  xnor_4 g07220(.A(new_n2607), .B(new_n4431), .Y(new_n9569));
  nor_5  g07221(.A(new_n2611), .B(new_n4435), .Y(new_n9570));
  xnor_4 g07222(.A(new_n2611), .B(new_n4435), .Y(new_n9571));
  nor_5  g07223(.A(new_n2647), .B(new_n4442), .Y(new_n9572));
  nor_5  g07224(.A(new_n2615), .B(n11011), .Y(new_n9573));
  xnor_4 g07225(.A(new_n2615), .B(n11011), .Y(new_n9574));
  nor_5  g07226(.A(new_n2618), .B(n16029), .Y(new_n9575));
  xnor_4 g07227(.A(new_n2618), .B(new_n3939), .Y(new_n9576));
  nor_5  g07228(.A(new_n2623), .B(new_n3943), .Y(new_n9577));
  xnor_4 g07229(.A(new_n2623), .B(new_n3943), .Y(new_n9578));
  nor_5  g07230(.A(new_n2636), .B(new_n3947), .Y(new_n9579));
  nor_5  g07231(.A(new_n2627), .B(n22433), .Y(new_n9580));
  nor_5  g07232(.A(new_n2630), .B(new_n3952_1), .Y(new_n9581));
  xnor_4 g07233(.A(new_n2627), .B(n22433), .Y(new_n9582));
  nor_5  g07234(.A(new_n9582), .B(new_n9581), .Y(new_n9583));
  nor_5  g07235(.A(new_n9583), .B(new_n9580), .Y(new_n9584));
  xnor_4 g07236(.A(new_n2636), .B(n11615), .Y(new_n9585));
  and_5  g07237(.A(new_n9585), .B(new_n9584), .Y(new_n9586));
  nor_5  g07238(.A(new_n9586), .B(new_n9579), .Y(new_n9587));
  nor_5  g07239(.A(new_n9587), .B(new_n9578), .Y(new_n9588));
  nor_5  g07240(.A(new_n9588), .B(new_n9577), .Y(new_n9589));
  and_5  g07241(.A(new_n9589), .B(new_n9576), .Y(new_n9590));
  nor_5  g07242(.A(new_n9590), .B(new_n9575), .Y(new_n9591));
  nor_5  g07243(.A(new_n9591), .B(new_n9574), .Y(new_n9592));
  or_5   g07244(.A(new_n9592), .B(new_n9573), .Y(new_n9593));
  xnor_4 g07245(.A(new_n2647), .B(new_n4442), .Y(new_n9594));
  nor_5  g07246(.A(new_n9594), .B(new_n9593), .Y(new_n9595));
  nor_5  g07247(.A(new_n9595), .B(new_n9572), .Y(new_n9596));
  nor_5  g07248(.A(new_n9596), .B(new_n9571), .Y(new_n9597));
  nor_5  g07249(.A(new_n9597), .B(new_n9570), .Y(new_n9598_1));
  xor_4  g07250(.A(new_n9598_1), .B(new_n9569), .Y(new_n9599));
  not_8  g07251(.A(new_n9599), .Y(new_n9600));
  not_8  g07252(.A(new_n9412), .Y(new_n9601));
  nor_5  g07253(.A(new_n9601), .B(n25074), .Y(new_n9602));
  not_8  g07254(.A(new_n9602), .Y(new_n9603));
  nor_5  g07255(.A(new_n9603), .B(n8006), .Y(new_n9604));
  not_8  g07256(.A(new_n9604), .Y(new_n9605));
  nor_5  g07257(.A(new_n9605), .B(n20929), .Y(new_n9606));
  not_8  g07258(.A(new_n9606), .Y(new_n9607));
  nor_5  g07259(.A(new_n9607), .B(n10710), .Y(new_n9608));
  not_8  g07260(.A(new_n9608), .Y(new_n9609));
  nor_5  g07261(.A(new_n9609), .B(n11841), .Y(new_n9610));
  xnor_4 g07262(.A(new_n9610), .B(n27089), .Y(new_n9611));
  xnor_4 g07263(.A(new_n9611), .B(new_n2725), .Y(new_n9612));
  xnor_4 g07264(.A(new_n9608), .B(n11841), .Y(new_n9613));
  and_5  g07265(.A(new_n9613), .B(new_n2729), .Y(new_n9614));
  not_8  g07266(.A(new_n2729), .Y(new_n9615));
  xnor_4 g07267(.A(new_n9613), .B(new_n9615), .Y(new_n9616_1));
  xnor_4 g07268(.A(new_n9606), .B(n10710), .Y(new_n9617));
  nor_5  g07269(.A(new_n9617), .B(new_n2733), .Y(new_n9618));
  xnor_4 g07270(.A(new_n9617), .B(new_n2733), .Y(new_n9619));
  xnor_4 g07271(.A(new_n9604), .B(n20929), .Y(new_n9620));
  nor_5  g07272(.A(new_n9620), .B(new_n2738), .Y(new_n9621));
  xnor_4 g07273(.A(new_n9620), .B(new_n2740), .Y(new_n9622_1));
  xnor_4 g07274(.A(new_n9602), .B(n8006), .Y(new_n9623));
  nor_5  g07275(.A(new_n9623), .B(new_n2744), .Y(new_n9624));
  nor_5  g07276(.A(new_n9413), .B(new_n2748), .Y(new_n9625));
  not_8  g07277(.A(new_n2748), .Y(new_n9626_1));
  xnor_4 g07278(.A(new_n9413), .B(new_n9626_1), .Y(new_n9627));
  nor_5  g07279(.A(new_n9415), .B(new_n2753), .Y(new_n9628));
  not_8  g07280(.A(new_n2753), .Y(new_n9629));
  xnor_4 g07281(.A(new_n9415), .B(new_n9629), .Y(new_n9630));
  nor_5  g07282(.A(new_n5781), .B(new_n2759), .Y(new_n9631));
  nor_5  g07283(.A(new_n2761_1), .B(n2088), .Y(new_n9632));
  xnor_4 g07284(.A(new_n5781), .B(new_n2763), .Y(new_n9633_1));
  and_5  g07285(.A(new_n9633_1), .B(new_n9632), .Y(new_n9634));
  or_5   g07286(.A(new_n9634), .B(new_n9631), .Y(new_n9635_1));
  and_5  g07287(.A(new_n9635_1), .B(new_n9630), .Y(new_n9636));
  or_5   g07288(.A(new_n9636), .B(new_n9628), .Y(new_n9637));
  and_5  g07289(.A(new_n9637), .B(new_n9627), .Y(new_n9638));
  or_5   g07290(.A(new_n9638), .B(new_n9625), .Y(new_n9639));
  xnor_4 g07291(.A(new_n9623), .B(new_n2771), .Y(new_n9640));
  and_5  g07292(.A(new_n9640), .B(new_n9639), .Y(new_n9641));
  or_5   g07293(.A(new_n9641), .B(new_n9624), .Y(new_n9642));
  and_5  g07294(.A(new_n9642), .B(new_n9622_1), .Y(new_n9643));
  nor_5  g07295(.A(new_n9643), .B(new_n9621), .Y(new_n9644));
  nor_5  g07296(.A(new_n9644), .B(new_n9619), .Y(new_n9645));
  nor_5  g07297(.A(new_n9645), .B(new_n9618), .Y(new_n9646_1));
  and_5  g07298(.A(new_n9646_1), .B(new_n9616_1), .Y(new_n9647));
  or_5   g07299(.A(new_n9647), .B(new_n9614), .Y(new_n9648_1));
  xor_4  g07300(.A(new_n9648_1), .B(new_n9612), .Y(new_n9649));
  xnor_4 g07301(.A(new_n9649), .B(new_n9600), .Y(new_n9650));
  xor_4  g07302(.A(new_n9596), .B(new_n9571), .Y(new_n9651));
  not_8  g07303(.A(new_n9651), .Y(new_n9652));
  xnor_4 g07304(.A(new_n9646_1), .B(new_n9616_1), .Y(new_n9653));
  nor_5  g07305(.A(new_n9653), .B(new_n9652), .Y(new_n9654));
  xnor_4 g07306(.A(new_n9653), .B(new_n9651), .Y(new_n9655_1));
  nor_5  g07307(.A(new_n9592), .B(new_n9573), .Y(new_n9656));
  xnor_4 g07308(.A(new_n9594), .B(new_n9656), .Y(new_n9657));
  xnor_4 g07309(.A(new_n9644), .B(new_n9619), .Y(new_n9658));
  nor_5  g07310(.A(new_n9658), .B(new_n9657), .Y(new_n9659));
  not_8  g07311(.A(new_n9657), .Y(new_n9660));
  xnor_4 g07312(.A(new_n9658), .B(new_n9660), .Y(new_n9661));
  xnor_4 g07313(.A(new_n9591), .B(new_n9574), .Y(new_n9662));
  not_8  g07314(.A(new_n9662), .Y(new_n9663));
  xor_4  g07315(.A(new_n9642), .B(new_n9622_1), .Y(new_n9664));
  nor_5  g07316(.A(new_n9664), .B(new_n9663), .Y(new_n9665));
  xnor_4 g07317(.A(new_n9664), .B(new_n9662), .Y(new_n9666));
  xnor_4 g07318(.A(new_n9589), .B(new_n9576), .Y(new_n9667));
  not_8  g07319(.A(new_n9667), .Y(new_n9668));
  xor_4  g07320(.A(new_n9640), .B(new_n9639), .Y(new_n9669));
  nor_5  g07321(.A(new_n9669), .B(new_n9668), .Y(new_n9670));
  xnor_4 g07322(.A(new_n9669), .B(new_n9667), .Y(new_n9671));
  xor_4  g07323(.A(new_n9637), .B(new_n9627), .Y(new_n9672));
  xnor_4 g07324(.A(new_n9587), .B(new_n9578), .Y(new_n9673));
  nor_5  g07325(.A(new_n9673), .B(new_n9672), .Y(new_n9674));
  not_8  g07326(.A(new_n9673), .Y(new_n9675));
  xnor_4 g07327(.A(new_n9675), .B(new_n9672), .Y(new_n9676));
  xor_4  g07328(.A(new_n9635_1), .B(new_n9630), .Y(new_n9677));
  xnor_4 g07329(.A(new_n9585), .B(new_n9584), .Y(new_n9678));
  nor_5  g07330(.A(new_n9678), .B(new_n9677), .Y(new_n9679));
  not_8  g07331(.A(new_n9678), .Y(new_n9680));
  xnor_4 g07332(.A(new_n9680), .B(new_n9677), .Y(new_n9681));
  xnor_4 g07333(.A(new_n9633_1), .B(new_n9632), .Y(new_n9682));
  xnor_4 g07334(.A(new_n9582), .B(new_n9581), .Y(new_n9683));
  nor_5  g07335(.A(new_n9683), .B(new_n9682), .Y(new_n9684));
  xnor_4 g07336(.A(new_n2630), .B(n14090), .Y(new_n9685));
  not_8  g07337(.A(new_n9685), .Y(new_n9686));
  xnor_4 g07338(.A(new_n2761_1), .B(new_n2951), .Y(new_n9687));
  nor_5  g07339(.A(new_n9687), .B(new_n9686), .Y(new_n9688));
  xnor_4 g07340(.A(new_n9683), .B(new_n9682), .Y(new_n9689_1));
  nor_5  g07341(.A(new_n9689_1), .B(new_n9688), .Y(new_n9690));
  nor_5  g07342(.A(new_n9690), .B(new_n9684), .Y(new_n9691));
  and_5  g07343(.A(new_n9691), .B(new_n9681), .Y(new_n9692));
  or_5   g07344(.A(new_n9692), .B(new_n9679), .Y(new_n9693));
  and_5  g07345(.A(new_n9693), .B(new_n9676), .Y(new_n9694));
  or_5   g07346(.A(new_n9694), .B(new_n9674), .Y(new_n9695_1));
  and_5  g07347(.A(new_n9695_1), .B(new_n9671), .Y(new_n9696));
  or_5   g07348(.A(new_n9696), .B(new_n9670), .Y(new_n9697));
  and_5  g07349(.A(new_n9697), .B(new_n9666), .Y(new_n9698));
  nor_5  g07350(.A(new_n9698), .B(new_n9665), .Y(new_n9699_1));
  and_5  g07351(.A(new_n9699_1), .B(new_n9661), .Y(new_n9700));
  nor_5  g07352(.A(new_n9700), .B(new_n9659), .Y(new_n9701));
  and_5  g07353(.A(new_n9701), .B(new_n9655_1), .Y(new_n9702));
  nor_5  g07354(.A(new_n9702), .B(new_n9654), .Y(new_n9703));
  xnor_4 g07355(.A(new_n9703), .B(new_n9650), .Y(n1119));
  xnor_4 g07356(.A(new_n7877), .B(new_n7879), .Y(new_n9705));
  xnor_4 g07357(.A(new_n9705), .B(new_n7902), .Y(n1120));
  xnor_4 g07358(.A(n9246), .B(n3925), .Y(new_n9707));
  xnor_4 g07359(.A(new_n9707), .B(new_n7749), .Y(new_n9708));
  not_8  g07360(.A(new_n9708), .Y(new_n9709));
  xnor_4 g07361(.A(n12495), .B(n7428), .Y(new_n9710));
  xnor_4 g07362(.A(new_n9710), .B(new_n9709), .Y(n1196));
  xnor_4 g07363(.A(n16223), .B(n15636), .Y(new_n9712));
  nor_5  g07364(.A(new_n2444_1), .B(n19494), .Y(new_n9713));
  or_5   g07365(.A(n20077), .B(new_n2365), .Y(new_n9714));
  nor_5  g07366(.A(new_n2447), .B(n2387), .Y(new_n9715));
  and_5  g07367(.A(new_n9715), .B(new_n9714), .Y(new_n9716));
  or_5   g07368(.A(new_n9716), .B(new_n9713), .Y(new_n9717));
  xor_4  g07369(.A(new_n9717), .B(new_n9712), .Y(new_n9718));
  xnor_4 g07370(.A(new_n9718), .B(new_n7882), .Y(new_n9719));
  xnor_4 g07371(.A(n6794), .B(n2387), .Y(new_n9720));
  nor_5  g07372(.A(new_n9720), .B(new_n7890), .Y(new_n9721));
  xnor_4 g07373(.A(n20077), .B(n19494), .Y(new_n9722));
  xnor_4 g07374(.A(new_n9722), .B(new_n9715), .Y(new_n9723));
  nor_5  g07375(.A(new_n9723), .B(new_n9721), .Y(new_n9724));
  xnor_4 g07376(.A(new_n9723), .B(new_n9721), .Y(new_n9725));
  nor_5  g07377(.A(new_n9725), .B(new_n7884_1), .Y(new_n9726_1));
  nor_5  g07378(.A(new_n9726_1), .B(new_n9724), .Y(new_n9727));
  xnor_4 g07379(.A(new_n9727), .B(new_n9719), .Y(n1237));
  xnor_4 g07380(.A(new_n5702), .B(new_n5498), .Y(new_n9729));
  xnor_4 g07381(.A(new_n9729), .B(new_n5765_1), .Y(n1239));
  xnor_4 g07382(.A(n22764), .B(n1536), .Y(new_n9731));
  nor_5  g07383(.A(n26264), .B(n19454), .Y(new_n9732));
  xnor_4 g07384(.A(n26264), .B(n19454), .Y(new_n9733));
  nor_5  g07385(.A(n9445), .B(n7841), .Y(new_n9734));
  xnor_4 g07386(.A(n9445), .B(n7841), .Y(new_n9735));
  nor_5  g07387(.A(n16812), .B(n1279), .Y(new_n9736));
  xnor_4 g07388(.A(n16812), .B(n1279), .Y(new_n9737));
  nor_5  g07389(.A(n25068), .B(n8324), .Y(new_n9738));
  xnor_4 g07390(.A(n25068), .B(n8324), .Y(new_n9739));
  nor_5  g07391(.A(n12546), .B(n2331), .Y(new_n9740));
  xnor_4 g07392(.A(n12546), .B(n2331), .Y(new_n9741));
  nor_5  g07393(.A(n22631), .B(n21078), .Y(new_n9742));
  xnor_4 g07394(.A(n22631), .B(n21078), .Y(new_n9743));
  nor_5  g07395(.A(n24485), .B(n16743), .Y(new_n9744));
  xnor_4 g07396(.A(n24485), .B(n16743), .Y(new_n9745));
  nor_5  g07397(.A(n15258), .B(n2420), .Y(new_n9746));
  nor_5  g07398(.A(new_n8110), .B(new_n2542), .Y(new_n9747));
  xnor_4 g07399(.A(n15258), .B(n2420), .Y(new_n9748));
  nor_5  g07400(.A(new_n9748), .B(new_n9747), .Y(new_n9749));
  nor_5  g07401(.A(new_n9749), .B(new_n9746), .Y(new_n9750));
  nor_5  g07402(.A(new_n9750), .B(new_n9745), .Y(new_n9751));
  nor_5  g07403(.A(new_n9751), .B(new_n9744), .Y(new_n9752));
  nor_5  g07404(.A(new_n9752), .B(new_n9743), .Y(new_n9753_1));
  nor_5  g07405(.A(new_n9753_1), .B(new_n9742), .Y(new_n9754));
  nor_5  g07406(.A(new_n9754), .B(new_n9741), .Y(new_n9755));
  nor_5  g07407(.A(new_n9755), .B(new_n9740), .Y(new_n9756));
  nor_5  g07408(.A(new_n9756), .B(new_n9739), .Y(new_n9757));
  nor_5  g07409(.A(new_n9757), .B(new_n9738), .Y(new_n9758));
  nor_5  g07410(.A(new_n9758), .B(new_n9737), .Y(new_n9759));
  nor_5  g07411(.A(new_n9759), .B(new_n9736), .Y(new_n9760));
  nor_5  g07412(.A(new_n9760), .B(new_n9735), .Y(new_n9761_1));
  nor_5  g07413(.A(new_n9761_1), .B(new_n9734), .Y(new_n9762));
  nor_5  g07414(.A(new_n9762), .B(new_n9733), .Y(new_n9763_1));
  nor_5  g07415(.A(new_n9763_1), .B(new_n9732), .Y(new_n9764));
  xnor_4 g07416(.A(new_n9764), .B(new_n9731), .Y(new_n9765));
  nor_5  g07417(.A(new_n9765), .B(n2416), .Y(new_n9766));
  xnor_4 g07418(.A(new_n9765), .B(n2416), .Y(new_n9767_1));
  xnor_4 g07419(.A(new_n9762), .B(new_n9733), .Y(new_n9768));
  nor_5  g07420(.A(new_n9768), .B(n21905), .Y(new_n9769));
  xnor_4 g07421(.A(new_n9768), .B(n21905), .Y(new_n9770));
  xnor_4 g07422(.A(new_n9760), .B(new_n9735), .Y(new_n9771_1));
  nor_5  g07423(.A(new_n9771_1), .B(n22918), .Y(new_n9772));
  xnor_4 g07424(.A(new_n9771_1), .B(n22918), .Y(new_n9773));
  xnor_4 g07425(.A(new_n9758), .B(new_n9737), .Y(new_n9774));
  nor_5  g07426(.A(new_n9774), .B(n25923), .Y(new_n9775));
  xnor_4 g07427(.A(new_n9774), .B(n25923), .Y(new_n9776));
  xnor_4 g07428(.A(new_n9756), .B(new_n9739), .Y(new_n9777));
  nor_5  g07429(.A(new_n9777), .B(n6790), .Y(new_n9778_1));
  xnor_4 g07430(.A(new_n9777), .B(n6790), .Y(new_n9779));
  xnor_4 g07431(.A(new_n9754), .B(new_n9741), .Y(new_n9780));
  nor_5  g07432(.A(new_n9780), .B(n22879), .Y(new_n9781));
  xnor_4 g07433(.A(new_n9780), .B(n22879), .Y(new_n9782));
  xnor_4 g07434(.A(new_n9752), .B(new_n9743), .Y(new_n9783_1));
  nor_5  g07435(.A(new_n9783_1), .B(n2117), .Y(new_n9784));
  xnor_4 g07436(.A(new_n9783_1), .B(n2117), .Y(new_n9785));
  xnor_4 g07437(.A(new_n9750), .B(new_n9745), .Y(new_n9786));
  nor_5  g07438(.A(new_n9786), .B(n5882), .Y(new_n9787));
  xnor_4 g07439(.A(new_n9748), .B(new_n9747), .Y(new_n9788));
  nor_5  g07440(.A(new_n9788), .B(n11775), .Y(new_n9789));
  not_8  g07441(.A(n27134), .Y(new_n9790));
  xnor_4 g07442(.A(n22201), .B(n4588), .Y(new_n9791));
  or_5   g07443(.A(new_n9791), .B(new_n9790), .Y(new_n9792));
  not_8  g07444(.A(n11775), .Y(new_n9793));
  xnor_4 g07445(.A(new_n9788), .B(new_n9793), .Y(new_n9794));
  and_5  g07446(.A(new_n9794), .B(new_n9792), .Y(new_n9795));
  nor_5  g07447(.A(new_n9795), .B(new_n9789), .Y(new_n9796));
  xnor_4 g07448(.A(new_n9786), .B(n5882), .Y(new_n9797));
  nor_5  g07449(.A(new_n9797), .B(new_n9796), .Y(new_n9798));
  nor_5  g07450(.A(new_n9798), .B(new_n9787), .Y(new_n9799));
  nor_5  g07451(.A(new_n9799), .B(new_n9785), .Y(new_n9800));
  nor_5  g07452(.A(new_n9800), .B(new_n9784), .Y(new_n9801));
  nor_5  g07453(.A(new_n9801), .B(new_n9782), .Y(new_n9802));
  nor_5  g07454(.A(new_n9802), .B(new_n9781), .Y(new_n9803_1));
  nor_5  g07455(.A(new_n9803_1), .B(new_n9779), .Y(new_n9804));
  nor_5  g07456(.A(new_n9804), .B(new_n9778_1), .Y(new_n9805));
  nor_5  g07457(.A(new_n9805), .B(new_n9776), .Y(new_n9806));
  nor_5  g07458(.A(new_n9806), .B(new_n9775), .Y(new_n9807));
  nor_5  g07459(.A(new_n9807), .B(new_n9773), .Y(new_n9808));
  nor_5  g07460(.A(new_n9808), .B(new_n9772), .Y(new_n9809));
  nor_5  g07461(.A(new_n9809), .B(new_n9770), .Y(new_n9810));
  nor_5  g07462(.A(new_n9810), .B(new_n9769), .Y(new_n9811));
  nor_5  g07463(.A(new_n9811), .B(new_n9767_1), .Y(new_n9812));
  nor_5  g07464(.A(new_n9812), .B(new_n9766), .Y(new_n9813));
  nor_5  g07465(.A(n22764), .B(n1536), .Y(new_n9814));
  nor_5  g07466(.A(new_n9764), .B(new_n9731), .Y(new_n9815));
  nor_5  g07467(.A(new_n9815), .B(new_n9814), .Y(new_n9816));
  and_5  g07468(.A(new_n9816), .B(new_n9813), .Y(new_n9817));
  nor_5  g07469(.A(n23493), .B(n8405), .Y(new_n9818));
  nor_5  g07470(.A(n22359), .B(n10275), .Y(new_n9819));
  nor_5  g07471(.A(n15146), .B(n5532), .Y(new_n9820));
  nor_5  g07472(.A(n11579), .B(n3962), .Y(new_n9821));
  nor_5  g07473(.A(n23513), .B(n21), .Y(new_n9822));
  xnor_4 g07474(.A(n23513), .B(n21), .Y(new_n9823));
  nor_5  g07475(.A(n6427), .B(n1682), .Y(new_n9824));
  and_5  g07476(.A(n6427), .B(n1682), .Y(new_n9825));
  nor_5  g07477(.A(n7963), .B(n6590), .Y(new_n9826));
  nor_5  g07478(.A(n20349), .B(n10017), .Y(new_n9827));
  not_8  g07479(.A(n15936), .Y(new_n9828));
  nor_5  g07480(.A(new_n9828), .B(new_n7939), .Y(new_n9829));
  not_8  g07481(.A(n20349), .Y(new_n9830));
  nor_5  g07482(.A(new_n9830), .B(new_n7941), .Y(new_n9831));
  nor_5  g07483(.A(new_n9831), .B(new_n9829), .Y(new_n9832_1));
  nor_5  g07484(.A(new_n9832_1), .B(new_n9827), .Y(new_n9833_1));
  not_8  g07485(.A(n6590), .Y(new_n9834));
  not_8  g07486(.A(n7963), .Y(new_n9835));
  nor_5  g07487(.A(new_n9835), .B(new_n9834), .Y(new_n9836));
  nor_5  g07488(.A(new_n9836), .B(new_n9833_1), .Y(new_n9837));
  nor_5  g07489(.A(new_n9837), .B(new_n9826), .Y(new_n9838_1));
  nor_5  g07490(.A(new_n9838_1), .B(new_n9825), .Y(new_n9839));
  nor_5  g07491(.A(new_n9839), .B(new_n9824), .Y(new_n9840));
  nor_5  g07492(.A(new_n9840), .B(new_n9823), .Y(new_n9841));
  nor_5  g07493(.A(new_n9841), .B(new_n9822), .Y(new_n9842));
  xnor_4 g07494(.A(n11579), .B(n3962), .Y(new_n9843));
  nor_5  g07495(.A(new_n9843), .B(new_n9842), .Y(new_n9844));
  nor_5  g07496(.A(new_n9844), .B(new_n9821), .Y(new_n9845));
  xnor_4 g07497(.A(n15146), .B(n5532), .Y(new_n9846));
  nor_5  g07498(.A(new_n9846), .B(new_n9845), .Y(new_n9847));
  nor_5  g07499(.A(new_n9847), .B(new_n9820), .Y(new_n9848));
  xnor_4 g07500(.A(n22359), .B(n10275), .Y(new_n9849));
  nor_5  g07501(.A(new_n9849), .B(new_n9848), .Y(new_n9850));
  nor_5  g07502(.A(new_n9850), .B(new_n9819), .Y(new_n9851));
  xnor_4 g07503(.A(n23493), .B(n8405), .Y(new_n9852));
  nor_5  g07504(.A(new_n9852), .B(new_n9851), .Y(new_n9853));
  nor_5  g07505(.A(new_n9853), .B(new_n9818), .Y(new_n9854));
  xnor_4 g07506(.A(n14826), .B(n13549), .Y(new_n9855));
  xnor_4 g07507(.A(new_n9855), .B(new_n9854), .Y(new_n9856));
  nor_5  g07508(.A(new_n9856), .B(n18105), .Y(new_n9857));
  xnor_4 g07509(.A(new_n9856), .B(n18105), .Y(new_n9858));
  xnor_4 g07510(.A(new_n9852), .B(new_n9851), .Y(new_n9859));
  nor_5  g07511(.A(new_n9859), .B(n24196), .Y(new_n9860));
  xnor_4 g07512(.A(new_n9859), .B(n24196), .Y(new_n9861));
  xnor_4 g07513(.A(new_n9849), .B(new_n9848), .Y(new_n9862));
  nor_5  g07514(.A(new_n9862), .B(n16376), .Y(new_n9863));
  xnor_4 g07515(.A(new_n9862), .B(n16376), .Y(new_n9864));
  xnor_4 g07516(.A(new_n9846), .B(new_n9845), .Y(new_n9865));
  nor_5  g07517(.A(new_n9865), .B(n25381), .Y(new_n9866));
  xnor_4 g07518(.A(new_n9865), .B(n25381), .Y(new_n9867_1));
  xnor_4 g07519(.A(new_n9843), .B(new_n9842), .Y(new_n9868));
  nor_5  g07520(.A(new_n9868), .B(n12587), .Y(new_n9869));
  xnor_4 g07521(.A(new_n9868), .B(n12587), .Y(new_n9870));
  xnor_4 g07522(.A(new_n9840), .B(new_n9823), .Y(new_n9871));
  nor_5  g07523(.A(new_n9871), .B(n268), .Y(new_n9872_1));
  xnor_4 g07524(.A(new_n9871), .B(n268), .Y(new_n9873));
  xnor_4 g07525(.A(n6427), .B(new_n7934), .Y(new_n9874));
  not_8  g07526(.A(new_n9874), .Y(new_n9875));
  xnor_4 g07527(.A(new_n9875), .B(new_n9838_1), .Y(new_n9876));
  nor_5  g07528(.A(new_n9876), .B(n24879), .Y(new_n9877));
  xnor_4 g07529(.A(new_n9876), .B(n24879), .Y(new_n9878));
  xnor_4 g07530(.A(n7963), .B(n6590), .Y(new_n9879));
  xnor_4 g07531(.A(new_n9879), .B(new_n9833_1), .Y(new_n9880));
  nor_5  g07532(.A(new_n9880), .B(n6785), .Y(new_n9881));
  xnor_4 g07533(.A(n20349), .B(n10017), .Y(new_n9882));
  xnor_4 g07534(.A(new_n9882), .B(new_n9829), .Y(new_n9883));
  nor_5  g07535(.A(new_n9883), .B(n24032), .Y(new_n9884));
  xnor_4 g07536(.A(n15936), .B(n3618), .Y(new_n9885));
  or_5   g07537(.A(new_n9885), .B(new_n4507), .Y(new_n9886));
  xnor_4 g07538(.A(new_n9883), .B(new_n8052_1), .Y(new_n9887));
  and_5  g07539(.A(new_n9887), .B(new_n9886), .Y(new_n9888));
  nor_5  g07540(.A(new_n9888), .B(new_n9884), .Y(new_n9889));
  xnor_4 g07541(.A(new_n9880), .B(n6785), .Y(new_n9890_1));
  nor_5  g07542(.A(new_n9890_1), .B(new_n9889), .Y(new_n9891));
  nor_5  g07543(.A(new_n9891), .B(new_n9881), .Y(new_n9892));
  nor_5  g07544(.A(new_n9892), .B(new_n9878), .Y(new_n9893));
  nor_5  g07545(.A(new_n9893), .B(new_n9877), .Y(new_n9894));
  nor_5  g07546(.A(new_n9894), .B(new_n9873), .Y(new_n9895));
  nor_5  g07547(.A(new_n9895), .B(new_n9872_1), .Y(new_n9896));
  nor_5  g07548(.A(new_n9896), .B(new_n9870), .Y(new_n9897));
  nor_5  g07549(.A(new_n9897), .B(new_n9869), .Y(new_n9898));
  nor_5  g07550(.A(new_n9898), .B(new_n9867_1), .Y(new_n9899));
  nor_5  g07551(.A(new_n9899), .B(new_n9866), .Y(new_n9900));
  nor_5  g07552(.A(new_n9900), .B(new_n9864), .Y(new_n9901));
  nor_5  g07553(.A(new_n9901), .B(new_n9863), .Y(new_n9902));
  nor_5  g07554(.A(new_n9902), .B(new_n9861), .Y(new_n9903));
  nor_5  g07555(.A(new_n9903), .B(new_n9860), .Y(new_n9904));
  nor_5  g07556(.A(new_n9904), .B(new_n9858), .Y(new_n9905));
  nor_5  g07557(.A(new_n9905), .B(new_n9857), .Y(new_n9906));
  nor_5  g07558(.A(new_n9855), .B(new_n9854), .Y(new_n9907));
  nor_5  g07559(.A(n14826), .B(n13549), .Y(new_n9908));
  nor_5  g07560(.A(new_n9908), .B(new_n9907), .Y(new_n9909));
  nand_5 g07561(.A(new_n9909), .B(new_n9906), .Y(new_n9910));
  xnor_4 g07562(.A(new_n9910), .B(new_n9817), .Y(new_n9911));
  xnor_4 g07563(.A(new_n9816), .B(new_n9813), .Y(new_n9912));
  xnor_4 g07564(.A(new_n9909), .B(new_n9906), .Y(new_n9913));
  not_8  g07565(.A(new_n9913), .Y(new_n9914));
  and_5  g07566(.A(new_n9914), .B(new_n9912), .Y(new_n9915));
  xnor_4 g07567(.A(new_n9914), .B(new_n9912), .Y(new_n9916));
  xnor_4 g07568(.A(new_n9811), .B(new_n9767_1), .Y(new_n9917_1));
  xnor_4 g07569(.A(new_n9904), .B(new_n9858), .Y(new_n9918));
  not_8  g07570(.A(new_n9918), .Y(new_n9919_1));
  nor_5  g07571(.A(new_n9919_1), .B(new_n9917_1), .Y(new_n9920));
  xnor_4 g07572(.A(new_n9919_1), .B(new_n9917_1), .Y(new_n9921));
  xnor_4 g07573(.A(new_n9809), .B(new_n9770), .Y(new_n9922));
  xnor_4 g07574(.A(new_n9902), .B(new_n9861), .Y(new_n9923));
  not_8  g07575(.A(new_n9923), .Y(new_n9924));
  nor_5  g07576(.A(new_n9924), .B(new_n9922), .Y(new_n9925));
  xnor_4 g07577(.A(new_n9924), .B(new_n9922), .Y(new_n9926_1));
  xnor_4 g07578(.A(new_n9807), .B(new_n9773), .Y(new_n9927));
  xnor_4 g07579(.A(new_n9900), .B(new_n9864), .Y(new_n9928));
  not_8  g07580(.A(new_n9928), .Y(new_n9929));
  nor_5  g07581(.A(new_n9929), .B(new_n9927), .Y(new_n9930));
  xnor_4 g07582(.A(new_n9929), .B(new_n9927), .Y(new_n9931));
  xnor_4 g07583(.A(new_n9805), .B(new_n9776), .Y(new_n9932));
  xnor_4 g07584(.A(new_n9898), .B(new_n9867_1), .Y(new_n9933));
  not_8  g07585(.A(new_n9933), .Y(new_n9934_1));
  nor_5  g07586(.A(new_n9934_1), .B(new_n9932), .Y(new_n9935));
  xnor_4 g07587(.A(new_n9934_1), .B(new_n9932), .Y(new_n9936));
  xnor_4 g07588(.A(new_n9803_1), .B(new_n9779), .Y(new_n9937));
  xnor_4 g07589(.A(new_n9896), .B(new_n9870), .Y(new_n9938_1));
  not_8  g07590(.A(new_n9938_1), .Y(new_n9939));
  nor_5  g07591(.A(new_n9939), .B(new_n9937), .Y(new_n9940));
  xnor_4 g07592(.A(new_n9939), .B(new_n9937), .Y(new_n9941));
  xnor_4 g07593(.A(new_n9801), .B(new_n9782), .Y(new_n9942_1));
  xor_4  g07594(.A(new_n9894), .B(new_n9873), .Y(new_n9943));
  nor_5  g07595(.A(new_n9943), .B(new_n9942_1), .Y(new_n9944));
  xnor_4 g07596(.A(new_n9943), .B(new_n9942_1), .Y(new_n9945));
  xnor_4 g07597(.A(new_n9799), .B(new_n9785), .Y(new_n9946_1));
  xnor_4 g07598(.A(new_n9892), .B(new_n9878), .Y(new_n9947));
  not_8  g07599(.A(new_n9947), .Y(new_n9948));
  nor_5  g07600(.A(new_n9948), .B(new_n9946_1), .Y(new_n9949));
  xnor_4 g07601(.A(new_n9948), .B(new_n9946_1), .Y(new_n9950));
  xnor_4 g07602(.A(new_n9797), .B(new_n9796), .Y(new_n9951));
  xnor_4 g07603(.A(new_n9890_1), .B(new_n9889), .Y(new_n9952));
  not_8  g07604(.A(new_n9952), .Y(new_n9953));
  nor_5  g07605(.A(new_n9953), .B(new_n9951), .Y(new_n9954));
  xnor_4 g07606(.A(new_n9953), .B(new_n9951), .Y(new_n9955));
  xor_4  g07607(.A(new_n9794), .B(new_n9792), .Y(new_n9956));
  not_8  g07608(.A(new_n9956), .Y(new_n9957));
  nor_5  g07609(.A(new_n9885), .B(new_n4507), .Y(new_n9958));
  xnor_4 g07610(.A(new_n9887), .B(new_n9958), .Y(new_n9959));
  nor_5  g07611(.A(new_n9959), .B(new_n9957), .Y(new_n9960));
  xnor_4 g07612(.A(new_n9791), .B(n27134), .Y(new_n9961));
  xnor_4 g07613(.A(new_n9885), .B(n22843), .Y(new_n9962));
  not_8  g07614(.A(new_n9962), .Y(new_n9963));
  nor_5  g07615(.A(new_n9963), .B(new_n9961), .Y(new_n9964));
  not_8  g07616(.A(new_n9959), .Y(new_n9965));
  xnor_4 g07617(.A(new_n9965), .B(new_n9957), .Y(new_n9966));
  and_5  g07618(.A(new_n9966), .B(new_n9964), .Y(new_n9967_1));
  nor_5  g07619(.A(new_n9967_1), .B(new_n9960), .Y(new_n9968_1));
  nor_5  g07620(.A(new_n9968_1), .B(new_n9955), .Y(new_n9969));
  nor_5  g07621(.A(new_n9969), .B(new_n9954), .Y(new_n9970));
  nor_5  g07622(.A(new_n9970), .B(new_n9950), .Y(new_n9971));
  nor_5  g07623(.A(new_n9971), .B(new_n9949), .Y(new_n9972));
  nor_5  g07624(.A(new_n9972), .B(new_n9945), .Y(new_n9973));
  nor_5  g07625(.A(new_n9973), .B(new_n9944), .Y(new_n9974));
  nor_5  g07626(.A(new_n9974), .B(new_n9941), .Y(new_n9975));
  nor_5  g07627(.A(new_n9975), .B(new_n9940), .Y(new_n9976));
  nor_5  g07628(.A(new_n9976), .B(new_n9936), .Y(new_n9977));
  nor_5  g07629(.A(new_n9977), .B(new_n9935), .Y(new_n9978));
  nor_5  g07630(.A(new_n9978), .B(new_n9931), .Y(new_n9979));
  nor_5  g07631(.A(new_n9979), .B(new_n9930), .Y(new_n9980));
  nor_5  g07632(.A(new_n9980), .B(new_n9926_1), .Y(new_n9981));
  nor_5  g07633(.A(new_n9981), .B(new_n9925), .Y(new_n9982));
  nor_5  g07634(.A(new_n9982), .B(new_n9921), .Y(new_n9983));
  nor_5  g07635(.A(new_n9983), .B(new_n9920), .Y(new_n9984));
  nor_5  g07636(.A(new_n9984), .B(new_n9916), .Y(new_n9985));
  nor_5  g07637(.A(new_n9985), .B(new_n9915), .Y(new_n9986));
  xnor_4 g07638(.A(new_n9986), .B(new_n9911), .Y(n1302));
  nor_5  g07639(.A(n13951), .B(new_n8719), .Y(new_n9988));
  xnor_4 g07640(.A(n13951), .B(n12507), .Y(new_n9989));
  nor_5  g07641(.A(n22793), .B(new_n8789), .Y(new_n9990));
  xnor_4 g07642(.A(n22793), .B(n15077), .Y(new_n9991));
  not_8  g07643(.A(n3710), .Y(new_n9992));
  nor_5  g07644(.A(n8439), .B(new_n9992), .Y(new_n9993));
  xnor_4 g07645(.A(n8439), .B(n3710), .Y(new_n9994));
  nor_5  g07646(.A(new_n8745_1), .B(n25523), .Y(new_n9995));
  xnor_4 g07647(.A(n26318), .B(n25523), .Y(new_n9996));
  nor_5  g07648(.A(new_n8749), .B(n5579), .Y(new_n9997));
  xnor_4 g07649(.A(n26054), .B(n5579), .Y(new_n9998));
  nor_5  g07650(.A(n23430), .B(new_n8753), .Y(new_n9999));
  xnor_4 g07651(.A(n23430), .B(n19081), .Y(new_n10000));
  nor_5  g07652(.A(n10411), .B(new_n8771), .Y(new_n10001));
  xnor_4 g07653(.A(n10411), .B(n8309), .Y(new_n10002));
  not_8  g07654(.A(n16971), .Y(new_n10003));
  nor_5  g07655(.A(n19144), .B(new_n10003), .Y(new_n10004));
  nor_5  g07656(.A(new_n8759), .B(n16971), .Y(new_n10005));
  nor_5  g07657(.A(n12593), .B(new_n2756), .Y(new_n10006));
  not_8  g07658(.A(n12593), .Y(new_n10007));
  nor_5  g07659(.A(new_n10007), .B(n11503), .Y(new_n10008));
  nor_5  g07660(.A(new_n2828), .B(n13714), .Y(new_n10009_1));
  not_8  g07661(.A(new_n10009_1), .Y(new_n10010_1));
  nor_5  g07662(.A(new_n10010_1), .B(new_n10008), .Y(new_n10011));
  nor_5  g07663(.A(new_n10011), .B(new_n10006), .Y(new_n10012));
  nor_5  g07664(.A(new_n10012), .B(new_n10005), .Y(new_n10013));
  nor_5  g07665(.A(new_n10013), .B(new_n10004), .Y(new_n10014));
  and_5  g07666(.A(new_n10014), .B(new_n10002), .Y(new_n10015));
  or_5   g07667(.A(new_n10015), .B(new_n10001), .Y(new_n10016));
  and_5  g07668(.A(new_n10016), .B(new_n10000), .Y(new_n10017_1));
  or_5   g07669(.A(new_n10017_1), .B(new_n9999), .Y(new_n10018_1));
  and_5  g07670(.A(new_n10018_1), .B(new_n9998), .Y(new_n10019_1));
  or_5   g07671(.A(new_n10019_1), .B(new_n9997), .Y(new_n10020));
  and_5  g07672(.A(new_n10020), .B(new_n9996), .Y(new_n10021_1));
  or_5   g07673(.A(new_n10021_1), .B(new_n9995), .Y(new_n10022));
  and_5  g07674(.A(new_n10022), .B(new_n9994), .Y(new_n10023));
  or_5   g07675(.A(new_n10023), .B(new_n9993), .Y(new_n10024));
  and_5  g07676(.A(new_n10024), .B(new_n9991), .Y(new_n10025));
  or_5   g07677(.A(new_n10025), .B(new_n9990), .Y(new_n10026));
  and_5  g07678(.A(new_n10026), .B(new_n9989), .Y(new_n10027));
  nor_5  g07679(.A(new_n10027), .B(new_n9988), .Y(new_n10028));
  nor_5  g07680(.A(n12650), .B(n11220), .Y(new_n10029));
  not_8  g07681(.A(n11220), .Y(new_n10030));
  xnor_4 g07682(.A(n12650), .B(new_n10030), .Y(new_n10031));
  nor_5  g07683(.A(n22379), .B(n10201), .Y(new_n10032));
  xnor_4 g07684(.A(n22379), .B(new_n5560), .Y(new_n10033));
  nor_5  g07685(.A(n10593), .B(n1662), .Y(new_n10034));
  xnor_4 g07686(.A(n10593), .B(new_n2850), .Y(new_n10035));
  nor_5  g07687(.A(n18290), .B(n12875), .Y(new_n10036));
  and_5  g07688(.A(new_n9247), .B(new_n9226), .Y(new_n10037));
  or_5   g07689(.A(new_n10037), .B(new_n10036), .Y(new_n10038));
  and_5  g07690(.A(new_n10038), .B(new_n10035), .Y(new_n10039));
  or_5   g07691(.A(new_n10039), .B(new_n10034), .Y(new_n10040));
  and_5  g07692(.A(new_n10040), .B(new_n10033), .Y(new_n10041));
  or_5   g07693(.A(new_n10041), .B(new_n10032), .Y(new_n10042));
  and_5  g07694(.A(new_n10042), .B(new_n10031), .Y(new_n10043));
  nor_5  g07695(.A(new_n10043), .B(new_n10029), .Y(new_n10044));
  not_8  g07696(.A(new_n10044), .Y(new_n10045));
  nor_5  g07697(.A(n22270), .B(n2944), .Y(new_n10046));
  or_5   g07698(.A(new_n2717), .B(new_n2676), .Y(new_n10047));
  and_5  g07699(.A(new_n10047), .B(new_n2675), .Y(new_n10048));
  nor_5  g07700(.A(new_n10048), .B(new_n10046), .Y(new_n10049));
  not_8  g07701(.A(new_n10049), .Y(new_n10050));
  xnor_4 g07702(.A(new_n10050), .B(new_n10045), .Y(new_n10051));
  not_8  g07703(.A(new_n2719), .Y(new_n10052));
  nor_5  g07704(.A(new_n10041), .B(new_n10032), .Y(new_n10053_1));
  xnor_4 g07705(.A(new_n10053_1), .B(new_n10031), .Y(new_n10054));
  nor_5  g07706(.A(new_n10054), .B(new_n10052), .Y(new_n10055_1));
  nor_5  g07707(.A(new_n10039), .B(new_n10034), .Y(new_n10056));
  xnor_4 g07708(.A(new_n10056), .B(new_n10033), .Y(new_n10057_1));
  not_8  g07709(.A(new_n10057_1), .Y(new_n10058));
  nor_5  g07710(.A(new_n10058), .B(new_n2723), .Y(new_n10059));
  xnor_4 g07711(.A(new_n10057_1), .B(new_n2725), .Y(new_n10060));
  nor_5  g07712(.A(new_n10037), .B(new_n10036), .Y(new_n10061));
  xnor_4 g07713(.A(new_n10061), .B(new_n10035), .Y(new_n10062));
  not_8  g07714(.A(new_n10062), .Y(new_n10063));
  nor_5  g07715(.A(new_n10063), .B(new_n2729), .Y(new_n10064));
  xnor_4 g07716(.A(new_n10062), .B(new_n9615), .Y(new_n10065));
  nor_5  g07717(.A(new_n9249), .B(new_n2733), .Y(new_n10066));
  nor_5  g07718(.A(new_n9251_1), .B(new_n2738), .Y(new_n10067));
  xnor_4 g07719(.A(new_n9251_1), .B(new_n2740), .Y(new_n10068));
  nor_5  g07720(.A(new_n9255), .B(new_n2771), .Y(new_n10069));
  nor_5  g07721(.A(new_n9261_1), .B(new_n2748), .Y(new_n10070));
  xnor_4 g07722(.A(new_n9261_1), .B(new_n9626_1), .Y(new_n10071));
  nor_5  g07723(.A(new_n9266), .B(new_n2753), .Y(new_n10072));
  xnor_4 g07724(.A(new_n9266), .B(new_n9629), .Y(new_n10073));
  nor_5  g07725(.A(new_n9274), .B(new_n2759), .Y(new_n10074));
  nor_5  g07726(.A(new_n9271), .B(new_n2761_1), .Y(new_n10075));
  xnor_4 g07727(.A(new_n9274), .B(new_n2763), .Y(new_n10076));
  and_5  g07728(.A(new_n10076), .B(new_n10075), .Y(new_n10077));
  or_5   g07729(.A(new_n10077), .B(new_n10074), .Y(new_n10078));
  and_5  g07730(.A(new_n10078), .B(new_n10073), .Y(new_n10079));
  or_5   g07731(.A(new_n10079), .B(new_n10072), .Y(new_n10080));
  and_5  g07732(.A(new_n10080), .B(new_n10071), .Y(new_n10081));
  nor_5  g07733(.A(new_n10081), .B(new_n10070), .Y(new_n10082));
  xnor_4 g07734(.A(new_n9256), .B(new_n2771), .Y(new_n10083));
  and_5  g07735(.A(new_n10083), .B(new_n10082), .Y(new_n10084));
  nor_5  g07736(.A(new_n10084), .B(new_n10069), .Y(new_n10085));
  and_5  g07737(.A(new_n10085), .B(new_n10068), .Y(new_n10086));
  nor_5  g07738(.A(new_n10086), .B(new_n10067), .Y(new_n10087));
  xnor_4 g07739(.A(new_n9249), .B(new_n2733), .Y(new_n10088));
  nor_5  g07740(.A(new_n10088), .B(new_n10087), .Y(new_n10089));
  nor_5  g07741(.A(new_n10089), .B(new_n10066), .Y(new_n10090));
  nor_5  g07742(.A(new_n10090), .B(new_n10065), .Y(new_n10091));
  nor_5  g07743(.A(new_n10091), .B(new_n10064), .Y(new_n10092));
  nor_5  g07744(.A(new_n10092), .B(new_n10060), .Y(new_n10093));
  nor_5  g07745(.A(new_n10093), .B(new_n10059), .Y(new_n10094));
  not_8  g07746(.A(new_n10054), .Y(new_n10095));
  xnor_4 g07747(.A(new_n10095), .B(new_n10052), .Y(new_n10096_1));
  and_5  g07748(.A(new_n10096_1), .B(new_n10094), .Y(new_n10097));
  or_5   g07749(.A(new_n10097), .B(new_n10055_1), .Y(new_n10098));
  xor_4  g07750(.A(new_n10098), .B(new_n10051), .Y(new_n10099));
  xnor_4 g07751(.A(new_n10099), .B(new_n10028), .Y(new_n10100));
  xor_4  g07752(.A(new_n10026), .B(new_n9989), .Y(new_n10101_1));
  xor_4  g07753(.A(new_n10096_1), .B(new_n10094), .Y(new_n10102));
  nor_5  g07754(.A(new_n10102), .B(new_n10101_1), .Y(new_n10103));
  xnor_4 g07755(.A(new_n10102), .B(new_n10101_1), .Y(new_n10104));
  xor_4  g07756(.A(new_n10024), .B(new_n9991), .Y(new_n10105));
  xnor_4 g07757(.A(new_n10092), .B(new_n10060), .Y(new_n10106));
  nor_5  g07758(.A(new_n10106), .B(new_n10105), .Y(new_n10107));
  xnor_4 g07759(.A(new_n10106), .B(new_n10105), .Y(new_n10108));
  xor_4  g07760(.A(new_n10022), .B(new_n9994), .Y(new_n10109));
  xnor_4 g07761(.A(new_n10090), .B(new_n10065), .Y(new_n10110));
  nor_5  g07762(.A(new_n10110), .B(new_n10109), .Y(new_n10111_1));
  xnor_4 g07763(.A(new_n10110), .B(new_n10109), .Y(new_n10112));
  xor_4  g07764(.A(new_n10020), .B(new_n9996), .Y(new_n10113));
  xnor_4 g07765(.A(new_n10088), .B(new_n10087), .Y(new_n10114));
  nor_5  g07766(.A(new_n10114), .B(new_n10113), .Y(new_n10115));
  xnor_4 g07767(.A(new_n10114), .B(new_n10113), .Y(new_n10116));
  xor_4  g07768(.A(new_n10018_1), .B(new_n9998), .Y(new_n10117_1));
  xnor_4 g07769(.A(new_n10085), .B(new_n10068), .Y(new_n10118));
  nor_5  g07770(.A(new_n10118), .B(new_n10117_1), .Y(new_n10119));
  xor_4  g07771(.A(new_n10016), .B(new_n10000), .Y(new_n10120));
  xor_4  g07772(.A(new_n10083), .B(new_n10082), .Y(new_n10121));
  nor_5  g07773(.A(new_n10121), .B(new_n10120), .Y(new_n10122));
  xnor_4 g07774(.A(new_n10121), .B(new_n10120), .Y(new_n10123));
  xor_4  g07775(.A(new_n10080), .B(new_n10071), .Y(new_n10124));
  xnor_4 g07776(.A(new_n10014), .B(new_n10002), .Y(new_n10125_1));
  and_5  g07777(.A(new_n10125_1), .B(new_n10124), .Y(new_n10126));
  nor_5  g07778(.A(new_n10077), .B(new_n10074), .Y(new_n10127));
  xnor_4 g07779(.A(new_n10127), .B(new_n10073), .Y(new_n10128));
  xnor_4 g07780(.A(n19144), .B(n16971), .Y(new_n10129));
  xnor_4 g07781(.A(new_n10129), .B(new_n10012), .Y(new_n10130));
  and_5  g07782(.A(new_n10130), .B(new_n10128), .Y(new_n10131));
  not_8  g07783(.A(new_n10128), .Y(new_n10132));
  xnor_4 g07784(.A(new_n10130), .B(new_n10132), .Y(new_n10133));
  xnor_4 g07785(.A(new_n9272), .B(new_n2761_1), .Y(new_n10134));
  xnor_4 g07786(.A(n18151), .B(n13714), .Y(new_n10135));
  nor_5  g07787(.A(new_n10135), .B(new_n10134), .Y(new_n10136));
  xnor_4 g07788(.A(n12593), .B(n11503), .Y(new_n10137));
  xnor_4 g07789(.A(new_n10137), .B(new_n10010_1), .Y(new_n10138));
  not_8  g07790(.A(new_n10138), .Y(new_n10139));
  and_5  g07791(.A(new_n10139), .B(new_n10136), .Y(new_n10140));
  xnor_4 g07792(.A(new_n10076), .B(new_n10075), .Y(new_n10141));
  not_8  g07793(.A(new_n10141), .Y(new_n10142));
  xnor_4 g07794(.A(new_n10139), .B(new_n10136), .Y(new_n10143));
  nor_5  g07795(.A(new_n10143), .B(new_n10142), .Y(new_n10144));
  nor_5  g07796(.A(new_n10144), .B(new_n10140), .Y(new_n10145));
  and_5  g07797(.A(new_n10145), .B(new_n10133), .Y(new_n10146));
  nor_5  g07798(.A(new_n10146), .B(new_n10131), .Y(new_n10147));
  xnor_4 g07799(.A(new_n10125_1), .B(new_n10124), .Y(new_n10148));
  nor_5  g07800(.A(new_n10148), .B(new_n10147), .Y(new_n10149));
  nor_5  g07801(.A(new_n10149), .B(new_n10126), .Y(new_n10150));
  nor_5  g07802(.A(new_n10150), .B(new_n10123), .Y(new_n10151));
  nor_5  g07803(.A(new_n10151), .B(new_n10122), .Y(new_n10152));
  xnor_4 g07804(.A(new_n10118), .B(new_n10117_1), .Y(new_n10153));
  nor_5  g07805(.A(new_n10153), .B(new_n10152), .Y(new_n10154));
  nor_5  g07806(.A(new_n10154), .B(new_n10119), .Y(new_n10155));
  nor_5  g07807(.A(new_n10155), .B(new_n10116), .Y(new_n10156));
  nor_5  g07808(.A(new_n10156), .B(new_n10115), .Y(new_n10157));
  nor_5  g07809(.A(new_n10157), .B(new_n10112), .Y(new_n10158_1));
  nor_5  g07810(.A(new_n10158_1), .B(new_n10111_1), .Y(new_n10159));
  nor_5  g07811(.A(new_n10159), .B(new_n10108), .Y(new_n10160));
  nor_5  g07812(.A(new_n10160), .B(new_n10107), .Y(new_n10161));
  nor_5  g07813(.A(new_n10161), .B(new_n10104), .Y(new_n10162));
  nor_5  g07814(.A(new_n10162), .B(new_n10103), .Y(new_n10163));
  xnor_4 g07815(.A(new_n10163), .B(new_n10100), .Y(n1332));
  not_8  g07816(.A(new_n5542), .Y(new_n10165_1));
  nor_5  g07817(.A(new_n5544), .B(n14692), .Y(new_n10166));
  not_8  g07818(.A(new_n5544), .Y(new_n10167));
  xnor_4 g07819(.A(new_n10167), .B(n14692), .Y(new_n10168));
  nor_5  g07820(.A(new_n5619), .B(n4100), .Y(new_n10169));
  not_8  g07821(.A(n4100), .Y(new_n10170));
  xnor_4 g07822(.A(new_n5620), .B(new_n10170), .Y(new_n10171));
  nor_5  g07823(.A(new_n5625), .B(n21957), .Y(new_n10172));
  not_8  g07824(.A(n21957), .Y(new_n10173));
  xnor_4 g07825(.A(new_n5626), .B(new_n10173), .Y(new_n10174));
  nor_5  g07826(.A(new_n5631), .B(n15761), .Y(new_n10175));
  not_8  g07827(.A(n15761), .Y(new_n10176));
  xnor_4 g07828(.A(new_n5632), .B(new_n10176), .Y(new_n10177));
  nor_5  g07829(.A(new_n5637), .B(n11201), .Y(new_n10178));
  not_8  g07830(.A(n11201), .Y(new_n10179));
  xnor_4 g07831(.A(new_n5638), .B(new_n10179), .Y(new_n10180));
  nor_5  g07832(.A(new_n5643_1), .B(n18690), .Y(new_n10181));
  not_8  g07833(.A(n18690), .Y(new_n10182));
  xnor_4 g07834(.A(new_n5644), .B(new_n10182), .Y(new_n10183));
  nor_5  g07835(.A(new_n5648), .B(n12153), .Y(new_n10184));
  xnor_4 g07836(.A(new_n5649), .B(n12153), .Y(new_n10185));
  not_8  g07837(.A(n13044), .Y(new_n10186));
  nor_5  g07838(.A(new_n5655), .B(new_n10186), .Y(new_n10187));
  nand_5 g07839(.A(new_n5655), .B(new_n10186), .Y(new_n10188));
  nor_5  g07840(.A(new_n5666), .B(n18745), .Y(new_n10189));
  and_5  g07841(.A(new_n5808), .B(new_n5806), .Y(new_n10190));
  nor_5  g07842(.A(new_n10190), .B(new_n10189), .Y(new_n10191));
  and_5  g07843(.A(new_n10191), .B(new_n10188), .Y(new_n10192));
  nor_5  g07844(.A(new_n10192), .B(new_n10187), .Y(new_n10193));
  and_5  g07845(.A(new_n10193), .B(new_n10185), .Y(new_n10194));
  nor_5  g07846(.A(new_n10194), .B(new_n10184), .Y(new_n10195));
  nor_5  g07847(.A(new_n10195), .B(new_n10183), .Y(new_n10196));
  nor_5  g07848(.A(new_n10196), .B(new_n10181), .Y(new_n10197));
  nor_5  g07849(.A(new_n10197), .B(new_n10180), .Y(new_n10198));
  nor_5  g07850(.A(new_n10198), .B(new_n10178), .Y(new_n10199));
  nor_5  g07851(.A(new_n10199), .B(new_n10177), .Y(new_n10200));
  nor_5  g07852(.A(new_n10200), .B(new_n10175), .Y(new_n10201_1));
  nor_5  g07853(.A(new_n10201_1), .B(new_n10174), .Y(new_n10202));
  nor_5  g07854(.A(new_n10202), .B(new_n10172), .Y(new_n10203));
  nor_5  g07855(.A(new_n10203), .B(new_n10171), .Y(new_n10204));
  or_5   g07856(.A(new_n10204), .B(new_n10169), .Y(new_n10205));
  and_5  g07857(.A(new_n10205), .B(new_n10168), .Y(new_n10206));
  nor_5  g07858(.A(new_n10206), .B(new_n10166), .Y(new_n10207));
  not_8  g07859(.A(new_n10207), .Y(new_n10208));
  nor_5  g07860(.A(new_n10208), .B(new_n10165_1), .Y(new_n10209));
  not_8  g07861(.A(new_n10209), .Y(new_n10210));
  not_8  g07862(.A(new_n5817), .Y(new_n10211));
  nor_5  g07863(.A(new_n10211), .B(n11302), .Y(new_n10212));
  not_8  g07864(.A(new_n10212), .Y(new_n10213));
  nor_5  g07865(.A(new_n10213), .B(n10405), .Y(new_n10214));
  not_8  g07866(.A(new_n10214), .Y(new_n10215));
  nor_5  g07867(.A(new_n10215), .B(n7693), .Y(new_n10216));
  not_8  g07868(.A(new_n10216), .Y(new_n10217));
  nor_5  g07869(.A(new_n10217), .B(n20151), .Y(new_n10218));
  not_8  g07870(.A(new_n10218), .Y(new_n10219));
  nor_5  g07871(.A(new_n10219), .B(n8964), .Y(new_n10220));
  not_8  g07872(.A(new_n10220), .Y(new_n10221));
  nor_5  g07873(.A(new_n10221), .B(n27037), .Y(new_n10222));
  and_5  g07874(.A(new_n10222), .B(new_n6215), .Y(new_n10223));
  and_5  g07875(.A(new_n10223), .B(new_n6198), .Y(new_n10224));
  nor_5  g07876(.A(n25926), .B(n7657), .Y(new_n10225));
  not_8  g07877(.A(new_n10225), .Y(new_n10226));
  nor_5  g07878(.A(new_n10226), .B(n5330), .Y(new_n10227));
  not_8  g07879(.A(new_n10227), .Y(new_n10228));
  nor_5  g07880(.A(new_n10228), .B(n5451), .Y(new_n10229));
  not_8  g07881(.A(new_n10229), .Y(new_n10230));
  nor_5  g07882(.A(new_n10230), .B(n18926), .Y(new_n10231));
  not_8  g07883(.A(new_n10231), .Y(new_n10232));
  nor_5  g07884(.A(new_n10232), .B(n13677), .Y(new_n10233));
  not_8  g07885(.A(new_n10233), .Y(new_n10234));
  nor_5  g07886(.A(new_n10234), .B(n23039), .Y(new_n10235));
  not_8  g07887(.A(new_n10235), .Y(new_n10236_1));
  nor_5  g07888(.A(new_n10236_1), .B(n7692), .Y(new_n10237));
  not_8  g07889(.A(new_n10237), .Y(new_n10238));
  nor_5  g07890(.A(new_n10238), .B(n25629), .Y(new_n10239_1));
  and_5  g07891(.A(new_n10239_1), .B(new_n6320), .Y(new_n10240));
  xnor_4 g07892(.A(new_n10239_1), .B(n15766), .Y(new_n10241));
  nor_5  g07893(.A(new_n10241), .B(n23895), .Y(new_n10242));
  xnor_4 g07894(.A(new_n10237), .B(n25629), .Y(new_n10243));
  nor_5  g07895(.A(new_n10243), .B(n17351), .Y(new_n10244_1));
  xnor_4 g07896(.A(new_n10243), .B(new_n5456), .Y(new_n10245));
  xnor_4 g07897(.A(new_n10235), .B(n7692), .Y(new_n10246));
  nor_5  g07898(.A(new_n10246), .B(n11736), .Y(new_n10247));
  xnor_4 g07899(.A(new_n10246), .B(new_n5459), .Y(new_n10248));
  xnor_4 g07900(.A(new_n10233), .B(n23039), .Y(new_n10249));
  nor_5  g07901(.A(new_n10249), .B(n23200), .Y(new_n10250_1));
  xnor_4 g07902(.A(new_n10249), .B(new_n5462), .Y(new_n10251));
  xnor_4 g07903(.A(new_n10231), .B(n13677), .Y(new_n10252));
  nor_5  g07904(.A(new_n10252), .B(n17959), .Y(new_n10253));
  xnor_4 g07905(.A(new_n10229), .B(n18926), .Y(new_n10254));
  nor_5  g07906(.A(new_n10254), .B(n7566), .Y(new_n10255));
  xnor_4 g07907(.A(new_n10254), .B(new_n5468), .Y(new_n10256));
  xnor_4 g07908(.A(new_n10227), .B(n5451), .Y(new_n10257));
  and_5  g07909(.A(new_n10257), .B(n7731), .Y(new_n10258));
  nor_5  g07910(.A(new_n10257), .B(n7731), .Y(new_n10259));
  xnor_4 g07911(.A(new_n10225), .B(n5330), .Y(new_n10260));
  and_5  g07912(.A(new_n10260), .B(n12341), .Y(new_n10261_1));
  xnor_4 g07913(.A(new_n10260), .B(new_n5475), .Y(new_n10262_1));
  nor_5  g07914(.A(new_n5811), .B(new_n5478), .Y(new_n10263));
  and_5  g07915(.A(new_n5812), .B(new_n5810), .Y(new_n10264));
  or_5   g07916(.A(new_n10264), .B(new_n10263), .Y(new_n10265));
  and_5  g07917(.A(new_n10265), .B(new_n10262_1), .Y(new_n10266));
  nor_5  g07918(.A(new_n10266), .B(new_n10261_1), .Y(new_n10267));
  nor_5  g07919(.A(new_n10267), .B(new_n10259), .Y(new_n10268));
  nor_5  g07920(.A(new_n10268), .B(new_n10258), .Y(new_n10269));
  and_5  g07921(.A(new_n10269), .B(new_n10256), .Y(new_n10270));
  or_5   g07922(.A(new_n10270), .B(new_n10255), .Y(new_n10271));
  xnor_4 g07923(.A(new_n10252), .B(new_n5465), .Y(new_n10272));
  and_5  g07924(.A(new_n10272), .B(new_n10271), .Y(new_n10273));
  or_5   g07925(.A(new_n10273), .B(new_n10253), .Y(new_n10274));
  and_5  g07926(.A(new_n10274), .B(new_n10251), .Y(new_n10275_1));
  or_5   g07927(.A(new_n10275_1), .B(new_n10250_1), .Y(new_n10276));
  and_5  g07928(.A(new_n10276), .B(new_n10248), .Y(new_n10277));
  or_5   g07929(.A(new_n10277), .B(new_n10247), .Y(new_n10278));
  and_5  g07930(.A(new_n10278), .B(new_n10245), .Y(new_n10279));
  nor_5  g07931(.A(new_n10279), .B(new_n10244_1), .Y(new_n10280));
  not_8  g07932(.A(new_n10241), .Y(new_n10281));
  nor_5  g07933(.A(new_n10281), .B(new_n5453), .Y(new_n10282));
  nor_5  g07934(.A(new_n10282), .B(new_n10280), .Y(new_n10283));
  nor_5  g07935(.A(new_n10283), .B(new_n10242), .Y(new_n10284));
  nor_5  g07936(.A(new_n10284), .B(new_n10240), .Y(new_n10285));
  nor_5  g07937(.A(new_n10285), .B(new_n10224), .Y(new_n10286));
  xnor_4 g07938(.A(new_n10223), .B(n8614), .Y(new_n10287_1));
  not_8  g07939(.A(new_n10287_1), .Y(new_n10288));
  xnor_4 g07940(.A(new_n10281), .B(n23895), .Y(new_n10289));
  xnor_4 g07941(.A(new_n10289), .B(new_n10280), .Y(new_n10290));
  nor_5  g07942(.A(new_n10290), .B(new_n10288), .Y(new_n10291));
  xnor_4 g07943(.A(new_n10222), .B(n15182), .Y(new_n10292));
  nor_5  g07944(.A(new_n10277), .B(new_n10247), .Y(new_n10293));
  xnor_4 g07945(.A(new_n10293), .B(new_n10245), .Y(new_n10294));
  not_8  g07946(.A(new_n10294), .Y(new_n10295_1));
  nor_5  g07947(.A(new_n10295_1), .B(new_n10292), .Y(new_n10296));
  xnor_4 g07948(.A(new_n10294), .B(new_n10292), .Y(new_n10297));
  xnor_4 g07949(.A(new_n10220), .B(n27037), .Y(new_n10298));
  xor_4  g07950(.A(new_n10276), .B(new_n10248), .Y(new_n10299));
  not_8  g07951(.A(new_n10299), .Y(new_n10300));
  nor_5  g07952(.A(new_n10300), .B(new_n10298), .Y(new_n10301));
  xnor_4 g07953(.A(new_n10300), .B(new_n10298), .Y(new_n10302));
  xnor_4 g07954(.A(new_n10218), .B(n8964), .Y(new_n10303));
  xor_4  g07955(.A(new_n10274), .B(new_n10251), .Y(new_n10304));
  not_8  g07956(.A(new_n10304), .Y(new_n10305));
  nor_5  g07957(.A(new_n10305), .B(new_n10303), .Y(new_n10306));
  xnor_4 g07958(.A(new_n10304), .B(new_n10303), .Y(new_n10307));
  xnor_4 g07959(.A(new_n10216), .B(n20151), .Y(new_n10308));
  xor_4  g07960(.A(new_n10272), .B(new_n10271), .Y(new_n10309));
  not_8  g07961(.A(new_n10309), .Y(new_n10310));
  nor_5  g07962(.A(new_n10310), .B(new_n10308), .Y(new_n10311));
  xnor_4 g07963(.A(new_n10310), .B(new_n10308), .Y(new_n10312));
  xnor_4 g07964(.A(new_n10214), .B(n7693), .Y(new_n10313));
  xnor_4 g07965(.A(new_n10269), .B(new_n10256), .Y(new_n10314));
  nor_5  g07966(.A(new_n10314), .B(new_n10313), .Y(new_n10315));
  xor_4  g07967(.A(new_n10314), .B(new_n10313), .Y(new_n10316));
  xnor_4 g07968(.A(new_n10212), .B(n10405), .Y(new_n10317));
  xnor_4 g07969(.A(new_n10257), .B(new_n5471), .Y(new_n10318));
  xnor_4 g07970(.A(new_n10318), .B(new_n10267), .Y(new_n10319));
  nor_5  g07971(.A(new_n10319), .B(new_n10317), .Y(new_n10320));
  xnor_4 g07972(.A(new_n10319), .B(new_n10317), .Y(new_n10321_1));
  xor_4  g07973(.A(new_n10265), .B(new_n10262_1), .Y(new_n10322));
  xnor_4 g07974(.A(new_n5817), .B(n11302), .Y(new_n10323));
  nor_5  g07975(.A(new_n10323), .B(new_n10322), .Y(new_n10324));
  xnor_4 g07976(.A(new_n10323), .B(new_n10322), .Y(new_n10325));
  and_5  g07977(.A(new_n5821), .B(new_n5813), .Y(new_n10326_1));
  nor_5  g07978(.A(new_n10326_1), .B(new_n5820), .Y(new_n10327_1));
  nor_5  g07979(.A(new_n10327_1), .B(new_n10325), .Y(new_n10328));
  nor_5  g07980(.A(new_n10328), .B(new_n10324), .Y(new_n10329));
  nor_5  g07981(.A(new_n10329), .B(new_n10321_1), .Y(new_n10330_1));
  or_5   g07982(.A(new_n10330_1), .B(new_n10320), .Y(new_n10331));
  and_5  g07983(.A(new_n10331), .B(new_n10316), .Y(new_n10332));
  nor_5  g07984(.A(new_n10332), .B(new_n10315), .Y(new_n10333));
  nor_5  g07985(.A(new_n10333), .B(new_n10312), .Y(new_n10334));
  or_5   g07986(.A(new_n10334), .B(new_n10311), .Y(new_n10335));
  and_5  g07987(.A(new_n10335), .B(new_n10307), .Y(new_n10336));
  nor_5  g07988(.A(new_n10336), .B(new_n10306), .Y(new_n10337));
  nor_5  g07989(.A(new_n10337), .B(new_n10302), .Y(new_n10338));
  or_5   g07990(.A(new_n10338), .B(new_n10301), .Y(new_n10339));
  and_5  g07991(.A(new_n10339), .B(new_n10297), .Y(new_n10340_1));
  nor_5  g07992(.A(new_n10340_1), .B(new_n10296), .Y(new_n10341));
  not_8  g07993(.A(new_n10290), .Y(new_n10342));
  xnor_4 g07994(.A(new_n10342), .B(new_n10288), .Y(new_n10343));
  and_5  g07995(.A(new_n10343), .B(new_n10341), .Y(new_n10344));
  nor_5  g07996(.A(new_n10344), .B(new_n10291), .Y(new_n10345_1));
  and_5  g07997(.A(new_n10345_1), .B(new_n10286), .Y(new_n10346));
  xnor_4 g07998(.A(new_n10346), .B(new_n10210), .Y(new_n10347));
  xnor_4 g07999(.A(new_n10208), .B(new_n5542), .Y(new_n10348));
  xnor_4 g08000(.A(new_n10285), .B(new_n10224), .Y(new_n10349));
  xnor_4 g08001(.A(new_n10349), .B(new_n10345_1), .Y(new_n10350));
  nor_5  g08002(.A(new_n10350), .B(new_n10348), .Y(new_n10351));
  not_8  g08003(.A(new_n10348), .Y(new_n10352));
  xnor_4 g08004(.A(new_n10350), .B(new_n10352), .Y(new_n10353));
  xor_4  g08005(.A(new_n10205), .B(new_n10168), .Y(new_n10354));
  xnor_4 g08006(.A(new_n10343), .B(new_n10341), .Y(new_n10355));
  nor_5  g08007(.A(new_n10355), .B(new_n10354), .Y(new_n10356_1));
  xor_4  g08008(.A(new_n10355), .B(new_n10354), .Y(new_n10357));
  xnor_4 g08009(.A(new_n10339), .B(new_n10297), .Y(new_n10358));
  xnor_4 g08010(.A(new_n10203), .B(new_n10171), .Y(new_n10359));
  and_5  g08011(.A(new_n10359), .B(new_n10358), .Y(new_n10360));
  xnor_4 g08012(.A(new_n10337), .B(new_n10302), .Y(new_n10361));
  xnor_4 g08013(.A(new_n10201_1), .B(new_n10174), .Y(new_n10362));
  nor_5  g08014(.A(new_n10362), .B(new_n10361), .Y(new_n10363));
  xnor_4 g08015(.A(new_n10362), .B(new_n10361), .Y(new_n10364));
  not_8  g08016(.A(new_n10364), .Y(new_n10365));
  xnor_4 g08017(.A(new_n10335), .B(new_n10307), .Y(new_n10366));
  xnor_4 g08018(.A(new_n10199), .B(new_n10177), .Y(new_n10367));
  and_5  g08019(.A(new_n10367), .B(new_n10366), .Y(new_n10368));
  xnor_4 g08020(.A(new_n10333), .B(new_n10312), .Y(new_n10369));
  xnor_4 g08021(.A(new_n10197), .B(new_n10180), .Y(new_n10370));
  nor_5  g08022(.A(new_n10370), .B(new_n10369), .Y(new_n10371));
  xnor_4 g08023(.A(new_n10370), .B(new_n10369), .Y(new_n10372_1));
  not_8  g08024(.A(new_n10372_1), .Y(new_n10373));
  xnor_4 g08025(.A(new_n10331), .B(new_n10316), .Y(new_n10374));
  xnor_4 g08026(.A(new_n10195), .B(new_n10183), .Y(new_n10375));
  and_5  g08027(.A(new_n10375), .B(new_n10374), .Y(new_n10376));
  xor_4  g08028(.A(new_n10375), .B(new_n10374), .Y(new_n10377));
  xnor_4 g08029(.A(new_n10329), .B(new_n10321_1), .Y(new_n10378));
  xnor_4 g08030(.A(new_n10193), .B(new_n10185), .Y(new_n10379));
  nor_5  g08031(.A(new_n10379), .B(new_n10378), .Y(new_n10380));
  xnor_4 g08032(.A(new_n10379), .B(new_n10378), .Y(new_n10381));
  xnor_4 g08033(.A(new_n10327_1), .B(new_n10325), .Y(new_n10382));
  xnor_4 g08034(.A(new_n5655), .B(new_n10186), .Y(new_n10383));
  xnor_4 g08035(.A(new_n10383), .B(new_n10191), .Y(new_n10384));
  nor_5  g08036(.A(new_n10384), .B(new_n10382), .Y(new_n10385_1));
  and_5  g08037(.A(new_n5822_1), .B(new_n5809), .Y(new_n10386));
  nor_5  g08038(.A(new_n5823), .B(new_n5804), .Y(new_n10387_1));
  nor_5  g08039(.A(new_n10387_1), .B(new_n10386), .Y(new_n10388_1));
  xnor_4 g08040(.A(new_n10384), .B(new_n10382), .Y(new_n10389));
  nor_5  g08041(.A(new_n10389), .B(new_n10388_1), .Y(new_n10390_1));
  nor_5  g08042(.A(new_n10390_1), .B(new_n10385_1), .Y(new_n10391));
  nor_5  g08043(.A(new_n10391), .B(new_n10381), .Y(new_n10392));
  nor_5  g08044(.A(new_n10392), .B(new_n10380), .Y(new_n10393));
  and_5  g08045(.A(new_n10393), .B(new_n10377), .Y(new_n10394));
  nor_5  g08046(.A(new_n10394), .B(new_n10376), .Y(new_n10395));
  and_5  g08047(.A(new_n10395), .B(new_n10373), .Y(new_n10396));
  nor_5  g08048(.A(new_n10396), .B(new_n10371), .Y(new_n10397));
  xor_4  g08049(.A(new_n10367), .B(new_n10366), .Y(new_n10398));
  and_5  g08050(.A(new_n10398), .B(new_n10397), .Y(new_n10399));
  nor_5  g08051(.A(new_n10399), .B(new_n10368), .Y(new_n10400));
  and_5  g08052(.A(new_n10400), .B(new_n10365), .Y(new_n10401));
  nor_5  g08053(.A(new_n10401), .B(new_n10363), .Y(new_n10402));
  xor_4  g08054(.A(new_n10359), .B(new_n10358), .Y(new_n10403));
  and_5  g08055(.A(new_n10403), .B(new_n10402), .Y(new_n10404_1));
  or_5   g08056(.A(new_n10404_1), .B(new_n10360), .Y(new_n10405_1));
  and_5  g08057(.A(new_n10405_1), .B(new_n10357), .Y(new_n10406));
  nor_5  g08058(.A(new_n10406), .B(new_n10356_1), .Y(new_n10407));
  and_5  g08059(.A(new_n10407), .B(new_n10353), .Y(new_n10408));
  nor_5  g08060(.A(new_n10408), .B(new_n10351), .Y(new_n10409_1));
  not_8  g08061(.A(new_n10409_1), .Y(new_n10410));
  xnor_4 g08062(.A(new_n10410), .B(new_n10347), .Y(n1357));
  xnor_4 g08063(.A(new_n7971), .B(n25240), .Y(new_n10412));
  nor_5  g08064(.A(new_n7976), .B(n10125), .Y(new_n10413));
  not_8  g08065(.A(n10125), .Y(new_n10414));
  xnor_4 g08066(.A(new_n7976), .B(new_n10414), .Y(new_n10415));
  nor_5  g08067(.A(new_n7981), .B(n8067), .Y(new_n10416));
  xnor_4 g08068(.A(new_n7981), .B(n8067), .Y(new_n10417));
  nor_5  g08069(.A(new_n7986), .B(n20923), .Y(new_n10418));
  xnor_4 g08070(.A(new_n7986), .B(n20923), .Y(new_n10419));
  nor_5  g08071(.A(new_n7991), .B(n18157), .Y(new_n10420_1));
  or_5   g08072(.A(new_n8441), .B(new_n8434), .Y(new_n10421));
  and_5  g08073(.A(new_n10421), .B(new_n8433), .Y(new_n10422));
  nor_5  g08074(.A(new_n10422), .B(new_n10420_1), .Y(new_n10423));
  nor_5  g08075(.A(new_n10423), .B(new_n10419), .Y(new_n10424));
  nor_5  g08076(.A(new_n10424), .B(new_n10418), .Y(new_n10425));
  nor_5  g08077(.A(new_n10425), .B(new_n10417), .Y(new_n10426));
  or_5   g08078(.A(new_n10426), .B(new_n10416), .Y(new_n10427));
  and_5  g08079(.A(new_n10427), .B(new_n10415), .Y(new_n10428));
  nor_5  g08080(.A(new_n10428), .B(new_n10413), .Y(new_n10429));
  xnor_4 g08081(.A(new_n10429), .B(new_n10412), .Y(new_n10430));
  not_8  g08082(.A(n5077), .Y(new_n10431));
  xnor_4 g08083(.A(n6381), .B(n1099), .Y(new_n10432_1));
  nor_5  g08084(.A(n14345), .B(n2113), .Y(new_n10433));
  not_8  g08085(.A(n2113), .Y(new_n10434));
  xnor_4 g08086(.A(n14345), .B(new_n10434), .Y(new_n10435));
  nor_5  g08087(.A(n21134), .B(n11356), .Y(new_n10436));
  xnor_4 g08088(.A(n21134), .B(new_n9088), .Y(new_n10437));
  nor_5  g08089(.A(new_n4165_1), .B(new_n9091), .Y(new_n10438));
  or_5   g08090(.A(n6369), .B(n3164), .Y(new_n10439));
  nor_5  g08091(.A(n25797), .B(n10611), .Y(new_n10440));
  or_5   g08092(.A(new_n6601), .B(new_n6592), .Y(new_n10441));
  and_5  g08093(.A(new_n10441), .B(new_n6591), .Y(new_n10442));
  nor_5  g08094(.A(new_n10442), .B(new_n10440), .Y(new_n10443));
  and_5  g08095(.A(new_n10443), .B(new_n10439), .Y(new_n10444));
  nor_5  g08096(.A(new_n10444), .B(new_n10438), .Y(new_n10445));
  and_5  g08097(.A(new_n10445), .B(new_n10437), .Y(new_n10446));
  or_5   g08098(.A(new_n10446), .B(new_n10436), .Y(new_n10447));
  and_5  g08099(.A(new_n10447), .B(new_n10435), .Y(new_n10448));
  nor_5  g08100(.A(new_n10448), .B(new_n10433), .Y(new_n10449));
  xnor_4 g08101(.A(new_n10449), .B(new_n10432_1), .Y(new_n10450));
  xnor_4 g08102(.A(new_n10450), .B(new_n10431), .Y(new_n10451));
  not_8  g08103(.A(n15546), .Y(new_n10452));
  nor_5  g08104(.A(new_n10446), .B(new_n10436), .Y(new_n10453));
  xnor_4 g08105(.A(new_n10453), .B(new_n10435), .Y(new_n10454));
  nor_5  g08106(.A(new_n10454), .B(new_n10452), .Y(new_n10455));
  not_8  g08107(.A(new_n10454), .Y(new_n10456));
  xnor_4 g08108(.A(new_n10456), .B(new_n10452), .Y(new_n10457));
  xnor_4 g08109(.A(new_n10445), .B(new_n10437), .Y(new_n10458));
  nor_5  g08110(.A(new_n10458), .B(n26452), .Y(new_n10459));
  not_8  g08111(.A(n19905), .Y(new_n10460));
  xnor_4 g08112(.A(n6369), .B(new_n9091), .Y(new_n10461));
  xnor_4 g08113(.A(new_n10461), .B(new_n10443), .Y(new_n10462));
  nor_5  g08114(.A(new_n10462), .B(new_n10460), .Y(new_n10463));
  not_8  g08115(.A(new_n10462), .Y(new_n10464));
  xnor_4 g08116(.A(new_n10464), .B(new_n10460), .Y(new_n10465));
  nor_5  g08117(.A(new_n6603), .B(new_n8469), .Y(new_n10466));
  and_5  g08118(.A(new_n8473), .B(new_n8470), .Y(new_n10467));
  or_5   g08119(.A(new_n10467), .B(new_n10466), .Y(new_n10468));
  and_5  g08120(.A(new_n10468), .B(new_n10465), .Y(new_n10469));
  nor_5  g08121(.A(new_n10469), .B(new_n10463), .Y(new_n10470));
  not_8  g08122(.A(new_n10458), .Y(new_n10471));
  xnor_4 g08123(.A(new_n10471), .B(n26452), .Y(new_n10472));
  and_5  g08124(.A(new_n10472), .B(new_n10470), .Y(new_n10473));
  nor_5  g08125(.A(new_n10473), .B(new_n10459), .Y(new_n10474));
  and_5  g08126(.A(new_n10474), .B(new_n10457), .Y(new_n10475));
  nor_5  g08127(.A(new_n10475), .B(new_n10455), .Y(new_n10476));
  xor_4  g08128(.A(new_n10476), .B(new_n10451), .Y(new_n10477));
  xnor_4 g08129(.A(new_n10477), .B(new_n10430), .Y(new_n10478));
  xor_4  g08130(.A(new_n10427), .B(new_n10415), .Y(new_n10479));
  xnor_4 g08131(.A(new_n10474), .B(new_n10457), .Y(new_n10480));
  not_8  g08132(.A(new_n10480), .Y(new_n10481));
  and_5  g08133(.A(new_n10481), .B(new_n10479), .Y(new_n10482));
  xnor_4 g08134(.A(new_n10481), .B(new_n10479), .Y(new_n10483));
  xnor_4 g08135(.A(new_n10425), .B(new_n10417), .Y(new_n10484_1));
  xor_4  g08136(.A(new_n10472), .B(new_n10470), .Y(new_n10485));
  nor_5  g08137(.A(new_n10485), .B(new_n10484_1), .Y(new_n10486));
  xnor_4 g08138(.A(new_n10485), .B(new_n10484_1), .Y(new_n10487));
  xnor_4 g08139(.A(new_n10423), .B(new_n10419), .Y(new_n10488));
  nor_5  g08140(.A(new_n10467), .B(new_n10466), .Y(new_n10489_1));
  xnor_4 g08141(.A(new_n10489_1), .B(new_n10465), .Y(new_n10490));
  not_8  g08142(.A(new_n10490), .Y(new_n10491));
  nor_5  g08143(.A(new_n10491), .B(new_n10488), .Y(new_n10492));
  xnor_4 g08144(.A(new_n10490), .B(new_n10488), .Y(new_n10493));
  not_8  g08145(.A(new_n8467), .Y(new_n10494));
  nor_5  g08146(.A(new_n10494), .B(new_n8443), .Y(new_n10495));
  and_5  g08147(.A(new_n8474), .B(new_n8468), .Y(new_n10496));
  nor_5  g08148(.A(new_n10496), .B(new_n10495), .Y(new_n10497));
  and_5  g08149(.A(new_n10497), .B(new_n10493), .Y(new_n10498));
  nor_5  g08150(.A(new_n10498), .B(new_n10492), .Y(new_n10499));
  nor_5  g08151(.A(new_n10499), .B(new_n10487), .Y(new_n10500));
  nor_5  g08152(.A(new_n10500), .B(new_n10486), .Y(new_n10501));
  nor_5  g08153(.A(new_n10501), .B(new_n10483), .Y(new_n10502));
  nor_5  g08154(.A(new_n10502), .B(new_n10482), .Y(new_n10503));
  xnor_4 g08155(.A(new_n10503), .B(new_n10478), .Y(n1371));
  xnor_4 g08156(.A(n17250), .B(n15241), .Y(new_n10505));
  not_8  g08157(.A(n23160), .Y(new_n10506));
  nor_5  g08158(.A(new_n10506), .B(n7678), .Y(new_n10507));
  and_5  g08159(.A(n16524), .B(new_n4377), .Y(new_n10508));
  xnor_4 g08160(.A(n16524), .B(n3785), .Y(new_n10509));
  nor_5  g08161(.A(new_n4382), .B(n11056), .Y(new_n10510));
  nor_5  g08162(.A(n15271), .B(new_n4384), .Y(new_n10511));
  xnor_4 g08163(.A(n15271), .B(n5822), .Y(new_n10512));
  nor_5  g08164(.A(new_n6644), .B(n25877), .Y(new_n10513));
  and_5  g08165(.A(new_n5778), .B(new_n5777), .Y(new_n10514_1));
  or_5   g08166(.A(new_n10514_1), .B(new_n10513), .Y(new_n10515));
  and_5  g08167(.A(new_n10515), .B(new_n10512), .Y(new_n10516));
  or_5   g08168(.A(new_n10516), .B(new_n10511), .Y(new_n10517));
  xnor_4 g08169(.A(n20250), .B(n11056), .Y(new_n10518));
  and_5  g08170(.A(new_n10518), .B(new_n10517), .Y(new_n10519));
  nor_5  g08171(.A(new_n10519), .B(new_n10510), .Y(new_n10520));
  and_5  g08172(.A(new_n10520), .B(new_n10509), .Y(new_n10521));
  or_5   g08173(.A(new_n10521), .B(new_n10508), .Y(new_n10522));
  xnor_4 g08174(.A(n23160), .B(n7678), .Y(new_n10523));
  and_5  g08175(.A(new_n10523), .B(new_n10522), .Y(new_n10524));
  or_5   g08176(.A(new_n10524), .B(new_n10507), .Y(new_n10525_1));
  xor_4  g08177(.A(new_n10525_1), .B(new_n10505), .Y(new_n10526));
  xnor_4 g08178(.A(new_n9617), .B(new_n2425), .Y(new_n10527));
  not_8  g08179(.A(new_n10527), .Y(new_n10528));
  nor_5  g08180(.A(new_n9620), .B(n26660), .Y(new_n10529));
  xnor_4 g08181(.A(new_n9620), .B(new_n7618), .Y(new_n10530));
  and_5  g08182(.A(new_n9623), .B(n3018), .Y(new_n10531));
  nor_5  g08183(.A(new_n9623), .B(n3018), .Y(new_n10532));
  and_5  g08184(.A(new_n9413), .B(n3480), .Y(new_n10533));
  not_8  g08185(.A(new_n9414), .Y(new_n10534));
  nor_5  g08186(.A(new_n9422), .B(new_n10534), .Y(new_n10535));
  nor_5  g08187(.A(new_n10535), .B(new_n10533), .Y(new_n10536));
  nor_5  g08188(.A(new_n10536), .B(new_n10532), .Y(new_n10537));
  nor_5  g08189(.A(new_n10537), .B(new_n10531), .Y(new_n10538));
  and_5  g08190(.A(new_n10538), .B(new_n10530), .Y(new_n10539));
  nor_5  g08191(.A(new_n10539), .B(new_n10529), .Y(new_n10540_1));
  xnor_4 g08192(.A(new_n10540_1), .B(new_n10528), .Y(new_n10541));
  xnor_4 g08193(.A(new_n10541), .B(new_n10526), .Y(new_n10542));
  xnor_4 g08194(.A(new_n10538), .B(new_n10530), .Y(new_n10543));
  xor_4  g08195(.A(new_n10523), .B(new_n10522), .Y(new_n10544));
  and_5  g08196(.A(new_n10544), .B(new_n10543), .Y(new_n10545));
  not_8  g08197(.A(new_n10543), .Y(new_n10546));
  xnor_4 g08198(.A(new_n10544), .B(new_n10546), .Y(new_n10547));
  xnor_4 g08199(.A(new_n10520), .B(new_n10509), .Y(new_n10548));
  not_8  g08200(.A(new_n10548), .Y(new_n10549));
  not_8  g08201(.A(n3018), .Y(new_n10550));
  xnor_4 g08202(.A(new_n9623), .B(new_n10550), .Y(new_n10551));
  xnor_4 g08203(.A(new_n10551), .B(new_n10536), .Y(new_n10552));
  nor_5  g08204(.A(new_n10552), .B(new_n10549), .Y(new_n10553));
  not_8  g08205(.A(new_n10552), .Y(new_n10554));
  xnor_4 g08206(.A(new_n10554), .B(new_n10548), .Y(new_n10555));
  nor_5  g08207(.A(new_n10516), .B(new_n10511), .Y(new_n10556));
  xnor_4 g08208(.A(new_n10518), .B(new_n10556), .Y(new_n10557));
  not_8  g08209(.A(new_n10557), .Y(new_n10558));
  nor_5  g08210(.A(new_n10558), .B(new_n9423_1), .Y(new_n10559));
  xnor_4 g08211(.A(new_n10557), .B(new_n9423_1), .Y(new_n10560));
  xor_4  g08212(.A(new_n10515), .B(new_n10512), .Y(new_n10561_1));
  nor_5  g08213(.A(new_n10561_1), .B(new_n9425), .Y(new_n10562));
  xnor_4 g08214(.A(new_n10561_1), .B(new_n9425), .Y(new_n10563));
  and_5  g08215(.A(new_n5779), .B(new_n5776_1), .Y(new_n10564_1));
  nor_5  g08216(.A(new_n5788), .B(new_n5780), .Y(new_n10565));
  nor_5  g08217(.A(new_n10565), .B(new_n10564_1), .Y(new_n10566));
  nor_5  g08218(.A(new_n10566), .B(new_n10563), .Y(new_n10567));
  nor_5  g08219(.A(new_n10567), .B(new_n10562), .Y(new_n10568));
  and_5  g08220(.A(new_n10568), .B(new_n10560), .Y(new_n10569));
  nor_5  g08221(.A(new_n10569), .B(new_n10559), .Y(new_n10570));
  nor_5  g08222(.A(new_n10570), .B(new_n10555), .Y(new_n10571));
  nor_5  g08223(.A(new_n10571), .B(new_n10553), .Y(new_n10572));
  and_5  g08224(.A(new_n10572), .B(new_n10547), .Y(new_n10573));
  nor_5  g08225(.A(new_n10573), .B(new_n10545), .Y(new_n10574));
  xnor_4 g08226(.A(new_n10574), .B(new_n10542), .Y(new_n10575));
  not_8  g08227(.A(new_n10575), .Y(new_n10576));
  xnor_4 g08228(.A(new_n10576), .B(new_n5632), .Y(new_n10577_1));
  xor_4  g08229(.A(new_n10572), .B(new_n10547), .Y(new_n10578));
  nor_5  g08230(.A(new_n10578), .B(new_n5637), .Y(new_n10579));
  xnor_4 g08231(.A(new_n10578), .B(new_n5637), .Y(new_n10580));
  not_8  g08232(.A(new_n10580), .Y(new_n10581));
  xor_4  g08233(.A(new_n10570), .B(new_n10555), .Y(new_n10582));
  nor_5  g08234(.A(new_n10582), .B(new_n5644), .Y(new_n10583));
  xnor_4 g08235(.A(new_n10568), .B(new_n10560), .Y(new_n10584));
  nor_5  g08236(.A(new_n10584), .B(new_n5648), .Y(new_n10585));
  xnor_4 g08237(.A(new_n10584), .B(new_n5648), .Y(new_n10586));
  not_8  g08238(.A(new_n10586), .Y(new_n10587));
  xor_4  g08239(.A(new_n10566), .B(new_n10563), .Y(new_n10588_1));
  not_8  g08240(.A(new_n10588_1), .Y(new_n10589));
  nor_5  g08241(.A(new_n10589), .B(new_n5655), .Y(new_n10590));
  and_5  g08242(.A(new_n5773), .B(new_n5666), .Y(new_n10591));
  not_8  g08243(.A(new_n5790), .Y(new_n10592));
  nor_5  g08244(.A(new_n10592), .B(new_n5774), .Y(new_n10593_1));
  nor_5  g08245(.A(new_n10593_1), .B(new_n10591), .Y(new_n10594));
  xnor_4 g08246(.A(new_n10589), .B(new_n5655), .Y(new_n10595_1));
  nor_5  g08247(.A(new_n10595_1), .B(new_n10594), .Y(new_n10596));
  nor_5  g08248(.A(new_n10596), .B(new_n10590), .Y(new_n10597));
  and_5  g08249(.A(new_n10597), .B(new_n10587), .Y(new_n10598));
  nor_5  g08250(.A(new_n10598), .B(new_n10585), .Y(new_n10599));
  not_8  g08251(.A(new_n10582), .Y(new_n10600));
  xnor_4 g08252(.A(new_n10600), .B(new_n5644), .Y(new_n10601));
  and_5  g08253(.A(new_n10601), .B(new_n10599), .Y(new_n10602));
  nor_5  g08254(.A(new_n10602), .B(new_n10583), .Y(new_n10603));
  and_5  g08255(.A(new_n10603), .B(new_n10581), .Y(new_n10604));
  nor_5  g08256(.A(new_n10604), .B(new_n10579), .Y(new_n10605));
  xor_4  g08257(.A(new_n10605), .B(new_n10577_1), .Y(n1385));
  xnor_4 g08258(.A(n26808), .B(n24732), .Y(new_n10607));
  not_8  g08259(.A(new_n10607), .Y(new_n10608));
  nor_5  g08260(.A(new_n9155), .B(new_n4183), .Y(new_n10609));
  xnor_4 g08261(.A(n7339), .B(n6631), .Y(new_n10610));
  xnor_4 g08262(.A(new_n10610), .B(new_n10609), .Y(new_n10611_1));
  nor_5  g08263(.A(new_n10611_1), .B(new_n10608), .Y(new_n10612));
  not_8  g08264(.A(new_n10612), .Y(new_n10613));
  not_8  g08265(.A(n1667), .Y(new_n10614_1));
  xnor_4 g08266(.A(n14684), .B(new_n10614_1), .Y(new_n10615));
  nor_5  g08267(.A(n7339), .B(n6631), .Y(new_n10616));
  nor_5  g08268(.A(new_n10610), .B(new_n10609), .Y(new_n10617_1));
  nor_5  g08269(.A(new_n10617_1), .B(new_n10616), .Y(new_n10618));
  xnor_4 g08270(.A(new_n10618), .B(new_n10615), .Y(new_n10619));
  not_8  g08271(.A(new_n10619), .Y(new_n10620));
  nor_5  g08272(.A(new_n10620), .B(new_n10613), .Y(new_n10621));
  not_8  g08273(.A(new_n10621), .Y(new_n10622));
  not_8  g08274(.A(n2680), .Y(new_n10623));
  xnor_4 g08275(.A(n17035), .B(new_n10623), .Y(new_n10624));
  nor_5  g08276(.A(n14684), .B(n1667), .Y(new_n10625));
  or_5   g08277(.A(new_n10617_1), .B(new_n10616), .Y(new_n10626));
  and_5  g08278(.A(new_n10626), .B(new_n10615), .Y(new_n10627));
  nor_5  g08279(.A(new_n10627), .B(new_n10625), .Y(new_n10628_1));
  xnor_4 g08280(.A(new_n10628_1), .B(new_n10624), .Y(new_n10629));
  not_8  g08281(.A(new_n10629), .Y(new_n10630));
  nor_5  g08282(.A(new_n10630), .B(new_n10622), .Y(new_n10631));
  not_8  g08283(.A(new_n10631), .Y(new_n10632));
  not_8  g08284(.A(n2547), .Y(new_n10633));
  xnor_4 g08285(.A(n19905), .B(new_n10633), .Y(new_n10634));
  nor_5  g08286(.A(n17035), .B(n2680), .Y(new_n10635));
  or_5   g08287(.A(new_n10627), .B(new_n10625), .Y(new_n10636));
  and_5  g08288(.A(new_n10636), .B(new_n10624), .Y(new_n10637));
  nor_5  g08289(.A(new_n10637), .B(new_n10635), .Y(new_n10638));
  xnor_4 g08290(.A(new_n10638), .B(new_n10634), .Y(new_n10639));
  not_8  g08291(.A(new_n10639), .Y(new_n10640));
  nor_5  g08292(.A(new_n10640), .B(new_n10632), .Y(new_n10641));
  not_8  g08293(.A(new_n10641), .Y(new_n10642));
  not_8  g08294(.A(n2999), .Y(new_n10643));
  xnor_4 g08295(.A(n26452), .B(new_n10643), .Y(new_n10644));
  nor_5  g08296(.A(n19905), .B(n2547), .Y(new_n10645));
  not_8  g08297(.A(new_n10634), .Y(new_n10646));
  nor_5  g08298(.A(new_n10638), .B(new_n10646), .Y(new_n10647_1));
  nor_5  g08299(.A(new_n10647_1), .B(new_n10645), .Y(new_n10648));
  xnor_4 g08300(.A(new_n10648), .B(new_n10644), .Y(new_n10649));
  not_8  g08301(.A(new_n10649), .Y(new_n10650_1));
  nor_5  g08302(.A(new_n10650_1), .B(new_n10642), .Y(new_n10651));
  not_8  g08303(.A(new_n10651), .Y(new_n10652));
  xnor_4 g08304(.A(new_n10452), .B(n14702), .Y(new_n10653_1));
  nor_5  g08305(.A(n26452), .B(n2999), .Y(new_n10654));
  not_8  g08306(.A(new_n10644), .Y(new_n10655));
  nor_5  g08307(.A(new_n10648), .B(new_n10655), .Y(new_n10656));
  nor_5  g08308(.A(new_n10656), .B(new_n10654), .Y(new_n10657));
  xnor_4 g08309(.A(new_n10657), .B(new_n10653_1), .Y(new_n10658));
  not_8  g08310(.A(new_n10658), .Y(new_n10659));
  nor_5  g08311(.A(new_n10659), .B(new_n10652), .Y(new_n10660));
  not_8  g08312(.A(new_n10660), .Y(new_n10661));
  xnor_4 g08313(.A(n13914), .B(new_n10431), .Y(new_n10662));
  nor_5  g08314(.A(n15546), .B(n14702), .Y(new_n10663));
  not_8  g08315(.A(new_n10653_1), .Y(new_n10664));
  nor_5  g08316(.A(new_n10657), .B(new_n10664), .Y(new_n10665));
  nor_5  g08317(.A(new_n10665), .B(new_n10663), .Y(new_n10666));
  xnor_4 g08318(.A(new_n10666), .B(new_n10662), .Y(new_n10667));
  not_8  g08319(.A(new_n10667), .Y(new_n10668));
  nor_5  g08320(.A(new_n10668), .B(new_n10661), .Y(new_n10669));
  not_8  g08321(.A(new_n10669), .Y(new_n10670));
  xnor_4 g08322(.A(n18035), .B(new_n9062), .Y(new_n10671));
  nor_5  g08323(.A(n13914), .B(n5077), .Y(new_n10672));
  not_8  g08324(.A(new_n10662), .Y(new_n10673));
  nor_5  g08325(.A(new_n10666), .B(new_n10673), .Y(new_n10674));
  nor_5  g08326(.A(new_n10674), .B(new_n10672), .Y(new_n10675));
  xnor_4 g08327(.A(new_n10675), .B(new_n10671), .Y(new_n10676));
  not_8  g08328(.A(new_n10676), .Y(new_n10677));
  nor_5  g08329(.A(new_n10677), .B(new_n10670), .Y(new_n10678));
  not_8  g08330(.A(n4306), .Y(new_n10679));
  xnor_4 g08331(.A(n8827), .B(new_n10679), .Y(new_n10680));
  nor_5  g08332(.A(n18035), .B(n3279), .Y(new_n10681));
  not_8  g08333(.A(new_n10671), .Y(new_n10682));
  nor_5  g08334(.A(new_n10675), .B(new_n10682), .Y(new_n10683));
  nor_5  g08335(.A(new_n10683), .B(new_n10681), .Y(new_n10684));
  xnor_4 g08336(.A(new_n10684), .B(new_n10680), .Y(new_n10685));
  xor_4  g08337(.A(new_n10685), .B(new_n10678), .Y(new_n10686));
  xnor_4 g08338(.A(new_n10686), .B(new_n7959_1), .Y(new_n10687));
  xnor_4 g08339(.A(new_n10677), .B(new_n10669), .Y(new_n10688));
  nor_5  g08340(.A(new_n10688), .B(new_n7966), .Y(new_n10689));
  xnor_4 g08341(.A(new_n10688), .B(new_n7964), .Y(new_n10690));
  xnor_4 g08342(.A(new_n10668), .B(new_n10660), .Y(new_n10691));
  nor_5  g08343(.A(new_n10691), .B(new_n7971), .Y(new_n10692_1));
  xnor_4 g08344(.A(new_n10691), .B(new_n7969), .Y(new_n10693));
  xnor_4 g08345(.A(new_n10659), .B(new_n10651), .Y(new_n10694_1));
  nor_5  g08346(.A(new_n10694_1), .B(new_n7976), .Y(new_n10695));
  xnor_4 g08347(.A(new_n10694_1), .B(new_n7974), .Y(new_n10696));
  xnor_4 g08348(.A(new_n10650_1), .B(new_n10641), .Y(new_n10697));
  nor_5  g08349(.A(new_n10697), .B(new_n7981), .Y(new_n10698));
  xnor_4 g08350(.A(new_n10697), .B(new_n7979), .Y(new_n10699));
  xnor_4 g08351(.A(new_n10640), .B(new_n10631), .Y(new_n10700));
  nor_5  g08352(.A(new_n10700), .B(new_n7986), .Y(new_n10701_1));
  xnor_4 g08353(.A(new_n10700), .B(new_n7984), .Y(new_n10702));
  xnor_4 g08354(.A(new_n10630), .B(new_n10621), .Y(new_n10703));
  nor_5  g08355(.A(new_n10703), .B(new_n7991), .Y(new_n10704));
  xnor_4 g08356(.A(new_n10703), .B(new_n7991), .Y(new_n10705));
  xnor_4 g08357(.A(new_n10620), .B(new_n10612), .Y(new_n10706));
  nor_5  g08358(.A(new_n10706), .B(new_n7995), .Y(new_n10707));
  xnor_4 g08359(.A(new_n10706), .B(new_n7995), .Y(new_n10708));
  nor_5  g08360(.A(new_n10607), .B(new_n2543), .Y(new_n10709));
  nor_5  g08361(.A(new_n10709), .B(new_n8003), .Y(new_n10710_1));
  nor_5  g08362(.A(new_n10610), .B(new_n10607), .Y(new_n10711));
  or_5   g08363(.A(new_n10711), .B(new_n10612), .Y(new_n10712_1));
  and_5  g08364(.A(new_n10709), .B(new_n7942), .Y(new_n10713));
  nor_5  g08365(.A(new_n10713), .B(new_n10710_1), .Y(new_n10714));
  and_5  g08366(.A(new_n10714), .B(new_n10712_1), .Y(new_n10715));
  nor_5  g08367(.A(new_n10715), .B(new_n10710_1), .Y(new_n10716));
  nor_5  g08368(.A(new_n10716), .B(new_n10708), .Y(new_n10717));
  nor_5  g08369(.A(new_n10717), .B(new_n10707), .Y(new_n10718));
  nor_5  g08370(.A(new_n10718), .B(new_n10705), .Y(new_n10719));
  or_5   g08371(.A(new_n10719), .B(new_n10704), .Y(new_n10720));
  and_5  g08372(.A(new_n10720), .B(new_n10702), .Y(new_n10721));
  or_5   g08373(.A(new_n10721), .B(new_n10701_1), .Y(new_n10722));
  and_5  g08374(.A(new_n10722), .B(new_n10699), .Y(new_n10723));
  or_5   g08375(.A(new_n10723), .B(new_n10698), .Y(new_n10724));
  and_5  g08376(.A(new_n10724), .B(new_n10696), .Y(new_n10725));
  or_5   g08377(.A(new_n10725), .B(new_n10695), .Y(new_n10726));
  and_5  g08378(.A(new_n10726), .B(new_n10693), .Y(new_n10727));
  or_5   g08379(.A(new_n10727), .B(new_n10692_1), .Y(new_n10728));
  and_5  g08380(.A(new_n10728), .B(new_n10690), .Y(new_n10729));
  or_5   g08381(.A(new_n10729), .B(new_n10689), .Y(new_n10730));
  xor_4  g08382(.A(new_n10730), .B(new_n10687), .Y(new_n10731));
  xnor_4 g08383(.A(new_n10731), .B(new_n9119), .Y(new_n10732));
  xor_4  g08384(.A(new_n10728), .B(new_n10690), .Y(new_n10733));
  and_5  g08385(.A(new_n10733), .B(new_n9123), .Y(new_n10734));
  xnor_4 g08386(.A(new_n10733), .B(new_n9123), .Y(new_n10735));
  xor_4  g08387(.A(new_n10726), .B(new_n10693), .Y(new_n10736));
  and_5  g08388(.A(new_n10736), .B(new_n9127), .Y(new_n10737));
  xnor_4 g08389(.A(new_n10736), .B(new_n9127), .Y(new_n10738));
  xor_4  g08390(.A(new_n10724), .B(new_n10696), .Y(new_n10739_1));
  and_5  g08391(.A(new_n10739_1), .B(new_n9131), .Y(new_n10740));
  xnor_4 g08392(.A(new_n10739_1), .B(new_n9131), .Y(new_n10741));
  xor_4  g08393(.A(new_n10722), .B(new_n10699), .Y(new_n10742));
  and_5  g08394(.A(new_n10742), .B(new_n9135), .Y(new_n10743));
  xnor_4 g08395(.A(new_n10742), .B(new_n9135), .Y(new_n10744));
  xor_4  g08396(.A(new_n10720), .B(new_n10702), .Y(new_n10745));
  and_5  g08397(.A(new_n10745), .B(new_n9138), .Y(new_n10746));
  xnor_4 g08398(.A(new_n10745), .B(new_n9138), .Y(new_n10747));
  xnor_4 g08399(.A(new_n10718), .B(new_n10705), .Y(new_n10748));
  nor_5  g08400(.A(new_n10748), .B(new_n9142), .Y(new_n10749));
  xnor_4 g08401(.A(new_n10716), .B(new_n10708), .Y(new_n10750));
  nor_5  g08402(.A(new_n10750), .B(new_n9147), .Y(new_n10751));
  xnor_4 g08403(.A(new_n10750), .B(new_n9147), .Y(new_n10752));
  xnor_4 g08404(.A(new_n10608), .B(new_n2543), .Y(new_n10753));
  nor_5  g08405(.A(new_n10753), .B(new_n9156), .Y(new_n10754));
  and_5  g08406(.A(new_n10754), .B(new_n9158), .Y(new_n10755));
  xnor_4 g08407(.A(new_n10754), .B(new_n9153), .Y(new_n10756_1));
  xnor_4 g08408(.A(new_n10714), .B(new_n10712_1), .Y(new_n10757));
  not_8  g08409(.A(new_n10757), .Y(new_n10758));
  and_5  g08410(.A(new_n10758), .B(new_n10756_1), .Y(new_n10759));
  nor_5  g08411(.A(new_n10759), .B(new_n10755), .Y(new_n10760));
  nor_5  g08412(.A(new_n10760), .B(new_n10752), .Y(new_n10761));
  nor_5  g08413(.A(new_n10761), .B(new_n10751), .Y(new_n10762));
  xnor_4 g08414(.A(new_n10748), .B(new_n9142), .Y(new_n10763_1));
  nor_5  g08415(.A(new_n10763_1), .B(new_n10762), .Y(new_n10764));
  nor_5  g08416(.A(new_n10764), .B(new_n10749), .Y(new_n10765));
  nor_5  g08417(.A(new_n10765), .B(new_n10747), .Y(new_n10766));
  nor_5  g08418(.A(new_n10766), .B(new_n10746), .Y(new_n10767));
  nor_5  g08419(.A(new_n10767), .B(new_n10744), .Y(new_n10768));
  nor_5  g08420(.A(new_n10768), .B(new_n10743), .Y(new_n10769));
  nor_5  g08421(.A(new_n10769), .B(new_n10741), .Y(new_n10770));
  nor_5  g08422(.A(new_n10770), .B(new_n10740), .Y(new_n10771));
  nor_5  g08423(.A(new_n10771), .B(new_n10738), .Y(new_n10772));
  nor_5  g08424(.A(new_n10772), .B(new_n10737), .Y(new_n10773));
  nor_5  g08425(.A(new_n10773), .B(new_n10735), .Y(new_n10774));
  nor_5  g08426(.A(new_n10774), .B(new_n10734), .Y(new_n10775_1));
  xnor_4 g08427(.A(new_n10775_1), .B(new_n10732), .Y(n1498));
  not_8  g08428(.A(new_n5956), .Y(new_n10777));
  xnor_4 g08429(.A(n20658), .B(n9090), .Y(new_n10778));
  xnor_4 g08430(.A(new_n10778), .B(new_n10777), .Y(new_n10779));
  xnor_4 g08431(.A(new_n10779), .B(new_n5004), .Y(n1501));
  nor_5  g08432(.A(n15506), .B(n11473), .Y(new_n10781));
  not_8  g08433(.A(new_n10781), .Y(new_n10782));
  nor_5  g08434(.A(new_n10782), .B(n5131), .Y(new_n10783));
  not_8  g08435(.A(new_n10783), .Y(new_n10784));
  nor_5  g08436(.A(new_n10784), .B(n21538), .Y(new_n10785));
  not_8  g08437(.A(new_n10785), .Y(new_n10786));
  nor_5  g08438(.A(new_n10786), .B(n25094), .Y(new_n10787));
  not_8  g08439(.A(new_n10787), .Y(new_n10788));
  nor_5  g08440(.A(new_n10788), .B(n1611), .Y(new_n10789));
  xnor_4 g08441(.A(new_n10789), .B(n752), .Y(new_n10790));
  xnor_4 g08442(.A(new_n10790), .B(new_n9660), .Y(new_n10791));
  xnor_4 g08443(.A(new_n10787), .B(n1611), .Y(new_n10792_1));
  nor_5  g08444(.A(new_n10792_1), .B(new_n9662), .Y(new_n10793));
  xnor_4 g08445(.A(new_n10792_1), .B(new_n9662), .Y(new_n10794));
  xnor_4 g08446(.A(new_n10785), .B(n25094), .Y(new_n10795));
  nor_5  g08447(.A(new_n10795), .B(new_n9667), .Y(new_n10796));
  xnor_4 g08448(.A(new_n10795), .B(new_n9667), .Y(new_n10797));
  xnor_4 g08449(.A(new_n10783), .B(n21538), .Y(new_n10798));
  and_5  g08450(.A(new_n10798), .B(new_n9675), .Y(new_n10799));
  xnor_4 g08451(.A(new_n10781), .B(n5131), .Y(new_n10800));
  nor_5  g08452(.A(new_n10800), .B(new_n9680), .Y(new_n10801));
  xnor_4 g08453(.A(new_n10800), .B(new_n9680), .Y(new_n10802));
  not_8  g08454(.A(n15506), .Y(new_n10803));
  nor_5  g08455(.A(new_n9686), .B(new_n10803), .Y(new_n10804));
  xnor_4 g08456(.A(n15506), .B(n11473), .Y(new_n10805));
  not_8  g08457(.A(new_n10805), .Y(new_n10806));
  nor_5  g08458(.A(new_n10806), .B(new_n10804), .Y(new_n10807));
  not_8  g08459(.A(new_n9683), .Y(new_n10808));
  not_8  g08460(.A(n11473), .Y(new_n10809));
  and_5  g08461(.A(new_n10804), .B(new_n10809), .Y(new_n10810));
  nor_5  g08462(.A(new_n10810), .B(new_n10807), .Y(new_n10811));
  and_5  g08463(.A(new_n10811), .B(new_n10808), .Y(new_n10812));
  nor_5  g08464(.A(new_n10812), .B(new_n10807), .Y(new_n10813));
  nor_5  g08465(.A(new_n10813), .B(new_n10802), .Y(new_n10814));
  nor_5  g08466(.A(new_n10814), .B(new_n10801), .Y(new_n10815));
  xnor_4 g08467(.A(new_n10798), .B(new_n9673), .Y(new_n10816));
  and_5  g08468(.A(new_n10816), .B(new_n10815), .Y(new_n10817_1));
  or_5   g08469(.A(new_n10817_1), .B(new_n10799), .Y(new_n10818));
  nor_5  g08470(.A(new_n10818), .B(new_n10797), .Y(new_n10819));
  nor_5  g08471(.A(new_n10819), .B(new_n10796), .Y(new_n10820));
  nor_5  g08472(.A(new_n10820), .B(new_n10794), .Y(new_n10821));
  nor_5  g08473(.A(new_n10821), .B(new_n10793), .Y(new_n10822));
  xor_4  g08474(.A(new_n10822), .B(new_n10791), .Y(new_n10823));
  not_8  g08475(.A(n20470), .Y(new_n10824));
  xnor_4 g08476(.A(new_n10824), .B(n3366), .Y(new_n10825));
  and_5  g08477(.A(n26565), .B(n21222), .Y(new_n10826));
  or_5   g08478(.A(n26565), .B(n21222), .Y(new_n10827));
  nor_5  g08479(.A(n9832), .B(n3959), .Y(new_n10828));
  or_5   g08480(.A(new_n9493_1), .B(new_n9478), .Y(new_n10829));
  and_5  g08481(.A(new_n10829), .B(new_n9477), .Y(new_n10830));
  nor_5  g08482(.A(new_n10830), .B(new_n10828), .Y(new_n10831));
  and_5  g08483(.A(new_n10831), .B(new_n10827), .Y(new_n10832));
  nor_5  g08484(.A(new_n10832), .B(new_n10826), .Y(new_n10833));
  xor_4  g08485(.A(new_n10833), .B(new_n10825), .Y(new_n10834_1));
  xnor_4 g08486(.A(new_n10834_1), .B(new_n10823), .Y(new_n10835));
  xor_4  g08487(.A(new_n10820), .B(new_n10794), .Y(new_n10836));
  not_8  g08488(.A(n21222), .Y(new_n10837));
  xnor_4 g08489(.A(n26565), .B(new_n10837), .Y(new_n10838));
  xnor_4 g08490(.A(new_n10838), .B(new_n10831), .Y(new_n10839));
  not_8  g08491(.A(new_n10839), .Y(new_n10840));
  and_5  g08492(.A(new_n10840), .B(new_n10836), .Y(new_n10841));
  xnor_4 g08493(.A(new_n10840), .B(new_n10836), .Y(new_n10842));
  not_8  g08494(.A(new_n9495), .Y(new_n10843));
  xor_4  g08495(.A(new_n10818), .B(new_n10797), .Y(new_n10844));
  and_5  g08496(.A(new_n10844), .B(new_n10843), .Y(new_n10845));
  xnor_4 g08497(.A(new_n10844), .B(new_n10843), .Y(new_n10846));
  xnor_4 g08498(.A(new_n10816), .B(new_n10815), .Y(new_n10847));
  not_8  g08499(.A(new_n10847), .Y(new_n10848));
  nor_5  g08500(.A(new_n10848), .B(new_n9546), .Y(new_n10849));
  xnor_4 g08501(.A(new_n10848), .B(new_n9546), .Y(new_n10850));
  xor_4  g08502(.A(new_n10813), .B(new_n10802), .Y(new_n10851_1));
  nor_5  g08503(.A(new_n10851_1), .B(new_n9551), .Y(new_n10852));
  xnor_4 g08504(.A(new_n10811), .B(new_n10808), .Y(new_n10853));
  nor_5  g08505(.A(new_n10853), .B(new_n9557_1), .Y(new_n10854));
  xnor_4 g08506(.A(new_n9686), .B(n15506), .Y(new_n10855));
  nor_5  g08507(.A(new_n10855), .B(new_n7198), .Y(new_n10856));
  xnor_4 g08508(.A(new_n10853), .B(new_n9560), .Y(new_n10857));
  and_5  g08509(.A(new_n10857), .B(new_n10856), .Y(new_n10858));
  nor_5  g08510(.A(new_n10858), .B(new_n10854), .Y(new_n10859));
  xor_4  g08511(.A(new_n10851_1), .B(new_n9551), .Y(new_n10860));
  and_5  g08512(.A(new_n10860), .B(new_n10859), .Y(new_n10861));
  or_5   g08513(.A(new_n10861), .B(new_n10852), .Y(new_n10862));
  nor_5  g08514(.A(new_n10862), .B(new_n10850), .Y(new_n10863));
  nor_5  g08515(.A(new_n10863), .B(new_n10849), .Y(new_n10864));
  nor_5  g08516(.A(new_n10864), .B(new_n10846), .Y(new_n10865));
  nor_5  g08517(.A(new_n10865), .B(new_n10845), .Y(new_n10866));
  nor_5  g08518(.A(new_n10866), .B(new_n10842), .Y(new_n10867));
  nor_5  g08519(.A(new_n10867), .B(new_n10841), .Y(new_n10868));
  xnor_4 g08520(.A(new_n10868), .B(new_n10835), .Y(n1518));
  not_8  g08521(.A(n17458), .Y(new_n10870));
  nor_5  g08522(.A(new_n10870), .B(n14826), .Y(new_n10871));
  xnor_4 g08523(.A(n17458), .B(n14826), .Y(new_n10872));
  not_8  g08524(.A(n1222), .Y(new_n10873));
  nor_5  g08525(.A(n23493), .B(new_n10873), .Y(new_n10874_1));
  xnor_4 g08526(.A(n23493), .B(n1222), .Y(new_n10875));
  not_8  g08527(.A(n25240), .Y(new_n10876));
  nor_5  g08528(.A(new_n10876), .B(n10275), .Y(new_n10877));
  xnor_4 g08529(.A(n25240), .B(n10275), .Y(new_n10878));
  nor_5  g08530(.A(n15146), .B(new_n10414), .Y(new_n10879));
  xnor_4 g08531(.A(n15146), .B(n10125), .Y(new_n10880));
  not_8  g08532(.A(n8067), .Y(new_n10881));
  nor_5  g08533(.A(n11579), .B(new_n10881), .Y(new_n10882));
  xnor_4 g08534(.A(n11579), .B(n8067), .Y(new_n10883));
  not_8  g08535(.A(n20923), .Y(new_n10884));
  nor_5  g08536(.A(new_n10884), .B(n21), .Y(new_n10885));
  xnor_4 g08537(.A(n20923), .B(n21), .Y(new_n10886));
  nor_5  g08538(.A(new_n8432_1), .B(n1682), .Y(new_n10887));
  xnor_4 g08539(.A(n18157), .B(n1682), .Y(new_n10888));
  nor_5  g08540(.A(n12161), .B(new_n9835), .Y(new_n10889));
  nor_5  g08541(.A(new_n7217), .B(n7963), .Y(new_n10890));
  nor_5  g08542(.A(new_n7941), .B(n5026), .Y(new_n10891));
  nor_5  g08543(.A(n10017), .B(new_n7220), .Y(new_n10892));
  nor_5  g08544(.A(n8581), .B(new_n7939), .Y(new_n10893));
  not_8  g08545(.A(new_n10893), .Y(new_n10894));
  nor_5  g08546(.A(new_n10894), .B(new_n10892), .Y(new_n10895));
  nor_5  g08547(.A(new_n10895), .B(new_n10891), .Y(new_n10896));
  nor_5  g08548(.A(new_n10896), .B(new_n10890), .Y(new_n10897));
  nor_5  g08549(.A(new_n10897), .B(new_n10889), .Y(new_n10898));
  and_5  g08550(.A(new_n10898), .B(new_n10888), .Y(new_n10899));
  or_5   g08551(.A(new_n10899), .B(new_n10887), .Y(new_n10900));
  and_5  g08552(.A(new_n10900), .B(new_n10886), .Y(new_n10901));
  or_5   g08553(.A(new_n10901), .B(new_n10885), .Y(new_n10902));
  and_5  g08554(.A(new_n10902), .B(new_n10883), .Y(new_n10903));
  or_5   g08555(.A(new_n10903), .B(new_n10882), .Y(new_n10904));
  and_5  g08556(.A(new_n10904), .B(new_n10880), .Y(new_n10905));
  or_5   g08557(.A(new_n10905), .B(new_n10879), .Y(new_n10906));
  and_5  g08558(.A(new_n10906), .B(new_n10878), .Y(new_n10907));
  or_5   g08559(.A(new_n10907), .B(new_n10877), .Y(new_n10908));
  and_5  g08560(.A(new_n10908), .B(new_n10875), .Y(new_n10909));
  or_5   g08561(.A(new_n10909), .B(new_n10874_1), .Y(new_n10910));
  and_5  g08562(.A(new_n10910), .B(new_n10872), .Y(new_n10911));
  nor_5  g08563(.A(new_n10911), .B(new_n10871), .Y(new_n10912));
  not_8  g08564(.A(new_n4200), .Y(new_n10913));
  nor_5  g08565(.A(new_n10913), .B(n3468), .Y(new_n10914));
  not_8  g08566(.A(new_n10914), .Y(new_n10915));
  nor_5  g08567(.A(new_n10915), .B(n12821), .Y(new_n10916));
  not_8  g08568(.A(new_n10916), .Y(new_n10917));
  nor_5  g08569(.A(new_n10917), .B(n22492), .Y(new_n10918));
  not_8  g08570(.A(new_n10918), .Y(new_n10919));
  nor_5  g08571(.A(new_n10919), .B(n7330), .Y(new_n10920));
  not_8  g08572(.A(new_n10920), .Y(new_n10921));
  nor_5  g08573(.A(new_n10921), .B(n767), .Y(new_n10922));
  xnor_4 g08574(.A(new_n10922), .B(n2944), .Y(new_n10923));
  and_5  g08575(.A(new_n10923), .B(n19282), .Y(new_n10924_1));
  and_5  g08576(.A(new_n10922), .B(new_n2674), .Y(new_n10925));
  xnor_4 g08577(.A(new_n10920), .B(n767), .Y(new_n10926));
  nor_5  g08578(.A(new_n10926), .B(n12657), .Y(new_n10927));
  xnor_4 g08579(.A(new_n10926), .B(new_n2926), .Y(new_n10928));
  xnor_4 g08580(.A(new_n10918), .B(n7330), .Y(new_n10929));
  and_5  g08581(.A(new_n10929), .B(n17077), .Y(new_n10930));
  xnor_4 g08582(.A(new_n10929), .B(n17077), .Y(new_n10931));
  xnor_4 g08583(.A(new_n10916), .B(n22492), .Y(new_n10932));
  not_8  g08584(.A(new_n10932), .Y(new_n10933));
  nor_5  g08585(.A(new_n10933), .B(new_n7251), .Y(new_n10934));
  xnor_4 g08586(.A(new_n10933), .B(n26510), .Y(new_n10935));
  xnor_4 g08587(.A(new_n10914), .B(n12821), .Y(new_n10936));
  not_8  g08588(.A(new_n10936), .Y(new_n10937));
  nor_5  g08589(.A(new_n10937), .B(new_n3815), .Y(new_n10938));
  nor_5  g08590(.A(new_n10936), .B(n23068), .Y(new_n10939));
  and_5  g08591(.A(new_n4201), .B(n19514), .Y(new_n10940));
  or_5   g08592(.A(new_n4219), .B(new_n4205_1), .Y(new_n10941));
  and_5  g08593(.A(new_n10941), .B(new_n4203), .Y(new_n10942));
  nor_5  g08594(.A(new_n10942), .B(new_n10940), .Y(new_n10943_1));
  nor_5  g08595(.A(new_n10943_1), .B(new_n10939), .Y(new_n10944));
  or_5   g08596(.A(new_n10944), .B(new_n10938), .Y(new_n10945));
  and_5  g08597(.A(new_n10945), .B(new_n10935), .Y(new_n10946));
  nor_5  g08598(.A(new_n10946), .B(new_n10934), .Y(new_n10947));
  nor_5  g08599(.A(new_n10947), .B(new_n10931), .Y(new_n10948));
  nor_5  g08600(.A(new_n10948), .B(new_n10930), .Y(new_n10949));
  and_5  g08601(.A(new_n10949), .B(new_n10928), .Y(new_n10950));
  nor_5  g08602(.A(new_n10950), .B(new_n10927), .Y(new_n10951));
  or_5   g08603(.A(new_n10923), .B(n19282), .Y(new_n10952));
  and_5  g08604(.A(new_n10952), .B(new_n10951), .Y(new_n10953));
  or_5   g08605(.A(new_n10953), .B(new_n10925), .Y(new_n10954));
  nor_5  g08606(.A(new_n10954), .B(new_n10924_1), .Y(new_n10955));
  nor_5  g08607(.A(new_n10955), .B(new_n10912), .Y(new_n10956));
  xor_4  g08608(.A(new_n10910), .B(new_n10872), .Y(new_n10957));
  not_8  g08609(.A(n19282), .Y(new_n10958));
  xnor_4 g08610(.A(new_n10923), .B(new_n10958), .Y(new_n10959));
  xnor_4 g08611(.A(new_n10959), .B(new_n10951), .Y(new_n10960));
  not_8  g08612(.A(new_n10960), .Y(new_n10961_1));
  nor_5  g08613(.A(new_n10961_1), .B(new_n10957), .Y(new_n10962));
  xnor_4 g08614(.A(new_n10961_1), .B(new_n10957), .Y(new_n10963));
  xor_4  g08615(.A(new_n10908), .B(new_n10875), .Y(new_n10964));
  xnor_4 g08616(.A(new_n10949), .B(new_n10928), .Y(new_n10965));
  nor_5  g08617(.A(new_n10965), .B(new_n10964), .Y(new_n10966));
  xnor_4 g08618(.A(new_n10965), .B(new_n10964), .Y(new_n10967));
  xor_4  g08619(.A(new_n10906), .B(new_n10878), .Y(new_n10968));
  xnor_4 g08620(.A(new_n10947), .B(new_n10931), .Y(new_n10969));
  not_8  g08621(.A(new_n10969), .Y(new_n10970));
  nor_5  g08622(.A(new_n10970), .B(new_n10968), .Y(new_n10971));
  xnor_4 g08623(.A(new_n10970), .B(new_n10968), .Y(new_n10972));
  xor_4  g08624(.A(new_n10904), .B(new_n10880), .Y(new_n10973));
  xor_4  g08625(.A(new_n10945), .B(new_n10935), .Y(new_n10974));
  nor_5  g08626(.A(new_n10974), .B(new_n10973), .Y(new_n10975));
  xnor_4 g08627(.A(new_n10974), .B(new_n10973), .Y(new_n10976));
  xor_4  g08628(.A(new_n10902), .B(new_n10883), .Y(new_n10977));
  xnor_4 g08629(.A(new_n10937), .B(n23068), .Y(new_n10978));
  xnor_4 g08630(.A(new_n10978), .B(new_n10943_1), .Y(new_n10979));
  nor_5  g08631(.A(new_n10979), .B(new_n10977), .Y(new_n10980));
  xnor_4 g08632(.A(new_n10979), .B(new_n10977), .Y(new_n10981));
  xor_4  g08633(.A(new_n10900), .B(new_n10886), .Y(new_n10982));
  nor_5  g08634(.A(new_n10982), .B(new_n4221_1), .Y(new_n10983));
  xnor_4 g08635(.A(new_n10898), .B(new_n10888), .Y(new_n10984));
  not_8  g08636(.A(new_n10984), .Y(new_n10985));
  nor_5  g08637(.A(new_n10985), .B(new_n4254), .Y(new_n10986));
  xnor_4 g08638(.A(new_n10984), .B(new_n4255), .Y(new_n10987));
  xnor_4 g08639(.A(n12161), .B(n7963), .Y(new_n10988));
  xnor_4 g08640(.A(new_n10988), .B(new_n10896), .Y(new_n10989));
  and_5  g08641(.A(new_n10989), .B(new_n4290), .Y(new_n10990));
  xnor_4 g08642(.A(new_n10989), .B(new_n4290), .Y(new_n10991));
  xnor_4 g08643(.A(n8581), .B(n3618), .Y(new_n10992));
  nor_5  g08644(.A(new_n10992), .B(new_n4268), .Y(new_n10993));
  xnor_4 g08645(.A(n10017), .B(n5026), .Y(new_n10994));
  xnor_4 g08646(.A(new_n10994), .B(new_n10894), .Y(new_n10995));
  not_8  g08647(.A(new_n10995), .Y(new_n10996));
  nor_5  g08648(.A(new_n10996), .B(new_n10993), .Y(new_n10997));
  xnor_4 g08649(.A(new_n10995), .B(new_n10993), .Y(new_n10998));
  and_5  g08650(.A(new_n10998), .B(new_n4262), .Y(new_n10999));
  nor_5  g08651(.A(new_n10999), .B(new_n10997), .Y(new_n11000));
  nor_5  g08652(.A(new_n11000), .B(new_n10991), .Y(new_n11001));
  nor_5  g08653(.A(new_n11001), .B(new_n10990), .Y(new_n11002));
  nor_5  g08654(.A(new_n11002), .B(new_n10987), .Y(new_n11003));
  nor_5  g08655(.A(new_n11003), .B(new_n10986), .Y(new_n11004));
  xnor_4 g08656(.A(new_n10982), .B(new_n4221_1), .Y(new_n11005_1));
  nor_5  g08657(.A(new_n11005_1), .B(new_n11004), .Y(new_n11006));
  nor_5  g08658(.A(new_n11006), .B(new_n10983), .Y(new_n11007));
  nor_5  g08659(.A(new_n11007), .B(new_n10981), .Y(new_n11008));
  nor_5  g08660(.A(new_n11008), .B(new_n10980), .Y(new_n11009));
  nor_5  g08661(.A(new_n11009), .B(new_n10976), .Y(new_n11010));
  nor_5  g08662(.A(new_n11010), .B(new_n10975), .Y(new_n11011_1));
  nor_5  g08663(.A(new_n11011_1), .B(new_n10972), .Y(new_n11012));
  nor_5  g08664(.A(new_n11012), .B(new_n10971), .Y(new_n11013));
  nor_5  g08665(.A(new_n11013), .B(new_n10967), .Y(new_n11014));
  nor_5  g08666(.A(new_n11014), .B(new_n10966), .Y(new_n11015));
  nor_5  g08667(.A(new_n11015), .B(new_n10963), .Y(new_n11016));
  nor_5  g08668(.A(new_n11016), .B(new_n10962), .Y(new_n11017));
  not_8  g08669(.A(new_n10912), .Y(new_n11018));
  xnor_4 g08670(.A(new_n10955), .B(new_n11018), .Y(new_n11019));
  and_5  g08671(.A(new_n11019), .B(new_n11017), .Y(new_n11020));
  nor_5  g08672(.A(new_n11020), .B(new_n10956), .Y(new_n11021));
  nor_5  g08673(.A(n20040), .B(new_n7429), .Y(new_n11022));
  or_5   g08674(.A(new_n8716_1), .B(new_n8683), .Y(new_n11023_1));
  and_5  g08675(.A(new_n11023_1), .B(new_n8682), .Y(new_n11024));
  nor_5  g08676(.A(new_n11024), .B(new_n11022), .Y(new_n11025_1));
  not_8  g08677(.A(new_n11025_1), .Y(new_n11026));
  xnor_4 g08678(.A(new_n11026), .B(new_n11021), .Y(new_n11027));
  xor_4  g08679(.A(new_n11019), .B(new_n11017), .Y(new_n11028));
  nor_5  g08680(.A(new_n11028), .B(new_n11025_1), .Y(new_n11029));
  xnor_4 g08681(.A(new_n11015), .B(new_n10963), .Y(new_n11030));
  nor_5  g08682(.A(new_n11030), .B(new_n8718), .Y(new_n11031));
  not_8  g08683(.A(new_n8718), .Y(new_n11032));
  not_8  g08684(.A(new_n11030), .Y(new_n11033));
  xnor_4 g08685(.A(new_n11033), .B(new_n11032), .Y(new_n11034));
  xnor_4 g08686(.A(new_n11013), .B(new_n10967), .Y(new_n11035));
  nor_5  g08687(.A(new_n11035), .B(new_n8788), .Y(new_n11036));
  not_8  g08688(.A(new_n11035), .Y(new_n11037));
  xnor_4 g08689(.A(new_n11037), .B(new_n8793), .Y(new_n11038));
  xnor_4 g08690(.A(new_n11011_1), .B(new_n10972), .Y(new_n11039));
  nor_5  g08691(.A(new_n11039), .B(new_n8795), .Y(new_n11040));
  xnor_4 g08692(.A(new_n11039), .B(new_n8795), .Y(new_n11041));
  xnor_4 g08693(.A(new_n11009), .B(new_n10976), .Y(new_n11042));
  nor_5  g08694(.A(new_n11042), .B(new_n8801), .Y(new_n11043));
  not_8  g08695(.A(new_n11042), .Y(new_n11044_1));
  xnor_4 g08696(.A(new_n11044_1), .B(new_n8802), .Y(new_n11045));
  xnor_4 g08697(.A(new_n11007), .B(new_n10981), .Y(new_n11046));
  nor_5  g08698(.A(new_n11046), .B(new_n8807), .Y(new_n11047));
  not_8  g08699(.A(new_n11046), .Y(new_n11048));
  xnor_4 g08700(.A(new_n11048), .B(new_n8807), .Y(new_n11049));
  xnor_4 g08701(.A(new_n11005_1), .B(new_n11004), .Y(new_n11050));
  not_8  g08702(.A(new_n11050), .Y(new_n11051));
  nor_5  g08703(.A(new_n11051), .B(new_n8814), .Y(new_n11052));
  xnor_4 g08704(.A(new_n11002), .B(new_n10987), .Y(new_n11053));
  nor_5  g08705(.A(new_n11053), .B(new_n8821_1), .Y(new_n11054));
  not_8  g08706(.A(new_n11053), .Y(new_n11055));
  xnor_4 g08707(.A(new_n11055), .B(new_n8818), .Y(new_n11056_1));
  not_8  g08708(.A(new_n8825), .Y(new_n11057));
  xnor_4 g08709(.A(new_n11000), .B(new_n10991), .Y(new_n11058));
  nor_5  g08710(.A(new_n11058), .B(new_n11057), .Y(new_n11059));
  xnor_4 g08711(.A(new_n10992), .B(new_n4267), .Y(new_n11060));
  not_8  g08712(.A(new_n11060), .Y(new_n11061));
  nor_5  g08713(.A(new_n11061), .B(new_n8832), .Y(new_n11062));
  and_5  g08714(.A(new_n11062), .B(new_n8835), .Y(new_n11063_1));
  xnor_4 g08715(.A(new_n10998), .B(new_n4270), .Y(new_n11064));
  xnor_4 g08716(.A(new_n11062), .B(new_n8830), .Y(new_n11065));
  not_8  g08717(.A(new_n11065), .Y(new_n11066));
  nor_5  g08718(.A(new_n11066), .B(new_n11064), .Y(new_n11067));
  nor_5  g08719(.A(new_n11067), .B(new_n11063_1), .Y(new_n11068));
  not_8  g08720(.A(new_n11058), .Y(new_n11069));
  xnor_4 g08721(.A(new_n11069), .B(new_n11057), .Y(new_n11070));
  and_5  g08722(.A(new_n11070), .B(new_n11068), .Y(new_n11071));
  nor_5  g08723(.A(new_n11071), .B(new_n11059), .Y(new_n11072));
  nor_5  g08724(.A(new_n11072), .B(new_n11056_1), .Y(new_n11073));
  nor_5  g08725(.A(new_n11073), .B(new_n11054), .Y(new_n11074));
  xnor_4 g08726(.A(new_n11051), .B(new_n8813), .Y(new_n11075));
  and_5  g08727(.A(new_n11075), .B(new_n11074), .Y(new_n11076));
  nor_5  g08728(.A(new_n11076), .B(new_n11052), .Y(new_n11077));
  and_5  g08729(.A(new_n11077), .B(new_n11049), .Y(new_n11078_1));
  nor_5  g08730(.A(new_n11078_1), .B(new_n11047), .Y(new_n11079));
  nor_5  g08731(.A(new_n11079), .B(new_n11045), .Y(new_n11080_1));
  nor_5  g08732(.A(new_n11080_1), .B(new_n11043), .Y(new_n11081));
  nor_5  g08733(.A(new_n11081), .B(new_n11041), .Y(new_n11082));
  nor_5  g08734(.A(new_n11082), .B(new_n11040), .Y(new_n11083));
  nor_5  g08735(.A(new_n11083), .B(new_n11038), .Y(new_n11084));
  nor_5  g08736(.A(new_n11084), .B(new_n11036), .Y(new_n11085));
  nor_5  g08737(.A(new_n11085), .B(new_n11034), .Y(new_n11086));
  nor_5  g08738(.A(new_n11086), .B(new_n11031), .Y(new_n11087));
  xnor_4 g08739(.A(new_n11028), .B(new_n11025_1), .Y(new_n11088));
  nor_5  g08740(.A(new_n11088), .B(new_n11087), .Y(new_n11089));
  nor_5  g08741(.A(new_n11089), .B(new_n11029), .Y(new_n11090));
  xor_4  g08742(.A(new_n11090), .B(new_n11027), .Y(n1527));
  xnor_4 g08743(.A(n25345), .B(n23463), .Y(new_n11092));
  nor_5  g08744(.A(new_n3095), .B(n9655), .Y(new_n11093));
  xnor_4 g08745(.A(n13074), .B(n9655), .Y(new_n11094_1));
  nor_5  g08746(.A(n13490), .B(new_n3099), .Y(new_n11095));
  xnor_4 g08747(.A(n13490), .B(n10739), .Y(new_n11096));
  nor_5  g08748(.A(n22660), .B(new_n2350), .Y(new_n11097));
  xnor_4 g08749(.A(n22660), .B(n21753), .Y(new_n11098));
  nor_5  g08750(.A(new_n2353), .B(n1777), .Y(new_n11099));
  xnor_4 g08751(.A(n21832), .B(n1777), .Y(new_n11100));
  nor_5  g08752(.A(new_n2356), .B(n8745), .Y(new_n11101_1));
  nor_5  g08753(.A(n16223), .B(new_n2441), .Y(new_n11102));
  and_5  g08754(.A(new_n9717), .B(new_n9712), .Y(new_n11103_1));
  nor_5  g08755(.A(new_n11103_1), .B(new_n11102), .Y(new_n11104));
  xnor_4 g08756(.A(n26913), .B(n8745), .Y(new_n11105));
  and_5  g08757(.A(new_n11105), .B(new_n11104), .Y(new_n11106));
  or_5   g08758(.A(new_n11106), .B(new_n11101_1), .Y(new_n11107));
  and_5  g08759(.A(new_n11107), .B(new_n11100), .Y(new_n11108));
  or_5   g08760(.A(new_n11108), .B(new_n11099), .Y(new_n11109));
  and_5  g08761(.A(new_n11109), .B(new_n11098), .Y(new_n11110));
  or_5   g08762(.A(new_n11110), .B(new_n11097), .Y(new_n11111));
  and_5  g08763(.A(new_n11111), .B(new_n11096), .Y(new_n11112));
  or_5   g08764(.A(new_n11112), .B(new_n11095), .Y(new_n11113));
  and_5  g08765(.A(new_n11113), .B(new_n11094_1), .Y(new_n11114));
  or_5   g08766(.A(new_n11114), .B(new_n11093), .Y(new_n11115));
  xor_4  g08767(.A(new_n11115), .B(new_n11092), .Y(new_n11116));
  xnor_4 g08768(.A(new_n11116), .B(new_n7845), .Y(new_n11117));
  xor_4  g08769(.A(new_n11113), .B(new_n11094_1), .Y(new_n11118));
  nor_5  g08770(.A(new_n11118), .B(new_n7851), .Y(new_n11119));
  xnor_4 g08771(.A(new_n11118), .B(new_n7851), .Y(new_n11120_1));
  xor_4  g08772(.A(new_n11111), .B(new_n11096), .Y(new_n11121_1));
  nor_5  g08773(.A(new_n11121_1), .B(new_n7858), .Y(new_n11122));
  xnor_4 g08774(.A(new_n11121_1), .B(new_n7858), .Y(new_n11123));
  xor_4  g08775(.A(new_n11109), .B(new_n11098), .Y(new_n11124));
  nor_5  g08776(.A(new_n11124), .B(new_n7864), .Y(new_n11125));
  xnor_4 g08777(.A(new_n11124), .B(new_n7864), .Y(new_n11126));
  xor_4  g08778(.A(new_n11107), .B(new_n11100), .Y(new_n11127_1));
  nor_5  g08779(.A(new_n11127_1), .B(new_n7871), .Y(new_n11128));
  xnor_4 g08780(.A(new_n11127_1), .B(new_n7871), .Y(new_n11129));
  xnor_4 g08781(.A(new_n11105), .B(new_n11104), .Y(new_n11130));
  and_5  g08782(.A(new_n11130), .B(new_n7879), .Y(new_n11131));
  and_5  g08783(.A(new_n9718), .B(new_n7882), .Y(new_n11132_1));
  nor_5  g08784(.A(new_n9727), .B(new_n9719), .Y(new_n11133));
  nor_5  g08785(.A(new_n11133), .B(new_n11132_1), .Y(new_n11134_1));
  xnor_4 g08786(.A(new_n11130), .B(new_n7879), .Y(new_n11135));
  nor_5  g08787(.A(new_n11135), .B(new_n11134_1), .Y(new_n11136));
  nor_5  g08788(.A(new_n11136), .B(new_n11131), .Y(new_n11137));
  nor_5  g08789(.A(new_n11137), .B(new_n11129), .Y(new_n11138_1));
  nor_5  g08790(.A(new_n11138_1), .B(new_n11128), .Y(new_n11139));
  nor_5  g08791(.A(new_n11139), .B(new_n11126), .Y(new_n11140));
  nor_5  g08792(.A(new_n11140), .B(new_n11125), .Y(new_n11141));
  nor_5  g08793(.A(new_n11141), .B(new_n11123), .Y(new_n11142));
  nor_5  g08794(.A(new_n11142), .B(new_n11122), .Y(new_n11143));
  nor_5  g08795(.A(new_n11143), .B(new_n11120_1), .Y(new_n11144));
  nor_5  g08796(.A(new_n11144), .B(new_n11119), .Y(new_n11145));
  xor_4  g08797(.A(new_n11145), .B(new_n11117), .Y(n1580));
  xnor_4 g08798(.A(n18962), .B(n12315), .Y(new_n11147));
  nor_5  g08799(.A(new_n11147), .B(new_n7401), .Y(new_n11148));
  nor_5  g08800(.A(new_n6771), .B(n12315), .Y(new_n11149));
  xnor_4 g08801(.A(n10158), .B(n3952), .Y(new_n11150));
  xnor_4 g08802(.A(new_n11150), .B(new_n11149), .Y(new_n11151));
  xnor_4 g08803(.A(new_n11151), .B(new_n11148), .Y(new_n11152));
  xnor_4 g08804(.A(new_n11152), .B(new_n7407), .Y(n1586));
  xnor_4 g08805(.A(n19539), .B(n1483), .Y(new_n11154));
  not_8  g08806(.A(n8194), .Y(new_n11155));
  nor_5  g08807(.A(n24093), .B(new_n11155), .Y(new_n11156));
  xnor_4 g08808(.A(n24093), .B(n8194), .Y(new_n11157));
  not_8  g08809(.A(n23657), .Y(new_n11158));
  nor_5  g08810(.A(new_n11158), .B(n23035), .Y(new_n11159));
  xnor_4 g08811(.A(n23657), .B(n23035), .Y(new_n11160));
  not_8  g08812(.A(n16911), .Y(new_n11161));
  nor_5  g08813(.A(new_n11161), .B(n7773), .Y(new_n11162));
  and_5  g08814(.A(new_n6460), .B(new_n6432), .Y(new_n11163));
  or_5   g08815(.A(new_n11163), .B(new_n11162), .Y(new_n11164));
  and_5  g08816(.A(new_n11164), .B(new_n11160), .Y(new_n11165));
  or_5   g08817(.A(new_n11165), .B(new_n11159), .Y(new_n11166));
  and_5  g08818(.A(new_n11166), .B(new_n11157), .Y(new_n11167));
  or_5   g08819(.A(new_n11167), .B(new_n11156), .Y(new_n11168));
  xor_4  g08820(.A(new_n11168), .B(new_n11154), .Y(new_n11169));
  xnor_4 g08821(.A(n25494), .B(n1314), .Y(new_n11170));
  and_5  g08822(.A(new_n3424), .B(n3306), .Y(new_n11171));
  xnor_4 g08823(.A(n10117), .B(n3306), .Y(new_n11172));
  nor_5  g08824(.A(new_n8230), .B(n13460), .Y(new_n11173));
  xnor_4 g08825(.A(n22335), .B(n13460), .Y(new_n11174));
  nor_5  g08826(.A(new_n8234), .B(n6104), .Y(new_n11175));
  nor_5  g08827(.A(n4119), .B(new_n8238), .Y(new_n11176));
  and_5  g08828(.A(new_n4659), .B(new_n4637), .Y(new_n11177));
  or_5   g08829(.A(new_n11177), .B(new_n11176), .Y(new_n11178));
  xnor_4 g08830(.A(n24048), .B(n6104), .Y(new_n11179));
  and_5  g08831(.A(new_n11179), .B(new_n11178), .Y(new_n11180));
  or_5   g08832(.A(new_n11180), .B(new_n11175), .Y(new_n11181));
  and_5  g08833(.A(new_n11181), .B(new_n11174), .Y(new_n11182_1));
  or_5   g08834(.A(new_n11182_1), .B(new_n11173), .Y(new_n11183));
  and_5  g08835(.A(new_n11183), .B(new_n11172), .Y(new_n11184_1));
  or_5   g08836(.A(new_n11184_1), .B(new_n11171), .Y(new_n11185));
  xor_4  g08837(.A(new_n11185), .B(new_n11170), .Y(new_n11186));
  xnor_4 g08838(.A(n25296), .B(n23717), .Y(new_n11187));
  not_8  g08839(.A(n7788), .Y(new_n11188));
  nor_5  g08840(.A(n20013), .B(new_n11188), .Y(new_n11189));
  xnor_4 g08841(.A(n20013), .B(n7788), .Y(new_n11190));
  not_8  g08842(.A(n5443), .Y(new_n11191));
  nor_5  g08843(.A(new_n11191), .B(n1320), .Y(new_n11192_1));
  xnor_4 g08844(.A(n5443), .B(n1320), .Y(new_n11193));
  not_8  g08845(.A(n18584), .Y(new_n11194));
  nor_5  g08846(.A(n19803), .B(new_n11194), .Y(new_n11195));
  or_5   g08847(.A(new_n6428), .B(new_n6427_1), .Y(new_n11196));
  and_5  g08848(.A(new_n11196), .B(new_n6425), .Y(new_n11197));
  or_5   g08849(.A(new_n11197), .B(new_n11195), .Y(new_n11198));
  and_5  g08850(.A(new_n11198), .B(new_n11193), .Y(new_n11199));
  or_5   g08851(.A(new_n11199), .B(new_n11192_1), .Y(new_n11200));
  and_5  g08852(.A(new_n11200), .B(new_n11190), .Y(new_n11201_1));
  or_5   g08853(.A(new_n11201_1), .B(new_n11189), .Y(new_n11202));
  xor_4  g08854(.A(new_n11202), .B(new_n11187), .Y(new_n11203));
  xnor_4 g08855(.A(new_n11203), .B(new_n11186), .Y(new_n11204));
  xor_4  g08856(.A(new_n11183), .B(new_n11172), .Y(new_n11205));
  xor_4  g08857(.A(new_n11200), .B(new_n11190), .Y(new_n11206));
  and_5  g08858(.A(new_n11206), .B(new_n11205), .Y(new_n11207));
  xor_4  g08859(.A(new_n11206), .B(new_n11205), .Y(new_n11208));
  xor_4  g08860(.A(new_n11181), .B(new_n11174), .Y(new_n11209));
  xor_4  g08861(.A(new_n11198), .B(new_n11193), .Y(new_n11210));
  nor_5  g08862(.A(new_n11210), .B(new_n11209), .Y(new_n11211));
  xnor_4 g08863(.A(new_n11210), .B(new_n11209), .Y(new_n11212));
  not_8  g08864(.A(new_n11212), .Y(new_n11213));
  xor_4  g08865(.A(new_n11179), .B(new_n11178), .Y(new_n11214));
  and_5  g08866(.A(new_n11214), .B(new_n6430), .Y(new_n11215));
  xnor_4 g08867(.A(new_n11214), .B(new_n6430), .Y(new_n11216));
  and_5  g08868(.A(new_n4685), .B(new_n4660), .Y(new_n11217));
  nor_5  g08869(.A(new_n4722_1), .B(new_n4686), .Y(new_n11218));
  nor_5  g08870(.A(new_n11218), .B(new_n11217), .Y(new_n11219));
  nor_5  g08871(.A(new_n11219), .B(new_n11216), .Y(new_n11220_1));
  nor_5  g08872(.A(new_n11220_1), .B(new_n11215), .Y(new_n11221));
  and_5  g08873(.A(new_n11221), .B(new_n11213), .Y(new_n11222));
  nor_5  g08874(.A(new_n11222), .B(new_n11211), .Y(new_n11223_1));
  and_5  g08875(.A(new_n11223_1), .B(new_n11208), .Y(new_n11224));
  nor_5  g08876(.A(new_n11224), .B(new_n11207), .Y(new_n11225));
  xnor_4 g08877(.A(new_n11225), .B(new_n11204), .Y(new_n11226));
  xnor_4 g08878(.A(new_n11226), .B(new_n11169), .Y(new_n11227));
  xor_4  g08879(.A(new_n11166), .B(new_n11157), .Y(new_n11228));
  xor_4  g08880(.A(new_n11223_1), .B(new_n11208), .Y(new_n11229));
  nor_5  g08881(.A(new_n11229), .B(new_n11228), .Y(new_n11230));
  xnor_4 g08882(.A(new_n11229), .B(new_n11228), .Y(new_n11231));
  xor_4  g08883(.A(new_n11164), .B(new_n11160), .Y(new_n11232));
  xnor_4 g08884(.A(new_n11221), .B(new_n11213), .Y(new_n11233));
  nor_5  g08885(.A(new_n11233), .B(new_n11232), .Y(new_n11234_1));
  xnor_4 g08886(.A(new_n11233), .B(new_n11232), .Y(new_n11235));
  xnor_4 g08887(.A(new_n11219), .B(new_n11216), .Y(new_n11236));
  not_8  g08888(.A(new_n11236), .Y(new_n11237));
  nor_5  g08889(.A(new_n11237), .B(new_n6461), .Y(new_n11238));
  xnor_4 g08890(.A(new_n11237), .B(new_n6461), .Y(new_n11239));
  not_8  g08891(.A(new_n4723), .Y(new_n11240));
  nor_5  g08892(.A(new_n6510), .B(new_n11240), .Y(new_n11241));
  nor_5  g08893(.A(new_n6520), .B(new_n4726), .Y(new_n11242));
  xnor_4 g08894(.A(new_n6520), .B(new_n4726), .Y(new_n11243));
  and_5  g08895(.A(new_n6522), .B(new_n4730), .Y(new_n11244));
  and_5  g08896(.A(new_n6528), .B(new_n4734), .Y(new_n11245_1));
  xnor_4 g08897(.A(new_n6528), .B(new_n4734), .Y(new_n11246));
  nor_5  g08898(.A(new_n6532), .B(new_n4740), .Y(new_n11247));
  nor_5  g08899(.A(new_n11247), .B(new_n6536), .Y(new_n11248));
  xnor_4 g08900(.A(new_n11247), .B(new_n6535), .Y(new_n11249));
  and_5  g08901(.A(new_n11249), .B(new_n4745_1), .Y(new_n11250));
  nor_5  g08902(.A(new_n11250), .B(new_n11248), .Y(new_n11251));
  nor_5  g08903(.A(new_n11251), .B(new_n11246), .Y(new_n11252));
  nor_5  g08904(.A(new_n11252), .B(new_n11245_1), .Y(new_n11253));
  xnor_4 g08905(.A(new_n6522), .B(new_n4730), .Y(new_n11254));
  nor_5  g08906(.A(new_n11254), .B(new_n11253), .Y(new_n11255));
  nor_5  g08907(.A(new_n11255), .B(new_n11244), .Y(new_n11256));
  nor_5  g08908(.A(new_n11256), .B(new_n11243), .Y(new_n11257));
  nor_5  g08909(.A(new_n11257), .B(new_n11242), .Y(new_n11258));
  xnor_4 g08910(.A(new_n6510), .B(new_n11240), .Y(new_n11259));
  nor_5  g08911(.A(new_n11259), .B(new_n11258), .Y(new_n11260));
  nor_5  g08912(.A(new_n11260), .B(new_n11241), .Y(new_n11261_1));
  nor_5  g08913(.A(new_n11261_1), .B(new_n11239), .Y(new_n11262));
  nor_5  g08914(.A(new_n11262), .B(new_n11238), .Y(new_n11263));
  nor_5  g08915(.A(new_n11263), .B(new_n11235), .Y(new_n11264));
  nor_5  g08916(.A(new_n11264), .B(new_n11234_1), .Y(new_n11265));
  nor_5  g08917(.A(new_n11265), .B(new_n11231), .Y(new_n11266_1));
  nor_5  g08918(.A(new_n11266_1), .B(new_n11230), .Y(new_n11267));
  xor_4  g08919(.A(new_n11267), .B(new_n11227), .Y(n1590));
  xnor_4 g08920(.A(new_n7590), .B(new_n7576), .Y(n1602));
  xor_4  g08921(.A(new_n2845), .B(new_n2790), .Y(n1634));
  xnor_4 g08922(.A(new_n11265), .B(new_n11231), .Y(n1636));
  nor_5  g08923(.A(n10514), .B(n4514), .Y(new_n11272));
  not_8  g08924(.A(n4514), .Y(new_n11273_1));
  xnor_4 g08925(.A(n10514), .B(new_n11273_1), .Y(new_n11274));
  nor_5  g08926(.A(n18649), .B(n3984), .Y(new_n11275_1));
  not_8  g08927(.A(n18649), .Y(new_n11276));
  xnor_4 g08928(.A(new_n11276), .B(n3984), .Y(new_n11277));
  and_5  g08929(.A(n19652), .B(n6218), .Y(new_n11278));
  or_5   g08930(.A(n19652), .B(n6218), .Y(new_n11279));
  nor_5  g08931(.A(n20470), .B(n3366), .Y(new_n11280));
  and_5  g08932(.A(new_n10833), .B(new_n10825), .Y(new_n11281));
  nor_5  g08933(.A(new_n11281), .B(new_n11280), .Y(new_n11282));
  and_5  g08934(.A(new_n11282), .B(new_n11279), .Y(new_n11283));
  nor_5  g08935(.A(new_n11283), .B(new_n11278), .Y(new_n11284));
  and_5  g08936(.A(new_n11284), .B(new_n11277), .Y(new_n11285));
  or_5   g08937(.A(new_n11285), .B(new_n11275_1), .Y(new_n11286));
  and_5  g08938(.A(new_n11286), .B(new_n11274), .Y(new_n11287));
  nor_5  g08939(.A(new_n11287), .B(new_n11272), .Y(new_n11288));
  not_8  g08940(.A(n20040), .Y(new_n11289));
  xnor_4 g08941(.A(n18880), .B(new_n7429), .Y(new_n11290_1));
  not_8  g08942(.A(new_n11290_1), .Y(new_n11291));
  nor_5  g08943(.A(n25475), .B(n23697), .Y(new_n11292));
  nor_5  g08944(.A(new_n6787), .B(new_n6746), .Y(new_n11293));
  nor_5  g08945(.A(new_n11293), .B(new_n11292), .Y(new_n11294));
  xnor_4 g08946(.A(new_n11294), .B(new_n11291), .Y(new_n11295));
  not_8  g08947(.A(new_n11295), .Y(new_n11296));
  nor_5  g08948(.A(new_n11296), .B(new_n11289), .Y(new_n11297));
  xnor_4 g08949(.A(new_n11296), .B(new_n11289), .Y(new_n11298));
  nor_5  g08950(.A(new_n6789), .B(new_n2558), .Y(new_n11299));
  xnor_4 g08951(.A(new_n6789), .B(new_n2558), .Y(new_n11300));
  nor_5  g08952(.A(new_n6791_1), .B(n18345), .Y(new_n11301));
  xnor_4 g08953(.A(new_n6791_1), .B(n18345), .Y(new_n11302_1));
  nor_5  g08954(.A(new_n6794_1), .B(n13190), .Y(new_n11303));
  xnor_4 g08955(.A(new_n6794_1), .B(new_n2566), .Y(new_n11304));
  not_8  g08956(.A(n3460), .Y(new_n11305));
  nor_5  g08957(.A(new_n6798), .B(new_n11305), .Y(new_n11306));
  nor_5  g08958(.A(new_n6802_1), .B(new_n9502), .Y(new_n11307));
  nor_5  g08959(.A(new_n9516), .B(new_n9503), .Y(new_n11308));
  nor_5  g08960(.A(new_n11308), .B(new_n11307), .Y(new_n11309));
  xnor_4 g08961(.A(new_n6798), .B(new_n11305), .Y(new_n11310));
  nor_5  g08962(.A(new_n11310), .B(new_n11309), .Y(new_n11311));
  nor_5  g08963(.A(new_n11311), .B(new_n11306), .Y(new_n11312));
  and_5  g08964(.A(new_n11312), .B(new_n11304), .Y(new_n11313_1));
  nor_5  g08965(.A(new_n11313_1), .B(new_n11303), .Y(new_n11314));
  nor_5  g08966(.A(new_n11314), .B(new_n11302_1), .Y(new_n11315));
  or_5   g08967(.A(new_n11315), .B(new_n11301), .Y(new_n11316));
  nor_5  g08968(.A(new_n11316), .B(new_n11300), .Y(new_n11317));
  nor_5  g08969(.A(new_n11317), .B(new_n11299), .Y(new_n11318));
  nor_5  g08970(.A(new_n11318), .B(new_n11298), .Y(new_n11319));
  nor_5  g08971(.A(new_n11319), .B(new_n11297), .Y(new_n11320));
  nor_5  g08972(.A(n18880), .B(n2978), .Y(new_n11321));
  nor_5  g08973(.A(new_n11294), .B(new_n11291), .Y(new_n11322));
  nor_5  g08974(.A(new_n11322), .B(new_n11321), .Y(new_n11323));
  xnor_4 g08975(.A(new_n11323), .B(new_n11320), .Y(new_n11324));
  not_8  g08976(.A(n7569), .Y(new_n11325_1));
  not_8  g08977(.A(n17037), .Y(new_n11326_1));
  not_8  g08978(.A(new_n9500), .Y(new_n11327));
  nor_5  g08979(.A(new_n11327), .B(n19575), .Y(new_n11328));
  not_8  g08980(.A(new_n11328), .Y(new_n11329));
  nor_5  g08981(.A(new_n11329), .B(n26512), .Y(new_n11330_1));
  not_8  g08982(.A(new_n11330_1), .Y(new_n11331));
  nor_5  g08983(.A(new_n11331), .B(n26191), .Y(new_n11332));
  not_8  g08984(.A(new_n11332), .Y(new_n11333));
  nor_5  g08985(.A(new_n11333), .B(n5386), .Y(new_n11334));
  and_5  g08986(.A(new_n11334), .B(new_n11326_1), .Y(new_n11335));
  and_5  g08987(.A(new_n11335), .B(new_n11325_1), .Y(new_n11336));
  xnor_4 g08988(.A(new_n11336), .B(new_n11324), .Y(new_n11337));
  xnor_4 g08989(.A(new_n11318), .B(new_n11298), .Y(new_n11338));
  not_8  g08990(.A(new_n11338), .Y(new_n11339));
  xnor_4 g08991(.A(new_n11335), .B(n7569), .Y(new_n11340));
  nor_5  g08992(.A(new_n11340), .B(new_n11339), .Y(new_n11341));
  xnor_4 g08993(.A(new_n11340), .B(new_n11339), .Y(new_n11342));
  nor_5  g08994(.A(new_n11315), .B(new_n11301), .Y(new_n11343));
  xnor_4 g08995(.A(new_n11343), .B(new_n11300), .Y(new_n11344));
  xnor_4 g08996(.A(new_n11334), .B(n17037), .Y(new_n11345));
  nor_5  g08997(.A(new_n11345), .B(new_n11344), .Y(new_n11346));
  xnor_4 g08998(.A(new_n11345), .B(new_n11344), .Y(new_n11347_1));
  xnor_4 g08999(.A(new_n11314), .B(new_n11302_1), .Y(new_n11348_1));
  xnor_4 g09000(.A(new_n11332), .B(n5386), .Y(new_n11349));
  nor_5  g09001(.A(new_n11349), .B(new_n11348_1), .Y(new_n11350));
  xnor_4 g09002(.A(new_n11349), .B(new_n11348_1), .Y(new_n11351));
  xnor_4 g09003(.A(new_n11312), .B(new_n11304), .Y(new_n11352_1));
  xnor_4 g09004(.A(new_n11330_1), .B(n26191), .Y(new_n11353));
  nor_5  g09005(.A(new_n11353), .B(new_n11352_1), .Y(new_n11354));
  xnor_4 g09006(.A(new_n11328), .B(n26512), .Y(new_n11355));
  not_8  g09007(.A(new_n11355), .Y(new_n11356_1));
  xor_4  g09008(.A(new_n11310), .B(new_n11309), .Y(new_n11357));
  not_8  g09009(.A(new_n11357), .Y(new_n11358));
  nor_5  g09010(.A(new_n11358), .B(new_n11356_1), .Y(new_n11359));
  xnor_4 g09011(.A(new_n11358), .B(new_n11356_1), .Y(new_n11360));
  nor_5  g09012(.A(new_n9517), .B(new_n9501), .Y(new_n11361));
  and_5  g09013(.A(new_n9542), .B(new_n9519), .Y(new_n11362));
  or_5   g09014(.A(new_n11362), .B(new_n11361), .Y(new_n11363));
  nor_5  g09015(.A(new_n11363), .B(new_n11360), .Y(new_n11364));
  nor_5  g09016(.A(new_n11364), .B(new_n11359), .Y(new_n11365));
  not_8  g09017(.A(new_n11352_1), .Y(new_n11366));
  xnor_4 g09018(.A(new_n11353), .B(new_n11366), .Y(new_n11367));
  and_5  g09019(.A(new_n11367), .B(new_n11365), .Y(new_n11368));
  nor_5  g09020(.A(new_n11368), .B(new_n11354), .Y(new_n11369));
  nor_5  g09021(.A(new_n11369), .B(new_n11351), .Y(new_n11370));
  nor_5  g09022(.A(new_n11370), .B(new_n11350), .Y(new_n11371));
  nor_5  g09023(.A(new_n11371), .B(new_n11347_1), .Y(new_n11372));
  nor_5  g09024(.A(new_n11372), .B(new_n11346), .Y(new_n11373));
  nor_5  g09025(.A(new_n11373), .B(new_n11342), .Y(new_n11374));
  nor_5  g09026(.A(new_n11374), .B(new_n11341), .Y(new_n11375_1));
  xnor_4 g09027(.A(new_n11375_1), .B(new_n11337), .Y(new_n11376));
  xnor_4 g09028(.A(new_n11376), .B(new_n11288), .Y(new_n11377));
  xor_4  g09029(.A(new_n11373), .B(new_n11342), .Y(new_n11378));
  xor_4  g09030(.A(new_n11286), .B(new_n11274), .Y(new_n11379_1));
  not_8  g09031(.A(new_n11379_1), .Y(new_n11380));
  and_5  g09032(.A(new_n11380), .B(new_n11378), .Y(new_n11381));
  xnor_4 g09033(.A(new_n11380), .B(new_n11378), .Y(new_n11382));
  xnor_4 g09034(.A(new_n11371), .B(new_n11347_1), .Y(new_n11383));
  xnor_4 g09035(.A(new_n11284), .B(new_n11277), .Y(new_n11384));
  not_8  g09036(.A(new_n11384), .Y(new_n11385));
  nor_5  g09037(.A(new_n11385), .B(new_n11383), .Y(new_n11386_1));
  xnor_4 g09038(.A(new_n11385), .B(new_n11383), .Y(new_n11387));
  xor_4  g09039(.A(new_n11369), .B(new_n11351), .Y(new_n11388));
  not_8  g09040(.A(n6218), .Y(new_n11389));
  xnor_4 g09041(.A(n19652), .B(new_n11389), .Y(new_n11390));
  xnor_4 g09042(.A(new_n11390), .B(new_n11282), .Y(new_n11391_1));
  not_8  g09043(.A(new_n11391_1), .Y(new_n11392));
  and_5  g09044(.A(new_n11392), .B(new_n11388), .Y(new_n11393));
  xnor_4 g09045(.A(new_n11392), .B(new_n11388), .Y(new_n11394));
  xnor_4 g09046(.A(new_n11367), .B(new_n11365), .Y(new_n11395));
  nor_5  g09047(.A(new_n11395), .B(new_n10834_1), .Y(new_n11396));
  xnor_4 g09048(.A(new_n11395), .B(new_n10834_1), .Y(new_n11397));
  xor_4  g09049(.A(new_n11363), .B(new_n11360), .Y(new_n11398_1));
  and_5  g09050(.A(new_n11398_1), .B(new_n10839), .Y(new_n11399));
  nor_5  g09051(.A(new_n11398_1), .B(new_n10839), .Y(new_n11400));
  nor_5  g09052(.A(new_n9543), .B(new_n10843), .Y(new_n11401));
  and_5  g09053(.A(new_n9567), .B(new_n9544), .Y(new_n11402));
  nor_5  g09054(.A(new_n11402), .B(new_n11401), .Y(new_n11403_1));
  nor_5  g09055(.A(new_n11403_1), .B(new_n11400), .Y(new_n11404));
  or_5   g09056(.A(new_n11404), .B(new_n11399), .Y(new_n11405));
  nor_5  g09057(.A(new_n11405), .B(new_n11397), .Y(new_n11406));
  nor_5  g09058(.A(new_n11406), .B(new_n11396), .Y(new_n11407));
  nor_5  g09059(.A(new_n11407), .B(new_n11394), .Y(new_n11408));
  nor_5  g09060(.A(new_n11408), .B(new_n11393), .Y(new_n11409));
  nor_5  g09061(.A(new_n11409), .B(new_n11387), .Y(new_n11410));
  nor_5  g09062(.A(new_n11410), .B(new_n11386_1), .Y(new_n11411));
  nor_5  g09063(.A(new_n11411), .B(new_n11382), .Y(new_n11412));
  nor_5  g09064(.A(new_n11412), .B(new_n11381), .Y(new_n11413));
  xnor_4 g09065(.A(new_n11413), .B(new_n11377), .Y(n1684));
  xnor_4 g09066(.A(new_n6216), .B(n3984), .Y(new_n11415));
  nor_5  g09067(.A(new_n6218_1), .B(n19652), .Y(new_n11416));
  xnor_4 g09068(.A(new_n6220), .B(n19652), .Y(new_n11417));
  nor_5  g09069(.A(new_n6223_1), .B(n3366), .Y(new_n11418));
  xnor_4 g09070(.A(new_n6224), .B(n3366), .Y(new_n11419_1));
  nor_5  g09071(.A(new_n4012), .B(n26565), .Y(new_n11420));
  xnor_4 g09072(.A(new_n4013), .B(n26565), .Y(new_n11421));
  nor_5  g09073(.A(new_n4016), .B(n3959), .Y(new_n11422));
  xnor_4 g09074(.A(new_n4017), .B(n3959), .Y(new_n11423));
  nor_5  g09075(.A(new_n4019), .B(n11566), .Y(new_n11424_1));
  xor_4  g09076(.A(new_n4019), .B(n11566), .Y(new_n11425));
  nor_5  g09077(.A(new_n4023), .B(n26744), .Y(new_n11426));
  xnor_4 g09078(.A(new_n4025), .B(n26744), .Y(new_n11427));
  nor_5  g09079(.A(new_n4028), .B(n26625), .Y(new_n11428));
  or_5   g09080(.A(new_n4031), .B(new_n9484), .Y(new_n11429));
  xnor_4 g09081(.A(new_n4027), .B(n26625), .Y(new_n11430));
  and_5  g09082(.A(new_n11430), .B(new_n11429), .Y(new_n11431));
  or_5   g09083(.A(new_n11431), .B(new_n11428), .Y(new_n11432));
  and_5  g09084(.A(new_n11432), .B(new_n11427), .Y(new_n11433));
  or_5   g09085(.A(new_n11433), .B(new_n11426), .Y(new_n11434));
  and_5  g09086(.A(new_n11434), .B(new_n11425), .Y(new_n11435));
  or_5   g09087(.A(new_n11435), .B(new_n11424_1), .Y(new_n11436));
  and_5  g09088(.A(new_n11436), .B(new_n11423), .Y(new_n11437));
  or_5   g09089(.A(new_n11437), .B(new_n11422), .Y(new_n11438));
  and_5  g09090(.A(new_n11438), .B(new_n11421), .Y(new_n11439_1));
  or_5   g09091(.A(new_n11439_1), .B(new_n11420), .Y(new_n11440));
  and_5  g09092(.A(new_n11440), .B(new_n11419_1), .Y(new_n11441));
  or_5   g09093(.A(new_n11441), .B(new_n11418), .Y(new_n11442));
  and_5  g09094(.A(new_n11442), .B(new_n11417), .Y(new_n11443));
  or_5   g09095(.A(new_n11443), .B(new_n11416), .Y(new_n11444));
  xor_4  g09096(.A(new_n11444), .B(new_n11415), .Y(new_n11445));
  nor_5  g09097(.A(new_n11445), .B(n13026), .Y(new_n11446));
  xor_4  g09098(.A(new_n11445), .B(n13026), .Y(new_n11447));
  xor_4  g09099(.A(new_n11442), .B(new_n11417), .Y(new_n11448));
  nor_5  g09100(.A(new_n11448), .B(n2175), .Y(new_n11449));
  xor_4  g09101(.A(new_n11448), .B(n2175), .Y(new_n11450));
  xor_4  g09102(.A(new_n11440), .B(new_n11419_1), .Y(new_n11451));
  nor_5  g09103(.A(new_n11451), .B(n752), .Y(new_n11452));
  xnor_4 g09104(.A(new_n11451), .B(n752), .Y(new_n11453));
  xor_4  g09105(.A(new_n11438), .B(new_n11421), .Y(new_n11454));
  nor_5  g09106(.A(new_n11454), .B(n1611), .Y(new_n11455_1));
  xor_4  g09107(.A(new_n11436), .B(new_n11423), .Y(new_n11456));
  nor_5  g09108(.A(new_n11456), .B(n25094), .Y(new_n11457));
  xnor_4 g09109(.A(new_n11456), .B(n25094), .Y(new_n11458));
  xor_4  g09110(.A(new_n11434), .B(new_n11425), .Y(new_n11459));
  nor_5  g09111(.A(new_n11459), .B(n21538), .Y(new_n11460));
  xnor_4 g09112(.A(new_n11459), .B(n21538), .Y(new_n11461));
  xor_4  g09113(.A(new_n11432), .B(new_n11427), .Y(new_n11462_1));
  nor_5  g09114(.A(new_n11462_1), .B(n5131), .Y(new_n11463));
  xor_4  g09115(.A(new_n11430), .B(new_n11429), .Y(new_n11464));
  nor_5  g09116(.A(new_n11464), .B(n11473), .Y(new_n11465));
  xnor_4 g09117(.A(n19922), .B(new_n9484), .Y(new_n11466));
  or_5   g09118(.A(new_n11466), .B(new_n10803), .Y(new_n11467));
  xnor_4 g09119(.A(new_n11464), .B(new_n10809), .Y(new_n11468));
  and_5  g09120(.A(new_n11468), .B(new_n11467), .Y(new_n11469));
  nor_5  g09121(.A(new_n11469), .B(new_n11465), .Y(new_n11470_1));
  xnor_4 g09122(.A(new_n11462_1), .B(n5131), .Y(new_n11471));
  nor_5  g09123(.A(new_n11471), .B(new_n11470_1), .Y(new_n11472_1));
  nor_5  g09124(.A(new_n11472_1), .B(new_n11463), .Y(new_n11473_1));
  nor_5  g09125(.A(new_n11473_1), .B(new_n11461), .Y(new_n11474));
  nor_5  g09126(.A(new_n11474), .B(new_n11460), .Y(new_n11475));
  nor_5  g09127(.A(new_n11475), .B(new_n11458), .Y(new_n11476));
  nor_5  g09128(.A(new_n11476), .B(new_n11457), .Y(new_n11477));
  xnor_4 g09129(.A(new_n11454), .B(n1611), .Y(new_n11478));
  nor_5  g09130(.A(new_n11478), .B(new_n11477), .Y(new_n11479_1));
  nor_5  g09131(.A(new_n11479_1), .B(new_n11455_1), .Y(new_n11480));
  nor_5  g09132(.A(new_n11480), .B(new_n11453), .Y(new_n11481_1));
  or_5   g09133(.A(new_n11481_1), .B(new_n11452), .Y(new_n11482));
  and_5  g09134(.A(new_n11482), .B(new_n11450), .Y(new_n11483));
  or_5   g09135(.A(new_n11483), .B(new_n11449), .Y(new_n11484));
  and_5  g09136(.A(new_n11484), .B(new_n11447), .Y(new_n11485));
  nor_5  g09137(.A(new_n11485), .B(new_n11446), .Y(new_n11486_1));
  and_5  g09138(.A(new_n11486_1), .B(n23912), .Y(new_n11487));
  xnor_4 g09139(.A(new_n11486_1), .B(n23912), .Y(new_n11488));
  nor_5  g09140(.A(new_n6213), .B(n3984), .Y(new_n11489));
  and_5  g09141(.A(new_n11444), .B(new_n11415), .Y(new_n11490));
  nor_5  g09142(.A(new_n11490), .B(new_n11489), .Y(new_n11491));
  not_8  g09143(.A(new_n11491), .Y(new_n11492));
  xnor_4 g09144(.A(new_n6208), .B(n4514), .Y(new_n11493));
  xnor_4 g09145(.A(new_n11493), .B(new_n11492), .Y(new_n11494));
  nor_5  g09146(.A(new_n11494), .B(new_n11488), .Y(new_n11495));
  nor_5  g09147(.A(new_n11495), .B(new_n11487), .Y(new_n11496_1));
  nor_5  g09148(.A(new_n6208), .B(new_n11273_1), .Y(new_n11497));
  nor_5  g09149(.A(new_n6207), .B(n4514), .Y(new_n11498));
  nor_5  g09150(.A(new_n11498), .B(new_n11492), .Y(new_n11499));
  or_5   g09151(.A(new_n11499), .B(new_n6211), .Y(new_n11500));
  or_5   g09152(.A(new_n11500), .B(new_n11497), .Y(new_n11501));
  and_5  g09153(.A(new_n11501), .B(new_n11496_1), .Y(new_n11502));
  nor_5  g09154(.A(new_n4477), .B(n15766), .Y(new_n11503_1));
  xnor_4 g09155(.A(new_n4477), .B(new_n6320), .Y(new_n11504));
  nor_5  g09156(.A(new_n4482), .B(n25629), .Y(new_n11505));
  xnor_4 g09157(.A(new_n4481), .B(n25629), .Y(new_n11506_1));
  nor_5  g09158(.A(new_n4488), .B(n7692), .Y(new_n11507));
  xnor_4 g09159(.A(new_n4488), .B(new_n6326), .Y(new_n11508));
  nor_5  g09160(.A(new_n4493), .B(n23039), .Y(new_n11509));
  xnor_4 g09161(.A(new_n4493), .B(n23039), .Y(new_n11510));
  nor_5  g09162(.A(new_n3963), .B(n13677), .Y(new_n11511));
  nor_5  g09163(.A(new_n3995), .B(new_n3964), .Y(new_n11512));
  nor_5  g09164(.A(new_n11512), .B(new_n11511), .Y(new_n11513));
  nor_5  g09165(.A(new_n11513), .B(new_n11510), .Y(new_n11514));
  or_5   g09166(.A(new_n11514), .B(new_n11509), .Y(new_n11515_1));
  and_5  g09167(.A(new_n11515_1), .B(new_n11508), .Y(new_n11516));
  or_5   g09168(.A(new_n11516), .B(new_n11507), .Y(new_n11517));
  and_5  g09169(.A(new_n11517), .B(new_n11506_1), .Y(new_n11518));
  or_5   g09170(.A(new_n11518), .B(new_n11505), .Y(new_n11519));
  and_5  g09171(.A(new_n11519), .B(new_n11504), .Y(new_n11520));
  nor_5  g09172(.A(new_n11520), .B(new_n11503_1), .Y(new_n11521));
  not_8  g09173(.A(new_n11521), .Y(new_n11522));
  nor_5  g09174(.A(new_n11522), .B(new_n4538), .Y(new_n11523));
  not_8  g09175(.A(new_n11523), .Y(new_n11524));
  xnor_4 g09176(.A(new_n11522), .B(new_n4453), .Y(new_n11525));
  xor_4  g09177(.A(new_n11501), .B(new_n11496_1), .Y(new_n11526));
  nor_5  g09178(.A(new_n11526), .B(new_n11525), .Y(new_n11527));
  xnor_4 g09179(.A(new_n11526), .B(new_n11525), .Y(new_n11528));
  xor_4  g09180(.A(new_n11519), .B(new_n11504), .Y(new_n11529));
  not_8  g09181(.A(new_n11529), .Y(new_n11530));
  xnor_4 g09182(.A(new_n11494), .B(new_n11488), .Y(new_n11531));
  nor_5  g09183(.A(new_n11531), .B(new_n11530), .Y(new_n11532));
  xor_4  g09184(.A(new_n11517), .B(new_n11506_1), .Y(new_n11533));
  not_8  g09185(.A(new_n11533), .Y(new_n11534));
  xor_4  g09186(.A(new_n11484), .B(new_n11447), .Y(new_n11535));
  nor_5  g09187(.A(new_n11535), .B(new_n11534), .Y(new_n11536));
  xnor_4 g09188(.A(new_n11535), .B(new_n11534), .Y(new_n11537));
  xor_4  g09189(.A(new_n11515_1), .B(new_n11508), .Y(new_n11538_1));
  not_8  g09190(.A(new_n11538_1), .Y(new_n11539));
  xor_4  g09191(.A(new_n11482), .B(new_n11450), .Y(new_n11540));
  nor_5  g09192(.A(new_n11540), .B(new_n11539), .Y(new_n11541));
  xnor_4 g09193(.A(new_n11540), .B(new_n11539), .Y(new_n11542));
  xnor_4 g09194(.A(new_n11513), .B(new_n11510), .Y(new_n11543));
  xor_4  g09195(.A(new_n11480), .B(new_n11453), .Y(new_n11544));
  nor_5  g09196(.A(new_n11544), .B(new_n11543), .Y(new_n11545));
  xnor_4 g09197(.A(new_n11544), .B(new_n11543), .Y(new_n11546));
  xor_4  g09198(.A(new_n11478), .B(new_n11477), .Y(new_n11547));
  nor_5  g09199(.A(new_n11547), .B(new_n3996), .Y(new_n11548_1));
  xnor_4 g09200(.A(new_n11547), .B(new_n3996), .Y(new_n11549));
  not_8  g09201(.A(new_n4080), .Y(new_n11550));
  xor_4  g09202(.A(new_n11475), .B(new_n11458), .Y(new_n11551));
  nor_5  g09203(.A(new_n11551), .B(new_n11550), .Y(new_n11552));
  xor_4  g09204(.A(new_n11473_1), .B(new_n11461), .Y(new_n11553));
  nor_5  g09205(.A(new_n11553), .B(new_n4084), .Y(new_n11554));
  xnor_4 g09206(.A(new_n11553), .B(new_n4084), .Y(new_n11555));
  xor_4  g09207(.A(new_n11471), .B(new_n11470_1), .Y(new_n11556));
  nor_5  g09208(.A(new_n11556), .B(new_n4087), .Y(new_n11557));
  xor_4  g09209(.A(new_n11468), .B(new_n11467), .Y(new_n11558));
  nor_5  g09210(.A(new_n11558), .B(new_n4092), .Y(new_n11559));
  xnor_4 g09211(.A(new_n11466), .B(n15506), .Y(new_n11560));
  nor_5  g09212(.A(new_n11560), .B(new_n4094), .Y(new_n11561));
  xnor_4 g09213(.A(new_n11558), .B(new_n4092), .Y(new_n11562));
  nor_5  g09214(.A(new_n11562), .B(new_n11561), .Y(new_n11563));
  nor_5  g09215(.A(new_n11563), .B(new_n11559), .Y(new_n11564_1));
  xnor_4 g09216(.A(new_n11556), .B(new_n4087), .Y(new_n11565));
  nor_5  g09217(.A(new_n11565), .B(new_n11564_1), .Y(new_n11566_1));
  nor_5  g09218(.A(new_n11566_1), .B(new_n11557), .Y(new_n11567));
  nor_5  g09219(.A(new_n11567), .B(new_n11555), .Y(new_n11568));
  nor_5  g09220(.A(new_n11568), .B(new_n11554), .Y(new_n11569));
  xnor_4 g09221(.A(new_n11551), .B(new_n11550), .Y(new_n11570));
  nor_5  g09222(.A(new_n11570), .B(new_n11569), .Y(new_n11571));
  nor_5  g09223(.A(new_n11571), .B(new_n11552), .Y(new_n11572));
  nor_5  g09224(.A(new_n11572), .B(new_n11549), .Y(new_n11573));
  nor_5  g09225(.A(new_n11573), .B(new_n11548_1), .Y(new_n11574));
  nor_5  g09226(.A(new_n11574), .B(new_n11546), .Y(new_n11575));
  nor_5  g09227(.A(new_n11575), .B(new_n11545), .Y(new_n11576));
  nor_5  g09228(.A(new_n11576), .B(new_n11542), .Y(new_n11577));
  nor_5  g09229(.A(new_n11577), .B(new_n11541), .Y(new_n11578));
  nor_5  g09230(.A(new_n11578), .B(new_n11537), .Y(new_n11579_1));
  nor_5  g09231(.A(new_n11579_1), .B(new_n11536), .Y(new_n11580_1));
  xnor_4 g09232(.A(new_n11531), .B(new_n11530), .Y(new_n11581));
  nor_5  g09233(.A(new_n11581), .B(new_n11580_1), .Y(new_n11582));
  nor_5  g09234(.A(new_n11582), .B(new_n11532), .Y(new_n11583));
  nor_5  g09235(.A(new_n11583), .B(new_n11528), .Y(new_n11584));
  nor_5  g09236(.A(new_n11584), .B(new_n11527), .Y(new_n11585));
  xnor_4 g09237(.A(new_n11585), .B(new_n11524), .Y(new_n11586));
  xnor_4 g09238(.A(new_n11586), .B(new_n11502), .Y(n1701));
  xnor_4 g09239(.A(new_n3924), .B(new_n3894), .Y(n1703));
  xnor_4 g09240(.A(new_n4604), .B(new_n4551), .Y(n1721));
  nor_5  g09241(.A(new_n7694), .B(new_n4353), .Y(new_n11590));
  and_5  g09242(.A(new_n8952), .B(new_n8951), .Y(new_n11591_1));
  nor_5  g09243(.A(new_n11591_1), .B(new_n11590), .Y(new_n11592));
  not_8  g09244(.A(new_n11592), .Y(new_n11593));
  and_5  g09245(.A(new_n11593), .B(new_n8996), .Y(new_n11594));
  nor_5  g09246(.A(new_n8996), .B(new_n8953), .Y(new_n11595));
  nor_5  g09247(.A(new_n9059), .B(new_n8997), .Y(new_n11596));
  nor_5  g09248(.A(new_n11596), .B(new_n11595), .Y(new_n11597));
  nor_5  g09249(.A(new_n11597), .B(new_n11594), .Y(new_n11598));
  nor_5  g09250(.A(new_n11593), .B(new_n8996), .Y(new_n11599));
  nor_5  g09251(.A(new_n11599), .B(new_n11596), .Y(new_n11600));
  nor_5  g09252(.A(new_n11600), .B(new_n11598), .Y(n1760));
  xnor_4 g09253(.A(new_n4098), .B(new_n4090), .Y(n1791));
  xnor_4 g09254(.A(n23333), .B(n16502), .Y(new_n11603));
  xnor_4 g09255(.A(new_n3368), .B(new_n11603), .Y(n1808));
  nor_5  g09256(.A(new_n7695), .B(new_n7650), .Y(new_n11605));
  nor_5  g09257(.A(new_n7769_1), .B(new_n7696), .Y(new_n11606));
  nor_5  g09258(.A(new_n11606), .B(new_n11605), .Y(new_n11607_1));
  nor_5  g09259(.A(n13494), .B(new_n3087), .Y(new_n11608));
  xnor_4 g09260(.A(n13494), .B(n4319), .Y(new_n11609));
  not_8  g09261(.A(n23463), .Y(new_n11610));
  nor_5  g09262(.A(n25345), .B(new_n11610), .Y(new_n11611));
  and_5  g09263(.A(new_n11115), .B(new_n11092), .Y(new_n11612));
  or_5   g09264(.A(new_n11612), .B(new_n11611), .Y(new_n11613));
  and_5  g09265(.A(new_n11613), .B(new_n11609), .Y(new_n11614));
  nor_5  g09266(.A(new_n11614), .B(new_n11608), .Y(new_n11615_1));
  and_5  g09267(.A(new_n11615_1), .B(new_n11607_1), .Y(new_n11616));
  nor_5  g09268(.A(new_n11615_1), .B(new_n7770), .Y(new_n11617));
  xnor_4 g09269(.A(new_n11615_1), .B(new_n7771), .Y(new_n11618));
  xor_4  g09270(.A(new_n11613), .B(new_n11609), .Y(new_n11619));
  and_5  g09271(.A(new_n11619), .B(new_n7837), .Y(new_n11620));
  xnor_4 g09272(.A(new_n11619), .B(new_n7842), .Y(new_n11621));
  and_5  g09273(.A(new_n11116), .B(new_n7844), .Y(new_n11622));
  and_5  g09274(.A(new_n11145), .B(new_n11117), .Y(new_n11623));
  or_5   g09275(.A(new_n11623), .B(new_n11622), .Y(new_n11624));
  and_5  g09276(.A(new_n11624), .B(new_n11621), .Y(new_n11625));
  nor_5  g09277(.A(new_n11625), .B(new_n11620), .Y(new_n11626));
  and_5  g09278(.A(new_n11626), .B(new_n11618), .Y(new_n11627));
  nor_5  g09279(.A(new_n11627), .B(new_n11617), .Y(new_n11628));
  nor_5  g09280(.A(new_n11628), .B(new_n11616), .Y(new_n11629));
  nor_5  g09281(.A(new_n11615_1), .B(new_n11607_1), .Y(new_n11630_1));
  nor_5  g09282(.A(new_n11630_1), .B(new_n11627), .Y(new_n11631));
  nor_5  g09283(.A(new_n11631), .B(new_n11629), .Y(n1821));
  xnor_4 g09284(.A(new_n6948), .B(new_n6947), .Y(n1832));
  xnor_4 g09285(.A(n9934), .B(new_n7179), .Y(new_n11634));
  nor_5  g09286(.A(n25331), .B(n18496), .Y(new_n11635));
  not_8  g09287(.A(n18496), .Y(new_n11636));
  xnor_4 g09288(.A(n25331), .B(new_n11636), .Y(new_n11637));
  nor_5  g09289(.A(n26224), .B(n18483), .Y(new_n11638));
  xnor_4 g09290(.A(n26224), .B(n18483), .Y(new_n11639));
  nor_5  g09291(.A(n21934), .B(n19327), .Y(new_n11640));
  xnor_4 g09292(.A(n21934), .B(n19327), .Y(new_n11641));
  nor_5  g09293(.A(n22597), .B(n18901), .Y(new_n11642));
  xnor_4 g09294(.A(n22597), .B(n18901), .Y(new_n11643));
  nor_5  g09295(.A(n26107), .B(n4376), .Y(new_n11644));
  xnor_4 g09296(.A(n26107), .B(n4376), .Y(new_n11645));
  nor_5  g09297(.A(n14570), .B(n342), .Y(new_n11646));
  xnor_4 g09298(.A(n14570), .B(n342), .Y(new_n11647_1));
  nor_5  g09299(.A(n26553), .B(n23775), .Y(new_n11648));
  xnor_4 g09300(.A(n26553), .B(n23775), .Y(new_n11649));
  nor_5  g09301(.A(n8259), .B(n4964), .Y(new_n11650));
  not_8  g09302(.A(n11479), .Y(new_n11651));
  or_5   g09303(.A(new_n11651), .B(new_n3755_1), .Y(new_n11652));
  xnor_4 g09304(.A(n8259), .B(new_n4776), .Y(new_n11653));
  and_5  g09305(.A(new_n11653), .B(new_n11652), .Y(new_n11654));
  nor_5  g09306(.A(new_n11654), .B(new_n11650), .Y(new_n11655));
  nor_5  g09307(.A(new_n11655), .B(new_n11649), .Y(new_n11656));
  nor_5  g09308(.A(new_n11656), .B(new_n11648), .Y(new_n11657));
  nor_5  g09309(.A(new_n11657), .B(new_n11647_1), .Y(new_n11658));
  nor_5  g09310(.A(new_n11658), .B(new_n11646), .Y(new_n11659));
  nor_5  g09311(.A(new_n11659), .B(new_n11645), .Y(new_n11660));
  nor_5  g09312(.A(new_n11660), .B(new_n11644), .Y(new_n11661));
  nor_5  g09313(.A(new_n11661), .B(new_n11643), .Y(new_n11662));
  nor_5  g09314(.A(new_n11662), .B(new_n11642), .Y(new_n11663));
  nor_5  g09315(.A(new_n11663), .B(new_n11641), .Y(new_n11664));
  nor_5  g09316(.A(new_n11664), .B(new_n11640), .Y(new_n11665));
  nor_5  g09317(.A(new_n11665), .B(new_n11639), .Y(new_n11666));
  or_5   g09318(.A(new_n11666), .B(new_n11638), .Y(new_n11667_1));
  and_5  g09319(.A(new_n11667_1), .B(new_n11637), .Y(new_n11668));
  or_5   g09320(.A(new_n11668), .B(new_n11635), .Y(new_n11669));
  xor_4  g09321(.A(new_n11669), .B(new_n11634), .Y(new_n11670));
  xnor_4 g09322(.A(new_n11670), .B(n2160), .Y(new_n11671));
  xor_4  g09323(.A(new_n11667_1), .B(new_n11637), .Y(new_n11672));
  nor_5  g09324(.A(new_n11672), .B(n10763), .Y(new_n11673));
  not_8  g09325(.A(n10763), .Y(new_n11674_1));
  xnor_4 g09326(.A(new_n11672), .B(new_n11674_1), .Y(new_n11675));
  xnor_4 g09327(.A(new_n11665), .B(new_n11639), .Y(new_n11676));
  nor_5  g09328(.A(new_n11676), .B(new_n2890), .Y(new_n11677));
  xnor_4 g09329(.A(new_n11676), .B(new_n2890), .Y(new_n11678));
  xnor_4 g09330(.A(new_n11663), .B(new_n11641), .Y(new_n11679));
  nor_5  g09331(.A(new_n11679), .B(new_n2893), .Y(new_n11680));
  xnor_4 g09332(.A(new_n11679), .B(new_n2893), .Y(new_n11681));
  xnor_4 g09333(.A(new_n11661), .B(new_n11643), .Y(new_n11682_1));
  nor_5  g09334(.A(new_n11682_1), .B(new_n2896), .Y(new_n11683));
  xnor_4 g09335(.A(new_n11682_1), .B(new_n2896), .Y(new_n11684));
  not_8  g09336(.A(n12811), .Y(new_n11685));
  xnor_4 g09337(.A(new_n11659), .B(new_n11645), .Y(new_n11686));
  nor_5  g09338(.A(new_n11686), .B(new_n11685), .Y(new_n11687));
  xnor_4 g09339(.A(new_n11686), .B(new_n11685), .Y(new_n11688));
  not_8  g09340(.A(n1118), .Y(new_n11689));
  xnor_4 g09341(.A(new_n11657), .B(new_n11647_1), .Y(new_n11690));
  nor_5  g09342(.A(new_n11690), .B(new_n11689), .Y(new_n11691));
  xnor_4 g09343(.A(new_n11690), .B(new_n11689), .Y(new_n11692));
  not_8  g09344(.A(n25974), .Y(new_n11693));
  xnor_4 g09345(.A(new_n11655), .B(new_n11649), .Y(new_n11694));
  nor_5  g09346(.A(new_n11694), .B(new_n11693), .Y(new_n11695));
  xnor_4 g09347(.A(new_n11694), .B(n25974), .Y(new_n11696));
  xnor_4 g09348(.A(n11479), .B(new_n3755_1), .Y(new_n11697));
  nor_5  g09349(.A(new_n11697), .B(new_n2906), .Y(new_n11698));
  nor_5  g09350(.A(new_n11698), .B(n1630), .Y(new_n11699));
  xor_4  g09351(.A(new_n11653), .B(new_n11652), .Y(new_n11700));
  xnor_4 g09352(.A(new_n11698), .B(new_n2909), .Y(new_n11701));
  not_8  g09353(.A(new_n11701), .Y(new_n11702));
  nor_5  g09354(.A(new_n11702), .B(new_n11700), .Y(new_n11703));
  nor_5  g09355(.A(new_n11703), .B(new_n11699), .Y(new_n11704));
  and_5  g09356(.A(new_n11704), .B(new_n11696), .Y(new_n11705));
  nor_5  g09357(.A(new_n11705), .B(new_n11695), .Y(new_n11706));
  nor_5  g09358(.A(new_n11706), .B(new_n11692), .Y(new_n11707));
  nor_5  g09359(.A(new_n11707), .B(new_n11691), .Y(new_n11708));
  nor_5  g09360(.A(new_n11708), .B(new_n11688), .Y(new_n11709));
  nor_5  g09361(.A(new_n11709), .B(new_n11687), .Y(new_n11710_1));
  nor_5  g09362(.A(new_n11710_1), .B(new_n11684), .Y(new_n11711));
  nor_5  g09363(.A(new_n11711), .B(new_n11683), .Y(new_n11712_1));
  nor_5  g09364(.A(new_n11712_1), .B(new_n11681), .Y(new_n11713));
  nor_5  g09365(.A(new_n11713), .B(new_n11680), .Y(new_n11714));
  nor_5  g09366(.A(new_n11714), .B(new_n11678), .Y(new_n11715));
  nor_5  g09367(.A(new_n11715), .B(new_n11677), .Y(new_n11716));
  and_5  g09368(.A(new_n11716), .B(new_n11675), .Y(new_n11717));
  nor_5  g09369(.A(new_n11717), .B(new_n11673), .Y(new_n11718));
  xnor_4 g09370(.A(new_n11718), .B(new_n11671), .Y(new_n11719));
  not_8  g09371(.A(new_n3849), .Y(new_n11720));
  nor_5  g09372(.A(new_n11720), .B(n4325), .Y(new_n11721));
  not_8  g09373(.A(new_n11721), .Y(new_n11722));
  nor_5  g09374(.A(new_n11722), .B(n11926), .Y(new_n11723));
  not_8  g09375(.A(new_n11723), .Y(new_n11724_1));
  nor_5  g09376(.A(new_n11724_1), .B(n5521), .Y(new_n11725));
  xnor_4 g09377(.A(new_n11725), .B(n21784), .Y(new_n11726));
  xnor_4 g09378(.A(new_n11726), .B(new_n7264), .Y(new_n11727));
  xnor_4 g09379(.A(new_n11723), .B(n5521), .Y(new_n11728));
  nor_5  g09380(.A(new_n11728), .B(new_n7270), .Y(new_n11729));
  xnor_4 g09381(.A(new_n11728), .B(new_n7270), .Y(new_n11730));
  xnor_4 g09382(.A(new_n11721), .B(n11926), .Y(new_n11731));
  nor_5  g09383(.A(new_n11731), .B(new_n7275), .Y(new_n11732));
  xnor_4 g09384(.A(new_n11731), .B(new_n7275), .Y(new_n11733));
  nor_5  g09385(.A(new_n3850_1), .B(new_n3840), .Y(new_n11734));
  nor_5  g09386(.A(new_n3888), .B(new_n3851), .Y(new_n11735));
  nor_5  g09387(.A(new_n11735), .B(new_n11734), .Y(new_n11736_1));
  nor_5  g09388(.A(new_n11736_1), .B(new_n11733), .Y(new_n11737));
  nor_5  g09389(.A(new_n11737), .B(new_n11732), .Y(new_n11738));
  nor_5  g09390(.A(new_n11738), .B(new_n11730), .Y(new_n11739));
  nor_5  g09391(.A(new_n11739), .B(new_n11729), .Y(new_n11740));
  xnor_4 g09392(.A(new_n11740), .B(new_n11727), .Y(new_n11741_1));
  not_8  g09393(.A(new_n11741_1), .Y(new_n11742));
  xnor_4 g09394(.A(new_n11742), .B(new_n11719), .Y(new_n11743));
  xnor_4 g09395(.A(new_n11716), .B(new_n11675), .Y(new_n11744));
  xnor_4 g09396(.A(new_n11738), .B(new_n11730), .Y(new_n11745));
  not_8  g09397(.A(new_n11745), .Y(new_n11746));
  and_5  g09398(.A(new_n11746), .B(new_n11744), .Y(new_n11747));
  xnor_4 g09399(.A(new_n11746), .B(new_n11744), .Y(new_n11748));
  xnor_4 g09400(.A(new_n11714), .B(new_n11678), .Y(new_n11749_1));
  xnor_4 g09401(.A(new_n11736_1), .B(new_n11733), .Y(new_n11750));
  nor_5  g09402(.A(new_n11750), .B(new_n11749_1), .Y(new_n11751));
  xnor_4 g09403(.A(new_n11750), .B(new_n11749_1), .Y(new_n11752));
  xnor_4 g09404(.A(new_n11712_1), .B(new_n11681), .Y(new_n11753));
  nor_5  g09405(.A(new_n11753), .B(new_n3889), .Y(new_n11754));
  xnor_4 g09406(.A(new_n11753), .B(new_n3889), .Y(new_n11755));
  xnor_4 g09407(.A(new_n11710_1), .B(new_n11684), .Y(new_n11756));
  nor_5  g09408(.A(new_n11756), .B(new_n3891_1), .Y(new_n11757));
  xnor_4 g09409(.A(new_n11756), .B(new_n3891_1), .Y(new_n11758));
  xnor_4 g09410(.A(new_n11708), .B(new_n11688), .Y(new_n11759));
  nor_5  g09411(.A(new_n11759), .B(new_n3895), .Y(new_n11760));
  xnor_4 g09412(.A(new_n11759), .B(new_n3895), .Y(new_n11761));
  xnor_4 g09413(.A(new_n11706), .B(new_n11692), .Y(new_n11762));
  nor_5  g09414(.A(new_n11762), .B(new_n3900), .Y(new_n11763));
  xnor_4 g09415(.A(new_n11762), .B(new_n3900), .Y(new_n11764));
  xnor_4 g09416(.A(new_n11704), .B(new_n11696), .Y(new_n11765));
  nor_5  g09417(.A(new_n11765), .B(new_n3904), .Y(new_n11766));
  xnor_4 g09418(.A(new_n11765), .B(new_n3904), .Y(new_n11767));
  not_8  g09419(.A(new_n11767), .Y(new_n11768));
  xnor_4 g09420(.A(new_n11697), .B(n1451), .Y(new_n11769));
  nor_5  g09421(.A(new_n11769), .B(new_n3914), .Y(new_n11770_1));
  xnor_4 g09422(.A(new_n11701), .B(new_n11700), .Y(new_n11771_1));
  and_5  g09423(.A(new_n11771_1), .B(new_n11770_1), .Y(new_n11772));
  xnor_4 g09424(.A(new_n11771_1), .B(new_n11770_1), .Y(new_n11773));
  nor_5  g09425(.A(new_n11773), .B(new_n3908), .Y(new_n11774));
  nor_5  g09426(.A(new_n11774), .B(new_n11772), .Y(new_n11775_1));
  and_5  g09427(.A(new_n11775_1), .B(new_n11768), .Y(new_n11776));
  nor_5  g09428(.A(new_n11776), .B(new_n11766), .Y(new_n11777));
  nor_5  g09429(.A(new_n11777), .B(new_n11764), .Y(new_n11778));
  nor_5  g09430(.A(new_n11778), .B(new_n11763), .Y(new_n11779));
  nor_5  g09431(.A(new_n11779), .B(new_n11761), .Y(new_n11780));
  nor_5  g09432(.A(new_n11780), .B(new_n11760), .Y(new_n11781));
  nor_5  g09433(.A(new_n11781), .B(new_n11758), .Y(new_n11782));
  nor_5  g09434(.A(new_n11782), .B(new_n11757), .Y(new_n11783));
  nor_5  g09435(.A(new_n11783), .B(new_n11755), .Y(new_n11784));
  nor_5  g09436(.A(new_n11784), .B(new_n11754), .Y(new_n11785));
  nor_5  g09437(.A(new_n11785), .B(new_n11752), .Y(new_n11786));
  nor_5  g09438(.A(new_n11786), .B(new_n11751), .Y(new_n11787));
  nor_5  g09439(.A(new_n11787), .B(new_n11748), .Y(new_n11788));
  nor_5  g09440(.A(new_n11788), .B(new_n11747), .Y(new_n11789));
  xnor_4 g09441(.A(new_n11789), .B(new_n11743), .Y(n1859));
  xnor_4 g09442(.A(new_n5215), .B(new_n5189), .Y(n1860));
  not_8  g09443(.A(new_n11323), .Y(new_n11792));
  nor_5  g09444(.A(new_n11792), .B(new_n11320), .Y(new_n11793));
  not_8  g09445(.A(new_n11793), .Y(new_n11794));
  not_8  g09446(.A(n10250), .Y(new_n11795));
  nor_5  g09447(.A(n21915), .B(n15182), .Y(new_n11796));
  or_5   g09448(.A(new_n6861_1), .B(new_n6835_1), .Y(new_n11797));
  and_5  g09449(.A(new_n11797), .B(new_n6834), .Y(new_n11798));
  nor_5  g09450(.A(new_n11798), .B(new_n11796), .Y(new_n11799));
  not_8  g09451(.A(new_n11799), .Y(new_n11800));
  xnor_4 g09452(.A(n25972), .B(new_n6198), .Y(new_n11801));
  xnor_4 g09453(.A(new_n11801), .B(new_n11800), .Y(new_n11802));
  not_8  g09454(.A(new_n11802), .Y(new_n11803));
  nor_5  g09455(.A(new_n11803), .B(new_n11795), .Y(new_n11804));
  xnor_4 g09456(.A(new_n11802), .B(new_n11795), .Y(new_n11805));
  nor_5  g09457(.A(new_n6863_1), .B(new_n6155), .Y(new_n11806));
  xnor_4 g09458(.A(new_n6864), .B(new_n6155), .Y(new_n11807));
  nor_5  g09459(.A(new_n6867_1), .B(new_n6158), .Y(new_n11808));
  xnor_4 g09460(.A(new_n6869), .B(new_n6158), .Y(new_n11809));
  nor_5  g09461(.A(new_n6872), .B(new_n6161), .Y(new_n11810));
  xnor_4 g09462(.A(new_n6874), .B(new_n6161), .Y(new_n11811));
  not_8  g09463(.A(n23586), .Y(new_n11812));
  nor_5  g09464(.A(new_n6877), .B(new_n11812), .Y(new_n11813));
  nor_5  g09465(.A(new_n6881), .B(n21226), .Y(new_n11814));
  xnor_4 g09466(.A(new_n6882), .B(n21226), .Y(new_n11815));
  nor_5  g09467(.A(new_n6886), .B(new_n6170), .Y(new_n11816));
  xnor_4 g09468(.A(new_n6888), .B(new_n6170), .Y(new_n11817));
  nor_5  g09469(.A(new_n4116), .B(n20036), .Y(new_n11818_1));
  nor_5  g09470(.A(new_n4130), .B(new_n4120), .Y(new_n11819));
  nor_5  g09471(.A(new_n4135), .B(new_n6176), .Y(new_n11820));
  xnor_4 g09472(.A(new_n4138), .B(new_n4120), .Y(new_n11821));
  and_5  g09473(.A(new_n11821), .B(new_n11820), .Y(new_n11822));
  nor_5  g09474(.A(new_n11822), .B(new_n11819), .Y(new_n11823));
  xnor_4 g09475(.A(new_n4116), .B(new_n8659), .Y(new_n11824));
  and_5  g09476(.A(new_n11824), .B(new_n11823), .Y(new_n11825));
  nor_5  g09477(.A(new_n11825), .B(new_n11818_1), .Y(new_n11826));
  and_5  g09478(.A(new_n11826), .B(new_n11817), .Y(new_n11827));
  nor_5  g09479(.A(new_n11827), .B(new_n11816), .Y(new_n11828));
  and_5  g09480(.A(new_n11828), .B(new_n11815), .Y(new_n11829));
  nor_5  g09481(.A(new_n11829), .B(new_n11814), .Y(new_n11830));
  xnor_4 g09482(.A(new_n6879), .B(new_n11812), .Y(new_n11831));
  and_5  g09483(.A(new_n11831), .B(new_n11830), .Y(new_n11832));
  or_5   g09484(.A(new_n11832), .B(new_n11813), .Y(new_n11833));
  and_5  g09485(.A(new_n11833), .B(new_n11811), .Y(new_n11834));
  or_5   g09486(.A(new_n11834), .B(new_n11810), .Y(new_n11835));
  and_5  g09487(.A(new_n11835), .B(new_n11809), .Y(new_n11836));
  or_5   g09488(.A(new_n11836), .B(new_n11808), .Y(new_n11837_1));
  and_5  g09489(.A(new_n11837_1), .B(new_n11807), .Y(new_n11838));
  or_5   g09490(.A(new_n11838), .B(new_n11806), .Y(new_n11839));
  and_5  g09491(.A(new_n11839), .B(new_n11805), .Y(new_n11840));
  nor_5  g09492(.A(new_n11840), .B(new_n11804), .Y(new_n11841_1));
  not_8  g09493(.A(n25972), .Y(new_n11842_1));
  nor_5  g09494(.A(new_n11842_1), .B(new_n6198), .Y(new_n11843_1));
  nor_5  g09495(.A(n25972), .B(n8614), .Y(new_n11844));
  nor_5  g09496(.A(new_n11844), .B(new_n11800), .Y(new_n11845));
  nor_5  g09497(.A(new_n11845), .B(new_n11843_1), .Y(new_n11846));
  nor_5  g09498(.A(new_n11846), .B(new_n11841_1), .Y(new_n11847));
  nor_5  g09499(.A(new_n11847), .B(new_n11794), .Y(new_n11848));
  xnor_4 g09500(.A(new_n11847), .B(new_n11794), .Y(new_n11849));
  not_8  g09501(.A(new_n11324), .Y(new_n11850));
  not_8  g09502(.A(new_n11846), .Y(new_n11851));
  xnor_4 g09503(.A(new_n11851), .B(new_n11841_1), .Y(new_n11852));
  nor_5  g09504(.A(new_n11852), .B(new_n11850), .Y(new_n11853));
  xnor_4 g09505(.A(new_n11852), .B(new_n11850), .Y(new_n11854));
  xor_4  g09506(.A(new_n11839), .B(new_n11805), .Y(new_n11855));
  nor_5  g09507(.A(new_n11855), .B(new_n11338), .Y(new_n11856));
  xnor_4 g09508(.A(new_n11855), .B(new_n11338), .Y(new_n11857));
  not_8  g09509(.A(new_n11344), .Y(new_n11858));
  xor_4  g09510(.A(new_n11837_1), .B(new_n11807), .Y(new_n11859));
  nor_5  g09511(.A(new_n11859), .B(new_n11858), .Y(new_n11860));
  xnor_4 g09512(.A(new_n11859), .B(new_n11858), .Y(new_n11861));
  not_8  g09513(.A(new_n11348_1), .Y(new_n11862));
  xor_4  g09514(.A(new_n11835), .B(new_n11809), .Y(new_n11863));
  nor_5  g09515(.A(new_n11863), .B(new_n11862), .Y(new_n11864));
  xnor_4 g09516(.A(new_n11863), .B(new_n11862), .Y(new_n11865));
  xor_4  g09517(.A(new_n11833), .B(new_n11811), .Y(new_n11866));
  nor_5  g09518(.A(new_n11866), .B(new_n11366), .Y(new_n11867));
  xnor_4 g09519(.A(new_n11866), .B(new_n11366), .Y(new_n11868));
  xor_4  g09520(.A(new_n11831), .B(new_n11830), .Y(new_n11869));
  nor_5  g09521(.A(new_n11869), .B(new_n11358), .Y(new_n11870));
  xnor_4 g09522(.A(new_n11869), .B(new_n11358), .Y(new_n11871));
  xnor_4 g09523(.A(new_n11828), .B(new_n11815), .Y(new_n11872));
  nor_5  g09524(.A(new_n11872), .B(new_n9518), .Y(new_n11873));
  xnor_4 g09525(.A(new_n11872), .B(new_n9518), .Y(new_n11874));
  not_8  g09526(.A(new_n9520), .Y(new_n11875));
  xor_4  g09527(.A(new_n11826), .B(new_n11817), .Y(new_n11876));
  nor_5  g09528(.A(new_n11876), .B(new_n11875), .Y(new_n11877));
  xnor_4 g09529(.A(new_n11876), .B(new_n11875), .Y(new_n11878));
  xnor_4 g09530(.A(new_n11824), .B(new_n11823), .Y(new_n11879));
  nor_5  g09531(.A(new_n11879), .B(new_n9528), .Y(new_n11880));
  xnor_4 g09532(.A(new_n11879), .B(new_n9528), .Y(new_n11881));
  xor_4  g09533(.A(new_n11821), .B(new_n11820), .Y(new_n11882));
  nor_5  g09534(.A(new_n11882), .B(new_n9554_1), .Y(new_n11883));
  xnor_4 g09535(.A(new_n4135), .B(n9380), .Y(new_n11884));
  nor_5  g09536(.A(new_n11884), .B(new_n7200), .Y(new_n11885));
  xnor_4 g09537(.A(new_n11882), .B(new_n9530), .Y(new_n11886));
  and_5  g09538(.A(new_n11886), .B(new_n11885), .Y(new_n11887));
  nor_5  g09539(.A(new_n11887), .B(new_n11883), .Y(new_n11888));
  nor_5  g09540(.A(new_n11888), .B(new_n11881), .Y(new_n11889));
  nor_5  g09541(.A(new_n11889), .B(new_n11880), .Y(new_n11890));
  nor_5  g09542(.A(new_n11890), .B(new_n11878), .Y(new_n11891));
  nor_5  g09543(.A(new_n11891), .B(new_n11877), .Y(new_n11892));
  nor_5  g09544(.A(new_n11892), .B(new_n11874), .Y(new_n11893));
  nor_5  g09545(.A(new_n11893), .B(new_n11873), .Y(new_n11894));
  nor_5  g09546(.A(new_n11894), .B(new_n11871), .Y(new_n11895));
  nor_5  g09547(.A(new_n11895), .B(new_n11870), .Y(new_n11896));
  nor_5  g09548(.A(new_n11896), .B(new_n11868), .Y(new_n11897));
  nor_5  g09549(.A(new_n11897), .B(new_n11867), .Y(new_n11898_1));
  nor_5  g09550(.A(new_n11898_1), .B(new_n11865), .Y(new_n11899));
  nor_5  g09551(.A(new_n11899), .B(new_n11864), .Y(new_n11900));
  nor_5  g09552(.A(new_n11900), .B(new_n11861), .Y(new_n11901));
  nor_5  g09553(.A(new_n11901), .B(new_n11860), .Y(new_n11902));
  nor_5  g09554(.A(new_n11902), .B(new_n11857), .Y(new_n11903));
  nor_5  g09555(.A(new_n11903), .B(new_n11856), .Y(new_n11904));
  nor_5  g09556(.A(new_n11904), .B(new_n11854), .Y(new_n11905_1));
  nor_5  g09557(.A(new_n11905_1), .B(new_n11853), .Y(new_n11906));
  nor_5  g09558(.A(new_n11906), .B(new_n11849), .Y(new_n11907));
  or_5   g09559(.A(new_n11907), .B(new_n11848), .Y(n1861));
  nor_5  g09560(.A(n13714), .B(n12593), .Y(new_n11909));
  not_8  g09561(.A(new_n11909), .Y(new_n11910));
  nor_5  g09562(.A(new_n11910), .B(n19144), .Y(new_n11911));
  not_8  g09563(.A(new_n11911), .Y(new_n11912));
  nor_5  g09564(.A(new_n11912), .B(n8309), .Y(new_n11913));
  not_8  g09565(.A(new_n11913), .Y(new_n11914));
  nor_5  g09566(.A(new_n11914), .B(n19081), .Y(new_n11915));
  not_8  g09567(.A(new_n11915), .Y(new_n11916));
  nor_5  g09568(.A(new_n11916), .B(n26054), .Y(new_n11917));
  xnor_4 g09569(.A(new_n11917), .B(n26318), .Y(new_n11918));
  xnor_4 g09570(.A(new_n11918), .B(new_n5348), .Y(new_n11919));
  xnor_4 g09571(.A(new_n11915), .B(n26054), .Y(new_n11920));
  nor_5  g09572(.A(new_n11920), .B(new_n5391), .Y(new_n11921));
  xnor_4 g09573(.A(new_n11913), .B(n19081), .Y(new_n11922));
  nor_5  g09574(.A(new_n11922), .B(new_n5388), .Y(new_n11923));
  xnor_4 g09575(.A(new_n11922), .B(new_n5388), .Y(new_n11924));
  xnor_4 g09576(.A(new_n11911), .B(n8309), .Y(new_n11925));
  nor_5  g09577(.A(new_n11925), .B(new_n5358), .Y(new_n11926_1));
  xnor_4 g09578(.A(new_n11909), .B(n19144), .Y(new_n11927));
  nor_5  g09579(.A(new_n11927), .B(new_n5376_1), .Y(new_n11928));
  xnor_4 g09580(.A(new_n11927), .B(new_n5362), .Y(new_n11929));
  nor_5  g09581(.A(new_n5368), .B(new_n8763), .Y(new_n11930));
  xnor_4 g09582(.A(new_n11930), .B(n12593), .Y(new_n11931));
  nor_5  g09583(.A(new_n11931), .B(new_n5365), .Y(new_n11932));
  or_5   g09584(.A(new_n5369), .B(new_n8763), .Y(new_n11933));
  nor_5  g09585(.A(new_n11933), .B(n12593), .Y(new_n11934));
  nor_5  g09586(.A(new_n11934), .B(new_n11932), .Y(new_n11935));
  and_5  g09587(.A(new_n11935), .B(new_n11929), .Y(new_n11936));
  nor_5  g09588(.A(new_n11936), .B(new_n11928), .Y(new_n11937));
  xnor_4 g09589(.A(new_n11925), .B(new_n5358), .Y(new_n11938));
  nor_5  g09590(.A(new_n11938), .B(new_n11937), .Y(new_n11939));
  nor_5  g09591(.A(new_n11939), .B(new_n11926_1), .Y(new_n11940));
  nor_5  g09592(.A(new_n11940), .B(new_n11924), .Y(new_n11941));
  nor_5  g09593(.A(new_n11941), .B(new_n11923), .Y(new_n11942));
  xnor_4 g09594(.A(new_n11920), .B(new_n5391), .Y(new_n11943));
  nor_5  g09595(.A(new_n11943), .B(new_n11942), .Y(new_n11944));
  nor_5  g09596(.A(new_n11944), .B(new_n11921), .Y(new_n11945));
  xnor_4 g09597(.A(new_n11945), .B(new_n11919), .Y(new_n11946));
  not_8  g09598(.A(new_n8577), .Y(new_n11947));
  nor_5  g09599(.A(new_n11947), .B(n19228), .Y(new_n11948));
  not_8  g09600(.A(new_n11948), .Y(new_n11949));
  nor_5  g09601(.A(new_n11949), .B(n20179), .Y(new_n11950));
  xnor_4 g09602(.A(new_n11950), .B(n1112), .Y(new_n11951));
  xnor_4 g09603(.A(new_n11951), .B(new_n7278), .Y(new_n11952));
  not_8  g09604(.A(new_n7282), .Y(new_n11953));
  xnor_4 g09605(.A(new_n11948), .B(n20179), .Y(new_n11954));
  not_8  g09606(.A(new_n11954), .Y(new_n11955));
  nor_5  g09607(.A(new_n11955), .B(new_n11953), .Y(new_n11956));
  xnor_4 g09608(.A(new_n11955), .B(new_n11953), .Y(new_n11957));
  nor_5  g09609(.A(new_n8578), .B(new_n7285), .Y(new_n11958));
  xnor_4 g09610(.A(new_n8578), .B(new_n7285), .Y(new_n11959));
  nor_5  g09611(.A(new_n8580), .B(new_n7288), .Y(new_n11960));
  xnor_4 g09612(.A(new_n8580), .B(new_n7288), .Y(new_n11961));
  nor_5  g09613(.A(new_n8584), .B(new_n7295), .Y(new_n11962));
  or_5   g09614(.A(new_n8583), .B(new_n7293), .Y(new_n11963));
  nor_5  g09615(.A(new_n8588), .B(new_n7302), .Y(new_n11964));
  nor_5  g09616(.A(new_n7300), .B(new_n6771), .Y(new_n11965_1));
  xnor_4 g09617(.A(new_n8588), .B(new_n7302), .Y(new_n11966));
  nor_5  g09618(.A(new_n11966), .B(new_n11965_1), .Y(new_n11967));
  nor_5  g09619(.A(new_n11967), .B(new_n11964), .Y(new_n11968));
  and_5  g09620(.A(new_n11968), .B(new_n11963), .Y(new_n11969));
  or_5   g09621(.A(new_n11969), .B(new_n11962), .Y(new_n11970));
  nor_5  g09622(.A(new_n11970), .B(new_n11961), .Y(new_n11971));
  nor_5  g09623(.A(new_n11971), .B(new_n11960), .Y(new_n11972));
  nor_5  g09624(.A(new_n11972), .B(new_n11959), .Y(new_n11973));
  or_5   g09625(.A(new_n11973), .B(new_n11958), .Y(new_n11974));
  nor_5  g09626(.A(new_n11974), .B(new_n11957), .Y(new_n11975));
  nor_5  g09627(.A(new_n11975), .B(new_n11956), .Y(new_n11976));
  xor_4  g09628(.A(new_n11976), .B(new_n11952), .Y(new_n11977));
  xnor_4 g09629(.A(new_n11977), .B(new_n11946), .Y(new_n11978));
  xnor_4 g09630(.A(new_n11974), .B(new_n11957), .Y(new_n11979));
  xnor_4 g09631(.A(new_n11943), .B(new_n11942), .Y(new_n11980_1));
  not_8  g09632(.A(new_n11980_1), .Y(new_n11981));
  and_5  g09633(.A(new_n11981), .B(new_n11979), .Y(new_n11982));
  xnor_4 g09634(.A(new_n11981), .B(new_n11979), .Y(new_n11983));
  xnor_4 g09635(.A(new_n11940), .B(new_n11924), .Y(new_n11984));
  xnor_4 g09636(.A(new_n11972), .B(new_n11959), .Y(new_n11985));
  nor_5  g09637(.A(new_n11985), .B(new_n11984), .Y(new_n11986));
  xnor_4 g09638(.A(new_n11985), .B(new_n11984), .Y(new_n11987));
  xnor_4 g09639(.A(new_n11938), .B(new_n11937), .Y(new_n11988));
  xnor_4 g09640(.A(new_n11970), .B(new_n11961), .Y(new_n11989));
  nor_5  g09641(.A(new_n11989), .B(new_n11988), .Y(new_n11990));
  xnor_4 g09642(.A(new_n11989), .B(new_n11988), .Y(new_n11991));
  xnor_4 g09643(.A(new_n11935), .B(new_n11929), .Y(new_n11992));
  xnor_4 g09644(.A(new_n8584), .B(new_n7295), .Y(new_n11993));
  xnor_4 g09645(.A(new_n11993), .B(new_n11968), .Y(new_n11994));
  nor_5  g09646(.A(new_n11994), .B(new_n11992), .Y(new_n11995));
  xnor_4 g09647(.A(new_n11994), .B(new_n11992), .Y(new_n11996));
  xnor_4 g09648(.A(new_n11966), .B(new_n11965_1), .Y(new_n11997));
  xnor_4 g09649(.A(new_n11931), .B(new_n5372), .Y(new_n11998));
  nor_5  g09650(.A(new_n11998), .B(new_n11997), .Y(new_n11999));
  xnor_4 g09651(.A(new_n7300), .B(n18962), .Y(new_n12000_1));
  not_8  g09652(.A(new_n12000_1), .Y(new_n12001));
  xnor_4 g09653(.A(new_n5369), .B(new_n8763), .Y(new_n12002));
  nor_5  g09654(.A(new_n12002), .B(new_n12001), .Y(new_n12003_1));
  xnor_4 g09655(.A(new_n11998), .B(new_n11997), .Y(new_n12004));
  nor_5  g09656(.A(new_n12004), .B(new_n12003_1), .Y(new_n12005));
  nor_5  g09657(.A(new_n12005), .B(new_n11999), .Y(new_n12006));
  nor_5  g09658(.A(new_n12006), .B(new_n11996), .Y(new_n12007));
  nor_5  g09659(.A(new_n12007), .B(new_n11995), .Y(new_n12008));
  nor_5  g09660(.A(new_n12008), .B(new_n11991), .Y(new_n12009));
  nor_5  g09661(.A(new_n12009), .B(new_n11990), .Y(new_n12010));
  nor_5  g09662(.A(new_n12010), .B(new_n11987), .Y(new_n12011_1));
  nor_5  g09663(.A(new_n12011_1), .B(new_n11986), .Y(new_n12012));
  nor_5  g09664(.A(new_n12012), .B(new_n11983), .Y(new_n12013));
  nor_5  g09665(.A(new_n12013), .B(new_n11982), .Y(new_n12014));
  xnor_4 g09666(.A(new_n12014), .B(new_n11978), .Y(n1891));
  xnor_4 g09667(.A(n20169), .B(n1949), .Y(new_n12016));
  and_5  g09668(.A(n9323), .B(new_n6173), .Y(new_n12017));
  nor_5  g09669(.A(n9323), .B(new_n6173), .Y(new_n12018));
  and_5  g09670(.A(n10792), .B(new_n6178), .Y(new_n12019));
  or_5   g09671(.A(n10792), .B(new_n6178), .Y(new_n12020));
  nor_5  g09672(.A(n21687), .B(new_n4031), .Y(new_n12021));
  and_5  g09673(.A(new_n12021), .B(new_n12020), .Y(new_n12022));
  nor_5  g09674(.A(new_n12022), .B(new_n12019), .Y(new_n12023));
  nor_5  g09675(.A(new_n12023), .B(new_n12018), .Y(new_n12024));
  or_5   g09676(.A(new_n12024), .B(new_n12017), .Y(new_n12025));
  xor_4  g09677(.A(new_n12025), .B(new_n12016), .Y(new_n12026));
  xnor_4 g09678(.A(new_n12026), .B(new_n6560_1), .Y(new_n12027));
  xnor_4 g09679(.A(n9323), .B(n8285), .Y(new_n12028));
  xnor_4 g09680(.A(new_n12028), .B(new_n12023), .Y(new_n12029));
  and_5  g09681(.A(new_n12029), .B(new_n6566), .Y(new_n12030));
  xnor_4 g09682(.A(new_n12029), .B(new_n6566), .Y(new_n12031));
  xnor_4 g09683(.A(n21687), .B(n19922), .Y(new_n12032));
  nor_5  g09684(.A(new_n12032), .B(new_n6568), .Y(new_n12033));
  xnor_4 g09685(.A(n10792), .B(n6729), .Y(new_n12034));
  xnor_4 g09686(.A(new_n12034), .B(new_n12021), .Y(new_n12035));
  nor_5  g09687(.A(new_n12035), .B(new_n12033), .Y(new_n12036));
  xnor_4 g09688(.A(new_n12035), .B(new_n12033), .Y(new_n12037));
  nor_5  g09689(.A(new_n12037), .B(new_n6571), .Y(new_n12038));
  nor_5  g09690(.A(new_n12038), .B(new_n12036), .Y(new_n12039));
  nor_5  g09691(.A(new_n12039), .B(new_n12031), .Y(new_n12040));
  nor_5  g09692(.A(new_n12040), .B(new_n12030), .Y(new_n12041));
  xnor_4 g09693(.A(new_n12041), .B(new_n12027), .Y(n1925));
  xnor_4 g09694(.A(new_n7594), .B(new_n7570), .Y(n1942));
  xnor_4 g09695(.A(new_n6419), .B(new_n6365), .Y(n1972));
  and_5  g09696(.A(new_n8785), .B(new_n8718), .Y(new_n12045));
  nor_5  g09697(.A(new_n8852), .B(new_n8786), .Y(new_n12046));
  nor_5  g09698(.A(new_n12046), .B(new_n12045), .Y(new_n12047));
  not_8  g09699(.A(n22764), .Y(new_n12048));
  and_5  g09700(.A(new_n8734), .B(new_n12048), .Y(new_n12049));
  and_5  g09701(.A(new_n8735), .B(n12507), .Y(new_n12050));
  nor_5  g09702(.A(new_n8735), .B(n12507), .Y(new_n12051));
  nor_5  g09703(.A(new_n8784), .B(new_n12051), .Y(new_n12052));
  or_5   g09704(.A(new_n12052), .B(new_n12050), .Y(new_n12053));
  nor_5  g09705(.A(new_n12053), .B(new_n12049), .Y(new_n12054));
  and_5  g09706(.A(new_n12054), .B(new_n11026), .Y(new_n12055));
  and_5  g09707(.A(new_n12055), .B(new_n12047), .Y(new_n12056));
  or_5   g09708(.A(new_n12054), .B(new_n11026), .Y(new_n12057));
  nor_5  g09709(.A(new_n12057), .B(new_n12047), .Y(new_n12058));
  nor_5  g09710(.A(new_n12058), .B(new_n12056), .Y(new_n12059));
  and_5  g09711(.A(new_n12059), .B(new_n11018), .Y(new_n12060));
  xnor_4 g09712(.A(new_n12059), .B(new_n10912), .Y(new_n12061));
  xnor_4 g09713(.A(new_n12054), .B(new_n11025_1), .Y(new_n12062));
  xnor_4 g09714(.A(new_n12062), .B(new_n12047), .Y(new_n12063));
  not_8  g09715(.A(new_n12063), .Y(new_n12064));
  nor_5  g09716(.A(new_n12064), .B(new_n10912), .Y(new_n12065));
  xnor_4 g09717(.A(new_n12064), .B(new_n10912), .Y(new_n12066));
  not_8  g09718(.A(new_n8853), .Y(new_n12067));
  nor_5  g09719(.A(new_n10957), .B(new_n12067), .Y(new_n12068));
  nor_5  g09720(.A(new_n10964), .B(new_n8856_1), .Y(new_n12069));
  xnor_4 g09721(.A(new_n10964), .B(new_n8856_1), .Y(new_n12070));
  nor_5  g09722(.A(new_n10968), .B(new_n8860), .Y(new_n12071));
  xnor_4 g09723(.A(new_n10968), .B(new_n8860), .Y(new_n12072_1));
  nor_5  g09724(.A(new_n10973), .B(new_n8864), .Y(new_n12073));
  xnor_4 g09725(.A(new_n10973), .B(new_n8864), .Y(new_n12074));
  nor_5  g09726(.A(new_n10977), .B(new_n8868), .Y(new_n12075));
  xnor_4 g09727(.A(new_n10977), .B(new_n8868), .Y(new_n12076));
  nor_5  g09728(.A(new_n10982), .B(new_n8872), .Y(new_n12077));
  xnor_4 g09729(.A(new_n10982), .B(new_n8872), .Y(new_n12078));
  nor_5  g09730(.A(new_n10985), .B(new_n8875), .Y(new_n12079));
  xnor_4 g09731(.A(new_n10984), .B(new_n8876), .Y(new_n12080));
  and_5  g09732(.A(new_n10989), .B(new_n8880), .Y(new_n12081));
  xnor_4 g09733(.A(new_n10989), .B(new_n8880), .Y(new_n12082));
  nor_5  g09734(.A(new_n10992), .B(new_n8886), .Y(new_n12083));
  nor_5  g09735(.A(new_n12083), .B(new_n10996), .Y(new_n12084));
  xnor_4 g09736(.A(new_n12083), .B(new_n10995), .Y(new_n12085));
  and_5  g09737(.A(new_n12085), .B(new_n8891), .Y(new_n12086));
  nor_5  g09738(.A(new_n12086), .B(new_n12084), .Y(new_n12087));
  nor_5  g09739(.A(new_n12087), .B(new_n12082), .Y(new_n12088));
  nor_5  g09740(.A(new_n12088), .B(new_n12081), .Y(new_n12089));
  nor_5  g09741(.A(new_n12089), .B(new_n12080), .Y(new_n12090));
  nor_5  g09742(.A(new_n12090), .B(new_n12079), .Y(new_n12091));
  nor_5  g09743(.A(new_n12091), .B(new_n12078), .Y(new_n12092));
  nor_5  g09744(.A(new_n12092), .B(new_n12077), .Y(new_n12093));
  nor_5  g09745(.A(new_n12093), .B(new_n12076), .Y(new_n12094));
  nor_5  g09746(.A(new_n12094), .B(new_n12075), .Y(new_n12095));
  nor_5  g09747(.A(new_n12095), .B(new_n12074), .Y(new_n12096));
  nor_5  g09748(.A(new_n12096), .B(new_n12073), .Y(new_n12097));
  nor_5  g09749(.A(new_n12097), .B(new_n12072_1), .Y(new_n12098));
  nor_5  g09750(.A(new_n12098), .B(new_n12071), .Y(new_n12099));
  nor_5  g09751(.A(new_n12099), .B(new_n12070), .Y(new_n12100));
  nor_5  g09752(.A(new_n12100), .B(new_n12069), .Y(new_n12101));
  xnor_4 g09753(.A(new_n10957), .B(new_n12067), .Y(new_n12102));
  nor_5  g09754(.A(new_n12102), .B(new_n12101), .Y(new_n12103));
  nor_5  g09755(.A(new_n12103), .B(new_n12068), .Y(new_n12104));
  nor_5  g09756(.A(new_n12104), .B(new_n12066), .Y(new_n12105));
  nor_5  g09757(.A(new_n12105), .B(new_n12065), .Y(new_n12106));
  and_5  g09758(.A(new_n12106), .B(new_n12061), .Y(new_n12107));
  nor_5  g09759(.A(new_n12107), .B(new_n12060), .Y(n1981));
  xnor_4 g09760(.A(new_n12102), .B(new_n12101), .Y(n2004));
  not_8  g09761(.A(n5140), .Y(new_n12110));
  nor_5  g09762(.A(n6105), .B(new_n12110), .Y(new_n12111));
  xnor_4 g09763(.A(n6105), .B(n5140), .Y(new_n12112));
  not_8  g09764(.A(n6204), .Y(new_n12113_1));
  nor_5  g09765(.A(new_n12113_1), .B(n3795), .Y(new_n12114));
  xnor_4 g09766(.A(n6204), .B(n3795), .Y(new_n12115));
  not_8  g09767(.A(n3349), .Y(new_n12116));
  nor_5  g09768(.A(n25464), .B(new_n12116), .Y(new_n12117));
  xnor_4 g09769(.A(n25464), .B(n3349), .Y(new_n12118));
  not_8  g09770(.A(n1742), .Y(new_n12119));
  nor_5  g09771(.A(n4590), .B(new_n12119), .Y(new_n12120));
  xnor_4 g09772(.A(n4590), .B(n1742), .Y(new_n12121_1));
  not_8  g09773(.A(n4858), .Y(new_n12122));
  nor_5  g09774(.A(n26752), .B(new_n12122), .Y(new_n12123));
  xnor_4 g09775(.A(n26752), .B(n4858), .Y(new_n12124));
  not_8  g09776(.A(n8244), .Y(new_n12125));
  nor_5  g09777(.A(new_n12125), .B(n6513), .Y(new_n12126));
  xnor_4 g09778(.A(n8244), .B(n6513), .Y(new_n12127));
  not_8  g09779(.A(n9493), .Y(new_n12128));
  nor_5  g09780(.A(new_n12128), .B(n3918), .Y(new_n12129));
  xnor_4 g09781(.A(n9493), .B(n3918), .Y(new_n12130));
  nor_5  g09782(.A(n15167), .B(new_n4143), .Y(new_n12131_1));
  not_8  g09783(.A(n15167), .Y(new_n12132));
  nor_5  g09784(.A(new_n12132), .B(n919), .Y(new_n12133));
  not_8  g09785(.A(n21095), .Y(new_n12134));
  and_5  g09786(.A(n25316), .B(new_n12134), .Y(new_n12135));
  nor_5  g09787(.A(n25316), .B(new_n12134), .Y(new_n12136));
  nor_5  g09788(.A(new_n4146_1), .B(n8656), .Y(new_n12137));
  not_8  g09789(.A(new_n12137), .Y(new_n12138));
  nor_5  g09790(.A(new_n12138), .B(new_n12136), .Y(new_n12139));
  nor_5  g09791(.A(new_n12139), .B(new_n12135), .Y(new_n12140));
  nor_5  g09792(.A(new_n12140), .B(new_n12133), .Y(new_n12141));
  nor_5  g09793(.A(new_n12141), .B(new_n12131_1), .Y(new_n12142));
  and_5  g09794(.A(new_n12142), .B(new_n12130), .Y(new_n12143));
  or_5   g09795(.A(new_n12143), .B(new_n12129), .Y(new_n12144));
  and_5  g09796(.A(new_n12144), .B(new_n12127), .Y(new_n12145));
  or_5   g09797(.A(new_n12145), .B(new_n12126), .Y(new_n12146_1));
  and_5  g09798(.A(new_n12146_1), .B(new_n12124), .Y(new_n12147));
  or_5   g09799(.A(new_n12147), .B(new_n12123), .Y(new_n12148));
  and_5  g09800(.A(new_n12148), .B(new_n12121_1), .Y(new_n12149));
  or_5   g09801(.A(new_n12149), .B(new_n12120), .Y(new_n12150));
  and_5  g09802(.A(new_n12150), .B(new_n12118), .Y(new_n12151));
  or_5   g09803(.A(new_n12151), .B(new_n12117), .Y(new_n12152_1));
  and_5  g09804(.A(new_n12152_1), .B(new_n12115), .Y(new_n12153_1));
  or_5   g09805(.A(new_n12153_1), .B(new_n12114), .Y(new_n12154));
  and_5  g09806(.A(new_n12154), .B(new_n12112), .Y(new_n12155));
  nor_5  g09807(.A(new_n12155), .B(new_n12111), .Y(new_n12156));
  nor_5  g09808(.A(new_n6208), .B(n10018), .Y(new_n12157_1));
  not_8  g09809(.A(n10018), .Y(new_n12158_1));
  nor_5  g09810(.A(new_n6207), .B(new_n12158_1), .Y(new_n12159));
  nor_5  g09811(.A(new_n6216), .B(n2184), .Y(new_n12160));
  xnor_4 g09812(.A(new_n6213), .B(n2184), .Y(new_n12161_1));
  nor_5  g09813(.A(new_n6220), .B(n3541), .Y(new_n12162));
  xnor_4 g09814(.A(new_n6218_1), .B(n3541), .Y(new_n12163));
  nor_5  g09815(.A(new_n6224), .B(n16818), .Y(new_n12164));
  xnor_4 g09816(.A(new_n6223_1), .B(n16818), .Y(new_n12165));
  nor_5  g09817(.A(new_n4013), .B(n1269), .Y(new_n12166));
  xnor_4 g09818(.A(new_n4012), .B(n1269), .Y(new_n12167));
  nor_5  g09819(.A(new_n4017), .B(n14576), .Y(new_n12168));
  xnor_4 g09820(.A(new_n4016), .B(n14576), .Y(new_n12169));
  not_8  g09821(.A(n2985), .Y(new_n12170));
  nor_5  g09822(.A(new_n4019), .B(new_n12170), .Y(new_n12171));
  xnor_4 g09823(.A(new_n4019), .B(n2985), .Y(new_n12172));
  nor_5  g09824(.A(new_n4025), .B(n5605), .Y(new_n12173));
  and_5  g09825(.A(new_n4027), .B(n15652), .Y(new_n12174));
  nor_5  g09826(.A(n19922), .B(new_n6491), .Y(new_n12175));
  xnor_4 g09827(.A(new_n4028), .B(n15652), .Y(new_n12176));
  and_5  g09828(.A(new_n12176), .B(new_n12175), .Y(new_n12177));
  nor_5  g09829(.A(new_n12177), .B(new_n12174), .Y(new_n12178));
  xnor_4 g09830(.A(new_n4023), .B(n5605), .Y(new_n12179_1));
  and_5  g09831(.A(new_n12179_1), .B(new_n12178), .Y(new_n12180));
  nor_5  g09832(.A(new_n12180), .B(new_n12173), .Y(new_n12181));
  and_5  g09833(.A(new_n12181), .B(new_n12172), .Y(new_n12182));
  nor_5  g09834(.A(new_n12182), .B(new_n12171), .Y(new_n12183));
  and_5  g09835(.A(new_n12183), .B(new_n12169), .Y(new_n12184));
  or_5   g09836(.A(new_n12184), .B(new_n12168), .Y(new_n12185));
  and_5  g09837(.A(new_n12185), .B(new_n12167), .Y(new_n12186));
  or_5   g09838(.A(new_n12186), .B(new_n12166), .Y(new_n12187));
  and_5  g09839(.A(new_n12187), .B(new_n12165), .Y(new_n12188));
  or_5   g09840(.A(new_n12188), .B(new_n12164), .Y(new_n12189));
  and_5  g09841(.A(new_n12189), .B(new_n12163), .Y(new_n12190));
  or_5   g09842(.A(new_n12190), .B(new_n12162), .Y(new_n12191));
  and_5  g09843(.A(new_n12191), .B(new_n12161_1), .Y(new_n12192_1));
  nor_5  g09844(.A(new_n12192_1), .B(new_n12160), .Y(new_n12193));
  nor_5  g09845(.A(new_n12193), .B(new_n12159), .Y(new_n12194));
  xor_4  g09846(.A(new_n12194), .B(new_n6211), .Y(new_n12195));
  nor_5  g09847(.A(new_n12195), .B(new_n12157_1), .Y(new_n12196));
  xnor_4 g09848(.A(new_n12196), .B(new_n6242), .Y(new_n12197));
  xnor_4 g09849(.A(new_n6208), .B(new_n12158_1), .Y(new_n12198));
  xnor_4 g09850(.A(new_n12198), .B(new_n12193), .Y(new_n12199));
  not_8  g09851(.A(new_n12199), .Y(new_n12200));
  and_5  g09852(.A(new_n12200), .B(new_n6244), .Y(new_n12201));
  xnor_4 g09853(.A(new_n12200), .B(new_n6244), .Y(new_n12202));
  xor_4  g09854(.A(new_n12191), .B(new_n12161_1), .Y(new_n12203));
  nor_5  g09855(.A(new_n12203), .B(new_n6251), .Y(new_n12204));
  xnor_4 g09856(.A(new_n12203), .B(new_n6251), .Y(new_n12205));
  xor_4  g09857(.A(new_n12189), .B(new_n12163), .Y(new_n12206));
  nor_5  g09858(.A(new_n12206), .B(new_n6257), .Y(new_n12207));
  xnor_4 g09859(.A(new_n12206), .B(new_n6257), .Y(new_n12208));
  xor_4  g09860(.A(new_n12187), .B(new_n12165), .Y(new_n12209_1));
  nor_5  g09861(.A(new_n12209_1), .B(new_n6304), .Y(new_n12210));
  xor_4  g09862(.A(new_n12185), .B(new_n12167), .Y(new_n12211));
  nor_5  g09863(.A(new_n12211), .B(new_n6269), .Y(new_n12212));
  xnor_4 g09864(.A(new_n12211), .B(new_n6269), .Y(new_n12213));
  xor_4  g09865(.A(new_n12183), .B(new_n12169), .Y(new_n12214));
  nor_5  g09866(.A(new_n12214), .B(new_n6274), .Y(new_n12215));
  xnor_4 g09867(.A(new_n12214), .B(new_n6274), .Y(new_n12216));
  xnor_4 g09868(.A(new_n12181), .B(new_n12172), .Y(new_n12217));
  nor_5  g09869(.A(new_n12217), .B(new_n6277), .Y(new_n12218));
  xnor_4 g09870(.A(new_n12179_1), .B(new_n12178), .Y(new_n12219));
  nor_5  g09871(.A(new_n12219), .B(new_n6280), .Y(new_n12220));
  xnor_4 g09872(.A(new_n12219), .B(new_n6280), .Y(new_n12221));
  xor_4  g09873(.A(new_n12176), .B(new_n12175), .Y(new_n12222));
  nor_5  g09874(.A(new_n12222), .B(new_n6285), .Y(new_n12223_1));
  xnor_4 g09875(.A(n19922), .B(n4939), .Y(new_n12224));
  nor_5  g09876(.A(new_n12224), .B(new_n6288), .Y(new_n12225_1));
  not_8  g09877(.A(new_n6285), .Y(new_n12226));
  xnor_4 g09878(.A(new_n12222), .B(new_n12226), .Y(new_n12227));
  and_5  g09879(.A(new_n12227), .B(new_n12225_1), .Y(new_n12228_1));
  nor_5  g09880(.A(new_n12228_1), .B(new_n12223_1), .Y(new_n12229));
  nor_5  g09881(.A(new_n12229), .B(new_n12221), .Y(new_n12230));
  nor_5  g09882(.A(new_n12230), .B(new_n12220), .Y(new_n12231));
  xnor_4 g09883(.A(new_n12217), .B(new_n6276_1), .Y(new_n12232));
  and_5  g09884(.A(new_n12232), .B(new_n12231), .Y(new_n12233));
  nor_5  g09885(.A(new_n12233), .B(new_n12218), .Y(new_n12234));
  nor_5  g09886(.A(new_n12234), .B(new_n12216), .Y(new_n12235_1));
  nor_5  g09887(.A(new_n12235_1), .B(new_n12215), .Y(new_n12236));
  nor_5  g09888(.A(new_n12236), .B(new_n12213), .Y(new_n12237));
  nor_5  g09889(.A(new_n12237), .B(new_n12212), .Y(new_n12238));
  xnor_4 g09890(.A(new_n12209_1), .B(new_n6304), .Y(new_n12239));
  nor_5  g09891(.A(new_n12239), .B(new_n12238), .Y(new_n12240));
  nor_5  g09892(.A(new_n12240), .B(new_n12210), .Y(new_n12241));
  nor_5  g09893(.A(new_n12241), .B(new_n12208), .Y(new_n12242));
  nor_5  g09894(.A(new_n12242), .B(new_n12207), .Y(new_n12243));
  nor_5  g09895(.A(new_n12243), .B(new_n12205), .Y(new_n12244));
  nor_5  g09896(.A(new_n12244), .B(new_n12204), .Y(new_n12245));
  nor_5  g09897(.A(new_n12245), .B(new_n12202), .Y(new_n12246));
  nor_5  g09898(.A(new_n12246), .B(new_n12201), .Y(new_n12247));
  xnor_4 g09899(.A(new_n12247), .B(new_n12197), .Y(new_n12248));
  nor_5  g09900(.A(new_n12248), .B(new_n12156), .Y(new_n12249));
  xnor_4 g09901(.A(new_n12248), .B(new_n12156), .Y(new_n12250));
  xor_4  g09902(.A(new_n12154), .B(new_n12112), .Y(new_n12251));
  xnor_4 g09903(.A(new_n12245), .B(new_n12202), .Y(new_n12252));
  nor_5  g09904(.A(new_n12252), .B(new_n12251), .Y(new_n12253));
  xnor_4 g09905(.A(new_n12252), .B(new_n12251), .Y(new_n12254));
  xor_4  g09906(.A(new_n12152_1), .B(new_n12115), .Y(new_n12255));
  xnor_4 g09907(.A(new_n12243), .B(new_n12205), .Y(new_n12256));
  nor_5  g09908(.A(new_n12256), .B(new_n12255), .Y(new_n12257));
  xnor_4 g09909(.A(new_n12256), .B(new_n12255), .Y(new_n12258));
  xor_4  g09910(.A(new_n12150), .B(new_n12118), .Y(new_n12259));
  xnor_4 g09911(.A(new_n12241), .B(new_n12208), .Y(new_n12260));
  nor_5  g09912(.A(new_n12260), .B(new_n12259), .Y(new_n12261));
  xnor_4 g09913(.A(new_n12260), .B(new_n12259), .Y(new_n12262));
  xor_4  g09914(.A(new_n12148), .B(new_n12121_1), .Y(new_n12263));
  xnor_4 g09915(.A(new_n12239), .B(new_n12238), .Y(new_n12264));
  nor_5  g09916(.A(new_n12264), .B(new_n12263), .Y(new_n12265));
  xnor_4 g09917(.A(new_n12264), .B(new_n12263), .Y(new_n12266));
  xor_4  g09918(.A(new_n12146_1), .B(new_n12124), .Y(new_n12267));
  xnor_4 g09919(.A(new_n12236), .B(new_n12213), .Y(new_n12268));
  nor_5  g09920(.A(new_n12268), .B(new_n12267), .Y(new_n12269));
  xnor_4 g09921(.A(new_n12268), .B(new_n12267), .Y(new_n12270));
  xor_4  g09922(.A(new_n12144), .B(new_n12127), .Y(new_n12271));
  xnor_4 g09923(.A(new_n12234), .B(new_n12216), .Y(new_n12272));
  nor_5  g09924(.A(new_n12272), .B(new_n12271), .Y(new_n12273));
  xnor_4 g09925(.A(new_n12272), .B(new_n12271), .Y(new_n12274));
  xnor_4 g09926(.A(new_n12142), .B(new_n12130), .Y(new_n12275));
  xnor_4 g09927(.A(new_n12232), .B(new_n12231), .Y(new_n12276));
  not_8  g09928(.A(new_n12276), .Y(new_n12277));
  and_5  g09929(.A(new_n12277), .B(new_n12275), .Y(new_n12278));
  xnor_4 g09930(.A(new_n12277), .B(new_n12275), .Y(new_n12279));
  xnor_4 g09931(.A(new_n12229), .B(new_n12221), .Y(new_n12280));
  xnor_4 g09932(.A(n15167), .B(n919), .Y(new_n12281));
  xnor_4 g09933(.A(new_n12281), .B(new_n12140), .Y(new_n12282));
  and_5  g09934(.A(new_n12282), .B(new_n12280), .Y(new_n12283));
  xnor_4 g09935(.A(new_n12282), .B(new_n12280), .Y(new_n12284));
  xnor_4 g09936(.A(new_n12224), .B(new_n6287), .Y(new_n12285));
  not_8  g09937(.A(new_n12285), .Y(new_n12286));
  xnor_4 g09938(.A(n20385), .B(n8656), .Y(new_n12287));
  nor_5  g09939(.A(new_n12287), .B(new_n12286), .Y(new_n12288));
  xnor_4 g09940(.A(n25316), .B(n21095), .Y(new_n12289));
  xnor_4 g09941(.A(new_n12289), .B(new_n12138), .Y(new_n12290));
  not_8  g09942(.A(new_n12290), .Y(new_n12291));
  nor_5  g09943(.A(new_n12291), .B(new_n12288), .Y(new_n12292));
  xnor_4 g09944(.A(new_n12227), .B(new_n12225_1), .Y(new_n12293));
  xnor_4 g09945(.A(new_n12290), .B(new_n12288), .Y(new_n12294));
  and_5  g09946(.A(new_n12294), .B(new_n12293), .Y(new_n12295));
  nor_5  g09947(.A(new_n12295), .B(new_n12292), .Y(new_n12296));
  nor_5  g09948(.A(new_n12296), .B(new_n12284), .Y(new_n12297));
  nor_5  g09949(.A(new_n12297), .B(new_n12283), .Y(new_n12298));
  nor_5  g09950(.A(new_n12298), .B(new_n12279), .Y(new_n12299));
  nor_5  g09951(.A(new_n12299), .B(new_n12278), .Y(new_n12300));
  nor_5  g09952(.A(new_n12300), .B(new_n12274), .Y(new_n12301));
  nor_5  g09953(.A(new_n12301), .B(new_n12273), .Y(new_n12302_1));
  nor_5  g09954(.A(new_n12302_1), .B(new_n12270), .Y(new_n12303));
  nor_5  g09955(.A(new_n12303), .B(new_n12269), .Y(new_n12304_1));
  nor_5  g09956(.A(new_n12304_1), .B(new_n12266), .Y(new_n12305));
  nor_5  g09957(.A(new_n12305), .B(new_n12265), .Y(new_n12306));
  nor_5  g09958(.A(new_n12306), .B(new_n12262), .Y(new_n12307));
  nor_5  g09959(.A(new_n12307), .B(new_n12261), .Y(new_n12308));
  nor_5  g09960(.A(new_n12308), .B(new_n12258), .Y(new_n12309));
  nor_5  g09961(.A(new_n12309), .B(new_n12257), .Y(new_n12310));
  nor_5  g09962(.A(new_n12310), .B(new_n12254), .Y(new_n12311));
  nor_5  g09963(.A(new_n12311), .B(new_n12253), .Y(new_n12312));
  nor_5  g09964(.A(new_n12312), .B(new_n12250), .Y(new_n12313));
  nor_5  g09965(.A(new_n12313), .B(new_n12249), .Y(new_n12314));
  not_8  g09966(.A(new_n12314), .Y(new_n12315_1));
  nor_5  g09967(.A(new_n12196), .B(new_n6242), .Y(new_n12316));
  and_5  g09968(.A(new_n12194), .B(new_n6211), .Y(new_n12317));
  nand_5 g09969(.A(new_n12196), .B(new_n6242), .Y(new_n12318));
  and_5  g09970(.A(new_n12247), .B(new_n12318), .Y(new_n12319));
  or_5   g09971(.A(new_n12319), .B(new_n12317), .Y(new_n12320));
  nor_5  g09972(.A(new_n12320), .B(new_n12316), .Y(new_n12321));
  and_5  g09973(.A(new_n12321), .B(new_n12315_1), .Y(n2007));
  xnor_4 g09974(.A(new_n8895), .B(new_n8884_1), .Y(n2061));
  xnor_4 g09975(.A(new_n11205), .B(new_n7122), .Y(new_n12324_1));
  nor_5  g09976(.A(new_n11209), .B(new_n7126), .Y(new_n12325_1));
  xnor_4 g09977(.A(new_n11209), .B(new_n7126), .Y(new_n12326));
  nor_5  g09978(.A(new_n11214), .B(new_n7130), .Y(new_n12327));
  nor_5  g09979(.A(new_n7134), .B(new_n4660), .Y(new_n12328));
  xnor_4 g09980(.A(new_n7134), .B(new_n4660), .Y(new_n12329_1));
  nor_5  g09981(.A(new_n7138), .B(new_n4687), .Y(new_n12330_1));
  xnor_4 g09982(.A(new_n7138), .B(new_n4687), .Y(new_n12331));
  and_5  g09983(.A(new_n7141), .B(new_n4691), .Y(new_n12332));
  nor_5  g09984(.A(new_n7144), .B(new_n4699), .Y(new_n12333));
  xnor_4 g09985(.A(new_n7145), .B(new_n4699), .Y(new_n12334));
  nor_5  g09986(.A(new_n7150), .B(new_n4710), .Y(new_n12335));
  and_5  g09987(.A(new_n12335), .B(new_n4713), .Y(new_n12336));
  xnor_4 g09988(.A(new_n12335), .B(new_n4706), .Y(new_n12337));
  and_5  g09989(.A(new_n12337), .B(new_n7157), .Y(new_n12338));
  nor_5  g09990(.A(new_n12338), .B(new_n12336), .Y(new_n12339));
  and_5  g09991(.A(new_n12339), .B(new_n12334), .Y(new_n12340));
  nor_5  g09992(.A(new_n12340), .B(new_n12333), .Y(new_n12341_1));
  xnor_4 g09993(.A(new_n7141), .B(new_n4691), .Y(new_n12342));
  nor_5  g09994(.A(new_n12342), .B(new_n12341_1), .Y(new_n12343));
  nor_5  g09995(.A(new_n12343), .B(new_n12332), .Y(new_n12344));
  nor_5  g09996(.A(new_n12344), .B(new_n12331), .Y(new_n12345));
  nor_5  g09997(.A(new_n12345), .B(new_n12330_1), .Y(new_n12346_1));
  nor_5  g09998(.A(new_n12346_1), .B(new_n12329_1), .Y(new_n12347));
  nor_5  g09999(.A(new_n12347), .B(new_n12328), .Y(new_n12348));
  xnor_4 g10000(.A(new_n11214), .B(new_n7130), .Y(new_n12349_1));
  nor_5  g10001(.A(new_n12349_1), .B(new_n12348), .Y(new_n12350));
  nor_5  g10002(.A(new_n12350), .B(new_n12327), .Y(new_n12351));
  nor_5  g10003(.A(new_n12351), .B(new_n12326), .Y(new_n12352));
  nor_5  g10004(.A(new_n12352), .B(new_n12325_1), .Y(new_n12353));
  xnor_4 g10005(.A(new_n12353), .B(new_n12324_1), .Y(n2092));
  xnor_4 g10006(.A(n22253), .B(n10650), .Y(new_n12355));
  nor_5  g10007(.A(n12900), .B(n1255), .Y(new_n12356));
  xnor_4 g10008(.A(n12900), .B(n1255), .Y(new_n12357));
  nor_5  g10009(.A(n20411), .B(n9512), .Y(new_n12358));
  xnor_4 g10010(.A(n20411), .B(n9512), .Y(new_n12359));
  nor_5  g10011(.A(n17069), .B(n16608), .Y(new_n12360));
  xnor_4 g10012(.A(n17069), .B(n16608), .Y(new_n12361));
  nor_5  g10013(.A(n21735), .B(n15918), .Y(new_n12362));
  xnor_4 g10014(.A(n21735), .B(n15918), .Y(new_n12363));
  nor_5  g10015(.A(n24085), .B(n17784), .Y(new_n12364_1));
  xnor_4 g10016(.A(n24085), .B(n17784), .Y(new_n12365));
  nor_5  g10017(.A(n14323), .B(n14071), .Y(new_n12366));
  xnor_4 g10018(.A(n14323), .B(n14071), .Y(new_n12367));
  nor_5  g10019(.A(n2886), .B(n1738), .Y(new_n12368));
  xnor_4 g10020(.A(n2886), .B(n1738), .Y(new_n12369));
  nor_5  g10021(.A(n12152), .B(n1040), .Y(new_n12370));
  not_8  g10022(.A(n9090), .Y(new_n12371));
  or_5   g10023(.A(new_n7025), .B(new_n12371), .Y(new_n12372));
  not_8  g10024(.A(n1040), .Y(new_n12373));
  xnor_4 g10025(.A(n12152), .B(new_n12373), .Y(new_n12374));
  and_5  g10026(.A(new_n12374), .B(new_n12372), .Y(new_n12375));
  nor_5  g10027(.A(new_n12375), .B(new_n12370), .Y(new_n12376));
  nor_5  g10028(.A(new_n12376), .B(new_n12369), .Y(new_n12377));
  nor_5  g10029(.A(new_n12377), .B(new_n12368), .Y(new_n12378));
  nor_5  g10030(.A(new_n12378), .B(new_n12367), .Y(new_n12379));
  nor_5  g10031(.A(new_n12379), .B(new_n12366), .Y(new_n12380_1));
  nor_5  g10032(.A(new_n12380_1), .B(new_n12365), .Y(new_n12381));
  nor_5  g10033(.A(new_n12381), .B(new_n12364_1), .Y(new_n12382));
  nor_5  g10034(.A(new_n12382), .B(new_n12363), .Y(new_n12383_1));
  nor_5  g10035(.A(new_n12383_1), .B(new_n12362), .Y(new_n12384_1));
  nor_5  g10036(.A(new_n12384_1), .B(new_n12361), .Y(new_n12385));
  nor_5  g10037(.A(new_n12385), .B(new_n12360), .Y(new_n12386));
  nor_5  g10038(.A(new_n12386), .B(new_n12359), .Y(new_n12387));
  nor_5  g10039(.A(new_n12387), .B(new_n12358), .Y(new_n12388));
  nor_5  g10040(.A(new_n12388), .B(new_n12357), .Y(new_n12389));
  nor_5  g10041(.A(new_n12389), .B(new_n12356), .Y(new_n12390));
  xnor_4 g10042(.A(new_n12390), .B(new_n12355), .Y(new_n12391));
  nor_5  g10043(.A(new_n12391), .B(new_n7179), .Y(new_n12392));
  xnor_4 g10044(.A(new_n12391), .B(new_n7179), .Y(new_n12393));
  xnor_4 g10045(.A(new_n12388), .B(new_n12357), .Y(new_n12394));
  nor_5  g10046(.A(new_n12394), .B(new_n6967_1), .Y(new_n12395));
  xnor_4 g10047(.A(new_n12394), .B(new_n6967_1), .Y(new_n12396));
  xnor_4 g10048(.A(new_n12386), .B(new_n12359), .Y(new_n12397_1));
  nor_5  g10049(.A(new_n12397_1), .B(new_n6970), .Y(new_n12398_1));
  xnor_4 g10050(.A(new_n12397_1), .B(new_n6970), .Y(new_n12399));
  xnor_4 g10051(.A(new_n12384_1), .B(new_n12361), .Y(new_n12400));
  nor_5  g10052(.A(new_n12400), .B(new_n6973), .Y(new_n12401));
  xnor_4 g10053(.A(new_n12400), .B(new_n6973), .Y(new_n12402));
  xnor_4 g10054(.A(new_n12382), .B(new_n12363), .Y(new_n12403));
  nor_5  g10055(.A(new_n12403), .B(new_n6976), .Y(new_n12404));
  xnor_4 g10056(.A(new_n12403), .B(new_n6976), .Y(new_n12405));
  xnor_4 g10057(.A(new_n12380_1), .B(new_n12365), .Y(new_n12406));
  nor_5  g10058(.A(new_n12406), .B(new_n6979), .Y(new_n12407));
  xnor_4 g10059(.A(new_n12406), .B(new_n6979), .Y(new_n12408_1));
  xnor_4 g10060(.A(new_n12378), .B(new_n12367), .Y(new_n12409));
  nor_5  g10061(.A(new_n12409), .B(new_n6982), .Y(new_n12410));
  xnor_4 g10062(.A(new_n12409), .B(new_n6982), .Y(new_n12411));
  xnor_4 g10063(.A(new_n12376), .B(new_n12369), .Y(new_n12412));
  nor_5  g10064(.A(new_n12412), .B(new_n6986), .Y(new_n12413));
  xnor_4 g10065(.A(new_n12412), .B(n23775), .Y(new_n12414));
  xnor_4 g10066(.A(n19107), .B(new_n12371), .Y(new_n12415));
  nor_5  g10067(.A(new_n12415), .B(new_n11651), .Y(new_n12416));
  nor_5  g10068(.A(new_n12416), .B(n8259), .Y(new_n12417));
  xor_4  g10069(.A(new_n12374), .B(new_n12372), .Y(new_n12418));
  xnor_4 g10070(.A(new_n12416), .B(new_n6989), .Y(new_n12419));
  not_8  g10071(.A(new_n12419), .Y(new_n12420));
  nor_5  g10072(.A(new_n12420), .B(new_n12418), .Y(new_n12421));
  nor_5  g10073(.A(new_n12421), .B(new_n12417), .Y(new_n12422));
  and_5  g10074(.A(new_n12422), .B(new_n12414), .Y(new_n12423));
  nor_5  g10075(.A(new_n12423), .B(new_n12413), .Y(new_n12424));
  nor_5  g10076(.A(new_n12424), .B(new_n12411), .Y(new_n12425));
  nor_5  g10077(.A(new_n12425), .B(new_n12410), .Y(new_n12426));
  nor_5  g10078(.A(new_n12426), .B(new_n12408_1), .Y(new_n12427));
  nor_5  g10079(.A(new_n12427), .B(new_n12407), .Y(new_n12428));
  nor_5  g10080(.A(new_n12428), .B(new_n12405), .Y(new_n12429));
  nor_5  g10081(.A(new_n12429), .B(new_n12404), .Y(new_n12430));
  nor_5  g10082(.A(new_n12430), .B(new_n12402), .Y(new_n12431));
  nor_5  g10083(.A(new_n12431), .B(new_n12401), .Y(new_n12432));
  nor_5  g10084(.A(new_n12432), .B(new_n12399), .Y(new_n12433));
  nor_5  g10085(.A(new_n12433), .B(new_n12398_1), .Y(new_n12434));
  nor_5  g10086(.A(new_n12434), .B(new_n12396), .Y(new_n12435));
  nor_5  g10087(.A(new_n12435), .B(new_n12395), .Y(new_n12436));
  nor_5  g10088(.A(new_n12436), .B(new_n12393), .Y(new_n12437));
  nor_5  g10089(.A(new_n12437), .B(new_n12392), .Y(new_n12438));
  nor_5  g10090(.A(n22253), .B(n10650), .Y(new_n12439));
  nor_5  g10091(.A(new_n12390), .B(new_n12355), .Y(new_n12440));
  nor_5  g10092(.A(new_n12440), .B(new_n12439), .Y(new_n12441));
  nor_5  g10093(.A(new_n12441), .B(new_n12438), .Y(new_n12442));
  not_8  g10094(.A(n9934), .Y(new_n12443));
  nor_5  g10095(.A(n7876), .B(n4964), .Y(new_n12444));
  not_8  g10096(.A(new_n12444), .Y(new_n12445));
  nor_5  g10097(.A(new_n12445), .B(n26553), .Y(new_n12446_1));
  not_8  g10098(.A(new_n12446_1), .Y(new_n12447));
  nor_5  g10099(.A(new_n12447), .B(n342), .Y(new_n12448));
  not_8  g10100(.A(new_n12448), .Y(new_n12449_1));
  nor_5  g10101(.A(new_n12449_1), .B(n26107), .Y(new_n12450));
  not_8  g10102(.A(new_n12450), .Y(new_n12451));
  nor_5  g10103(.A(new_n12451), .B(n22597), .Y(new_n12452));
  not_8  g10104(.A(new_n12452), .Y(new_n12453));
  nor_5  g10105(.A(new_n12453), .B(n19327), .Y(new_n12454));
  not_8  g10106(.A(new_n12454), .Y(new_n12455));
  nor_5  g10107(.A(new_n12455), .B(n26224), .Y(new_n12456));
  and_5  g10108(.A(new_n12456), .B(new_n11636), .Y(new_n12457));
  and_5  g10109(.A(new_n12457), .B(new_n12443), .Y(new_n12458));
  xnor_4 g10110(.A(new_n12457), .B(new_n12443), .Y(new_n12459));
  nor_5  g10111(.A(n18409), .B(n5704), .Y(new_n12460));
  not_8  g10112(.A(new_n12460), .Y(new_n12461_1));
  nor_5  g10113(.A(new_n12461_1), .B(n13708), .Y(new_n12462_1));
  not_8  g10114(.A(new_n12462_1), .Y(new_n12463));
  nor_5  g10115(.A(new_n12463), .B(n19911), .Y(new_n12464));
  not_8  g10116(.A(new_n12464), .Y(new_n12465));
  nor_5  g10117(.A(new_n12465), .B(n2731), .Y(new_n12466));
  not_8  g10118(.A(new_n12466), .Y(new_n12467_1));
  nor_5  g10119(.A(new_n12467_1), .B(n18907), .Y(new_n12468));
  not_8  g10120(.A(new_n12468), .Y(new_n12469_1));
  nor_5  g10121(.A(new_n12469_1), .B(n22332), .Y(new_n12470));
  not_8  g10122(.A(new_n12470), .Y(new_n12471));
  nor_5  g10123(.A(new_n12471), .B(n4256), .Y(new_n12472));
  xnor_4 g10124(.A(new_n12472), .B(n21287), .Y(new_n12473));
  nor_5  g10125(.A(new_n12473), .B(n12861), .Y(new_n12474));
  xnor_4 g10126(.A(new_n12473), .B(new_n7043), .Y(new_n12475));
  xnor_4 g10127(.A(new_n12470), .B(n4256), .Y(new_n12476));
  nor_5  g10128(.A(new_n12476), .B(n13333), .Y(new_n12477));
  xnor_4 g10129(.A(new_n12476), .B(new_n7046), .Y(new_n12478));
  xnor_4 g10130(.A(new_n12468), .B(n22332), .Y(new_n12479));
  nor_5  g10131(.A(new_n12479), .B(n2210), .Y(new_n12480));
  xnor_4 g10132(.A(new_n12479), .B(new_n7049), .Y(new_n12481));
  xnor_4 g10133(.A(new_n12466), .B(n18907), .Y(new_n12482));
  nor_5  g10134(.A(new_n12482), .B(n20604), .Y(new_n12483));
  xnor_4 g10135(.A(new_n12482), .B(new_n5125), .Y(new_n12484));
  xnor_4 g10136(.A(new_n12464), .B(n2731), .Y(new_n12485));
  nor_5  g10137(.A(new_n12485), .B(n16158), .Y(new_n12486));
  xnor_4 g10138(.A(new_n12485), .B(new_n4614), .Y(new_n12487));
  xnor_4 g10139(.A(new_n12462_1), .B(n19911), .Y(new_n12488));
  nor_5  g10140(.A(new_n12488), .B(n5752), .Y(new_n12489));
  xnor_4 g10141(.A(new_n12460), .B(n13708), .Y(new_n12490));
  nor_5  g10142(.A(new_n12490), .B(n18171), .Y(new_n12491));
  xnor_4 g10143(.A(new_n12490), .B(new_n4620), .Y(new_n12492));
  xnor_4 g10144(.A(n18409), .B(n5704), .Y(new_n12493));
  and_5  g10145(.A(new_n12493), .B(new_n4623), .Y(new_n12494));
  or_5   g10146(.A(new_n4626), .B(new_n2381), .Y(new_n12495_1));
  xnor_4 g10147(.A(new_n12493), .B(n25073), .Y(new_n12496));
  and_5  g10148(.A(new_n12496), .B(new_n12495_1), .Y(new_n12497));
  or_5   g10149(.A(new_n12497), .B(new_n12494), .Y(new_n12498));
  and_5  g10150(.A(new_n12498), .B(new_n12492), .Y(new_n12499));
  or_5   g10151(.A(new_n12499), .B(new_n12491), .Y(new_n12500));
  xnor_4 g10152(.A(new_n12488), .B(new_n4617), .Y(new_n12501));
  and_5  g10153(.A(new_n12501), .B(new_n12500), .Y(new_n12502));
  or_5   g10154(.A(new_n12502), .B(new_n12489), .Y(new_n12503));
  and_5  g10155(.A(new_n12503), .B(new_n12487), .Y(new_n12504));
  or_5   g10156(.A(new_n12504), .B(new_n12486), .Y(new_n12505));
  and_5  g10157(.A(new_n12505), .B(new_n12484), .Y(new_n12506));
  or_5   g10158(.A(new_n12506), .B(new_n12483), .Y(new_n12507_1));
  and_5  g10159(.A(new_n12507_1), .B(new_n12481), .Y(new_n12508));
  or_5   g10160(.A(new_n12508), .B(new_n12480), .Y(new_n12509));
  and_5  g10161(.A(new_n12509), .B(new_n12478), .Y(new_n12510));
  or_5   g10162(.A(new_n12510), .B(new_n12477), .Y(new_n12511));
  and_5  g10163(.A(new_n12511), .B(new_n12475), .Y(new_n12512));
  nor_5  g10164(.A(new_n12512), .B(new_n12474), .Y(new_n12513));
  not_8  g10165(.A(new_n12472), .Y(new_n12514));
  nor_5  g10166(.A(new_n12514), .B(n21287), .Y(new_n12515_1));
  xnor_4 g10167(.A(new_n12515_1), .B(n26986), .Y(new_n12516_1));
  xnor_4 g10168(.A(new_n12516_1), .B(new_n7110), .Y(new_n12517));
  xnor_4 g10169(.A(new_n12517), .B(new_n12513), .Y(new_n12518));
  nor_5  g10170(.A(new_n12518), .B(new_n12459), .Y(new_n12519));
  xnor_4 g10171(.A(new_n12518), .B(new_n12459), .Y(new_n12520));
  xnor_4 g10172(.A(new_n12456), .B(new_n11636), .Y(new_n12521));
  nor_5  g10173(.A(new_n12510), .B(new_n12477), .Y(new_n12522));
  xnor_4 g10174(.A(new_n12522), .B(new_n12475), .Y(new_n12523));
  nor_5  g10175(.A(new_n12523), .B(new_n12521), .Y(new_n12524));
  xnor_4 g10176(.A(new_n12523), .B(new_n12521), .Y(new_n12525));
  not_8  g10177(.A(n26224), .Y(new_n12526));
  xnor_4 g10178(.A(new_n12454), .B(new_n12526), .Y(new_n12527));
  xor_4  g10179(.A(new_n12509), .B(new_n12478), .Y(new_n12528));
  nor_5  g10180(.A(new_n12528), .B(new_n12527), .Y(new_n12529));
  xnor_4 g10181(.A(new_n12528), .B(new_n12527), .Y(new_n12530));
  xnor_4 g10182(.A(new_n12452), .B(new_n3726), .Y(new_n12531));
  nor_5  g10183(.A(new_n12506), .B(new_n12483), .Y(new_n12532));
  xnor_4 g10184(.A(new_n12532), .B(new_n12481), .Y(new_n12533));
  nor_5  g10185(.A(new_n12533), .B(new_n12531), .Y(new_n12534));
  xnor_4 g10186(.A(new_n12533), .B(new_n12531), .Y(new_n12535));
  xnor_4 g10187(.A(new_n12450), .B(new_n3740_1), .Y(new_n12536));
  xor_4  g10188(.A(new_n12505), .B(new_n12484), .Y(new_n12537));
  nor_5  g10189(.A(new_n12537), .B(new_n12536), .Y(new_n12538));
  xnor_4 g10190(.A(new_n12537), .B(new_n12536), .Y(new_n12539));
  xnor_4 g10191(.A(new_n12448), .B(n26107), .Y(new_n12540_1));
  not_8  g10192(.A(new_n12540_1), .Y(new_n12541));
  nor_5  g10193(.A(new_n12502), .B(new_n12489), .Y(new_n12542));
  xnor_4 g10194(.A(new_n12542), .B(new_n12487), .Y(new_n12543));
  nor_5  g10195(.A(new_n12543), .B(new_n12541), .Y(new_n12544));
  not_8  g10196(.A(new_n12543), .Y(new_n12545_1));
  xnor_4 g10197(.A(new_n12545_1), .B(new_n12541), .Y(new_n12546_1));
  xnor_4 g10198(.A(new_n12446_1), .B(n342), .Y(new_n12547));
  xnor_4 g10199(.A(new_n12501), .B(new_n12500), .Y(new_n12548));
  and_5  g10200(.A(new_n12548), .B(new_n12547), .Y(new_n12549));
  xor_4  g10201(.A(new_n12501), .B(new_n12500), .Y(new_n12550));
  xnor_4 g10202(.A(new_n12550), .B(new_n12547), .Y(new_n12551));
  nor_5  g10203(.A(new_n12497), .B(new_n12494), .Y(new_n12552_1));
  xnor_4 g10204(.A(new_n12552_1), .B(new_n12492), .Y(new_n12553));
  not_8  g10205(.A(new_n12553), .Y(new_n12554));
  xnor_4 g10206(.A(new_n12444), .B(n26553), .Y(new_n12555));
  and_5  g10207(.A(new_n12555), .B(new_n12554), .Y(new_n12556));
  xnor_4 g10208(.A(new_n12555), .B(new_n12553), .Y(new_n12557));
  xnor_4 g10209(.A(n7876), .B(n4964), .Y(new_n12558));
  nor_5  g10210(.A(new_n4626), .B(new_n2381), .Y(new_n12559));
  xnor_4 g10211(.A(new_n12496), .B(new_n12559), .Y(new_n12560));
  nor_5  g10212(.A(new_n12560), .B(new_n12558), .Y(new_n12561));
  xnor_4 g10213(.A(n22309), .B(new_n2381), .Y(new_n12562_1));
  not_8  g10214(.A(new_n12562_1), .Y(new_n12563));
  nor_5  g10215(.A(new_n12563), .B(new_n3755_1), .Y(new_n12564));
  not_8  g10216(.A(new_n12560), .Y(new_n12565));
  xnor_4 g10217(.A(new_n12565), .B(new_n12558), .Y(new_n12566_1));
  and_5  g10218(.A(new_n12566_1), .B(new_n12564), .Y(new_n12567));
  or_5   g10219(.A(new_n12567), .B(new_n12561), .Y(new_n12568));
  and_5  g10220(.A(new_n12568), .B(new_n12557), .Y(new_n12569_1));
  or_5   g10221(.A(new_n12569_1), .B(new_n12556), .Y(new_n12570));
  and_5  g10222(.A(new_n12570), .B(new_n12551), .Y(new_n12571));
  or_5   g10223(.A(new_n12571), .B(new_n12549), .Y(new_n12572));
  and_5  g10224(.A(new_n12572), .B(new_n12546_1), .Y(new_n12573));
  nor_5  g10225(.A(new_n12573), .B(new_n12544), .Y(new_n12574));
  nor_5  g10226(.A(new_n12574), .B(new_n12539), .Y(new_n12575));
  nor_5  g10227(.A(new_n12575), .B(new_n12538), .Y(new_n12576));
  nor_5  g10228(.A(new_n12576), .B(new_n12535), .Y(new_n12577));
  nor_5  g10229(.A(new_n12577), .B(new_n12534), .Y(new_n12578));
  nor_5  g10230(.A(new_n12578), .B(new_n12530), .Y(new_n12579));
  nor_5  g10231(.A(new_n12579), .B(new_n12529), .Y(new_n12580));
  nor_5  g10232(.A(new_n12580), .B(new_n12525), .Y(new_n12581));
  nor_5  g10233(.A(new_n12581), .B(new_n12524), .Y(new_n12582));
  nor_5  g10234(.A(new_n12582), .B(new_n12520), .Y(new_n12583));
  or_5   g10235(.A(new_n12583), .B(new_n12519), .Y(new_n12584));
  nor_5  g10236(.A(new_n12584), .B(new_n12458), .Y(new_n12585));
  and_5  g10237(.A(new_n12515_1), .B(new_n7243), .Y(new_n12586));
  nor_5  g10238(.A(new_n12516_1), .B(n8305), .Y(new_n12587_1));
  and_5  g10239(.A(new_n12516_1), .B(n8305), .Y(new_n12588));
  nor_5  g10240(.A(new_n12588), .B(new_n12513), .Y(new_n12589));
  nor_5  g10241(.A(new_n12589), .B(new_n12587_1), .Y(new_n12590));
  or_5   g10242(.A(new_n12590), .B(new_n12586), .Y(new_n12591));
  and_5  g10243(.A(new_n12591), .B(new_n12585), .Y(new_n12592));
  xnor_4 g10244(.A(new_n12592), .B(new_n12442), .Y(new_n12593_1));
  xnor_4 g10245(.A(new_n12441), .B(new_n12438), .Y(new_n12594));
  nor_5  g10246(.A(new_n12590), .B(new_n12586), .Y(new_n12595));
  xnor_4 g10247(.A(new_n12595), .B(new_n12585), .Y(new_n12596));
  not_8  g10248(.A(new_n12596), .Y(new_n12597));
  nor_5  g10249(.A(new_n12597), .B(new_n12594), .Y(new_n12598));
  xnor_4 g10250(.A(new_n12597), .B(new_n12594), .Y(new_n12599));
  xnor_4 g10251(.A(new_n12436), .B(new_n12393), .Y(new_n12600));
  xnor_4 g10252(.A(new_n12582), .B(new_n12520), .Y(new_n12601));
  not_8  g10253(.A(new_n12601), .Y(new_n12602));
  nor_5  g10254(.A(new_n12602), .B(new_n12600), .Y(new_n12603));
  xnor_4 g10255(.A(new_n12602), .B(new_n12600), .Y(new_n12604));
  xnor_4 g10256(.A(new_n12434), .B(new_n12396), .Y(new_n12605));
  xnor_4 g10257(.A(new_n12580), .B(new_n12525), .Y(new_n12606));
  not_8  g10258(.A(new_n12606), .Y(new_n12607_1));
  nor_5  g10259(.A(new_n12607_1), .B(new_n12605), .Y(new_n12608));
  xnor_4 g10260(.A(new_n12607_1), .B(new_n12605), .Y(new_n12609));
  xnor_4 g10261(.A(new_n12432), .B(new_n12399), .Y(new_n12610));
  xnor_4 g10262(.A(new_n12578), .B(new_n12530), .Y(new_n12611));
  not_8  g10263(.A(new_n12611), .Y(new_n12612));
  nor_5  g10264(.A(new_n12612), .B(new_n12610), .Y(new_n12613));
  xnor_4 g10265(.A(new_n12612), .B(new_n12610), .Y(new_n12614));
  xnor_4 g10266(.A(new_n12430), .B(new_n12402), .Y(new_n12615));
  xnor_4 g10267(.A(new_n12576), .B(new_n12535), .Y(new_n12616));
  not_8  g10268(.A(new_n12616), .Y(new_n12617));
  nor_5  g10269(.A(new_n12617), .B(new_n12615), .Y(new_n12618));
  xnor_4 g10270(.A(new_n12617), .B(new_n12615), .Y(new_n12619));
  xnor_4 g10271(.A(new_n12428), .B(new_n12405), .Y(new_n12620_1));
  xnor_4 g10272(.A(new_n12574), .B(new_n12539), .Y(new_n12621_1));
  not_8  g10273(.A(new_n12621_1), .Y(new_n12622));
  nor_5  g10274(.A(new_n12622), .B(new_n12620_1), .Y(new_n12623));
  xnor_4 g10275(.A(new_n12622), .B(new_n12620_1), .Y(new_n12624));
  xnor_4 g10276(.A(new_n12426), .B(new_n12408_1), .Y(new_n12625));
  xor_4  g10277(.A(new_n12572), .B(new_n12546_1), .Y(new_n12626_1));
  nor_5  g10278(.A(new_n12626_1), .B(new_n12625), .Y(new_n12627));
  xnor_4 g10279(.A(new_n12626_1), .B(new_n12625), .Y(new_n12628));
  xnor_4 g10280(.A(new_n12424), .B(new_n12411), .Y(new_n12629));
  xor_4  g10281(.A(new_n12570), .B(new_n12551), .Y(new_n12630));
  nor_5  g10282(.A(new_n12630), .B(new_n12629), .Y(new_n12631));
  xnor_4 g10283(.A(new_n12630), .B(new_n12629), .Y(new_n12632));
  xnor_4 g10284(.A(new_n12422), .B(new_n12414), .Y(new_n12633));
  nor_5  g10285(.A(new_n12567), .B(new_n12561), .Y(new_n12634));
  xnor_4 g10286(.A(new_n12634), .B(new_n12557), .Y(new_n12635));
  nor_5  g10287(.A(new_n12635), .B(new_n12633), .Y(new_n12636));
  not_8  g10288(.A(new_n12635), .Y(new_n12637));
  xnor_4 g10289(.A(new_n12637), .B(new_n12633), .Y(new_n12638));
  xnor_4 g10290(.A(new_n12566_1), .B(new_n12564), .Y(new_n12639));
  xnor_4 g10291(.A(new_n12419), .B(new_n12418), .Y(new_n12640));
  not_8  g10292(.A(new_n12640), .Y(new_n12641));
  nor_5  g10293(.A(new_n12641), .B(new_n12639), .Y(new_n12642));
  xnor_4 g10294(.A(new_n12415), .B(n11479), .Y(new_n12643));
  xnor_4 g10295(.A(new_n12563), .B(n7876), .Y(new_n12644));
  not_8  g10296(.A(new_n12644), .Y(new_n12645));
  nor_5  g10297(.A(new_n12645), .B(new_n12643), .Y(new_n12646));
  xnor_4 g10298(.A(new_n12640), .B(new_n12639), .Y(new_n12647));
  and_5  g10299(.A(new_n12647), .B(new_n12646), .Y(new_n12648));
  nor_5  g10300(.A(new_n12648), .B(new_n12642), .Y(new_n12649));
  and_5  g10301(.A(new_n12649), .B(new_n12638), .Y(new_n12650_1));
  nor_5  g10302(.A(new_n12650_1), .B(new_n12636), .Y(new_n12651));
  nor_5  g10303(.A(new_n12651), .B(new_n12632), .Y(new_n12652));
  nor_5  g10304(.A(new_n12652), .B(new_n12631), .Y(new_n12653));
  nor_5  g10305(.A(new_n12653), .B(new_n12628), .Y(new_n12654_1));
  nor_5  g10306(.A(new_n12654_1), .B(new_n12627), .Y(new_n12655));
  nor_5  g10307(.A(new_n12655), .B(new_n12624), .Y(new_n12656));
  nor_5  g10308(.A(new_n12656), .B(new_n12623), .Y(new_n12657_1));
  nor_5  g10309(.A(new_n12657_1), .B(new_n12619), .Y(new_n12658));
  nor_5  g10310(.A(new_n12658), .B(new_n12618), .Y(new_n12659));
  nor_5  g10311(.A(new_n12659), .B(new_n12614), .Y(new_n12660));
  nor_5  g10312(.A(new_n12660), .B(new_n12613), .Y(new_n12661));
  nor_5  g10313(.A(new_n12661), .B(new_n12609), .Y(new_n12662));
  nor_5  g10314(.A(new_n12662), .B(new_n12608), .Y(new_n12663));
  nor_5  g10315(.A(new_n12663), .B(new_n12604), .Y(new_n12664));
  nor_5  g10316(.A(new_n12664), .B(new_n12603), .Y(new_n12665_1));
  nor_5  g10317(.A(new_n12665_1), .B(new_n12599), .Y(new_n12666));
  nor_5  g10318(.A(new_n12666), .B(new_n12598), .Y(new_n12667));
  xnor_4 g10319(.A(new_n12667), .B(new_n12593_1), .Y(n2095));
  xnor_4 g10320(.A(new_n11259), .B(new_n11258), .Y(n2105));
  not_8  g10321(.A(new_n6088), .Y(new_n12670_1));
  not_8  g10322(.A(n11898), .Y(new_n12671));
  xnor_4 g10323(.A(n23166), .B(new_n12671), .Y(new_n12672));
  not_8  g10324(.A(n19941), .Y(new_n12673));
  nor_5  g10325(.A(new_n12673), .B(new_n9079), .Y(new_n12674));
  or_5   g10326(.A(n19941), .B(n10577), .Y(new_n12675));
  nor_5  g10327(.A(n6381), .B(n1099), .Y(new_n12676));
  nor_5  g10328(.A(new_n10449), .B(new_n10432_1), .Y(new_n12677));
  nor_5  g10329(.A(new_n12677), .B(new_n12676), .Y(new_n12678));
  and_5  g10330(.A(new_n12678), .B(new_n12675), .Y(new_n12679));
  nor_5  g10331(.A(new_n12679), .B(new_n12674), .Y(new_n12680));
  xor_4  g10332(.A(new_n12680), .B(new_n12672), .Y(new_n12681));
  xnor_4 g10333(.A(new_n12681), .B(n8827), .Y(new_n12682));
  not_8  g10334(.A(n18035), .Y(new_n12683));
  xnor_4 g10335(.A(n19941), .B(new_n9079), .Y(new_n12684));
  xnor_4 g10336(.A(new_n12684), .B(new_n12678), .Y(new_n12685));
  nor_5  g10337(.A(new_n12685), .B(new_n12683), .Y(new_n12686));
  not_8  g10338(.A(new_n12685), .Y(new_n12687));
  xnor_4 g10339(.A(new_n12687), .B(new_n12683), .Y(new_n12688));
  nor_5  g10340(.A(new_n10450), .B(n5077), .Y(new_n12689));
  and_5  g10341(.A(new_n10476), .B(new_n10451), .Y(new_n12690));
  nor_5  g10342(.A(new_n12690), .B(new_n12689), .Y(new_n12691));
  and_5  g10343(.A(new_n12691), .B(new_n12688), .Y(new_n12692));
  or_5   g10344(.A(new_n12692), .B(new_n12686), .Y(new_n12693));
  xor_4  g10345(.A(new_n12693), .B(new_n12682), .Y(new_n12694));
  xnor_4 g10346(.A(new_n12694), .B(new_n12670_1), .Y(new_n12695));
  xnor_4 g10347(.A(new_n12691), .B(new_n12688), .Y(new_n12696));
  nor_5  g10348(.A(new_n12696), .B(new_n6091), .Y(new_n12697));
  not_8  g10349(.A(new_n6091), .Y(new_n12698));
  not_8  g10350(.A(new_n12696), .Y(new_n12699));
  xnor_4 g10351(.A(new_n12699), .B(new_n12698), .Y(new_n12700));
  nor_5  g10352(.A(new_n10477), .B(new_n6097), .Y(new_n12701));
  xnor_4 g10353(.A(new_n10477), .B(new_n6097), .Y(new_n12702_1));
  nor_5  g10354(.A(new_n10480), .B(new_n6102), .Y(new_n12703));
  not_8  g10355(.A(new_n6102), .Y(new_n12704));
  xnor_4 g10356(.A(new_n10481), .B(new_n12704), .Y(new_n12705));
  nor_5  g10357(.A(new_n10485), .B(new_n6107), .Y(new_n12706));
  xnor_4 g10358(.A(new_n10485), .B(new_n6107), .Y(new_n12707_1));
  nor_5  g10359(.A(new_n10491), .B(new_n6112), .Y(new_n12708));
  xnor_4 g10360(.A(new_n10491), .B(new_n6112), .Y(new_n12709));
  nor_5  g10361(.A(new_n8474), .B(new_n6116), .Y(new_n12710));
  xnor_4 g10362(.A(new_n8474), .B(new_n6116), .Y(new_n12711));
  nor_5  g10363(.A(new_n8452), .B(new_n6122), .Y(new_n12712));
  xnor_4 g10364(.A(new_n8452), .B(new_n6122), .Y(new_n12713));
  nor_5  g10365(.A(new_n8455), .B(new_n6132), .Y(new_n12714));
  nor_5  g10366(.A(new_n8459), .B(new_n5793), .Y(new_n12715));
  xnor_4 g10367(.A(new_n8455), .B(new_n6126), .Y(new_n12716));
  and_5  g10368(.A(new_n12716), .B(new_n12715), .Y(new_n12717));
  nor_5  g10369(.A(new_n12717), .B(new_n12714), .Y(new_n12718));
  nor_5  g10370(.A(new_n12718), .B(new_n12713), .Y(new_n12719));
  nor_5  g10371(.A(new_n12719), .B(new_n12712), .Y(new_n12720));
  nor_5  g10372(.A(new_n12720), .B(new_n12711), .Y(new_n12721));
  nor_5  g10373(.A(new_n12721), .B(new_n12710), .Y(new_n12722));
  nor_5  g10374(.A(new_n12722), .B(new_n12709), .Y(new_n12723));
  nor_5  g10375(.A(new_n12723), .B(new_n12708), .Y(new_n12724));
  nor_5  g10376(.A(new_n12724), .B(new_n12707_1), .Y(new_n12725_1));
  nor_5  g10377(.A(new_n12725_1), .B(new_n12706), .Y(new_n12726));
  nor_5  g10378(.A(new_n12726), .B(new_n12705), .Y(new_n12727_1));
  nor_5  g10379(.A(new_n12727_1), .B(new_n12703), .Y(new_n12728));
  nor_5  g10380(.A(new_n12728), .B(new_n12702_1), .Y(new_n12729));
  nor_5  g10381(.A(new_n12729), .B(new_n12701), .Y(new_n12730));
  nor_5  g10382(.A(new_n12730), .B(new_n12700), .Y(new_n12731));
  nor_5  g10383(.A(new_n12731), .B(new_n12697), .Y(new_n12732));
  xnor_4 g10384(.A(new_n12732), .B(new_n12695), .Y(n2122));
  xnor_4 g10385(.A(new_n2837), .B(new_n2809_1), .Y(n2147));
  xnor_4 g10386(.A(new_n10400), .B(new_n10365), .Y(n2209));
  xnor_4 g10387(.A(new_n5771), .B(new_n5663), .Y(n2214));
  xnor_4 g10388(.A(new_n11051), .B(new_n4195), .Y(new_n12737));
  nor_5  g10389(.A(new_n11053), .B(new_n4285), .Y(new_n12738));
  xnor_4 g10390(.A(new_n11055), .B(new_n4285), .Y(new_n12739));
  nor_5  g10391(.A(new_n11069), .B(new_n4293), .Y(new_n12740_1));
  xnor_4 g10392(.A(new_n11058), .B(new_n4293), .Y(new_n12741));
  and_5  g10393(.A(new_n11064), .B(new_n4299), .Y(new_n12742_1));
  nor_5  g10394(.A(new_n11061), .B(new_n4301), .Y(new_n12743));
  xnor_4 g10395(.A(new_n11064), .B(new_n4299), .Y(new_n12744));
  nor_5  g10396(.A(new_n12744), .B(new_n12743), .Y(new_n12745));
  nor_5  g10397(.A(new_n12745), .B(new_n12742_1), .Y(new_n12746_1));
  and_5  g10398(.A(new_n12746_1), .B(new_n12741), .Y(new_n12747));
  nor_5  g10399(.A(new_n12747), .B(new_n12740_1), .Y(new_n12748));
  and_5  g10400(.A(new_n12748), .B(new_n12739), .Y(new_n12749));
  nor_5  g10401(.A(new_n12749), .B(new_n12738), .Y(new_n12750));
  xnor_4 g10402(.A(new_n12750), .B(new_n12737), .Y(n2238));
  xor_4  g10403(.A(new_n11075), .B(new_n11074), .Y(n2327));
  xnor_4 g10404(.A(new_n5755), .B(new_n5724), .Y(n2343));
  not_8  g10405(.A(n13453), .Y(new_n12754));
  xnor_4 g10406(.A(new_n10464), .B(new_n12754), .Y(new_n12755));
  nor_5  g10407(.A(new_n6603), .B(new_n6589), .Y(new_n12756_1));
  and_5  g10408(.A(new_n6621), .B(new_n6605), .Y(new_n12757));
  nor_5  g10409(.A(new_n12757), .B(new_n12756_1), .Y(new_n12758));
  xnor_4 g10410(.A(new_n12758), .B(new_n12755), .Y(new_n12759));
  xnor_4 g10411(.A(n20923), .B(n16524), .Y(new_n12760));
  nor_5  g10412(.A(n18157), .B(n11056), .Y(new_n12761));
  nor_5  g10413(.A(new_n6635), .B(new_n6624), .Y(new_n12762));
  nor_5  g10414(.A(new_n12762), .B(new_n12761), .Y(new_n12763));
  xnor_4 g10415(.A(new_n12763), .B(new_n12760), .Y(new_n12764));
  xnor_4 g10416(.A(new_n12764), .B(n3785), .Y(new_n12765));
  nor_5  g10417(.A(new_n6636), .B(n20250), .Y(new_n12766));
  nor_5  g10418(.A(new_n6650), .B(new_n6637), .Y(new_n12767));
  nor_5  g10419(.A(new_n12767), .B(new_n12766), .Y(new_n12768));
  xnor_4 g10420(.A(new_n12768), .B(new_n12765), .Y(new_n12769));
  not_8  g10421(.A(new_n12769), .Y(new_n12770));
  xnor_4 g10422(.A(new_n12770), .B(new_n12759), .Y(new_n12771));
  nor_5  g10423(.A(new_n6651), .B(new_n6623), .Y(new_n12772));
  and_5  g10424(.A(new_n6673_1), .B(new_n6653), .Y(new_n12773));
  nor_5  g10425(.A(new_n12773), .B(new_n12772), .Y(new_n12774));
  xnor_4 g10426(.A(new_n12774), .B(new_n12771), .Y(n2361));
  xnor_4 g10427(.A(new_n3705), .B(new_n8367), .Y(n2363));
  xnor_4 g10428(.A(new_n4598), .B(new_n4566), .Y(n2374));
  xnor_4 g10429(.A(n7305), .B(n1204), .Y(new_n12778));
  nor_5  g10430(.A(n25872), .B(n19618), .Y(new_n12779));
  and_5  g10431(.A(new_n5830), .B(new_n5825), .Y(new_n12780));
  nor_5  g10432(.A(new_n12780), .B(new_n12779), .Y(new_n12781));
  xnor_4 g10433(.A(new_n12781), .B(new_n12778), .Y(new_n12782));
  nor_5  g10434(.A(new_n12782), .B(new_n4864), .Y(new_n12783_1));
  xor_4  g10435(.A(new_n12782), .B(new_n4864), .Y(new_n12784));
  nor_5  g10436(.A(new_n5831), .B(new_n4880), .Y(new_n12785));
  nor_5  g10437(.A(new_n5841_1), .B(new_n5832), .Y(new_n12786));
  nor_5  g10438(.A(new_n12786), .B(new_n12785), .Y(new_n12787));
  and_5  g10439(.A(new_n12787), .B(new_n12784), .Y(new_n12788));
  nor_5  g10440(.A(new_n12788), .B(new_n12783_1), .Y(new_n12789));
  xnor_4 g10441(.A(n20826), .B(new_n4223), .Y(new_n12790));
  nor_5  g10442(.A(n7305), .B(n1204), .Y(new_n12791));
  nor_5  g10443(.A(new_n12781), .B(new_n12778), .Y(new_n12792));
  or_5   g10444(.A(new_n12792), .B(new_n12791), .Y(new_n12793));
  xor_4  g10445(.A(new_n12793), .B(new_n12790), .Y(new_n12794));
  not_8  g10446(.A(new_n12794), .Y(new_n12795));
  xnor_4 g10447(.A(new_n12795), .B(new_n12789), .Y(new_n12796));
  xnor_4 g10448(.A(new_n12796), .B(new_n4859), .Y(new_n12797));
  xnor_4 g10449(.A(new_n12797), .B(new_n3780), .Y(new_n12798));
  xor_4  g10450(.A(new_n12787), .B(new_n12784), .Y(new_n12799));
  nor_5  g10451(.A(new_n12799), .B(new_n3785_1), .Y(new_n12800));
  nor_5  g10452(.A(new_n5842_1), .B(new_n3790), .Y(new_n12801_1));
  and_5  g10453(.A(new_n5851), .B(new_n5843), .Y(new_n12802));
  nor_5  g10454(.A(new_n12802), .B(new_n12801_1), .Y(new_n12803));
  xnor_4 g10455(.A(new_n12799), .B(new_n3785_1), .Y(new_n12804));
  nor_5  g10456(.A(new_n12804), .B(new_n12803), .Y(new_n12805));
  or_5   g10457(.A(new_n12805), .B(new_n12800), .Y(new_n12806));
  xor_4  g10458(.A(new_n12806), .B(new_n12798), .Y(n2388));
  not_8  g10459(.A(n2160), .Y(new_n12808));
  xnor_4 g10460(.A(n7335), .B(new_n12808), .Y(new_n12809));
  nor_5  g10461(.A(n10763), .B(n5696), .Y(new_n12810));
  and_5  g10462(.A(new_n5334), .B(new_n5305), .Y(new_n12811_1));
  or_5   g10463(.A(new_n12811_1), .B(new_n12810), .Y(new_n12812_1));
  xor_4  g10464(.A(new_n12812_1), .B(new_n12809), .Y(new_n12813));
  xnor_4 g10465(.A(n11220), .B(n3425), .Y(new_n12814));
  nor_5  g10466(.A(n22379), .B(n9967), .Y(new_n12815));
  nor_5  g10467(.A(new_n5303), .B(new_n5271), .Y(new_n12816_1));
  nor_5  g10468(.A(new_n12816_1), .B(new_n12815), .Y(new_n12817));
  xnor_4 g10469(.A(new_n12817), .B(new_n12814), .Y(new_n12818));
  xnor_4 g10470(.A(new_n12818), .B(new_n12813), .Y(new_n12819));
  nor_5  g10471(.A(new_n5335), .B(new_n5304), .Y(new_n12820));
  nor_5  g10472(.A(new_n5398), .B(new_n5336), .Y(new_n12821_1));
  nor_5  g10473(.A(new_n12821_1), .B(new_n12820), .Y(new_n12822));
  xnor_4 g10474(.A(new_n12822), .B(new_n12819), .Y(new_n12823));
  not_8  g10475(.A(new_n12823), .Y(new_n12824));
  not_8  g10476(.A(new_n5231), .Y(new_n12825));
  nor_5  g10477(.A(new_n12825), .B(n337), .Y(new_n12826));
  xnor_4 g10478(.A(new_n12826), .B(n7593), .Y(new_n12827));
  xnor_4 g10479(.A(new_n12827), .B(new_n3086), .Y(new_n12828));
  nor_5  g10480(.A(new_n5232), .B(n6485), .Y(new_n12829));
  and_5  g10481(.A(new_n5269), .B(new_n5233), .Y(new_n12830));
  nor_5  g10482(.A(new_n12830), .B(new_n12829), .Y(new_n12831));
  xnor_4 g10483(.A(new_n12831), .B(new_n12828), .Y(new_n12832));
  xnor_4 g10484(.A(new_n12832), .B(new_n12824), .Y(new_n12833));
  nor_5  g10485(.A(new_n5399_1), .B(new_n5270), .Y(new_n12834));
  and_5  g10486(.A(new_n5451_1), .B(new_n5401), .Y(new_n12835));
  or_5   g10487(.A(new_n12835), .B(new_n12834), .Y(new_n12836));
  xor_4  g10488(.A(new_n12836), .B(new_n12833), .Y(n2440));
  xnor_4 g10489(.A(new_n11407), .B(new_n11394), .Y(n2444));
  xnor_4 g10490(.A(new_n5083), .B(new_n3257), .Y(n2513));
  xnor_4 g10491(.A(new_n5943_1), .B(n14323), .Y(new_n12840));
  not_8  g10492(.A(n2886), .Y(new_n12841));
  nor_5  g10493(.A(new_n5950), .B(new_n12841), .Y(new_n12842));
  xnor_4 g10494(.A(new_n5950), .B(n2886), .Y(new_n12843_1));
  nor_5  g10495(.A(new_n5961), .B(new_n12373), .Y(new_n12844));
  nor_5  g10496(.A(new_n3798), .B(new_n12371), .Y(new_n12845));
  xnor_4 g10497(.A(new_n5961), .B(n1040), .Y(new_n12846));
  and_5  g10498(.A(new_n12846), .B(new_n12845), .Y(new_n12847));
  or_5   g10499(.A(new_n12847), .B(new_n12844), .Y(new_n12848));
  and_5  g10500(.A(new_n12848), .B(new_n12843_1), .Y(new_n12849));
  nor_5  g10501(.A(new_n12849), .B(new_n12842), .Y(new_n12850));
  xnor_4 g10502(.A(new_n12850), .B(new_n12840), .Y(new_n12851));
  xnor_4 g10503(.A(new_n12851), .B(n12562), .Y(new_n12852));
  xor_4  g10504(.A(new_n12848), .B(new_n12843_1), .Y(new_n12853));
  nor_5  g10505(.A(new_n12853), .B(n7949), .Y(new_n12854));
  xnor_4 g10506(.A(new_n12853), .B(new_n5892), .Y(new_n12855));
  nor_5  g10507(.A(new_n10778), .B(new_n5895), .Y(new_n12856));
  nor_5  g10508(.A(new_n12856), .B(n24374), .Y(new_n12857));
  xnor_4 g10509(.A(new_n12846), .B(new_n12845), .Y(new_n12858));
  xor_4  g10510(.A(new_n12856), .B(n24374), .Y(new_n12859));
  and_5  g10511(.A(new_n12859), .B(new_n12858), .Y(new_n12860));
  or_5   g10512(.A(new_n12860), .B(new_n12857), .Y(new_n12861_1));
  and_5  g10513(.A(new_n12861_1), .B(new_n12855), .Y(new_n12862));
  nor_5  g10514(.A(new_n12862), .B(new_n12854), .Y(new_n12863));
  xor_4  g10515(.A(new_n12863), .B(new_n12852), .Y(new_n12864_1));
  xnor_4 g10516(.A(new_n12864_1), .B(new_n12630), .Y(new_n12865_1));
  xor_4  g10517(.A(new_n12861_1), .B(new_n12855), .Y(new_n12866));
  and_5  g10518(.A(new_n12866), .B(new_n12637), .Y(new_n12867));
  xnor_4 g10519(.A(new_n12866), .B(new_n12637), .Y(new_n12868));
  not_8  g10520(.A(new_n12858), .Y(new_n12869));
  xnor_4 g10521(.A(new_n12859), .B(new_n12869), .Y(new_n12870_1));
  and_5  g10522(.A(new_n12870_1), .B(new_n12639), .Y(new_n12871_1));
  xnor_4 g10523(.A(new_n10778), .B(n14575), .Y(new_n12872));
  and_5  g10524(.A(new_n12872), .B(new_n12644), .Y(new_n12873_1));
  xnor_4 g10525(.A(new_n12870_1), .B(new_n12639), .Y(new_n12874));
  nor_5  g10526(.A(new_n12874), .B(new_n12873_1), .Y(new_n12875_1));
  nor_5  g10527(.A(new_n12875_1), .B(new_n12871_1), .Y(new_n12876));
  nor_5  g10528(.A(new_n12876), .B(new_n12868), .Y(new_n12877));
  nor_5  g10529(.A(new_n12877), .B(new_n12867), .Y(new_n12878));
  xnor_4 g10530(.A(new_n12878), .B(new_n12865_1), .Y(n2515));
  xnor_4 g10531(.A(new_n10769), .B(new_n10741), .Y(n2533));
  nor_5  g10532(.A(n26986), .B(new_n3217), .Y(new_n12881));
  xnor_4 g10533(.A(n26986), .B(n3425), .Y(new_n12882));
  nor_5  g10534(.A(n21287), .B(new_n3198), .Y(new_n12883));
  xnor_4 g10535(.A(n21287), .B(n9967), .Y(new_n12884));
  nor_5  g10536(.A(new_n7508), .B(n4256), .Y(new_n12885));
  xnor_4 g10537(.A(n20946), .B(n4256), .Y(new_n12886));
  nor_5  g10538(.A(n22332), .B(new_n5275), .Y(new_n12887));
  xnor_4 g10539(.A(n22332), .B(n7751), .Y(new_n12888));
  not_8  g10540(.A(n26823), .Y(new_n12889));
  nor_5  g10541(.A(new_n12889), .B(n18907), .Y(new_n12890));
  xnor_4 g10542(.A(n26823), .B(n18907), .Y(new_n12891));
  nor_5  g10543(.A(new_n5280), .B(n2731), .Y(new_n12892_1));
  and_5  g10544(.A(new_n8409), .B(new_n8393), .Y(new_n12893));
  or_5   g10545(.A(new_n12893), .B(new_n12892_1), .Y(new_n12894));
  and_5  g10546(.A(new_n12894), .B(new_n12891), .Y(new_n12895));
  or_5   g10547(.A(new_n12895), .B(new_n12890), .Y(new_n12896));
  and_5  g10548(.A(new_n12896), .B(new_n12888), .Y(new_n12897));
  or_5   g10549(.A(new_n12897), .B(new_n12887), .Y(new_n12898));
  and_5  g10550(.A(new_n12898), .B(new_n12886), .Y(new_n12899));
  or_5   g10551(.A(new_n12899), .B(new_n12885), .Y(new_n12900_1));
  and_5  g10552(.A(new_n12900_1), .B(new_n12884), .Y(new_n12901));
  or_5   g10553(.A(new_n12901), .B(new_n12883), .Y(new_n12902));
  and_5  g10554(.A(new_n12902), .B(new_n12882), .Y(new_n12903));
  nor_5  g10555(.A(new_n12903), .B(new_n12881), .Y(new_n12904_1));
  not_8  g10556(.A(new_n7059), .Y(new_n12905));
  not_8  g10557(.A(new_n7064), .Y(new_n12906));
  not_8  g10558(.A(new_n5124), .Y(new_n12907));
  nor_5  g10559(.A(new_n5132), .B(new_n12907), .Y(new_n12908));
  not_8  g10560(.A(new_n12908), .Y(new_n12909));
  not_8  g10561(.A(new_n7068), .Y(new_n12910));
  nor_5  g10562(.A(new_n12910), .B(new_n12909), .Y(new_n12911));
  not_8  g10563(.A(new_n12911), .Y(new_n12912));
  nor_5  g10564(.A(new_n12912), .B(new_n12906), .Y(new_n12913));
  not_8  g10565(.A(new_n12913), .Y(new_n12914));
  nor_5  g10566(.A(new_n12914), .B(new_n12905), .Y(new_n12915));
  and_5  g10567(.A(new_n12915), .B(new_n7116), .Y(new_n12916));
  and_5  g10568(.A(new_n12916), .B(new_n7186), .Y(new_n12917_1));
  not_8  g10569(.A(new_n7189), .Y(new_n12918));
  nor_5  g10570(.A(new_n12916), .B(new_n12918), .Y(new_n12919));
  nor_5  g10571(.A(new_n12919), .B(new_n12917_1), .Y(new_n12920));
  nor_5  g10572(.A(new_n12920), .B(new_n3195), .Y(new_n12921));
  xor_4  g10573(.A(new_n12915), .B(new_n7116), .Y(new_n12922));
  nor_5  g10574(.A(new_n12922), .B(new_n3137), .Y(new_n12923));
  xnor_4 g10575(.A(new_n12922), .B(new_n3137), .Y(new_n12924));
  xnor_4 g10576(.A(new_n12913), .B(new_n12905), .Y(new_n12925));
  nor_5  g10577(.A(new_n12925), .B(new_n3141), .Y(new_n12926));
  xnor_4 g10578(.A(new_n12925), .B(new_n3141), .Y(new_n12927));
  xnor_4 g10579(.A(new_n12911), .B(new_n12906), .Y(new_n12928));
  nor_5  g10580(.A(new_n12928), .B(new_n3145), .Y(new_n12929));
  xnor_4 g10581(.A(new_n12928), .B(new_n3145), .Y(new_n12930));
  xnor_4 g10582(.A(new_n12910), .B(new_n12908), .Y(new_n12931));
  nor_5  g10583(.A(new_n12931), .B(new_n3149), .Y(new_n12932));
  xnor_4 g10584(.A(new_n12931), .B(new_n3149), .Y(new_n12933));
  nor_5  g10585(.A(new_n5133), .B(new_n3153), .Y(new_n12934));
  nor_5  g10586(.A(new_n5159), .B(new_n5134), .Y(new_n12935));
  nor_5  g10587(.A(new_n12935), .B(new_n12934), .Y(new_n12936));
  nor_5  g10588(.A(new_n12936), .B(new_n12933), .Y(new_n12937));
  nor_5  g10589(.A(new_n12937), .B(new_n12932), .Y(new_n12938));
  nor_5  g10590(.A(new_n12938), .B(new_n12930), .Y(new_n12939));
  nor_5  g10591(.A(new_n12939), .B(new_n12929), .Y(new_n12940));
  nor_5  g10592(.A(new_n12940), .B(new_n12927), .Y(new_n12941_1));
  nor_5  g10593(.A(new_n12941_1), .B(new_n12926), .Y(new_n12942_1));
  nor_5  g10594(.A(new_n12942_1), .B(new_n12924), .Y(new_n12943));
  nor_5  g10595(.A(new_n12943), .B(new_n12923), .Y(new_n12944));
  and_5  g10596(.A(new_n12920), .B(new_n3195), .Y(new_n12945));
  nor_5  g10597(.A(new_n12945), .B(new_n12944), .Y(new_n12946));
  nor_5  g10598(.A(new_n12946), .B(new_n12921), .Y(new_n12947));
  nor_5  g10599(.A(new_n12947), .B(new_n12917_1), .Y(new_n12948));
  xnor_4 g10600(.A(new_n12948), .B(new_n12904_1), .Y(new_n12949));
  xnor_4 g10601(.A(new_n12920), .B(new_n3196), .Y(new_n12950));
  xnor_4 g10602(.A(new_n12950), .B(new_n12944), .Y(new_n12951));
  not_8  g10603(.A(new_n12951), .Y(new_n12952));
  nor_5  g10604(.A(new_n12952), .B(new_n12904_1), .Y(new_n12953));
  xnor_4 g10605(.A(new_n12952), .B(new_n12904_1), .Y(new_n12954));
  xor_4  g10606(.A(new_n12902), .B(new_n12882), .Y(new_n12955));
  xnor_4 g10607(.A(new_n12942_1), .B(new_n12924), .Y(new_n12956_1));
  nor_5  g10608(.A(new_n12956_1), .B(new_n12955), .Y(new_n12957));
  xnor_4 g10609(.A(new_n12956_1), .B(new_n12955), .Y(new_n12958));
  xor_4  g10610(.A(new_n12900_1), .B(new_n12884), .Y(new_n12959));
  xnor_4 g10611(.A(new_n12940), .B(new_n12927), .Y(new_n12960));
  nor_5  g10612(.A(new_n12960), .B(new_n12959), .Y(new_n12961));
  xnor_4 g10613(.A(new_n12960), .B(new_n12959), .Y(new_n12962));
  xor_4  g10614(.A(new_n12898), .B(new_n12886), .Y(new_n12963));
  xnor_4 g10615(.A(new_n12938), .B(new_n12930), .Y(new_n12964));
  nor_5  g10616(.A(new_n12964), .B(new_n12963), .Y(new_n12965));
  xnor_4 g10617(.A(new_n12964), .B(new_n12963), .Y(new_n12966));
  xor_4  g10618(.A(new_n12896), .B(new_n12888), .Y(new_n12967));
  xnor_4 g10619(.A(new_n12936), .B(new_n12933), .Y(new_n12968));
  nor_5  g10620(.A(new_n12968), .B(new_n12967), .Y(new_n12969));
  not_8  g10621(.A(new_n12968), .Y(new_n12970));
  xnor_4 g10622(.A(new_n12970), .B(new_n12967), .Y(new_n12971));
  xor_4  g10623(.A(new_n12894), .B(new_n12891), .Y(new_n12972));
  and_5  g10624(.A(new_n12972), .B(new_n5160), .Y(new_n12973));
  xnor_4 g10625(.A(new_n12972), .B(new_n5161), .Y(new_n12974));
  and_5  g10626(.A(new_n8410), .B(new_n5187), .Y(new_n12975));
  and_5  g10627(.A(new_n8430), .B(new_n8411), .Y(new_n12976));
  or_5   g10628(.A(new_n12976), .B(new_n12975), .Y(new_n12977));
  and_5  g10629(.A(new_n12977), .B(new_n12974), .Y(new_n12978_1));
  nor_5  g10630(.A(new_n12978_1), .B(new_n12973), .Y(new_n12979));
  and_5  g10631(.A(new_n12979), .B(new_n12971), .Y(new_n12980_1));
  nor_5  g10632(.A(new_n12980_1), .B(new_n12969), .Y(new_n12981));
  nor_5  g10633(.A(new_n12981), .B(new_n12966), .Y(new_n12982));
  nor_5  g10634(.A(new_n12982), .B(new_n12965), .Y(new_n12983));
  nor_5  g10635(.A(new_n12983), .B(new_n12962), .Y(new_n12984));
  nor_5  g10636(.A(new_n12984), .B(new_n12961), .Y(new_n12985_1));
  nor_5  g10637(.A(new_n12985_1), .B(new_n12958), .Y(new_n12986));
  nor_5  g10638(.A(new_n12986), .B(new_n12957), .Y(new_n12987_1));
  nor_5  g10639(.A(new_n12987_1), .B(new_n12954), .Y(new_n12988));
  nor_5  g10640(.A(new_n12988), .B(new_n12953), .Y(new_n12989));
  xnor_4 g10641(.A(new_n12989), .B(new_n12949), .Y(n2535));
  nor_5  g10642(.A(n20259), .B(n3925), .Y(new_n12991));
  not_8  g10643(.A(new_n12991), .Y(new_n12992_1));
  nor_5  g10644(.A(new_n12992_1), .B(n25872), .Y(new_n12993));
  not_8  g10645(.A(new_n12993), .Y(new_n12994));
  nor_5  g10646(.A(new_n12994), .B(n7305), .Y(new_n12995));
  not_8  g10647(.A(new_n12995), .Y(new_n12996));
  nor_5  g10648(.A(new_n12996), .B(n20826), .Y(new_n12997));
  xnor_4 g10649(.A(new_n12997), .B(n22198), .Y(new_n12998));
  xnor_4 g10650(.A(new_n12998), .B(n21674), .Y(new_n12999));
  xnor_4 g10651(.A(new_n12995), .B(n20826), .Y(new_n13000));
  nor_5  g10652(.A(new_n13000), .B(n17251), .Y(new_n13001));
  xnor_4 g10653(.A(new_n13000), .B(n17251), .Y(new_n13002));
  xnor_4 g10654(.A(new_n12993), .B(n7305), .Y(new_n13003));
  nor_5  g10655(.A(new_n13003), .B(n14790), .Y(new_n13004));
  xnor_4 g10656(.A(new_n12991), .B(n25872), .Y(new_n13005_1));
  nor_5  g10657(.A(new_n13005_1), .B(n10096), .Y(new_n13006));
  xnor_4 g10658(.A(new_n13005_1), .B(new_n3555_1), .Y(new_n13007));
  xnor_4 g10659(.A(n20259), .B(n3925), .Y(new_n13008));
  and_5  g10660(.A(new_n13008), .B(new_n3558), .Y(new_n13009));
  or_5   g10661(.A(new_n3562), .B(new_n5002), .Y(new_n13010));
  xnor_4 g10662(.A(new_n13008), .B(n16994), .Y(new_n13011));
  and_5  g10663(.A(new_n13011), .B(new_n13010), .Y(new_n13012));
  or_5   g10664(.A(new_n13012), .B(new_n13009), .Y(new_n13013));
  and_5  g10665(.A(new_n13013), .B(new_n13007), .Y(new_n13014));
  nor_5  g10666(.A(new_n13014), .B(new_n13006), .Y(new_n13015));
  xnor_4 g10667(.A(new_n13003), .B(n14790), .Y(new_n13016));
  nor_5  g10668(.A(new_n13016), .B(new_n13015), .Y(new_n13017));
  nor_5  g10669(.A(new_n13017), .B(new_n13004), .Y(new_n13018));
  nor_5  g10670(.A(new_n13018), .B(new_n13002), .Y(new_n13019));
  nor_5  g10671(.A(new_n13019), .B(new_n13001), .Y(new_n13020));
  xnor_4 g10672(.A(new_n13020), .B(new_n12999), .Y(new_n13021));
  xnor_4 g10673(.A(new_n13021), .B(new_n7722), .Y(new_n13022));
  xnor_4 g10674(.A(new_n13018), .B(new_n13002), .Y(new_n13023));
  nor_5  g10675(.A(new_n13023), .B(new_n7726), .Y(new_n13024));
  xnor_4 g10676(.A(new_n13023), .B(new_n7726), .Y(new_n13025));
  xnor_4 g10677(.A(new_n13016), .B(new_n13015), .Y(new_n13026_1));
  nor_5  g10678(.A(new_n13026_1), .B(new_n7731_1), .Y(new_n13027));
  xor_4  g10679(.A(new_n13026_1), .B(new_n7731_1), .Y(new_n13028));
  xor_4  g10680(.A(new_n13013), .B(new_n13007), .Y(new_n13029));
  nor_5  g10681(.A(new_n13029), .B(new_n7737), .Y(new_n13030));
  xnor_4 g10682(.A(new_n13029), .B(new_n7737), .Y(new_n13031));
  xor_4  g10683(.A(new_n13011), .B(new_n13010), .Y(new_n13032));
  nor_5  g10684(.A(new_n13032), .B(new_n7745), .Y(new_n13033));
  nor_5  g10685(.A(new_n9707), .B(new_n7749), .Y(new_n13034));
  xnor_4 g10686(.A(new_n13032), .B(new_n7746), .Y(new_n13035));
  and_5  g10687(.A(new_n13035), .B(new_n13034), .Y(new_n13036));
  nor_5  g10688(.A(new_n13036), .B(new_n13033), .Y(new_n13037));
  nor_5  g10689(.A(new_n13037), .B(new_n13031), .Y(new_n13038));
  nor_5  g10690(.A(new_n13038), .B(new_n13030), .Y(new_n13039));
  and_5  g10691(.A(new_n13039), .B(new_n13028), .Y(new_n13040));
  nor_5  g10692(.A(new_n13040), .B(new_n13027), .Y(new_n13041));
  nor_5  g10693(.A(new_n13041), .B(new_n13025), .Y(new_n13042));
  nor_5  g10694(.A(new_n13042), .B(new_n13024), .Y(new_n13043_1));
  xnor_4 g10695(.A(new_n13043_1), .B(new_n13022), .Y(new_n13044_1));
  xnor_4 g10696(.A(n1163), .B(n329), .Y(new_n13045));
  not_8  g10697(.A(n24170), .Y(new_n13046));
  nor_5  g10698(.A(new_n13046), .B(n18537), .Y(new_n13047));
  xnor_4 g10699(.A(n24170), .B(n18537), .Y(new_n13048_1));
  not_8  g10700(.A(n2409), .Y(new_n13049));
  nor_5  g10701(.A(n7057), .B(new_n13049), .Y(new_n13050));
  xnor_4 g10702(.A(n7057), .B(n2409), .Y(new_n13051));
  nor_5  g10703(.A(n8869), .B(new_n8510_1), .Y(new_n13052));
  and_5  g10704(.A(n8869), .B(new_n8510_1), .Y(new_n13053));
  nor_5  g10705(.A(new_n5040), .B(n10372), .Y(new_n13054_1));
  nor_5  g10706(.A(new_n5080), .B(n7428), .Y(new_n13055));
  nand_5 g10707(.A(new_n5040), .B(n10372), .Y(new_n13056));
  and_5  g10708(.A(new_n13056), .B(new_n13055), .Y(new_n13057));
  nor_5  g10709(.A(new_n13057), .B(new_n13054_1), .Y(new_n13058));
  nor_5  g10710(.A(new_n13058), .B(new_n13053), .Y(new_n13059));
  nor_5  g10711(.A(new_n13059), .B(new_n13052), .Y(new_n13060));
  and_5  g10712(.A(new_n13060), .B(new_n13051), .Y(new_n13061));
  or_5   g10713(.A(new_n13061), .B(new_n13050), .Y(new_n13062));
  and_5  g10714(.A(new_n13062), .B(new_n13048_1), .Y(new_n13063));
  or_5   g10715(.A(new_n13063), .B(new_n13047), .Y(new_n13064));
  xor_4  g10716(.A(new_n13064), .B(new_n13045), .Y(new_n13065));
  xnor_4 g10717(.A(new_n13065), .B(new_n13044_1), .Y(new_n13066));
  xor_4  g10718(.A(new_n13062), .B(new_n13048_1), .Y(new_n13067));
  xnor_4 g10719(.A(new_n13041), .B(new_n13025), .Y(new_n13068));
  nor_5  g10720(.A(new_n13068), .B(new_n13067), .Y(new_n13069));
  xnor_4 g10721(.A(new_n13068), .B(new_n13067), .Y(new_n13070));
  xnor_4 g10722(.A(new_n13039), .B(new_n13028), .Y(new_n13071));
  not_8  g10723(.A(new_n13071), .Y(new_n13072));
  xnor_4 g10724(.A(new_n13060), .B(new_n13051), .Y(new_n13073));
  and_5  g10725(.A(new_n13073), .B(new_n13072), .Y(new_n13074_1));
  xnor_4 g10726(.A(new_n13073), .B(new_n13072), .Y(new_n13075));
  xnor_4 g10727(.A(new_n13037), .B(new_n13031), .Y(new_n13076));
  xnor_4 g10728(.A(n8869), .B(n8381), .Y(new_n13077));
  xnor_4 g10729(.A(new_n13077), .B(new_n13058), .Y(new_n13078));
  and_5  g10730(.A(new_n13078), .B(new_n13076), .Y(new_n13079));
  xnor_4 g10731(.A(new_n13078), .B(new_n13076), .Y(new_n13080));
  nor_5  g10732(.A(new_n9710), .B(new_n9708), .Y(new_n13081));
  xnor_4 g10733(.A(n20235), .B(n10372), .Y(new_n13082_1));
  xnor_4 g10734(.A(new_n13082_1), .B(new_n13055), .Y(new_n13083));
  nor_5  g10735(.A(new_n13083), .B(new_n13081), .Y(new_n13084));
  xnor_4 g10736(.A(new_n13035), .B(new_n13034), .Y(new_n13085));
  not_8  g10737(.A(new_n13085), .Y(new_n13086));
  xnor_4 g10738(.A(new_n13083), .B(new_n13081), .Y(new_n13087));
  nor_5  g10739(.A(new_n13087), .B(new_n13086), .Y(new_n13088));
  nor_5  g10740(.A(new_n13088), .B(new_n13084), .Y(new_n13089));
  nor_5  g10741(.A(new_n13089), .B(new_n13080), .Y(new_n13090));
  nor_5  g10742(.A(new_n13090), .B(new_n13079), .Y(new_n13091));
  nor_5  g10743(.A(new_n13091), .B(new_n13075), .Y(new_n13092));
  nor_5  g10744(.A(new_n13092), .B(new_n13074_1), .Y(new_n13093));
  nor_5  g10745(.A(new_n13093), .B(new_n13070), .Y(new_n13094));
  nor_5  g10746(.A(new_n13094), .B(new_n13069), .Y(new_n13095));
  xnor_4 g10747(.A(new_n13095), .B(new_n13066), .Y(n2537));
  not_8  g10748(.A(new_n2987), .Y(new_n13097));
  xnor_4 g10749(.A(new_n10936), .B(new_n13097), .Y(new_n13098));
  nor_5  g10750(.A(new_n4202), .B(new_n2994), .Y(new_n13099));
  xnor_4 g10751(.A(new_n4201), .B(new_n2994), .Y(new_n13100));
  nor_5  g10752(.A(new_n4204_1), .B(new_n2998), .Y(new_n13101));
  xnor_4 g10753(.A(new_n4204_1), .B(new_n3000), .Y(new_n13102));
  nor_5  g10754(.A(new_n4208), .B(new_n3004), .Y(new_n13103));
  xnor_4 g10755(.A(new_n4207), .B(new_n3004), .Y(new_n13104));
  and_5  g10756(.A(new_n4211), .B(new_n3010_1), .Y(new_n13105));
  nor_5  g10757(.A(new_n3015), .B(n1152), .Y(new_n13106));
  xnor_4 g10758(.A(new_n4211), .B(new_n3011), .Y(new_n13107));
  and_5  g10759(.A(new_n13107), .B(new_n13106), .Y(new_n13108));
  nor_5  g10760(.A(new_n13108), .B(new_n13105), .Y(new_n13109));
  and_5  g10761(.A(new_n13109), .B(new_n13104), .Y(new_n13110_1));
  nor_5  g10762(.A(new_n13110_1), .B(new_n13103), .Y(new_n13111));
  and_5  g10763(.A(new_n13111), .B(new_n13102), .Y(new_n13112));
  nor_5  g10764(.A(new_n13112), .B(new_n13101), .Y(new_n13113));
  and_5  g10765(.A(new_n13113), .B(new_n13100), .Y(new_n13114));
  or_5   g10766(.A(new_n13114), .B(new_n13099), .Y(new_n13115));
  xor_4  g10767(.A(new_n13115), .B(new_n13098), .Y(new_n13116_1));
  xnor_4 g10768(.A(new_n13116_1), .B(new_n11357), .Y(new_n13117));
  xor_4  g10769(.A(new_n13113), .B(new_n13100), .Y(new_n13118));
  nor_5  g10770(.A(new_n13118), .B(new_n9517), .Y(new_n13119));
  xnor_4 g10771(.A(new_n13118), .B(new_n9517), .Y(new_n13120));
  xnor_4 g10772(.A(new_n13111), .B(new_n13102), .Y(new_n13121));
  nor_5  g10773(.A(new_n13121), .B(new_n9520), .Y(new_n13122_1));
  xnor_4 g10774(.A(new_n13121), .B(new_n11875), .Y(new_n13123));
  xnor_4 g10775(.A(new_n13109), .B(new_n13104), .Y(new_n13124));
  nor_5  g10776(.A(new_n13124), .B(new_n9528), .Y(new_n13125));
  xnor_4 g10777(.A(new_n13124), .B(new_n9525), .Y(new_n13126));
  xnor_4 g10778(.A(new_n13107), .B(new_n13106), .Y(new_n13127));
  nor_5  g10779(.A(new_n13127), .B(new_n9530), .Y(new_n13128));
  xnor_4 g10780(.A(new_n3015), .B(new_n2698), .Y(new_n13129));
  nor_5  g10781(.A(new_n13129), .B(new_n7200), .Y(new_n13130));
  xnor_4 g10782(.A(new_n13127), .B(new_n9530), .Y(new_n13131));
  nor_5  g10783(.A(new_n13131), .B(new_n13130), .Y(new_n13132));
  nor_5  g10784(.A(new_n13132), .B(new_n13128), .Y(new_n13133));
  and_5  g10785(.A(new_n13133), .B(new_n13126), .Y(new_n13134));
  nor_5  g10786(.A(new_n13134), .B(new_n13125), .Y(new_n13135));
  and_5  g10787(.A(new_n13135), .B(new_n13123), .Y(new_n13136));
  nor_5  g10788(.A(new_n13136), .B(new_n13122_1), .Y(new_n13137_1));
  nor_5  g10789(.A(new_n13137_1), .B(new_n13120), .Y(new_n13138));
  nor_5  g10790(.A(new_n13138), .B(new_n13119), .Y(new_n13139));
  xnor_4 g10791(.A(new_n13139), .B(new_n13117), .Y(n2553));
  xnor_4 g10792(.A(new_n11779), .B(new_n11761), .Y(n2555));
  xnor_4 g10793(.A(new_n10607), .B(n12892), .Y(new_n13142));
  not_8  g10794(.A(new_n13142), .Y(new_n13143));
  nor_5  g10795(.A(new_n13143), .B(new_n9962), .Y(new_n13144_1));
  not_8  g10796(.A(n12892), .Y(new_n13145));
  nor_5  g10797(.A(new_n10607), .B(new_n13145), .Y(new_n13146));
  not_8  g10798(.A(new_n10611_1), .Y(new_n13147));
  xnor_4 g10799(.A(new_n13147), .B(n12209), .Y(new_n13148));
  xnor_4 g10800(.A(new_n13148), .B(new_n13146), .Y(new_n13149));
  not_8  g10801(.A(new_n13149), .Y(new_n13150));
  xnor_4 g10802(.A(new_n13150), .B(new_n9965), .Y(new_n13151));
  xnor_4 g10803(.A(new_n13151), .B(new_n13144_1), .Y(n2560));
  nor_5  g10804(.A(n26180), .B(n10650), .Y(new_n13153));
  xnor_4 g10805(.A(n26180), .B(n10650), .Y(new_n13154));
  nor_5  g10806(.A(n24004), .B(n12900), .Y(new_n13155));
  xnor_4 g10807(.A(n24004), .B(n12900), .Y(new_n13156));
  nor_5  g10808(.A(n20411), .B(n12871), .Y(new_n13157));
  xnor_4 g10809(.A(n20411), .B(n12871), .Y(new_n13158));
  nor_5  g10810(.A(n23304), .B(n17069), .Y(new_n13159));
  xnor_4 g10811(.A(n23304), .B(n17069), .Y(new_n13160));
  nor_5  g10812(.A(n19361), .B(n15918), .Y(new_n13161));
  xnor_4 g10813(.A(n19361), .B(n15918), .Y(new_n13162));
  nor_5  g10814(.A(n17784), .B(n1437), .Y(new_n13163));
  xnor_4 g10815(.A(n17784), .B(new_n3497), .Y(new_n13164));
  nor_5  g10816(.A(n14323), .B(n4722), .Y(new_n13165));
  xnor_4 g10817(.A(n14323), .B(new_n3503), .Y(new_n13166));
  nor_5  g10818(.A(n14633), .B(n2886), .Y(new_n13167));
  xnor_4 g10819(.A(n14633), .B(new_n12841), .Y(new_n13168_1));
  nor_5  g10820(.A(n8721), .B(n1040), .Y(new_n13169));
  or_5   g10821(.A(new_n3515), .B(new_n12371), .Y(new_n13170));
  xnor_4 g10822(.A(n8721), .B(new_n12373), .Y(new_n13171));
  and_5  g10823(.A(new_n13171), .B(new_n13170), .Y(new_n13172));
  or_5   g10824(.A(new_n13172), .B(new_n13169), .Y(new_n13173));
  and_5  g10825(.A(new_n13173), .B(new_n13168_1), .Y(new_n13174));
  or_5   g10826(.A(new_n13174), .B(new_n13167), .Y(new_n13175));
  and_5  g10827(.A(new_n13175), .B(new_n13166), .Y(new_n13176));
  or_5   g10828(.A(new_n13176), .B(new_n13165), .Y(new_n13177));
  and_5  g10829(.A(new_n13177), .B(new_n13164), .Y(new_n13178));
  nor_5  g10830(.A(new_n13178), .B(new_n13163), .Y(new_n13179));
  nor_5  g10831(.A(new_n13179), .B(new_n13162), .Y(new_n13180));
  nor_5  g10832(.A(new_n13180), .B(new_n13161), .Y(new_n13181));
  nor_5  g10833(.A(new_n13181), .B(new_n13160), .Y(new_n13182));
  nor_5  g10834(.A(new_n13182), .B(new_n13159), .Y(new_n13183));
  nor_5  g10835(.A(new_n13183), .B(new_n13158), .Y(new_n13184));
  nor_5  g10836(.A(new_n13184), .B(new_n13157), .Y(new_n13185));
  nor_5  g10837(.A(new_n13185), .B(new_n13156), .Y(new_n13186));
  nor_5  g10838(.A(new_n13186), .B(new_n13155), .Y(new_n13187));
  nor_5  g10839(.A(new_n13187), .B(new_n13154), .Y(new_n13188));
  nor_5  g10840(.A(new_n13188), .B(new_n13153), .Y(new_n13189));
  nor_5  g10841(.A(n9259), .B(n6456), .Y(new_n13190_1));
  or_5   g10842(.A(new_n5912), .B(new_n5874), .Y(new_n13191));
  and_5  g10843(.A(new_n13191), .B(new_n5873), .Y(new_n13192));
  nor_5  g10844(.A(new_n13192), .B(new_n13190_1), .Y(new_n13193));
  not_8  g10845(.A(new_n13193), .Y(new_n13194));
  nor_5  g10846(.A(new_n13194), .B(new_n13189), .Y(new_n13195));
  xnor_4 g10847(.A(new_n13194), .B(new_n13189), .Y(new_n13196));
  xnor_4 g10848(.A(new_n13187), .B(new_n13154), .Y(new_n13197));
  nor_5  g10849(.A(new_n13197), .B(new_n5914), .Y(new_n13198_1));
  xnor_4 g10850(.A(new_n13197), .B(new_n5914), .Y(new_n13199_1));
  xnor_4 g10851(.A(new_n13185), .B(new_n13156), .Y(new_n13200));
  nor_5  g10852(.A(new_n13200), .B(new_n5919), .Y(new_n13201));
  xnor_4 g10853(.A(new_n13200), .B(new_n5919), .Y(new_n13202));
  xnor_4 g10854(.A(new_n13183), .B(new_n13158), .Y(new_n13203));
  nor_5  g10855(.A(new_n13203), .B(new_n5925), .Y(new_n13204_1));
  xnor_4 g10856(.A(new_n13203), .B(new_n5925), .Y(new_n13205));
  xnor_4 g10857(.A(new_n13181), .B(new_n13160), .Y(new_n13206));
  nor_5  g10858(.A(new_n13206), .B(new_n5930), .Y(new_n13207));
  xnor_4 g10859(.A(new_n13206), .B(new_n5930), .Y(new_n13208));
  xnor_4 g10860(.A(new_n13179), .B(new_n13162), .Y(new_n13209_1));
  nor_5  g10861(.A(new_n13209_1), .B(new_n5935), .Y(new_n13210));
  not_8  g10862(.A(new_n5935), .Y(new_n13211));
  xnor_4 g10863(.A(new_n13209_1), .B(new_n13211), .Y(new_n13212));
  not_8  g10864(.A(new_n5940), .Y(new_n13213));
  xor_4  g10865(.A(new_n13177), .B(new_n13164), .Y(new_n13214));
  nor_5  g10866(.A(new_n13214), .B(new_n13213), .Y(new_n13215));
  xnor_4 g10867(.A(new_n13214), .B(new_n13213), .Y(new_n13216));
  nor_5  g10868(.A(new_n13174), .B(new_n13167), .Y(new_n13217));
  xnor_4 g10869(.A(new_n13217), .B(new_n13166), .Y(new_n13218));
  nor_5  g10870(.A(new_n13218), .B(new_n5947), .Y(new_n13219));
  xnor_4 g10871(.A(new_n13218), .B(new_n5945), .Y(new_n13220));
  nor_5  g10872(.A(new_n13172), .B(new_n13169), .Y(new_n13221));
  xnor_4 g10873(.A(new_n13221), .B(new_n13168_1), .Y(new_n13222));
  nor_5  g10874(.A(new_n13222), .B(new_n5953), .Y(new_n13223));
  xnor_4 g10875(.A(new_n13222), .B(new_n5952), .Y(new_n13224));
  xnor_4 g10876(.A(n18578), .B(new_n12371), .Y(new_n13225));
  nor_5  g10877(.A(new_n13225), .B(new_n5956), .Y(new_n13226));
  nor_5  g10878(.A(new_n13226), .B(new_n5959), .Y(new_n13227));
  xnor_4 g10879(.A(new_n13171), .B(new_n13170), .Y(new_n13228));
  not_8  g10880(.A(new_n13226), .Y(new_n13229));
  nor_5  g10881(.A(new_n13229), .B(new_n5897), .Y(new_n13230));
  nor_5  g10882(.A(new_n13230), .B(new_n13227), .Y(new_n13231));
  and_5  g10883(.A(new_n13231), .B(new_n13228), .Y(new_n13232));
  or_5   g10884(.A(new_n13232), .B(new_n13227), .Y(new_n13233));
  and_5  g10885(.A(new_n13233), .B(new_n13224), .Y(new_n13234));
  or_5   g10886(.A(new_n13234), .B(new_n13223), .Y(new_n13235));
  and_5  g10887(.A(new_n13235), .B(new_n13220), .Y(new_n13236));
  nor_5  g10888(.A(new_n13236), .B(new_n13219), .Y(new_n13237));
  nor_5  g10889(.A(new_n13237), .B(new_n13216), .Y(new_n13238));
  nor_5  g10890(.A(new_n13238), .B(new_n13215), .Y(new_n13239));
  and_5  g10891(.A(new_n13239), .B(new_n13212), .Y(new_n13240));
  nor_5  g10892(.A(new_n13240), .B(new_n13210), .Y(new_n13241));
  nor_5  g10893(.A(new_n13241), .B(new_n13208), .Y(new_n13242));
  nor_5  g10894(.A(new_n13242), .B(new_n13207), .Y(new_n13243));
  nor_5  g10895(.A(new_n13243), .B(new_n13205), .Y(new_n13244));
  nor_5  g10896(.A(new_n13244), .B(new_n13204_1), .Y(new_n13245));
  nor_5  g10897(.A(new_n13245), .B(new_n13202), .Y(new_n13246));
  nor_5  g10898(.A(new_n13246), .B(new_n13201), .Y(new_n13247));
  nor_5  g10899(.A(new_n13247), .B(new_n13199_1), .Y(new_n13248));
  nor_5  g10900(.A(new_n13248), .B(new_n13198_1), .Y(new_n13249));
  nor_5  g10901(.A(new_n13249), .B(new_n13196), .Y(new_n13250));
  nor_5  g10902(.A(new_n13250), .B(new_n13195), .Y(new_n13251));
  xnor_4 g10903(.A(new_n13249), .B(new_n13196), .Y(new_n13252));
  not_8  g10904(.A(new_n13252), .Y(new_n13253));
  not_8  g10905(.A(n2743), .Y(new_n13254));
  nor_5  g10906(.A(n3506), .B(new_n13254), .Y(new_n13255));
  and_5  g10907(.A(new_n3580), .B(new_n3536), .Y(new_n13256));
  nor_5  g10908(.A(new_n13256), .B(new_n13255), .Y(new_n13257));
  and_5  g10909(.A(new_n13257), .B(new_n13253), .Y(new_n13258));
  xnor_4 g10910(.A(new_n13257), .B(new_n13253), .Y(new_n13259));
  xnor_4 g10911(.A(new_n13247), .B(new_n13199_1), .Y(new_n13260));
  nor_5  g10912(.A(new_n13260), .B(new_n3582_1), .Y(new_n13261));
  xnor_4 g10913(.A(new_n13260), .B(new_n3582_1), .Y(new_n13262));
  xnor_4 g10914(.A(new_n13245), .B(new_n13202), .Y(new_n13263_1));
  nor_5  g10915(.A(new_n13263_1), .B(new_n3601), .Y(new_n13264));
  xnor_4 g10916(.A(new_n13263_1), .B(new_n3601), .Y(new_n13265));
  xnor_4 g10917(.A(new_n13243), .B(new_n13205), .Y(new_n13266));
  nor_5  g10918(.A(new_n13266), .B(new_n3610), .Y(new_n13267));
  xnor_4 g10919(.A(new_n13266), .B(new_n3610), .Y(new_n13268));
  xnor_4 g10920(.A(new_n13241), .B(new_n13208), .Y(new_n13269));
  not_8  g10921(.A(new_n13269), .Y(new_n13270_1));
  and_5  g10922(.A(new_n13270_1), .B(new_n3613), .Y(new_n13271));
  xnor_4 g10923(.A(new_n13270_1), .B(new_n3613), .Y(new_n13272));
  xnor_4 g10924(.A(new_n13239), .B(new_n13212), .Y(new_n13273_1));
  not_8  g10925(.A(new_n13273_1), .Y(new_n13274));
  and_5  g10926(.A(new_n13274), .B(new_n3617_1), .Y(new_n13275));
  xnor_4 g10927(.A(new_n13274), .B(new_n3617_1), .Y(new_n13276));
  xnor_4 g10928(.A(new_n13237), .B(new_n13216), .Y(new_n13277));
  and_5  g10929(.A(new_n13277), .B(new_n3622), .Y(new_n13278));
  xnor_4 g10930(.A(new_n13277), .B(new_n3622), .Y(new_n13279));
  xor_4  g10931(.A(new_n13235), .B(new_n13220), .Y(new_n13280));
  nor_5  g10932(.A(new_n13280), .B(new_n3627), .Y(new_n13281));
  xnor_4 g10933(.A(new_n13280), .B(new_n3627), .Y(new_n13282));
  xor_4  g10934(.A(new_n13233), .B(new_n13224), .Y(new_n13283));
  nor_5  g10935(.A(new_n13283), .B(new_n3632), .Y(new_n13284));
  xnor_4 g10936(.A(new_n13283), .B(new_n3632), .Y(new_n13285_1));
  xor_4  g10937(.A(new_n13231), .B(new_n13228), .Y(new_n13286));
  nor_5  g10938(.A(new_n13286), .B(new_n3638), .Y(new_n13287));
  xnor_4 g10939(.A(new_n13225), .B(new_n5956), .Y(new_n13288));
  nor_5  g10940(.A(new_n13288), .B(new_n3641), .Y(new_n13289));
  xnor_4 g10941(.A(new_n13286), .B(new_n3639), .Y(new_n13290));
  and_5  g10942(.A(new_n13290), .B(new_n13289), .Y(new_n13291));
  nor_5  g10943(.A(new_n13291), .B(new_n13287), .Y(new_n13292));
  nor_5  g10944(.A(new_n13292), .B(new_n13285_1), .Y(new_n13293));
  nor_5  g10945(.A(new_n13293), .B(new_n13284), .Y(new_n13294));
  nor_5  g10946(.A(new_n13294), .B(new_n13282), .Y(new_n13295));
  nor_5  g10947(.A(new_n13295), .B(new_n13281), .Y(new_n13296));
  nor_5  g10948(.A(new_n13296), .B(new_n13279), .Y(new_n13297));
  nor_5  g10949(.A(new_n13297), .B(new_n13278), .Y(new_n13298));
  nor_5  g10950(.A(new_n13298), .B(new_n13276), .Y(new_n13299));
  nor_5  g10951(.A(new_n13299), .B(new_n13275), .Y(new_n13300));
  nor_5  g10952(.A(new_n13300), .B(new_n13272), .Y(new_n13301));
  nor_5  g10953(.A(new_n13301), .B(new_n13271), .Y(new_n13302));
  nor_5  g10954(.A(new_n13302), .B(new_n13268), .Y(new_n13303));
  nor_5  g10955(.A(new_n13303), .B(new_n13267), .Y(new_n13304));
  nor_5  g10956(.A(new_n13304), .B(new_n13265), .Y(new_n13305));
  nor_5  g10957(.A(new_n13305), .B(new_n13264), .Y(new_n13306));
  nor_5  g10958(.A(new_n13306), .B(new_n13262), .Y(new_n13307));
  nor_5  g10959(.A(new_n13307), .B(new_n13261), .Y(new_n13308));
  nor_5  g10960(.A(new_n13308), .B(new_n13259), .Y(new_n13309));
  nor_5  g10961(.A(new_n13309), .B(new_n13258), .Y(new_n13310));
  xor_4  g10962(.A(new_n13310), .B(new_n13251), .Y(n2561));
  xor_4  g10963(.A(new_n8423), .B(new_n8421), .Y(n2573));
  xnor_4 g10964(.A(n18558), .B(n10411), .Y(new_n13313));
  nor_5  g10965(.A(new_n10003), .B(n7149), .Y(new_n13314));
  nor_5  g10966(.A(n16971), .B(new_n2695), .Y(new_n13315));
  nor_5  g10967(.A(n14148), .B(new_n2756), .Y(new_n13316));
  nor_5  g10968(.A(new_n2701), .B(n11503), .Y(new_n13317));
  nor_5  g10969(.A(new_n2828), .B(n1152), .Y(new_n13318));
  not_8  g10970(.A(new_n13318), .Y(new_n13319_1));
  nor_5  g10971(.A(new_n13319_1), .B(new_n13317), .Y(new_n13320));
  nor_5  g10972(.A(new_n13320), .B(new_n13316), .Y(new_n13321));
  nor_5  g10973(.A(new_n13321), .B(new_n13315), .Y(new_n13322));
  or_5   g10974(.A(new_n13322), .B(new_n13314), .Y(new_n13323));
  xor_4  g10975(.A(new_n13323), .B(new_n13313), .Y(new_n13324));
  nor_5  g10976(.A(n7963), .B(new_n9834), .Y(new_n13325));
  nor_5  g10977(.A(new_n9835), .B(n6590), .Y(new_n13326));
  nor_5  g10978(.A(new_n9830), .B(n10017), .Y(new_n13327));
  or_5   g10979(.A(n20349), .B(new_n7941), .Y(new_n13328));
  nor_5  g10980(.A(new_n9828), .B(n3618), .Y(new_n13329));
  and_5  g10981(.A(new_n13329), .B(new_n13328), .Y(new_n13330));
  nor_5  g10982(.A(new_n13330), .B(new_n13327), .Y(new_n13331));
  nor_5  g10983(.A(new_n13331), .B(new_n13326), .Y(new_n13332));
  nor_5  g10984(.A(new_n13332), .B(new_n13325), .Y(new_n13333_1));
  xnor_4 g10985(.A(new_n13333_1), .B(new_n9874), .Y(new_n13334));
  not_8  g10986(.A(new_n13334), .Y(new_n13335));
  xnor_4 g10987(.A(new_n13335), .B(new_n13324), .Y(new_n13336));
  xnor_4 g10988(.A(n16971), .B(n7149), .Y(new_n13337));
  xnor_4 g10989(.A(new_n13337), .B(new_n13321), .Y(new_n13338_1));
  xnor_4 g10990(.A(new_n13331), .B(new_n9879), .Y(new_n13339));
  nor_5  g10991(.A(new_n13339), .B(new_n13338_1), .Y(new_n13340));
  not_8  g10992(.A(new_n13339), .Y(new_n13341));
  xnor_4 g10993(.A(new_n13341), .B(new_n13338_1), .Y(new_n13342));
  xnor_4 g10994(.A(n18151), .B(n1152), .Y(new_n13343));
  or_5   g10995(.A(new_n13343), .B(new_n9885), .Y(new_n13344));
  xnor_4 g10996(.A(n14148), .B(n11503), .Y(new_n13345));
  xnor_4 g10997(.A(new_n13345), .B(new_n13319_1), .Y(new_n13346));
  and_5  g10998(.A(new_n13346), .B(new_n13344), .Y(new_n13347));
  nor_5  g10999(.A(new_n13343), .B(new_n9885), .Y(new_n13348));
  xnor_4 g11000(.A(new_n13346), .B(new_n13348), .Y(new_n13349));
  xor_4  g11001(.A(new_n13329), .B(new_n9882), .Y(new_n13350));
  and_5  g11002(.A(new_n13350), .B(new_n13349), .Y(new_n13351));
  nor_5  g11003(.A(new_n13351), .B(new_n13347), .Y(new_n13352));
  and_5  g11004(.A(new_n13352), .B(new_n13342), .Y(new_n13353));
  nor_5  g11005(.A(new_n13353), .B(new_n13340), .Y(new_n13354));
  xnor_4 g11006(.A(new_n13354), .B(new_n13336), .Y(new_n13355));
  not_8  g11007(.A(new_n13355), .Y(new_n13356));
  xnor_4 g11008(.A(n19515), .B(n17035), .Y(new_n13357));
  not_8  g11009(.A(n22588), .Y(new_n13358));
  nor_5  g11010(.A(new_n13358), .B(n14684), .Y(new_n13359));
  nor_5  g11011(.A(n22588), .B(new_n8445), .Y(new_n13360));
  and_5  g11012(.A(n12209), .B(new_n4180), .Y(new_n13361));
  nor_5  g11013(.A(n12209), .B(new_n4180), .Y(new_n13362));
  nor_5  g11014(.A(n24732), .B(new_n13145), .Y(new_n13363));
  not_8  g11015(.A(new_n13363), .Y(new_n13364));
  nor_5  g11016(.A(new_n13364), .B(new_n13362), .Y(new_n13365));
  nor_5  g11017(.A(new_n13365), .B(new_n13361), .Y(new_n13366));
  nor_5  g11018(.A(new_n13366), .B(new_n13360), .Y(new_n13367_1));
  nor_5  g11019(.A(new_n13367_1), .B(new_n13359), .Y(new_n13368));
  xnor_4 g11020(.A(new_n13368), .B(new_n13357), .Y(new_n13369));
  not_8  g11021(.A(new_n13369), .Y(new_n13370));
  xnor_4 g11022(.A(new_n13370), .B(new_n13356), .Y(new_n13371));
  xnor_4 g11023(.A(new_n13352), .B(new_n13342), .Y(new_n13372));
  xnor_4 g11024(.A(n22588), .B(n14684), .Y(new_n13373));
  xnor_4 g11025(.A(new_n13373), .B(new_n13366), .Y(new_n13374));
  and_5  g11026(.A(new_n13374), .B(new_n13372), .Y(new_n13375));
  xnor_4 g11027(.A(n24732), .B(n12892), .Y(new_n13376));
  xnor_4 g11028(.A(new_n13343), .B(new_n9885), .Y(new_n13377));
  nor_5  g11029(.A(new_n13377), .B(new_n13376), .Y(new_n13378));
  xnor_4 g11030(.A(n12209), .B(n6631), .Y(new_n13379));
  xnor_4 g11031(.A(new_n13379), .B(new_n13364), .Y(new_n13380));
  not_8  g11032(.A(new_n13380), .Y(new_n13381));
  nor_5  g11033(.A(new_n13381), .B(new_n13378), .Y(new_n13382));
  xnor_4 g11034(.A(new_n13380), .B(new_n13378), .Y(new_n13383));
  xnor_4 g11035(.A(new_n13329), .B(new_n9882), .Y(new_n13384));
  xnor_4 g11036(.A(new_n13384), .B(new_n13349), .Y(new_n13385));
  and_5  g11037(.A(new_n13385), .B(new_n13383), .Y(new_n13386));
  nor_5  g11038(.A(new_n13386), .B(new_n13382), .Y(new_n13387));
  xnor_4 g11039(.A(new_n13374), .B(new_n13372), .Y(new_n13388));
  nor_5  g11040(.A(new_n13388), .B(new_n13387), .Y(new_n13389));
  nor_5  g11041(.A(new_n13389), .B(new_n13375), .Y(new_n13390));
  xnor_4 g11042(.A(new_n13390), .B(new_n13371), .Y(n2578));
  not_8  g11043(.A(new_n11607_1), .Y(new_n13392));
  nor_5  g11044(.A(new_n13392), .B(new_n7835), .Y(new_n13393));
  not_8  g11045(.A(new_n7835), .Y(new_n13394));
  xnor_4 g11046(.A(new_n13392), .B(new_n13394), .Y(new_n13395));
  nor_5  g11047(.A(new_n13394), .B(new_n7771), .Y(new_n13396));
  and_5  g11048(.A(new_n7916), .B(new_n7836), .Y(new_n13397));
  or_5   g11049(.A(new_n13397), .B(new_n13396), .Y(new_n13398));
  and_5  g11050(.A(new_n13398), .B(new_n13395), .Y(new_n13399));
  nor_5  g11051(.A(new_n13399), .B(new_n13393), .Y(n2582));
  xor_4  g11052(.A(new_n4306_1), .B(new_n4295), .Y(n2602));
  nor_5  g11053(.A(n22201), .B(n2420), .Y(new_n13402));
  not_8  g11054(.A(new_n13402), .Y(new_n13403));
  nor_5  g11055(.A(new_n13403), .B(n24485), .Y(new_n13404));
  not_8  g11056(.A(new_n13404), .Y(new_n13405));
  nor_5  g11057(.A(new_n13405), .B(n21078), .Y(new_n13406));
  not_8  g11058(.A(new_n13406), .Y(new_n13407_1));
  nor_5  g11059(.A(new_n13407_1), .B(n12546), .Y(new_n13408));
  xnor_4 g11060(.A(new_n13408), .B(n8324), .Y(new_n13409_1));
  xnor_4 g11061(.A(new_n13409_1), .B(new_n3963), .Y(new_n13410));
  xnor_4 g11062(.A(new_n13406), .B(n12546), .Y(new_n13411));
  nor_5  g11063(.A(new_n13411), .B(new_n3965), .Y(new_n13412));
  xnor_4 g11064(.A(new_n13404), .B(n21078), .Y(new_n13413));
  nor_5  g11065(.A(new_n13413), .B(new_n3970), .Y(new_n13414));
  xnor_4 g11066(.A(new_n13413), .B(new_n3968), .Y(new_n13415));
  xnor_4 g11067(.A(new_n13402), .B(n24485), .Y(new_n13416));
  and_5  g11068(.A(new_n13416), .B(new_n3976), .Y(new_n13417));
  xnor_4 g11069(.A(new_n13416), .B(new_n3974), .Y(new_n13418));
  xnor_4 g11070(.A(n22201), .B(new_n8112), .Y(new_n13419_1));
  nor_5  g11071(.A(new_n13419_1), .B(new_n3984_1), .Y(new_n13420));
  or_5   g11072(.A(new_n2551), .B(new_n8110), .Y(new_n13421));
  xnor_4 g11073(.A(new_n13419_1), .B(new_n3980), .Y(new_n13422));
  and_5  g11074(.A(new_n13422), .B(new_n13421), .Y(new_n13423));
  nor_5  g11075(.A(new_n13423), .B(new_n13420), .Y(new_n13424_1));
  and_5  g11076(.A(new_n13424_1), .B(new_n13418), .Y(new_n13425));
  nor_5  g11077(.A(new_n13425), .B(new_n13417), .Y(new_n13426));
  and_5  g11078(.A(new_n13426), .B(new_n13415), .Y(new_n13427));
  nor_5  g11079(.A(new_n13427), .B(new_n13414), .Y(new_n13428));
  xnor_4 g11080(.A(new_n13411), .B(new_n3965), .Y(new_n13429));
  nor_5  g11081(.A(new_n13429), .B(new_n13428), .Y(new_n13430));
  nor_5  g11082(.A(new_n13430), .B(new_n13412), .Y(new_n13431));
  xnor_4 g11083(.A(new_n13431), .B(new_n13410), .Y(new_n13432));
  xnor_4 g11084(.A(new_n8093), .B(n7678), .Y(new_n13433));
  nor_5  g11085(.A(new_n8095_1), .B(n3785), .Y(new_n13434));
  xnor_4 g11086(.A(new_n8095_1), .B(new_n4377), .Y(new_n13435));
  nor_5  g11087(.A(new_n8099), .B(n20250), .Y(new_n13436));
  xnor_4 g11088(.A(new_n8099), .B(new_n4382), .Y(new_n13437));
  nor_5  g11089(.A(new_n8103_1), .B(new_n4384), .Y(new_n13438));
  or_5   g11090(.A(new_n8104), .B(n5822), .Y(new_n13439));
  nor_5  g11091(.A(new_n8108), .B(n26443), .Y(new_n13440));
  or_5   g11092(.A(new_n2545), .B(new_n4394), .Y(new_n13441));
  xnor_4 g11093(.A(new_n8108), .B(new_n6644), .Y(new_n13442));
  and_5  g11094(.A(new_n13442), .B(new_n13441), .Y(new_n13443));
  nor_5  g11095(.A(new_n13443), .B(new_n13440), .Y(new_n13444));
  and_5  g11096(.A(new_n13444), .B(new_n13439), .Y(new_n13445));
  nor_5  g11097(.A(new_n13445), .B(new_n13438), .Y(new_n13446));
  and_5  g11098(.A(new_n13446), .B(new_n13437), .Y(new_n13447));
  or_5   g11099(.A(new_n13447), .B(new_n13436), .Y(new_n13448));
  and_5  g11100(.A(new_n13448), .B(new_n13435), .Y(new_n13449));
  nor_5  g11101(.A(new_n13449), .B(new_n13434), .Y(new_n13450));
  xor_4  g11102(.A(new_n13450), .B(new_n13433), .Y(new_n13451));
  xnor_4 g11103(.A(new_n13451), .B(new_n13432), .Y(new_n13452));
  xor_4  g11104(.A(new_n13448), .B(new_n13435), .Y(new_n13453_1));
  xnor_4 g11105(.A(new_n13429), .B(new_n13428), .Y(new_n13454));
  not_8  g11106(.A(new_n13454), .Y(new_n13455));
  and_5  g11107(.A(new_n13455), .B(new_n13453_1), .Y(new_n13456_1));
  xnor_4 g11108(.A(new_n13455), .B(new_n13453_1), .Y(new_n13457_1));
  xnor_4 g11109(.A(new_n13426), .B(new_n13415), .Y(new_n13458));
  xnor_4 g11110(.A(new_n13446), .B(new_n13437), .Y(new_n13459));
  nor_5  g11111(.A(new_n13459), .B(new_n13458), .Y(new_n13460_1));
  xor_4  g11112(.A(new_n13459), .B(new_n13458), .Y(new_n13461));
  xnor_4 g11113(.A(new_n13424_1), .B(new_n13418), .Y(new_n13462));
  xnor_4 g11114(.A(new_n8104), .B(new_n4384), .Y(new_n13463));
  xnor_4 g11115(.A(new_n13463), .B(new_n13444), .Y(new_n13464));
  nor_5  g11116(.A(new_n13464), .B(new_n13462), .Y(new_n13465));
  xor_4  g11117(.A(new_n13422), .B(new_n13421), .Y(new_n13466));
  xor_4  g11118(.A(new_n13442), .B(new_n13441), .Y(new_n13467));
  and_5  g11119(.A(new_n13467), .B(new_n13466), .Y(new_n13468));
  xnor_4 g11120(.A(new_n2545), .B(new_n4394), .Y(new_n13469));
  xnor_4 g11121(.A(new_n2551), .B(n22201), .Y(new_n13470));
  not_8  g11122(.A(new_n13470), .Y(new_n13471));
  nor_5  g11123(.A(new_n13471), .B(new_n13469), .Y(new_n13472));
  xnor_4 g11124(.A(new_n13467), .B(new_n13466), .Y(new_n13473));
  nor_5  g11125(.A(new_n13473), .B(new_n13472), .Y(new_n13474));
  nor_5  g11126(.A(new_n13474), .B(new_n13468), .Y(new_n13475));
  xor_4  g11127(.A(new_n13464), .B(new_n13462), .Y(new_n13476));
  and_5  g11128(.A(new_n13476), .B(new_n13475), .Y(new_n13477_1));
  nor_5  g11129(.A(new_n13477_1), .B(new_n13465), .Y(new_n13478));
  and_5  g11130(.A(new_n13478), .B(new_n13461), .Y(new_n13479));
  nor_5  g11131(.A(new_n13479), .B(new_n13460_1), .Y(new_n13480));
  nor_5  g11132(.A(new_n13480), .B(new_n13457_1), .Y(new_n13481));
  nor_5  g11133(.A(new_n13481), .B(new_n13456_1), .Y(new_n13482));
  xnor_4 g11134(.A(new_n13482), .B(new_n13452), .Y(n2619));
  nor_5  g11135(.A(new_n5917), .B(n12900), .Y(new_n13484_1));
  xnor_4 g11136(.A(new_n5917), .B(n12900), .Y(new_n13485));
  nor_5  g11137(.A(new_n5923), .B(n20411), .Y(new_n13486_1));
  xnor_4 g11138(.A(new_n5923), .B(n20411), .Y(new_n13487_1));
  nor_5  g11139(.A(new_n5928), .B(n17069), .Y(new_n13488));
  xnor_4 g11140(.A(new_n5928), .B(n17069), .Y(new_n13489));
  nor_5  g11141(.A(new_n5933), .B(n15918), .Y(new_n13490_1));
  nor_5  g11142(.A(new_n5938), .B(n17784), .Y(new_n13491));
  xnor_4 g11143(.A(new_n5938), .B(n17784), .Y(new_n13492));
  and_5  g11144(.A(new_n5943_1), .B(n14323), .Y(new_n13493));
  nor_5  g11145(.A(new_n12850), .B(new_n12840), .Y(new_n13494_1));
  nor_5  g11146(.A(new_n13494_1), .B(new_n13493), .Y(new_n13495));
  not_8  g11147(.A(new_n13495), .Y(new_n13496));
  nor_5  g11148(.A(new_n13496), .B(new_n13492), .Y(new_n13497));
  nor_5  g11149(.A(new_n13497), .B(new_n13491), .Y(new_n13498));
  xnor_4 g11150(.A(new_n5933), .B(n15918), .Y(new_n13499));
  nor_5  g11151(.A(new_n13499), .B(new_n13498), .Y(new_n13500_1));
  nor_5  g11152(.A(new_n13500_1), .B(new_n13490_1), .Y(new_n13501_1));
  nor_5  g11153(.A(new_n13501_1), .B(new_n13489), .Y(new_n13502));
  nor_5  g11154(.A(new_n13502), .B(new_n13488), .Y(new_n13503));
  nor_5  g11155(.A(new_n13503), .B(new_n13487_1), .Y(new_n13504));
  nor_5  g11156(.A(new_n13504), .B(new_n13486_1), .Y(new_n13505));
  nor_5  g11157(.A(new_n13505), .B(new_n13485), .Y(new_n13506_1));
  nor_5  g11158(.A(new_n13506_1), .B(new_n13484_1), .Y(new_n13507));
  not_8  g11159(.A(new_n5871), .Y(new_n13508));
  xnor_4 g11160(.A(new_n13508), .B(n10650), .Y(new_n13509));
  xnor_4 g11161(.A(new_n13509), .B(new_n13507), .Y(new_n13510));
  not_8  g11162(.A(new_n13510), .Y(new_n13511));
  nor_5  g11163(.A(new_n13511), .B(n6456), .Y(new_n13512));
  xnor_4 g11164(.A(new_n13511), .B(new_n5872), .Y(new_n13513));
  xnor_4 g11165(.A(new_n13505), .B(new_n13485), .Y(new_n13514));
  nor_5  g11166(.A(new_n13514), .B(n4085), .Y(new_n13515));
  not_8  g11167(.A(new_n13514), .Y(new_n13516));
  xnor_4 g11168(.A(new_n13516), .B(n4085), .Y(new_n13517));
  xnor_4 g11169(.A(new_n13503), .B(new_n13487_1), .Y(new_n13518));
  nor_5  g11170(.A(new_n13518), .B(n26725), .Y(new_n13519));
  not_8  g11171(.A(new_n13518), .Y(new_n13520));
  xnor_4 g11172(.A(new_n13520), .B(n26725), .Y(new_n13521));
  xnor_4 g11173(.A(new_n13501_1), .B(new_n13489), .Y(new_n13522));
  nor_5  g11174(.A(new_n13522), .B(n11980), .Y(new_n13523));
  not_8  g11175(.A(new_n13522), .Y(new_n13524));
  xnor_4 g11176(.A(new_n13524), .B(n11980), .Y(new_n13525));
  xnor_4 g11177(.A(new_n13499), .B(new_n13498), .Y(new_n13526));
  nor_5  g11178(.A(new_n13526), .B(n3253), .Y(new_n13527));
  xnor_4 g11179(.A(new_n13526), .B(new_n5883), .Y(new_n13528));
  xnor_4 g11180(.A(new_n13495), .B(new_n13492), .Y(new_n13529));
  nor_5  g11181(.A(new_n13529), .B(new_n5886), .Y(new_n13530));
  not_8  g11182(.A(new_n13529), .Y(new_n13531));
  xnor_4 g11183(.A(new_n13531), .B(new_n5886), .Y(new_n13532));
  nor_5  g11184(.A(new_n12851), .B(new_n5889), .Y(new_n13533));
  and_5  g11185(.A(new_n12863), .B(new_n12852), .Y(new_n13534));
  or_5   g11186(.A(new_n13534), .B(new_n13533), .Y(new_n13535));
  and_5  g11187(.A(new_n13535), .B(new_n13532), .Y(new_n13536));
  nor_5  g11188(.A(new_n13536), .B(new_n13530), .Y(new_n13537));
  and_5  g11189(.A(new_n13537), .B(new_n13528), .Y(new_n13538));
  or_5   g11190(.A(new_n13538), .B(new_n13527), .Y(new_n13539));
  and_5  g11191(.A(new_n13539), .B(new_n13525), .Y(new_n13540));
  or_5   g11192(.A(new_n13540), .B(new_n13523), .Y(new_n13541));
  and_5  g11193(.A(new_n13541), .B(new_n13521), .Y(new_n13542));
  or_5   g11194(.A(new_n13542), .B(new_n13519), .Y(new_n13543));
  and_5  g11195(.A(new_n13543), .B(new_n13517), .Y(new_n13544));
  or_5   g11196(.A(new_n13544), .B(new_n13515), .Y(new_n13545));
  and_5  g11197(.A(new_n13545), .B(new_n13513), .Y(new_n13546));
  nor_5  g11198(.A(new_n13546), .B(new_n13512), .Y(new_n13547));
  or_5   g11199(.A(new_n5871), .B(n10650), .Y(new_n13548_1));
  and_5  g11200(.A(new_n13548_1), .B(new_n13507), .Y(new_n13549_1));
  and_5  g11201(.A(new_n5870), .B(new_n4798), .Y(new_n13550));
  and_5  g11202(.A(new_n5871), .B(n10650), .Y(new_n13551_1));
  or_5   g11203(.A(new_n13551_1), .B(new_n13550), .Y(new_n13552));
  nor_5  g11204(.A(new_n13552), .B(new_n13549_1), .Y(new_n13553));
  and_5  g11205(.A(new_n13553), .B(new_n13547), .Y(new_n13554));
  nor_5  g11206(.A(new_n13554), .B(new_n12592), .Y(new_n13555));
  xnor_4 g11207(.A(new_n13554), .B(new_n12592), .Y(new_n13556));
  xnor_4 g11208(.A(new_n13553), .B(new_n13547), .Y(new_n13557));
  and_5  g11209(.A(new_n13557), .B(new_n12596), .Y(new_n13558));
  xnor_4 g11210(.A(new_n13557), .B(new_n12596), .Y(new_n13559));
  xor_4  g11211(.A(new_n13545), .B(new_n13513), .Y(new_n13560));
  and_5  g11212(.A(new_n13560), .B(new_n12601), .Y(new_n13561));
  xnor_4 g11213(.A(new_n13560), .B(new_n12601), .Y(new_n13562));
  xor_4  g11214(.A(new_n13543), .B(new_n13517), .Y(new_n13563));
  and_5  g11215(.A(new_n13563), .B(new_n12606), .Y(new_n13564));
  xnor_4 g11216(.A(new_n13563), .B(new_n12606), .Y(new_n13565));
  xor_4  g11217(.A(new_n13541), .B(new_n13521), .Y(new_n13566));
  and_5  g11218(.A(new_n13566), .B(new_n12611), .Y(new_n13567));
  xnor_4 g11219(.A(new_n13566), .B(new_n12611), .Y(new_n13568));
  xor_4  g11220(.A(new_n13539), .B(new_n13525), .Y(new_n13569));
  and_5  g11221(.A(new_n13569), .B(new_n12616), .Y(new_n13570));
  xnor_4 g11222(.A(new_n13569), .B(new_n12616), .Y(new_n13571));
  xnor_4 g11223(.A(new_n13537), .B(new_n13528), .Y(new_n13572));
  nor_5  g11224(.A(new_n13572), .B(new_n12622), .Y(new_n13573));
  xnor_4 g11225(.A(new_n13572), .B(new_n12622), .Y(new_n13574));
  xor_4  g11226(.A(new_n13535), .B(new_n13532), .Y(new_n13575));
  nor_5  g11227(.A(new_n13575), .B(new_n12626_1), .Y(new_n13576));
  xnor_4 g11228(.A(new_n13575), .B(new_n12626_1), .Y(new_n13577));
  nor_5  g11229(.A(new_n12864_1), .B(new_n12630), .Y(new_n13578));
  nor_5  g11230(.A(new_n12878), .B(new_n12865_1), .Y(new_n13579));
  nor_5  g11231(.A(new_n13579), .B(new_n13578), .Y(new_n13580));
  nor_5  g11232(.A(new_n13580), .B(new_n13577), .Y(new_n13581));
  nor_5  g11233(.A(new_n13581), .B(new_n13576), .Y(new_n13582));
  nor_5  g11234(.A(new_n13582), .B(new_n13574), .Y(new_n13583));
  nor_5  g11235(.A(new_n13583), .B(new_n13573), .Y(new_n13584));
  nor_5  g11236(.A(new_n13584), .B(new_n13571), .Y(new_n13585));
  nor_5  g11237(.A(new_n13585), .B(new_n13570), .Y(new_n13586));
  nor_5  g11238(.A(new_n13586), .B(new_n13568), .Y(new_n13587));
  nor_5  g11239(.A(new_n13587), .B(new_n13567), .Y(new_n13588));
  nor_5  g11240(.A(new_n13588), .B(new_n13565), .Y(new_n13589));
  nor_5  g11241(.A(new_n13589), .B(new_n13564), .Y(new_n13590));
  nor_5  g11242(.A(new_n13590), .B(new_n13562), .Y(new_n13591));
  nor_5  g11243(.A(new_n13591), .B(new_n13561), .Y(new_n13592));
  nor_5  g11244(.A(new_n13592), .B(new_n13559), .Y(new_n13593));
  nor_5  g11245(.A(new_n13593), .B(new_n13558), .Y(new_n13594));
  nor_5  g11246(.A(new_n13594), .B(new_n13556), .Y(new_n13595));
  nor_5  g11247(.A(new_n13595), .B(new_n13555), .Y(n2661));
  xnor_4 g11248(.A(new_n11070), .B(new_n11068), .Y(n2693));
  xnor_4 g11249(.A(new_n13324), .B(new_n7288), .Y(new_n13598));
  nor_5  g11250(.A(new_n13338_1), .B(new_n7295), .Y(new_n13599));
  xnor_4 g11251(.A(new_n13338_1), .B(new_n7295), .Y(new_n13600));
  nor_5  g11252(.A(new_n13346), .B(new_n7298_1), .Y(new_n13601));
  nor_5  g11253(.A(new_n13343), .B(new_n7300), .Y(new_n13602_1));
  xnor_4 g11254(.A(new_n13346), .B(new_n7302), .Y(new_n13603));
  and_5  g11255(.A(new_n13603), .B(new_n13602_1), .Y(new_n13604));
  nor_5  g11256(.A(new_n13604), .B(new_n13601), .Y(new_n13605));
  nor_5  g11257(.A(new_n13605), .B(new_n13600), .Y(new_n13606));
  nor_5  g11258(.A(new_n13606), .B(new_n13599), .Y(new_n13607));
  xnor_4 g11259(.A(new_n13607), .B(new_n13598), .Y(new_n13608));
  not_8  g11260(.A(new_n13608), .Y(new_n13609));
  xnor_4 g11261(.A(n8309), .B(n4665), .Y(new_n13610));
  nor_5  g11262(.A(new_n8759), .B(n19005), .Y(new_n13611));
  nor_5  g11263(.A(n19144), .B(new_n2866), .Y(new_n13612));
  nor_5  g11264(.A(new_n10007), .B(n4326), .Y(new_n13613));
  or_5   g11265(.A(n12593), .B(new_n2869), .Y(new_n13614));
  nor_5  g11266(.A(new_n8763), .B(n5438), .Y(new_n13615));
  and_5  g11267(.A(new_n13615), .B(new_n13614), .Y(new_n13616));
  nor_5  g11268(.A(new_n13616), .B(new_n13613), .Y(new_n13617));
  nor_5  g11269(.A(new_n13617), .B(new_n13612), .Y(new_n13618));
  or_5   g11270(.A(new_n13618), .B(new_n13611), .Y(new_n13619));
  xor_4  g11271(.A(new_n13619), .B(new_n13610), .Y(new_n13620));
  xnor_4 g11272(.A(new_n13620), .B(new_n13609), .Y(new_n13621));
  xnor_4 g11273(.A(new_n13605), .B(new_n13600), .Y(new_n13622));
  xnor_4 g11274(.A(n19144), .B(n19005), .Y(new_n13623));
  xnor_4 g11275(.A(new_n13623), .B(new_n13617), .Y(new_n13624));
  and_5  g11276(.A(new_n13624), .B(new_n13622), .Y(new_n13625));
  xnor_4 g11277(.A(new_n13624), .B(new_n13622), .Y(new_n13626_1));
  xnor_4 g11278(.A(n13714), .B(n5438), .Y(new_n13627));
  xnor_4 g11279(.A(new_n13343), .B(new_n7399), .Y(new_n13628));
  not_8  g11280(.A(new_n13628), .Y(new_n13629));
  nor_5  g11281(.A(new_n13629), .B(new_n13627), .Y(new_n13630));
  xnor_4 g11282(.A(n12593), .B(n4326), .Y(new_n13631));
  xnor_4 g11283(.A(new_n13631), .B(new_n13615), .Y(new_n13632));
  nor_5  g11284(.A(new_n13632), .B(new_n13630), .Y(new_n13633));
  xnor_4 g11285(.A(new_n13603), .B(new_n13602_1), .Y(new_n13634));
  not_8  g11286(.A(new_n13634), .Y(new_n13635));
  xnor_4 g11287(.A(new_n13632), .B(new_n13630), .Y(new_n13636));
  nor_5  g11288(.A(new_n13636), .B(new_n13635), .Y(new_n13637));
  nor_5  g11289(.A(new_n13637), .B(new_n13633), .Y(new_n13638));
  nor_5  g11290(.A(new_n13638), .B(new_n13626_1), .Y(new_n13639));
  nor_5  g11291(.A(new_n13639), .B(new_n13625), .Y(new_n13640));
  xnor_4 g11292(.A(new_n13640), .B(new_n13621), .Y(n2703));
  xnor_4 g11293(.A(new_n12720), .B(new_n12711), .Y(n2706));
  nor_5  g11294(.A(n3320), .B(new_n6152), .Y(new_n13643));
  xnor_4 g11295(.A(n3320), .B(n1831), .Y(new_n13644));
  not_8  g11296(.A(n13137), .Y(new_n13645));
  nor_5  g11297(.A(new_n13645), .B(n1288), .Y(new_n13646));
  xnor_4 g11298(.A(n13137), .B(n1288), .Y(new_n13647));
  not_8  g11299(.A(n18452), .Y(new_n13648));
  nor_5  g11300(.A(new_n13648), .B(n1752), .Y(new_n13649));
  xnor_4 g11301(.A(n18452), .B(n1752), .Y(new_n13650));
  not_8  g11302(.A(n21317), .Y(new_n13651));
  nor_5  g11303(.A(new_n13651), .B(n13110), .Y(new_n13652));
  xnor_4 g11304(.A(n21317), .B(n13110), .Y(new_n13653));
  nor_5  g11305(.A(n25694), .B(new_n6164), .Y(new_n13654));
  xnor_4 g11306(.A(n25694), .B(n12398), .Y(new_n13655));
  nor_5  g11307(.A(new_n6167), .B(n15424), .Y(new_n13656));
  xnor_4 g11308(.A(n19789), .B(n15424), .Y(new_n13657));
  not_8  g11309(.A(n1949), .Y(new_n13658));
  nor_5  g11310(.A(n20169), .B(new_n13658), .Y(new_n13659));
  and_5  g11311(.A(new_n12025), .B(new_n12016), .Y(new_n13660));
  nor_5  g11312(.A(new_n13660), .B(new_n13659), .Y(new_n13661));
  and_5  g11313(.A(new_n13661), .B(new_n13657), .Y(new_n13662));
  or_5   g11314(.A(new_n13662), .B(new_n13656), .Y(new_n13663));
  and_5  g11315(.A(new_n13663), .B(new_n13655), .Y(new_n13664));
  or_5   g11316(.A(new_n13664), .B(new_n13654), .Y(new_n13665));
  and_5  g11317(.A(new_n13665), .B(new_n13653), .Y(new_n13666));
  or_5   g11318(.A(new_n13666), .B(new_n13652), .Y(new_n13667));
  and_5  g11319(.A(new_n13667), .B(new_n13650), .Y(new_n13668_1));
  or_5   g11320(.A(new_n13668_1), .B(new_n13649), .Y(new_n13669));
  and_5  g11321(.A(new_n13669), .B(new_n13647), .Y(new_n13670));
  or_5   g11322(.A(new_n13670), .B(new_n13646), .Y(new_n13671));
  and_5  g11323(.A(new_n13671), .B(new_n13644), .Y(new_n13672));
  nor_5  g11324(.A(new_n13672), .B(new_n13643), .Y(new_n13673));
  not_8  g11325(.A(new_n13673), .Y(new_n13674));
  not_8  g11326(.A(n1483), .Y(new_n13675));
  nor_5  g11327(.A(n19539), .B(new_n13675), .Y(new_n13676));
  and_5  g11328(.A(new_n11168), .B(new_n11154), .Y(new_n13677_1));
  nor_5  g11329(.A(new_n13677_1), .B(new_n13676), .Y(new_n13678));
  not_8  g11330(.A(new_n6470_1), .Y(new_n13679));
  nor_5  g11331(.A(new_n13679), .B(n16818), .Y(new_n13680));
  not_8  g11332(.A(new_n13680), .Y(new_n13681));
  nor_5  g11333(.A(new_n13681), .B(n3541), .Y(new_n13682));
  xnor_4 g11334(.A(new_n13682), .B(n2184), .Y(new_n13683_1));
  nor_5  g11335(.A(new_n13683_1), .B(n6204), .Y(new_n13684));
  not_8  g11336(.A(new_n13683_1), .Y(new_n13685));
  xnor_4 g11337(.A(new_n13685), .B(n6204), .Y(new_n13686));
  xnor_4 g11338(.A(new_n13680), .B(n3541), .Y(new_n13687));
  not_8  g11339(.A(new_n13687), .Y(new_n13688));
  nor_5  g11340(.A(new_n13688), .B(new_n12116), .Y(new_n13689));
  nor_5  g11341(.A(new_n13687), .B(n3349), .Y(new_n13690));
  nor_5  g11342(.A(new_n6472), .B(new_n12119), .Y(new_n13691));
  or_5   g11343(.A(new_n6471), .B(n1742), .Y(new_n13692));
  and_5  g11344(.A(new_n6506_1), .B(new_n13692), .Y(new_n13693));
  nor_5  g11345(.A(new_n13693), .B(new_n13691), .Y(new_n13694));
  nor_5  g11346(.A(new_n13694), .B(new_n13690), .Y(new_n13695));
  nor_5  g11347(.A(new_n13695), .B(new_n13689), .Y(new_n13696));
  and_5  g11348(.A(new_n13696), .B(new_n13686), .Y(new_n13697));
  nor_5  g11349(.A(new_n13697), .B(new_n13684), .Y(new_n13698));
  not_8  g11350(.A(new_n13682), .Y(new_n13699));
  nor_5  g11351(.A(new_n13699), .B(n2184), .Y(new_n13700));
  xnor_4 g11352(.A(new_n13700), .B(n10018), .Y(new_n13701));
  not_8  g11353(.A(new_n13701), .Y(new_n13702));
  xnor_4 g11354(.A(new_n13702), .B(new_n12110), .Y(new_n13703));
  xnor_4 g11355(.A(new_n13703), .B(new_n13698), .Y(new_n13704));
  nor_5  g11356(.A(new_n13704), .B(new_n11169), .Y(new_n13705));
  xnor_4 g11357(.A(new_n13704), .B(new_n11169), .Y(new_n13706));
  xnor_4 g11358(.A(new_n13696), .B(new_n13686), .Y(new_n13707));
  nor_5  g11359(.A(new_n13707), .B(new_n11228), .Y(new_n13708_1));
  xnor_4 g11360(.A(new_n13707), .B(new_n11228), .Y(new_n13709));
  not_8  g11361(.A(new_n13709), .Y(new_n13710_1));
  xnor_4 g11362(.A(new_n13688), .B(n3349), .Y(new_n13711));
  xnor_4 g11363(.A(new_n13711), .B(new_n13694), .Y(new_n13712));
  and_5  g11364(.A(new_n13712), .B(new_n11232), .Y(new_n13713));
  xnor_4 g11365(.A(new_n13712), .B(new_n11232), .Y(new_n13714_1));
  and_5  g11366(.A(new_n6508), .B(new_n6461), .Y(new_n13715));
  nor_5  g11367(.A(new_n6550), .B(new_n6509), .Y(new_n13716));
  nor_5  g11368(.A(new_n13716), .B(new_n13715), .Y(new_n13717));
  nor_5  g11369(.A(new_n13717), .B(new_n13714_1), .Y(new_n13718));
  nor_5  g11370(.A(new_n13718), .B(new_n13713), .Y(new_n13719_1));
  and_5  g11371(.A(new_n13719_1), .B(new_n13710_1), .Y(new_n13720));
  nor_5  g11372(.A(new_n13720), .B(new_n13708_1), .Y(new_n13721));
  nor_5  g11373(.A(new_n13721), .B(new_n13706), .Y(new_n13722_1));
  nor_5  g11374(.A(new_n13722_1), .B(new_n13705), .Y(new_n13723));
  and_5  g11375(.A(new_n13700), .B(new_n12158_1), .Y(new_n13724));
  nor_5  g11376(.A(new_n13701), .B(n5140), .Y(new_n13725));
  nor_5  g11377(.A(new_n13702), .B(new_n12110), .Y(new_n13726));
  nor_5  g11378(.A(new_n13726), .B(new_n13698), .Y(new_n13727));
  nor_5  g11379(.A(new_n13727), .B(new_n13725), .Y(new_n13728));
  nor_5  g11380(.A(new_n13728), .B(new_n13724), .Y(new_n13729));
  not_8  g11381(.A(new_n13729), .Y(new_n13730));
  and_5  g11382(.A(new_n13730), .B(new_n13723), .Y(new_n13731));
  and_5  g11383(.A(new_n13731), .B(new_n13678), .Y(new_n13732));
  or_5   g11384(.A(new_n13730), .B(new_n13723), .Y(new_n13733));
  nor_5  g11385(.A(new_n13733), .B(new_n13678), .Y(new_n13734));
  nor_5  g11386(.A(new_n13734), .B(new_n13732), .Y(new_n13735));
  not_8  g11387(.A(new_n13735), .Y(new_n13736));
  xnor_4 g11388(.A(new_n13736), .B(new_n13674), .Y(new_n13737));
  xnor_4 g11389(.A(new_n13729), .B(new_n13723), .Y(new_n13738));
  xnor_4 g11390(.A(new_n13738), .B(new_n13678), .Y(new_n13739));
  and_5  g11391(.A(new_n13739), .B(new_n13673), .Y(new_n13740));
  or_5   g11392(.A(new_n13739), .B(new_n13673), .Y(new_n13741));
  xor_4  g11393(.A(new_n13671), .B(new_n13644), .Y(new_n13742));
  xnor_4 g11394(.A(new_n13721), .B(new_n13706), .Y(new_n13743));
  nor_5  g11395(.A(new_n13743), .B(new_n13742), .Y(new_n13744));
  xnor_4 g11396(.A(new_n13743), .B(new_n13742), .Y(new_n13745));
  xor_4  g11397(.A(new_n13669), .B(new_n13647), .Y(new_n13746));
  xnor_4 g11398(.A(new_n13719_1), .B(new_n13710_1), .Y(new_n13747));
  nor_5  g11399(.A(new_n13747), .B(new_n13746), .Y(new_n13748));
  xnor_4 g11400(.A(new_n13747), .B(new_n13746), .Y(new_n13749));
  xor_4  g11401(.A(new_n13667), .B(new_n13650), .Y(new_n13750));
  xnor_4 g11402(.A(new_n13717), .B(new_n13714_1), .Y(new_n13751));
  not_8  g11403(.A(new_n13751), .Y(new_n13752));
  nor_5  g11404(.A(new_n13752), .B(new_n13750), .Y(new_n13753));
  xnor_4 g11405(.A(new_n13752), .B(new_n13750), .Y(new_n13754_1));
  xor_4  g11406(.A(new_n13665), .B(new_n13653), .Y(new_n13755));
  nor_5  g11407(.A(new_n13755), .B(new_n6552), .Y(new_n13756));
  xor_4  g11408(.A(new_n13663), .B(new_n13655), .Y(new_n13757));
  nor_5  g11409(.A(new_n13757), .B(new_n6554), .Y(new_n13758));
  xnor_4 g11410(.A(new_n13757), .B(new_n6554), .Y(new_n13759));
  not_8  g11411(.A(new_n6557), .Y(new_n13760));
  xnor_4 g11412(.A(new_n13661), .B(new_n13657), .Y(new_n13761));
  and_5  g11413(.A(new_n13761), .B(new_n13760), .Y(new_n13762));
  xnor_4 g11414(.A(new_n13761), .B(new_n13760), .Y(new_n13763));
  and_5  g11415(.A(new_n12026), .B(new_n6560_1), .Y(new_n13764_1));
  nor_5  g11416(.A(new_n12041), .B(new_n12027), .Y(new_n13765));
  nor_5  g11417(.A(new_n13765), .B(new_n13764_1), .Y(new_n13766));
  nor_5  g11418(.A(new_n13766), .B(new_n13763), .Y(new_n13767));
  nor_5  g11419(.A(new_n13767), .B(new_n13762), .Y(new_n13768));
  nor_5  g11420(.A(new_n13768), .B(new_n13759), .Y(new_n13769));
  nor_5  g11421(.A(new_n13769), .B(new_n13758), .Y(new_n13770));
  xnor_4 g11422(.A(new_n13755), .B(new_n6552), .Y(new_n13771));
  nor_5  g11423(.A(new_n13771), .B(new_n13770), .Y(new_n13772));
  nor_5  g11424(.A(new_n13772), .B(new_n13756), .Y(new_n13773));
  nor_5  g11425(.A(new_n13773), .B(new_n13754_1), .Y(new_n13774));
  nor_5  g11426(.A(new_n13774), .B(new_n13753), .Y(new_n13775_1));
  nor_5  g11427(.A(new_n13775_1), .B(new_n13749), .Y(new_n13776));
  nor_5  g11428(.A(new_n13776), .B(new_n13748), .Y(new_n13777));
  nor_5  g11429(.A(new_n13777), .B(new_n13745), .Y(new_n13778));
  nor_5  g11430(.A(new_n13778), .B(new_n13744), .Y(new_n13779));
  and_5  g11431(.A(new_n13779), .B(new_n13741), .Y(new_n13780));
  nor_5  g11432(.A(new_n13780), .B(new_n13740), .Y(new_n13781_1));
  xnor_4 g11433(.A(new_n13781_1), .B(new_n13737), .Y(n2711));
  xnor_4 g11434(.A(n10611), .B(n2680), .Y(new_n13783_1));
  nor_5  g11435(.A(n2783), .B(new_n10614_1), .Y(new_n13784));
  nor_5  g11436(.A(new_n6593), .B(n1667), .Y(new_n13785));
  and_5  g11437(.A(new_n9099), .B(n7339), .Y(new_n13786));
  or_5   g11438(.A(new_n9099), .B(n7339), .Y(new_n13787));
  nor_5  g11439(.A(new_n9155), .B(n18), .Y(new_n13788));
  and_5  g11440(.A(new_n13788), .B(new_n13787), .Y(new_n13789));
  nor_5  g11441(.A(new_n13789), .B(new_n13786), .Y(new_n13790));
  nor_5  g11442(.A(new_n13790), .B(new_n13785), .Y(new_n13791));
  or_5   g11443(.A(new_n13791), .B(new_n13784), .Y(new_n13792));
  xor_4  g11444(.A(new_n13792), .B(new_n13783_1), .Y(new_n13793));
  xnor_4 g11445(.A(new_n13793), .B(new_n9023), .Y(new_n13794));
  xnor_4 g11446(.A(n2783), .B(n1667), .Y(new_n13795));
  xnor_4 g11447(.A(new_n13795), .B(new_n13790), .Y(new_n13796));
  and_5  g11448(.A(new_n13796), .B(new_n9027), .Y(new_n13797));
  xnor_4 g11449(.A(new_n13796), .B(new_n9027), .Y(new_n13798_1));
  xnor_4 g11450(.A(n26808), .B(n18), .Y(new_n13799));
  nor_5  g11451(.A(new_n13799), .B(new_n9034), .Y(new_n13800));
  xnor_4 g11452(.A(n15490), .B(n7339), .Y(new_n13801));
  xnor_4 g11453(.A(new_n13801), .B(new_n13788), .Y(new_n13802));
  nor_5  g11454(.A(new_n13802), .B(new_n13800), .Y(new_n13803));
  xnor_4 g11455(.A(new_n13802), .B(new_n13800), .Y(new_n13804));
  nor_5  g11456(.A(new_n13804), .B(new_n9039), .Y(new_n13805));
  nor_5  g11457(.A(new_n13805), .B(new_n13803), .Y(new_n13806));
  nor_5  g11458(.A(new_n13806), .B(new_n13798_1), .Y(new_n13807));
  nor_5  g11459(.A(new_n13807), .B(new_n13797), .Y(new_n13808));
  xnor_4 g11460(.A(new_n13808), .B(new_n13794), .Y(n2761));
  xnor_4 g11461(.A(n25120), .B(n8526), .Y(new_n13810));
  nor_5  g11462(.A(n8363), .B(n2816), .Y(new_n13811));
  xnor_4 g11463(.A(n8363), .B(new_n6025), .Y(new_n13812));
  nor_5  g11464(.A(n20359), .B(n14680), .Y(new_n13813));
  xnor_4 g11465(.A(n20359), .B(n14680), .Y(new_n13814));
  nor_5  g11466(.A(n17250), .B(n4409), .Y(new_n13815));
  or_5   g11467(.A(new_n9309), .B(new_n9289), .Y(new_n13816));
  and_5  g11468(.A(new_n13816), .B(new_n9288), .Y(new_n13817));
  nor_5  g11469(.A(new_n13817), .B(new_n13815), .Y(new_n13818));
  nor_5  g11470(.A(new_n13818), .B(new_n13814), .Y(new_n13819));
  or_5   g11471(.A(new_n13819), .B(new_n13813), .Y(new_n13820));
  and_5  g11472(.A(new_n13820), .B(new_n13812), .Y(new_n13821));
  nor_5  g11473(.A(new_n13821), .B(new_n13811), .Y(new_n13822));
  xnor_4 g11474(.A(new_n13822), .B(new_n13810), .Y(new_n13823));
  nor_5  g11475(.A(new_n13823), .B(n17458), .Y(new_n13824));
  xnor_4 g11476(.A(new_n13823), .B(new_n10870), .Y(new_n13825));
  nor_5  g11477(.A(new_n13819), .B(new_n13813), .Y(new_n13826));
  xnor_4 g11478(.A(new_n13826), .B(new_n13812), .Y(new_n13827));
  nor_5  g11479(.A(new_n13827), .B(new_n10873), .Y(new_n13828));
  xnor_4 g11480(.A(new_n13818), .B(new_n13814), .Y(new_n13829));
  nor_5  g11481(.A(new_n13829), .B(n25240), .Y(new_n13830));
  xnor_4 g11482(.A(new_n13829), .B(new_n10876), .Y(new_n13831));
  nor_5  g11483(.A(new_n9311), .B(new_n10414), .Y(new_n13832));
  xnor_4 g11484(.A(new_n9312), .B(new_n10414), .Y(new_n13833));
  nor_5  g11485(.A(new_n9315), .B(new_n10881), .Y(new_n13834));
  xnor_4 g11486(.A(new_n9317), .B(new_n10881), .Y(new_n13835_1));
  nor_5  g11487(.A(new_n9320), .B(new_n10884), .Y(new_n13836));
  xnor_4 g11488(.A(new_n9322), .B(new_n10884), .Y(new_n13837));
  nor_5  g11489(.A(new_n9325), .B(new_n8432_1), .Y(new_n13838));
  xnor_4 g11490(.A(new_n9327), .B(new_n8432_1), .Y(new_n13839));
  nor_5  g11491(.A(new_n9330), .B(new_n7217), .Y(new_n13840));
  nor_5  g11492(.A(new_n9332), .B(n5026), .Y(new_n13841));
  or_5   g11493(.A(new_n9335), .B(new_n6628_1), .Y(new_n13842));
  xnor_4 g11494(.A(new_n9332), .B(new_n7220), .Y(new_n13843));
  and_5  g11495(.A(new_n13843), .B(new_n13842), .Y(new_n13844));
  nor_5  g11496(.A(new_n13844), .B(new_n13841), .Y(new_n13845));
  xnor_4 g11497(.A(new_n9340), .B(new_n7217), .Y(new_n13846));
  and_5  g11498(.A(new_n13846), .B(new_n13845), .Y(new_n13847));
  or_5   g11499(.A(new_n13847), .B(new_n13840), .Y(new_n13848));
  and_5  g11500(.A(new_n13848), .B(new_n13839), .Y(new_n13849));
  or_5   g11501(.A(new_n13849), .B(new_n13838), .Y(new_n13850_1));
  and_5  g11502(.A(new_n13850_1), .B(new_n13837), .Y(new_n13851_1));
  or_5   g11503(.A(new_n13851_1), .B(new_n13836), .Y(new_n13852));
  and_5  g11504(.A(new_n13852), .B(new_n13835_1), .Y(new_n13853));
  or_5   g11505(.A(new_n13853), .B(new_n13834), .Y(new_n13854));
  and_5  g11506(.A(new_n13854), .B(new_n13833), .Y(new_n13855));
  nor_5  g11507(.A(new_n13855), .B(new_n13832), .Y(new_n13856));
  and_5  g11508(.A(new_n13856), .B(new_n13831), .Y(new_n13857));
  nor_5  g11509(.A(new_n13857), .B(new_n13830), .Y(new_n13858));
  not_8  g11510(.A(new_n13827), .Y(new_n13859));
  xnor_4 g11511(.A(new_n13859), .B(new_n10873), .Y(new_n13860));
  and_5  g11512(.A(new_n13860), .B(new_n13858), .Y(new_n13861));
  nor_5  g11513(.A(new_n13861), .B(new_n13828), .Y(new_n13862));
  and_5  g11514(.A(new_n13862), .B(new_n13825), .Y(new_n13863));
  nor_5  g11515(.A(new_n13863), .B(new_n13824), .Y(new_n13864));
  not_8  g11516(.A(new_n13864), .Y(new_n13865));
  nor_5  g11517(.A(n25120), .B(n8526), .Y(new_n13866));
  nor_5  g11518(.A(new_n13822), .B(new_n13810), .Y(new_n13867));
  nor_5  g11519(.A(new_n13867), .B(new_n13866), .Y(new_n13868));
  not_8  g11520(.A(new_n13868), .Y(new_n13869));
  nor_5  g11521(.A(new_n13869), .B(new_n13865), .Y(new_n13870));
  not_8  g11522(.A(new_n3735), .Y(new_n13871));
  nor_5  g11523(.A(new_n13871), .B(n2113), .Y(new_n13872));
  not_8  g11524(.A(new_n13872), .Y(new_n13873));
  nor_5  g11525(.A(new_n13873), .B(n1099), .Y(new_n13874));
  not_8  g11526(.A(new_n13874), .Y(new_n13875));
  nor_5  g11527(.A(new_n13875), .B(n19941), .Y(new_n13876));
  xnor_4 g11528(.A(new_n13876), .B(n11898), .Y(new_n13877));
  nor_5  g11529(.A(new_n13877), .B(new_n4837), .Y(new_n13878));
  not_8  g11530(.A(new_n13877), .Y(new_n13879));
  xnor_4 g11531(.A(new_n13879), .B(new_n4839), .Y(new_n13880));
  xnor_4 g11532(.A(new_n13874), .B(n19941), .Y(new_n13881));
  nor_5  g11533(.A(new_n13881), .B(new_n4841), .Y(new_n13882));
  xnor_4 g11534(.A(new_n13881), .B(new_n4841), .Y(new_n13883));
  xnor_4 g11535(.A(new_n13872), .B(n1099), .Y(new_n13884));
  nor_5  g11536(.A(new_n13884), .B(new_n4845), .Y(new_n13885));
  xnor_4 g11537(.A(new_n13884), .B(new_n4845), .Y(new_n13886));
  nor_5  g11538(.A(new_n4850_1), .B(new_n3736), .Y(new_n13887));
  xnor_4 g11539(.A(new_n4850_1), .B(new_n3736), .Y(new_n13888));
  nor_5  g11540(.A(new_n4854), .B(new_n3738), .Y(new_n13889));
  xnor_4 g11541(.A(new_n4854), .B(new_n3738), .Y(new_n13890));
  nor_5  g11542(.A(new_n4859), .B(new_n3742), .Y(new_n13891));
  xnor_4 g11543(.A(new_n4859), .B(new_n3742), .Y(new_n13892));
  nor_5  g11544(.A(new_n4864), .B(new_n3746), .Y(new_n13893));
  xnor_4 g11545(.A(new_n4864), .B(new_n3746), .Y(new_n13894));
  nor_5  g11546(.A(new_n4869), .B(new_n3748), .Y(new_n13895));
  xnor_4 g11547(.A(new_n4880), .B(new_n3748), .Y(new_n13896));
  nor_5  g11548(.A(new_n4874), .B(n25435), .Y(new_n13897));
  and_5  g11549(.A(new_n13897), .B(new_n3752), .Y(new_n13898));
  nor_5  g11550(.A(new_n13897), .B(new_n3758_1), .Y(new_n13899));
  nor_5  g11551(.A(new_n13899), .B(new_n13898), .Y(new_n13900));
  and_5  g11552(.A(new_n13900), .B(new_n4872), .Y(new_n13901));
  or_5   g11553(.A(new_n13901), .B(new_n13898), .Y(new_n13902));
  and_5  g11554(.A(new_n13902), .B(new_n13896), .Y(new_n13903));
  nor_5  g11555(.A(new_n13903), .B(new_n13895), .Y(new_n13904));
  nor_5  g11556(.A(new_n13904), .B(new_n13894), .Y(new_n13905));
  nor_5  g11557(.A(new_n13905), .B(new_n13893), .Y(new_n13906));
  nor_5  g11558(.A(new_n13906), .B(new_n13892), .Y(new_n13907));
  nor_5  g11559(.A(new_n13907), .B(new_n13891), .Y(new_n13908));
  nor_5  g11560(.A(new_n13908), .B(new_n13890), .Y(new_n13909));
  nor_5  g11561(.A(new_n13909), .B(new_n13889), .Y(new_n13910));
  nor_5  g11562(.A(new_n13910), .B(new_n13888), .Y(new_n13911));
  nor_5  g11563(.A(new_n13911), .B(new_n13887), .Y(new_n13912_1));
  nor_5  g11564(.A(new_n13912_1), .B(new_n13886), .Y(new_n13913));
  nor_5  g11565(.A(new_n13913), .B(new_n13885), .Y(new_n13914_1));
  nor_5  g11566(.A(new_n13914_1), .B(new_n13883), .Y(new_n13915));
  nor_5  g11567(.A(new_n13915), .B(new_n13882), .Y(new_n13916));
  nor_5  g11568(.A(new_n13916), .B(new_n13880), .Y(new_n13917));
  nor_5  g11569(.A(new_n13917), .B(new_n13878), .Y(new_n13918));
  not_8  g11570(.A(new_n4901), .Y(new_n13919));
  and_5  g11571(.A(new_n13876), .B(new_n12671), .Y(new_n13920));
  and_5  g11572(.A(new_n13920), .B(new_n13919), .Y(new_n13921));
  and_5  g11573(.A(new_n13921), .B(new_n13918), .Y(new_n13922_1));
  or_5   g11574(.A(new_n13920), .B(new_n13919), .Y(new_n13923_1));
  nor_5  g11575(.A(new_n13923_1), .B(new_n13918), .Y(new_n13924));
  nor_5  g11576(.A(new_n13924), .B(new_n13922_1), .Y(new_n13925));
  and_5  g11577(.A(new_n13925), .B(new_n13870), .Y(new_n13926));
  or_5   g11578(.A(new_n13925), .B(new_n13870), .Y(new_n13927));
  xnor_4 g11579(.A(new_n13868), .B(new_n13865), .Y(new_n13928));
  xnor_4 g11580(.A(new_n13920), .B(new_n4901), .Y(new_n13929));
  xnor_4 g11581(.A(new_n13929), .B(new_n13918), .Y(new_n13930));
  nor_5  g11582(.A(new_n13930), .B(new_n13928), .Y(new_n13931));
  xnor_4 g11583(.A(new_n13930), .B(new_n13928), .Y(new_n13932));
  xnor_4 g11584(.A(new_n13862), .B(new_n13825), .Y(new_n13933));
  xnor_4 g11585(.A(new_n13916), .B(new_n13880), .Y(new_n13934));
  nor_5  g11586(.A(new_n13934), .B(new_n13933), .Y(new_n13935));
  xnor_4 g11587(.A(new_n13934), .B(new_n13933), .Y(new_n13936));
  xnor_4 g11588(.A(new_n13914_1), .B(new_n13883), .Y(new_n13937));
  xor_4  g11589(.A(new_n13860), .B(new_n13858), .Y(new_n13938));
  nor_5  g11590(.A(new_n13938), .B(new_n13937), .Y(new_n13939));
  xnor_4 g11591(.A(new_n13938), .B(new_n13937), .Y(new_n13940));
  xnor_4 g11592(.A(new_n13856), .B(new_n13831), .Y(new_n13941));
  xnor_4 g11593(.A(new_n13912_1), .B(new_n13886), .Y(new_n13942));
  nor_5  g11594(.A(new_n13942), .B(new_n13941), .Y(new_n13943));
  xnor_4 g11595(.A(new_n13942), .B(new_n13941), .Y(new_n13944));
  xnor_4 g11596(.A(new_n13910), .B(new_n13888), .Y(new_n13945));
  xor_4  g11597(.A(new_n13854), .B(new_n13833), .Y(new_n13946));
  nor_5  g11598(.A(new_n13946), .B(new_n13945), .Y(new_n13947));
  xnor_4 g11599(.A(new_n13946), .B(new_n13945), .Y(new_n13948));
  xnor_4 g11600(.A(new_n13908), .B(new_n13890), .Y(new_n13949));
  xor_4  g11601(.A(new_n13852), .B(new_n13835_1), .Y(new_n13950));
  nor_5  g11602(.A(new_n13950), .B(new_n13949), .Y(new_n13951_1));
  xnor_4 g11603(.A(new_n13950), .B(new_n13949), .Y(new_n13952));
  xnor_4 g11604(.A(new_n13906), .B(new_n13892), .Y(new_n13953));
  xor_4  g11605(.A(new_n13850_1), .B(new_n13837), .Y(new_n13954));
  nor_5  g11606(.A(new_n13954), .B(new_n13953), .Y(new_n13955));
  xnor_4 g11607(.A(new_n13954), .B(new_n13953), .Y(new_n13956));
  xnor_4 g11608(.A(new_n13904), .B(new_n13894), .Y(new_n13957));
  xor_4  g11609(.A(new_n13848), .B(new_n13839), .Y(new_n13958));
  nor_5  g11610(.A(new_n13958), .B(new_n13957), .Y(new_n13959));
  xnor_4 g11611(.A(new_n13958), .B(new_n13957), .Y(new_n13960));
  not_8  g11612(.A(new_n13960), .Y(new_n13961));
  xor_4  g11613(.A(new_n13902), .B(new_n13896), .Y(new_n13962));
  xnor_4 g11614(.A(new_n13846), .B(new_n13845), .Y(new_n13963));
  nor_5  g11615(.A(new_n13963), .B(new_n13962), .Y(new_n13964));
  xor_4  g11616(.A(new_n13963), .B(new_n13962), .Y(new_n13965));
  xor_4  g11617(.A(new_n13843), .B(new_n13842), .Y(new_n13966));
  xnor_4 g11618(.A(new_n13900), .B(new_n4871), .Y(new_n13967));
  and_5  g11619(.A(new_n13967), .B(new_n13966), .Y(new_n13968));
  xnor_4 g11620(.A(new_n9335), .B(n8581), .Y(new_n13969));
  xnor_4 g11621(.A(new_n4874), .B(n25435), .Y(new_n13970));
  and_5  g11622(.A(new_n13970), .B(new_n13969), .Y(new_n13971));
  xnor_4 g11623(.A(new_n13967), .B(new_n13966), .Y(new_n13972));
  nor_5  g11624(.A(new_n13972), .B(new_n13971), .Y(new_n13973));
  nor_5  g11625(.A(new_n13973), .B(new_n13968), .Y(new_n13974));
  and_5  g11626(.A(new_n13974), .B(new_n13965), .Y(new_n13975));
  nor_5  g11627(.A(new_n13975), .B(new_n13964), .Y(new_n13976));
  and_5  g11628(.A(new_n13976), .B(new_n13961), .Y(new_n13977));
  nor_5  g11629(.A(new_n13977), .B(new_n13959), .Y(new_n13978));
  nor_5  g11630(.A(new_n13978), .B(new_n13956), .Y(new_n13979));
  nor_5  g11631(.A(new_n13979), .B(new_n13955), .Y(new_n13980));
  nor_5  g11632(.A(new_n13980), .B(new_n13952), .Y(new_n13981));
  nor_5  g11633(.A(new_n13981), .B(new_n13951_1), .Y(new_n13982));
  nor_5  g11634(.A(new_n13982), .B(new_n13948), .Y(new_n13983));
  nor_5  g11635(.A(new_n13983), .B(new_n13947), .Y(new_n13984));
  nor_5  g11636(.A(new_n13984), .B(new_n13944), .Y(new_n13985));
  nor_5  g11637(.A(new_n13985), .B(new_n13943), .Y(new_n13986));
  nor_5  g11638(.A(new_n13986), .B(new_n13940), .Y(new_n13987));
  nor_5  g11639(.A(new_n13987), .B(new_n13939), .Y(new_n13988));
  nor_5  g11640(.A(new_n13988), .B(new_n13936), .Y(new_n13989));
  nor_5  g11641(.A(new_n13989), .B(new_n13935), .Y(new_n13990));
  nor_5  g11642(.A(new_n13990), .B(new_n13932), .Y(new_n13991));
  nor_5  g11643(.A(new_n13991), .B(new_n13931), .Y(new_n13992));
  and_5  g11644(.A(new_n13992), .B(new_n13927), .Y(new_n13993));
  or_5   g11645(.A(new_n13993), .B(new_n13922_1), .Y(new_n13994));
  nor_5  g11646(.A(new_n13994), .B(new_n13926), .Y(n2774));
  not_8  g11647(.A(new_n9395), .Y(new_n13996));
  nor_5  g11648(.A(new_n13996), .B(n20478), .Y(new_n13997));
  not_8  g11649(.A(new_n13997), .Y(new_n13998));
  nor_5  g11650(.A(new_n13998), .B(n987), .Y(new_n13999));
  not_8  g11651(.A(new_n13999), .Y(new_n14000));
  nor_5  g11652(.A(new_n14000), .B(n2421), .Y(new_n14001));
  not_8  g11653(.A(new_n14001), .Y(new_n14002));
  nor_5  g11654(.A(new_n14002), .B(n11044), .Y(new_n14003));
  not_8  g11655(.A(new_n14003), .Y(new_n14004_1));
  nor_5  g11656(.A(new_n14004_1), .B(n5031), .Y(new_n14005));
  xnor_4 g11657(.A(new_n14005), .B(n2145), .Y(new_n14006));
  xnor_4 g11658(.A(new_n14006), .B(new_n4909), .Y(new_n14007));
  xnor_4 g11659(.A(new_n14003), .B(n5031), .Y(new_n14008));
  nor_5  g11660(.A(new_n14008), .B(n2659), .Y(new_n14009));
  xnor_4 g11661(.A(new_n14008), .B(new_n4913_1), .Y(new_n14010));
  xnor_4 g11662(.A(new_n14001), .B(n11044), .Y(new_n14011));
  nor_5  g11663(.A(new_n14011), .B(n24327), .Y(new_n14012));
  xnor_4 g11664(.A(new_n14011), .B(new_n4917), .Y(new_n14013));
  xnor_4 g11665(.A(new_n13999), .B(n2421), .Y(new_n14014));
  nor_5  g11666(.A(new_n14014), .B(n22198), .Y(new_n14015));
  xnor_4 g11667(.A(new_n13997), .B(n987), .Y(new_n14016));
  and_5  g11668(.A(new_n14016), .B(n20826), .Y(new_n14017));
  xnor_4 g11669(.A(new_n14016), .B(new_n4927), .Y(new_n14018));
  and_5  g11670(.A(new_n9396_1), .B(n7305), .Y(new_n14019));
  or_5   g11671(.A(new_n9407), .B(new_n9399_1), .Y(new_n14020));
  and_5  g11672(.A(new_n14020), .B(new_n9397), .Y(new_n14021));
  or_5   g11673(.A(new_n14021), .B(new_n14019), .Y(new_n14022));
  and_5  g11674(.A(new_n14022), .B(new_n14018), .Y(new_n14023));
  nor_5  g11675(.A(new_n14023), .B(new_n14017), .Y(new_n14024));
  xnor_4 g11676(.A(new_n14014), .B(new_n4922), .Y(new_n14025));
  and_5  g11677(.A(new_n14025), .B(new_n14024), .Y(new_n14026));
  or_5   g11678(.A(new_n14026), .B(new_n14015), .Y(new_n14027));
  and_5  g11679(.A(new_n14027), .B(new_n14013), .Y(new_n14028));
  or_5   g11680(.A(new_n14028), .B(new_n14012), .Y(new_n14029));
  and_5  g11681(.A(new_n14029), .B(new_n14010), .Y(new_n14030));
  nor_5  g11682(.A(new_n14030), .B(new_n14009), .Y(new_n14031));
  xnor_4 g11683(.A(new_n14031), .B(new_n14007), .Y(new_n14032));
  xnor_4 g11684(.A(new_n14032), .B(new_n3476), .Y(new_n14033));
  nor_5  g11685(.A(new_n14028), .B(new_n14012), .Y(new_n14034));
  xnor_4 g11686(.A(new_n14034), .B(new_n14010), .Y(new_n14035));
  nor_5  g11687(.A(new_n14035), .B(new_n3480_1), .Y(new_n14036_1));
  xor_4  g11688(.A(new_n14027), .B(new_n14013), .Y(new_n14037));
  not_8  g11689(.A(new_n14037), .Y(new_n14038));
  nor_5  g11690(.A(new_n14038), .B(new_n3486), .Y(new_n14039));
  xnor_4 g11691(.A(new_n14038), .B(new_n3486), .Y(new_n14040));
  xnor_4 g11692(.A(new_n14025), .B(new_n14024), .Y(new_n14041));
  nor_5  g11693(.A(new_n14041), .B(new_n3491), .Y(new_n14042));
  not_8  g11694(.A(new_n14041), .Y(new_n14043));
  xnor_4 g11695(.A(new_n14043), .B(new_n3490), .Y(new_n14044));
  nor_5  g11696(.A(new_n14021), .B(new_n14019), .Y(new_n14045));
  xnor_4 g11697(.A(new_n14045), .B(new_n14018), .Y(new_n14046));
  nor_5  g11698(.A(new_n14046), .B(new_n3495), .Y(new_n14047));
  not_8  g11699(.A(new_n14046), .Y(new_n14048));
  xnor_4 g11700(.A(new_n14048), .B(new_n3495), .Y(new_n14049));
  not_8  g11701(.A(new_n9409), .Y(new_n14050));
  nor_5  g11702(.A(new_n14050), .B(new_n3500), .Y(new_n14051));
  xnor_4 g11703(.A(new_n14050), .B(new_n3501), .Y(new_n14052));
  nor_5  g11704(.A(new_n9428), .B(new_n3507), .Y(new_n14053));
  xnor_4 g11705(.A(new_n9428), .B(new_n3509), .Y(new_n14054));
  nor_5  g11706(.A(new_n9431), .B(new_n3513), .Y(new_n14055));
  nor_5  g11707(.A(new_n9434), .B(new_n3516_1), .Y(new_n14056));
  not_8  g11708(.A(new_n9431), .Y(new_n14057));
  xnor_4 g11709(.A(new_n14057), .B(new_n3513), .Y(new_n14058));
  and_5  g11710(.A(new_n14058), .B(new_n14056), .Y(new_n14059_1));
  or_5   g11711(.A(new_n14059_1), .B(new_n14055), .Y(new_n14060));
  and_5  g11712(.A(new_n14060), .B(new_n14054), .Y(new_n14061));
  or_5   g11713(.A(new_n14061), .B(new_n14053), .Y(new_n14062));
  and_5  g11714(.A(new_n14062), .B(new_n14052), .Y(new_n14063));
  nor_5  g11715(.A(new_n14063), .B(new_n14051), .Y(new_n14064));
  and_5  g11716(.A(new_n14064), .B(new_n14049), .Y(new_n14065));
  nor_5  g11717(.A(new_n14065), .B(new_n14047), .Y(new_n14066));
  nor_5  g11718(.A(new_n14066), .B(new_n14044), .Y(new_n14067));
  nor_5  g11719(.A(new_n14067), .B(new_n14042), .Y(new_n14068));
  nor_5  g11720(.A(new_n14068), .B(new_n14040), .Y(new_n14069));
  nor_5  g11721(.A(new_n14069), .B(new_n14039), .Y(new_n14070));
  xnor_4 g11722(.A(new_n14035), .B(new_n3481), .Y(new_n14071_1));
  and_5  g11723(.A(new_n14071_1), .B(new_n14070), .Y(new_n14072));
  nor_5  g11724(.A(new_n14072), .B(new_n14036_1), .Y(new_n14073));
  xnor_4 g11725(.A(new_n14073), .B(new_n14033), .Y(new_n14074));
  not_8  g11726(.A(new_n14074), .Y(new_n14075));
  xnor_4 g11727(.A(new_n3603), .B(n7026), .Y(new_n14076));
  nor_5  g11728(.A(new_n3611), .B(new_n3540), .Y(new_n14077));
  or_5   g11729(.A(new_n3608), .B(n13719), .Y(new_n14078));
  nor_5  g11730(.A(new_n3614), .B(n442), .Y(new_n14079));
  xnor_4 g11731(.A(new_n3614), .B(new_n3543), .Y(new_n14080));
  nor_5  g11732(.A(new_n3618_1), .B(n9172), .Y(new_n14081_1));
  xnor_4 g11733(.A(new_n3618_1), .B(n9172), .Y(new_n14082));
  nor_5  g11734(.A(new_n3621), .B(n4913), .Y(new_n14083));
  xnor_4 g11735(.A(new_n3621), .B(new_n3549), .Y(new_n14084));
  nor_5  g11736(.A(new_n3625), .B(n604), .Y(new_n14085));
  nor_5  g11737(.A(new_n3629), .B(n16824), .Y(new_n14086));
  xnor_4 g11738(.A(new_n3630), .B(n16824), .Y(new_n14087));
  nor_5  g11739(.A(new_n3636), .B(n16521), .Y(new_n14088));
  nand_5 g11740(.A(n21993), .B(n7139), .Y(new_n14089));
  xnor_4 g11741(.A(new_n3643), .B(n16521), .Y(new_n14090_1));
  and_5  g11742(.A(new_n14090_1), .B(new_n14089), .Y(new_n14091));
  or_5   g11743(.A(new_n14091), .B(new_n14088), .Y(new_n14092));
  and_5  g11744(.A(new_n14092), .B(new_n14087), .Y(new_n14093));
  or_5   g11745(.A(new_n14093), .B(new_n14086), .Y(new_n14094));
  xnor_4 g11746(.A(new_n3626), .B(n604), .Y(new_n14095_1));
  and_5  g11747(.A(new_n14095_1), .B(new_n14094), .Y(new_n14096));
  or_5   g11748(.A(new_n14096), .B(new_n14085), .Y(new_n14097));
  and_5  g11749(.A(new_n14097), .B(new_n14084), .Y(new_n14098));
  nor_5  g11750(.A(new_n14098), .B(new_n14083), .Y(new_n14099));
  nor_5  g11751(.A(new_n14099), .B(new_n14082), .Y(new_n14100));
  or_5   g11752(.A(new_n14100), .B(new_n14081_1), .Y(new_n14101));
  and_5  g11753(.A(new_n14101), .B(new_n14080), .Y(new_n14102));
  nor_5  g11754(.A(new_n14102), .B(new_n14079), .Y(new_n14103));
  and_5  g11755(.A(new_n14103), .B(new_n14078), .Y(new_n14104));
  nor_5  g11756(.A(new_n14104), .B(new_n14077), .Y(new_n14105));
  xnor_4 g11757(.A(new_n14105), .B(new_n14076), .Y(new_n14106));
  xnor_4 g11758(.A(new_n14106), .B(new_n14075), .Y(new_n14107_1));
  xnor_4 g11759(.A(new_n14071_1), .B(new_n14070), .Y(new_n14108));
  xnor_4 g11760(.A(new_n3611), .B(n13719), .Y(new_n14109));
  xnor_4 g11761(.A(new_n14109), .B(new_n14103), .Y(new_n14110));
  nor_5  g11762(.A(new_n14110), .B(new_n14108), .Y(new_n14111));
  not_8  g11763(.A(new_n14108), .Y(new_n14112));
  xnor_4 g11764(.A(new_n14110), .B(new_n14112), .Y(new_n14113));
  xor_4  g11765(.A(new_n14101), .B(new_n14080), .Y(new_n14114));
  xnor_4 g11766(.A(new_n14068), .B(new_n14040), .Y(new_n14115));
  not_8  g11767(.A(new_n14115), .Y(new_n14116));
  and_5  g11768(.A(new_n14116), .B(new_n14114), .Y(new_n14117));
  xnor_4 g11769(.A(new_n14116), .B(new_n14114), .Y(new_n14118));
  xnor_4 g11770(.A(new_n14099), .B(new_n14082), .Y(new_n14119));
  xnor_4 g11771(.A(new_n14066), .B(new_n14044), .Y(new_n14120));
  nor_5  g11772(.A(new_n14120), .B(new_n14119), .Y(new_n14121_1));
  not_8  g11773(.A(new_n14120), .Y(new_n14122));
  xnor_4 g11774(.A(new_n14122), .B(new_n14119), .Y(new_n14123));
  xor_4  g11775(.A(new_n14097), .B(new_n14084), .Y(new_n14124));
  xor_4  g11776(.A(new_n14064), .B(new_n14049), .Y(new_n14125));
  nor_5  g11777(.A(new_n14125), .B(new_n14124), .Y(new_n14126_1));
  xor_4  g11778(.A(new_n14095_1), .B(new_n14094), .Y(new_n14127));
  nor_5  g11779(.A(new_n14061), .B(new_n14053), .Y(new_n14128));
  xnor_4 g11780(.A(new_n14128), .B(new_n14052), .Y(new_n14129));
  not_8  g11781(.A(new_n14129), .Y(new_n14130_1));
  nor_5  g11782(.A(new_n14130_1), .B(new_n14127), .Y(new_n14131));
  xnor_4 g11783(.A(new_n14129), .B(new_n14127), .Y(new_n14132));
  xor_4  g11784(.A(new_n14092), .B(new_n14087), .Y(new_n14133));
  nor_5  g11785(.A(new_n14059_1), .B(new_n14055), .Y(new_n14134));
  xnor_4 g11786(.A(new_n14134), .B(new_n14054), .Y(new_n14135));
  not_8  g11787(.A(new_n14135), .Y(new_n14136_1));
  nor_5  g11788(.A(new_n14136_1), .B(new_n14133), .Y(new_n14137));
  xnor_4 g11789(.A(new_n14135), .B(new_n14133), .Y(new_n14138));
  xnor_4 g11790(.A(new_n14058), .B(new_n14056), .Y(new_n14139));
  not_8  g11791(.A(new_n14139), .Y(new_n14140));
  nor_5  g11792(.A(new_n14140), .B(new_n14090_1), .Y(new_n14141));
  xor_4  g11793(.A(new_n14090_1), .B(new_n14089), .Y(new_n14142));
  nor_5  g11794(.A(new_n14142), .B(new_n14139), .Y(new_n14143));
  xnor_4 g11795(.A(n21993), .B(n7139), .Y(new_n14144));
  xnor_4 g11796(.A(new_n9433), .B(new_n3516_1), .Y(new_n14145));
  not_8  g11797(.A(new_n14145), .Y(new_n14146));
  nor_5  g11798(.A(new_n14146), .B(new_n14144), .Y(new_n14147_1));
  nor_5  g11799(.A(new_n14147_1), .B(new_n14143), .Y(new_n14148_1));
  nor_5  g11800(.A(new_n14148_1), .B(new_n14141), .Y(new_n14149));
  and_5  g11801(.A(new_n14149), .B(new_n14138), .Y(new_n14150));
  or_5   g11802(.A(new_n14150), .B(new_n14137), .Y(new_n14151));
  and_5  g11803(.A(new_n14151), .B(new_n14132), .Y(new_n14152));
  nor_5  g11804(.A(new_n14152), .B(new_n14131), .Y(new_n14153));
  xnor_4 g11805(.A(new_n14125), .B(new_n14124), .Y(new_n14154));
  nor_5  g11806(.A(new_n14154), .B(new_n14153), .Y(new_n14155));
  nor_5  g11807(.A(new_n14155), .B(new_n14126_1), .Y(new_n14156));
  and_5  g11808(.A(new_n14156), .B(new_n14123), .Y(new_n14157));
  nor_5  g11809(.A(new_n14157), .B(new_n14121_1), .Y(new_n14158));
  nor_5  g11810(.A(new_n14158), .B(new_n14118), .Y(new_n14159));
  nor_5  g11811(.A(new_n14159), .B(new_n14117), .Y(new_n14160));
  and_5  g11812(.A(new_n14160), .B(new_n14113), .Y(new_n14161));
  nor_5  g11813(.A(new_n14161), .B(new_n14111), .Y(new_n14162));
  xnor_4 g11814(.A(new_n14162), .B(new_n14107_1), .Y(n2779));
  nor_5  g11815(.A(new_n10243), .B(n25751), .Y(new_n14164));
  not_8  g11816(.A(n25751), .Y(new_n14165));
  xnor_4 g11817(.A(new_n10243), .B(new_n14165), .Y(new_n14166));
  nor_5  g11818(.A(new_n10246), .B(n26053), .Y(new_n14167));
  not_8  g11819(.A(n26053), .Y(new_n14168));
  xnor_4 g11820(.A(new_n10246), .B(new_n14168), .Y(new_n14169));
  nor_5  g11821(.A(new_n10249), .B(n7917), .Y(new_n14170));
  not_8  g11822(.A(n7917), .Y(new_n14171));
  xnor_4 g11823(.A(new_n10249), .B(new_n14171), .Y(new_n14172));
  nor_5  g11824(.A(new_n10252), .B(n17302), .Y(new_n14173));
  not_8  g11825(.A(n17302), .Y(new_n14174_1));
  xnor_4 g11826(.A(new_n10252), .B(new_n14174_1), .Y(new_n14175));
  nor_5  g11827(.A(new_n10254), .B(n2013), .Y(new_n14176));
  not_8  g11828(.A(n2013), .Y(new_n14177));
  xnor_4 g11829(.A(new_n10254), .B(new_n14177), .Y(new_n14178));
  nor_5  g11830(.A(new_n10257), .B(n23755), .Y(new_n14179));
  nor_5  g11831(.A(new_n10260), .B(n19163), .Y(new_n14180));
  not_8  g11832(.A(n19163), .Y(new_n14181));
  xnor_4 g11833(.A(new_n10260), .B(new_n14181), .Y(new_n14182));
  not_8  g11834(.A(n22358), .Y(new_n14183));
  and_5  g11835(.A(new_n5811), .B(new_n14183), .Y(new_n14184));
  nor_5  g11836(.A(new_n3982), .B(new_n6585), .Y(new_n14185));
  xnor_4 g11837(.A(new_n5811), .B(new_n14183), .Y(new_n14186));
  nor_5  g11838(.A(new_n14186), .B(new_n14185), .Y(new_n14187));
  or_5   g11839(.A(new_n14187), .B(new_n14184), .Y(new_n14188));
  and_5  g11840(.A(new_n14188), .B(new_n14182), .Y(new_n14189));
  or_5   g11841(.A(new_n14189), .B(new_n14180), .Y(new_n14190_1));
  not_8  g11842(.A(n23755), .Y(new_n14191));
  xnor_4 g11843(.A(new_n10257), .B(new_n14191), .Y(new_n14192));
  and_5  g11844(.A(new_n14192), .B(new_n14190_1), .Y(new_n14193));
  or_5   g11845(.A(new_n14193), .B(new_n14179), .Y(new_n14194));
  and_5  g11846(.A(new_n14194), .B(new_n14178), .Y(new_n14195));
  or_5   g11847(.A(new_n14195), .B(new_n14176), .Y(new_n14196));
  and_5  g11848(.A(new_n14196), .B(new_n14175), .Y(new_n14197));
  or_5   g11849(.A(new_n14197), .B(new_n14173), .Y(new_n14198));
  and_5  g11850(.A(new_n14198), .B(new_n14172), .Y(new_n14199));
  or_5   g11851(.A(new_n14199), .B(new_n14170), .Y(new_n14200));
  and_5  g11852(.A(new_n14200), .B(new_n14169), .Y(new_n14201));
  or_5   g11853(.A(new_n14201), .B(new_n14167), .Y(new_n14202));
  and_5  g11854(.A(new_n14202), .B(new_n14166), .Y(new_n14203));
  nor_5  g11855(.A(new_n14203), .B(new_n14164), .Y(new_n14204));
  xnor_4 g11856(.A(new_n10281), .B(n25586), .Y(new_n14205));
  xnor_4 g11857(.A(new_n14205), .B(new_n14204), .Y(new_n14206));
  xnor_4 g11858(.A(new_n14206), .B(n4514), .Y(new_n14207));
  xor_4  g11859(.A(new_n14202), .B(new_n14166), .Y(new_n14208));
  nor_5  g11860(.A(new_n14208), .B(n3984), .Y(new_n14209));
  xnor_4 g11861(.A(new_n14208), .B(n3984), .Y(new_n14210));
  xor_4  g11862(.A(new_n14200), .B(new_n14169), .Y(new_n14211_1));
  nor_5  g11863(.A(new_n14211_1), .B(n19652), .Y(new_n14212));
  xnor_4 g11864(.A(new_n14211_1), .B(n19652), .Y(new_n14213));
  xor_4  g11865(.A(new_n14198), .B(new_n14172), .Y(new_n14214));
  nor_5  g11866(.A(new_n14214), .B(n3366), .Y(new_n14215));
  xor_4  g11867(.A(new_n14196), .B(new_n14175), .Y(new_n14216));
  nor_5  g11868(.A(new_n14216), .B(n26565), .Y(new_n14217));
  xnor_4 g11869(.A(new_n14216), .B(n26565), .Y(new_n14218));
  xor_4  g11870(.A(new_n14194), .B(new_n14178), .Y(new_n14219));
  nor_5  g11871(.A(new_n14219), .B(n3959), .Y(new_n14220));
  xnor_4 g11872(.A(new_n14219), .B(n3959), .Y(new_n14221));
  xor_4  g11873(.A(new_n14192), .B(new_n14190_1), .Y(new_n14222_1));
  nor_5  g11874(.A(new_n14222_1), .B(n11566), .Y(new_n14223));
  xnor_4 g11875(.A(new_n14222_1), .B(n11566), .Y(new_n14224));
  xor_4  g11876(.A(new_n14188), .B(new_n14182), .Y(new_n14225));
  nor_5  g11877(.A(new_n14225), .B(n26744), .Y(new_n14226));
  xor_4  g11878(.A(new_n14186), .B(new_n14185), .Y(new_n14227));
  nor_5  g11879(.A(new_n14227), .B(n26625), .Y(new_n14228));
  nor_5  g11880(.A(new_n6586), .B(new_n9484), .Y(new_n14229));
  xnor_4 g11881(.A(new_n14227), .B(n26625), .Y(new_n14230_1));
  nor_5  g11882(.A(new_n14230_1), .B(new_n14229), .Y(new_n14231));
  nor_5  g11883(.A(new_n14231), .B(new_n14228), .Y(new_n14232));
  xnor_4 g11884(.A(new_n14225), .B(n26744), .Y(new_n14233));
  nor_5  g11885(.A(new_n14233), .B(new_n14232), .Y(new_n14234));
  nor_5  g11886(.A(new_n14234), .B(new_n14226), .Y(new_n14235));
  nor_5  g11887(.A(new_n14235), .B(new_n14224), .Y(new_n14236));
  nor_5  g11888(.A(new_n14236), .B(new_n14223), .Y(new_n14237));
  nor_5  g11889(.A(new_n14237), .B(new_n14221), .Y(new_n14238));
  nor_5  g11890(.A(new_n14238), .B(new_n14220), .Y(new_n14239));
  nor_5  g11891(.A(new_n14239), .B(new_n14218), .Y(new_n14240));
  nor_5  g11892(.A(new_n14240), .B(new_n14217), .Y(new_n14241));
  xnor_4 g11893(.A(new_n14214), .B(n3366), .Y(new_n14242));
  nor_5  g11894(.A(new_n14242), .B(new_n14241), .Y(new_n14243));
  nor_5  g11895(.A(new_n14243), .B(new_n14215), .Y(new_n14244));
  nor_5  g11896(.A(new_n14244), .B(new_n14213), .Y(new_n14245));
  nor_5  g11897(.A(new_n14245), .B(new_n14212), .Y(new_n14246));
  nor_5  g11898(.A(new_n14246), .B(new_n14210), .Y(new_n14247));
  nor_5  g11899(.A(new_n14247), .B(new_n14209), .Y(new_n14248));
  xnor_4 g11900(.A(new_n14248), .B(new_n14207), .Y(new_n14249));
  and_5  g11901(.A(new_n14249), .B(new_n10354), .Y(new_n14250));
  xnor_4 g11902(.A(new_n14249), .B(new_n10354), .Y(new_n14251));
  xor_4  g11903(.A(new_n14246), .B(new_n14210), .Y(new_n14252));
  nor_5  g11904(.A(new_n14252), .B(new_n10359), .Y(new_n14253));
  xnor_4 g11905(.A(new_n14252), .B(new_n10359), .Y(new_n14254));
  xor_4  g11906(.A(new_n14244), .B(new_n14213), .Y(new_n14255));
  nor_5  g11907(.A(new_n14255), .B(new_n10362), .Y(new_n14256));
  xnor_4 g11908(.A(new_n14255), .B(new_n10362), .Y(new_n14257));
  xor_4  g11909(.A(new_n14242), .B(new_n14241), .Y(new_n14258));
  nor_5  g11910(.A(new_n14258), .B(new_n10367), .Y(new_n14259));
  xnor_4 g11911(.A(new_n14258), .B(new_n10367), .Y(new_n14260));
  xor_4  g11912(.A(new_n14239), .B(new_n14218), .Y(new_n14261));
  nor_5  g11913(.A(new_n14261), .B(new_n10370), .Y(new_n14262));
  xnor_4 g11914(.A(new_n14261), .B(new_n10370), .Y(new_n14263));
  xor_4  g11915(.A(new_n14237), .B(new_n14221), .Y(new_n14264));
  nor_5  g11916(.A(new_n14264), .B(new_n10375), .Y(new_n14265));
  xnor_4 g11917(.A(new_n14264), .B(new_n10375), .Y(new_n14266));
  xor_4  g11918(.A(new_n14235), .B(new_n14224), .Y(new_n14267_1));
  nor_5  g11919(.A(new_n14267_1), .B(new_n10379), .Y(new_n14268));
  xnor_4 g11920(.A(new_n14267_1), .B(new_n10379), .Y(new_n14269));
  xor_4  g11921(.A(new_n14233), .B(new_n14232), .Y(new_n14270));
  nor_5  g11922(.A(new_n14270), .B(new_n10384), .Y(new_n14271_1));
  xnor_4 g11923(.A(new_n14270), .B(new_n10384), .Y(new_n14272));
  xnor_4 g11924(.A(new_n14230_1), .B(new_n14229), .Y(new_n14273));
  not_8  g11925(.A(new_n14273), .Y(new_n14274));
  nor_5  g11926(.A(new_n14274), .B(new_n5808), .Y(new_n14275_1));
  nor_5  g11927(.A(new_n6587_1), .B(new_n5803), .Y(new_n14276));
  nor_5  g11928(.A(new_n14273), .B(new_n5809), .Y(new_n14277_1));
  nor_5  g11929(.A(new_n14277_1), .B(new_n14276), .Y(new_n14278));
  nor_5  g11930(.A(new_n14278), .B(new_n14275_1), .Y(new_n14279));
  nor_5  g11931(.A(new_n14279), .B(new_n14272), .Y(new_n14280));
  nor_5  g11932(.A(new_n14280), .B(new_n14271_1), .Y(new_n14281));
  nor_5  g11933(.A(new_n14281), .B(new_n14269), .Y(new_n14282));
  nor_5  g11934(.A(new_n14282), .B(new_n14268), .Y(new_n14283));
  nor_5  g11935(.A(new_n14283), .B(new_n14266), .Y(new_n14284));
  nor_5  g11936(.A(new_n14284), .B(new_n14265), .Y(new_n14285));
  nor_5  g11937(.A(new_n14285), .B(new_n14263), .Y(new_n14286));
  nor_5  g11938(.A(new_n14286), .B(new_n14262), .Y(new_n14287));
  nor_5  g11939(.A(new_n14287), .B(new_n14260), .Y(new_n14288));
  nor_5  g11940(.A(new_n14288), .B(new_n14259), .Y(new_n14289));
  nor_5  g11941(.A(new_n14289), .B(new_n14257), .Y(new_n14290));
  nor_5  g11942(.A(new_n14290), .B(new_n14256), .Y(new_n14291));
  nor_5  g11943(.A(new_n14291), .B(new_n14254), .Y(new_n14292));
  nor_5  g11944(.A(new_n14292), .B(new_n14253), .Y(new_n14293));
  nor_5  g11945(.A(new_n14293), .B(new_n14251), .Y(new_n14294_1));
  nor_5  g11946(.A(new_n14294_1), .B(new_n14250), .Y(new_n14295));
  xnor_4 g11947(.A(new_n14295), .B(new_n10352), .Y(new_n14296));
  and_5  g11948(.A(new_n14206), .B(n4514), .Y(new_n14297));
  not_8  g11949(.A(new_n14248), .Y(new_n14298));
  nor_5  g11950(.A(new_n14298), .B(new_n14207), .Y(new_n14299));
  or_5   g11951(.A(new_n14299), .B(new_n14297), .Y(new_n14300));
  or_5   g11952(.A(new_n10241), .B(n25586), .Y(new_n14301));
  and_5  g11953(.A(new_n14301), .B(new_n14204), .Y(new_n14302));
  not_8  g11954(.A(n25586), .Y(new_n14303));
  nor_5  g11955(.A(new_n10281), .B(new_n14303), .Y(new_n14304));
  or_5   g11956(.A(new_n14304), .B(new_n10240), .Y(new_n14305));
  nor_5  g11957(.A(new_n14305), .B(new_n14302), .Y(new_n14306));
  xnor_4 g11958(.A(new_n14306), .B(new_n14300), .Y(new_n14307));
  xnor_4 g11959(.A(new_n14307), .B(new_n14296), .Y(n2826));
  nor_5  g11960(.A(new_n6244), .B(new_n12110), .Y(new_n14309));
  xnor_4 g11961(.A(new_n6244), .B(n5140), .Y(new_n14310_1));
  nor_5  g11962(.A(new_n6250), .B(new_n12113_1), .Y(new_n14311));
  xnor_4 g11963(.A(new_n6251), .B(new_n12113_1), .Y(new_n14312));
  nor_5  g11964(.A(new_n6256_1), .B(new_n12116), .Y(new_n14313));
  xnor_4 g11965(.A(new_n6257), .B(new_n12116), .Y(new_n14314));
  nor_5  g11966(.A(new_n6262), .B(new_n12119), .Y(new_n14315));
  xnor_4 g11967(.A(new_n6304), .B(new_n12119), .Y(new_n14316));
  nor_5  g11968(.A(new_n6268), .B(new_n12122), .Y(new_n14317));
  nor_5  g11969(.A(new_n6274), .B(n8244), .Y(new_n14318));
  xnor_4 g11970(.A(new_n6274), .B(new_n12125), .Y(new_n14319));
  nor_5  g11971(.A(new_n6276_1), .B(new_n12128), .Y(new_n14320));
  xnor_4 g11972(.A(new_n6277), .B(new_n12128), .Y(new_n14321));
  nor_5  g11973(.A(new_n6282), .B(n15167), .Y(new_n14322));
  nor_5  g11974(.A(new_n6285), .B(new_n12134), .Y(new_n14323_1));
  nor_5  g11975(.A(new_n6288), .B(new_n6492), .Y(new_n14324));
  xnor_4 g11976(.A(new_n12226), .B(new_n12134), .Y(new_n14325));
  and_5  g11977(.A(new_n14325), .B(new_n14324), .Y(new_n14326_1));
  nor_5  g11978(.A(new_n14326_1), .B(new_n14323_1), .Y(new_n14327));
  xnor_4 g11979(.A(new_n6282), .B(new_n12132), .Y(new_n14328));
  and_5  g11980(.A(new_n14328), .B(new_n14327), .Y(new_n14329));
  nor_5  g11981(.A(new_n14329), .B(new_n14322), .Y(new_n14330));
  and_5  g11982(.A(new_n14330), .B(new_n14321), .Y(new_n14331));
  nor_5  g11983(.A(new_n14331), .B(new_n14320), .Y(new_n14332));
  and_5  g11984(.A(new_n14332), .B(new_n14319), .Y(new_n14333));
  nor_5  g11985(.A(new_n14333), .B(new_n14318), .Y(new_n14334));
  xnor_4 g11986(.A(new_n6269), .B(new_n12122), .Y(new_n14335));
  and_5  g11987(.A(new_n14335), .B(new_n14334), .Y(new_n14336));
  or_5   g11988(.A(new_n14336), .B(new_n14317), .Y(new_n14337));
  and_5  g11989(.A(new_n14337), .B(new_n14316), .Y(new_n14338));
  or_5   g11990(.A(new_n14338), .B(new_n14315), .Y(new_n14339));
  and_5  g11991(.A(new_n14339), .B(new_n14314), .Y(new_n14340));
  or_5   g11992(.A(new_n14340), .B(new_n14313), .Y(new_n14341));
  and_5  g11993(.A(new_n14341), .B(new_n14312), .Y(new_n14342_1));
  or_5   g11994(.A(new_n14342_1), .B(new_n14311), .Y(new_n14343));
  and_5  g11995(.A(new_n14343), .B(new_n14310_1), .Y(new_n14344));
  nor_5  g11996(.A(new_n14344), .B(new_n14309), .Y(new_n14345_1));
  nor_5  g11997(.A(new_n14345_1), .B(new_n6242), .Y(new_n14346));
  not_8  g11998(.A(n25365), .Y(new_n14347));
  nor_5  g11999(.A(new_n2603), .B(new_n14347), .Y(new_n14348));
  or_5   g12000(.A(new_n2653), .B(new_n2606), .Y(new_n14349));
  and_5  g12001(.A(new_n14349), .B(new_n2604), .Y(new_n14350));
  nor_5  g12002(.A(new_n14350), .B(new_n14348), .Y(new_n14351));
  nor_5  g12003(.A(n20040), .B(n9396), .Y(new_n14352));
  nor_5  g12004(.A(new_n2601), .B(new_n2556), .Y(new_n14353_1));
  nor_5  g12005(.A(new_n14353_1), .B(new_n14352), .Y(new_n14354));
  not_8  g12006(.A(new_n14354), .Y(new_n14355));
  nor_5  g12007(.A(new_n14355), .B(new_n14351), .Y(new_n14356));
  not_8  g12008(.A(new_n14356), .Y(new_n14357));
  xnor_4 g12009(.A(new_n14357), .B(new_n14346), .Y(new_n14358));
  xnor_4 g12010(.A(new_n14345_1), .B(new_n6197), .Y(new_n14359));
  not_8  g12011(.A(new_n14359), .Y(new_n14360));
  xnor_4 g12012(.A(new_n14354), .B(new_n14351), .Y(new_n14361));
  and_5  g12013(.A(new_n14361), .B(new_n14360), .Y(new_n14362));
  xnor_4 g12014(.A(new_n14361), .B(new_n14360), .Y(new_n14363));
  xor_4  g12015(.A(new_n14343), .B(new_n14310_1), .Y(new_n14364_1));
  nor_5  g12016(.A(new_n14364_1), .B(new_n2656), .Y(new_n14365));
  xnor_4 g12017(.A(new_n14364_1), .B(new_n2656), .Y(new_n14366));
  xor_4  g12018(.A(new_n14341), .B(new_n14312), .Y(new_n14367));
  nor_5  g12019(.A(new_n14367), .B(new_n2787), .Y(new_n14368));
  xnor_4 g12020(.A(new_n14367), .B(new_n2787), .Y(new_n14369));
  not_8  g12021(.A(new_n2792), .Y(new_n14370));
  xor_4  g12022(.A(new_n14339), .B(new_n14314), .Y(new_n14371));
  nor_5  g12023(.A(new_n14371), .B(new_n14370), .Y(new_n14372));
  xnor_4 g12024(.A(new_n14371), .B(new_n14370), .Y(new_n14373));
  xor_4  g12025(.A(new_n14337), .B(new_n14316), .Y(new_n14374));
  nor_5  g12026(.A(new_n14374), .B(new_n2796), .Y(new_n14375_1));
  xnor_4 g12027(.A(new_n14374), .B(new_n2796), .Y(new_n14376));
  xor_4  g12028(.A(new_n14335), .B(new_n14334), .Y(new_n14377));
  nor_5  g12029(.A(new_n14377), .B(new_n2802), .Y(new_n14378));
  xnor_4 g12030(.A(new_n14377), .B(new_n2802), .Y(new_n14379));
  xnor_4 g12031(.A(new_n14332), .B(new_n14319), .Y(new_n14380));
  nor_5  g12032(.A(new_n14380), .B(new_n2806), .Y(new_n14381));
  xnor_4 g12033(.A(new_n14380), .B(new_n2806), .Y(new_n14382));
  xor_4  g12034(.A(new_n14330), .B(new_n14321), .Y(new_n14383));
  nor_5  g12035(.A(new_n14383), .B(new_n2814), .Y(new_n14384));
  xnor_4 g12036(.A(new_n14383), .B(new_n2814), .Y(new_n14385));
  xnor_4 g12037(.A(new_n14328), .B(new_n14327), .Y(new_n14386));
  nor_5  g12038(.A(new_n14386), .B(new_n2817), .Y(new_n14387));
  xnor_4 g12039(.A(new_n14386), .B(new_n2817), .Y(new_n14388));
  xor_4  g12040(.A(new_n14325), .B(new_n14324), .Y(new_n14389));
  nor_5  g12041(.A(new_n14389), .B(new_n2823), .Y(new_n14390));
  xnor_4 g12042(.A(new_n6288), .B(n8656), .Y(new_n14391));
  nor_5  g12043(.A(new_n14391), .B(new_n2827), .Y(new_n14392));
  xnor_4 g12044(.A(new_n14389), .B(new_n2824), .Y(new_n14393));
  and_5  g12045(.A(new_n14393), .B(new_n14392), .Y(new_n14394));
  nor_5  g12046(.A(new_n14394), .B(new_n14390), .Y(new_n14395));
  nor_5  g12047(.A(new_n14395), .B(new_n14388), .Y(new_n14396));
  nor_5  g12048(.A(new_n14396), .B(new_n14387), .Y(new_n14397));
  nor_5  g12049(.A(new_n14397), .B(new_n14385), .Y(new_n14398));
  nor_5  g12050(.A(new_n14398), .B(new_n14384), .Y(new_n14399));
  nor_5  g12051(.A(new_n14399), .B(new_n14382), .Y(new_n14400));
  nor_5  g12052(.A(new_n14400), .B(new_n14381), .Y(new_n14401));
  nor_5  g12053(.A(new_n14401), .B(new_n14379), .Y(new_n14402));
  nor_5  g12054(.A(new_n14402), .B(new_n14378), .Y(new_n14403));
  nor_5  g12055(.A(new_n14403), .B(new_n14376), .Y(new_n14404));
  nor_5  g12056(.A(new_n14404), .B(new_n14375_1), .Y(new_n14405));
  nor_5  g12057(.A(new_n14405), .B(new_n14373), .Y(new_n14406));
  nor_5  g12058(.A(new_n14406), .B(new_n14372), .Y(new_n14407));
  nor_5  g12059(.A(new_n14407), .B(new_n14369), .Y(new_n14408));
  nor_5  g12060(.A(new_n14408), .B(new_n14368), .Y(new_n14409));
  nor_5  g12061(.A(new_n14409), .B(new_n14366), .Y(new_n14410));
  nor_5  g12062(.A(new_n14410), .B(new_n14365), .Y(new_n14411));
  nor_5  g12063(.A(new_n14411), .B(new_n14363), .Y(new_n14412_1));
  nor_5  g12064(.A(new_n14412_1), .B(new_n14362), .Y(new_n14413));
  xnor_4 g12065(.A(new_n14413), .B(new_n14358), .Y(n2853));
  xnor_4 g12066(.A(n7099), .B(n2035), .Y(new_n14415));
  nor_5  g12067(.A(new_n11685), .B(n5213), .Y(new_n14416));
  xnor_4 g12068(.A(n12811), .B(n5213), .Y(new_n14417));
  nor_5  g12069(.A(n4665), .B(new_n11689), .Y(new_n14418));
  xnor_4 g12070(.A(n4665), .B(n1118), .Y(new_n14419));
  nor_5  g12071(.A(n25974), .B(new_n2866), .Y(new_n14420));
  nor_5  g12072(.A(new_n11693), .B(n19005), .Y(new_n14421));
  nor_5  g12073(.A(new_n2869), .B(n1630), .Y(new_n14422));
  nor_5  g12074(.A(n4326), .B(new_n2909), .Y(new_n14423));
  nor_5  g12075(.A(new_n5287), .B(n1451), .Y(new_n14424));
  not_8  g12076(.A(new_n14424), .Y(new_n14425));
  nor_5  g12077(.A(new_n14425), .B(new_n14423), .Y(new_n14426));
  nor_5  g12078(.A(new_n14426), .B(new_n14422), .Y(new_n14427));
  nor_5  g12079(.A(new_n14427), .B(new_n14421), .Y(new_n14428));
  nor_5  g12080(.A(new_n14428), .B(new_n14420), .Y(new_n14429));
  and_5  g12081(.A(new_n14429), .B(new_n14419), .Y(new_n14430));
  or_5   g12082(.A(new_n14430), .B(new_n14418), .Y(new_n14431));
  and_5  g12083(.A(new_n14431), .B(new_n14417), .Y(new_n14432));
  or_5   g12084(.A(new_n14432), .B(new_n14416), .Y(new_n14433));
  xor_4  g12085(.A(new_n14433), .B(new_n14415), .Y(new_n14434));
  not_8  g12086(.A(n5337), .Y(new_n14435));
  not_8  g12087(.A(new_n4228), .Y(new_n14436));
  nor_5  g12088(.A(new_n14436), .B(n13668), .Y(new_n14437));
  xnor_4 g12089(.A(new_n14437), .B(n3570), .Y(new_n14438));
  xnor_4 g12090(.A(new_n14438), .B(new_n14435), .Y(new_n14439));
  and_5  g12091(.A(new_n4229), .B(n626), .Y(new_n14440_1));
  or_5   g12092(.A(new_n4249), .B(new_n4232), .Y(new_n14441));
  and_5  g12093(.A(new_n14441), .B(new_n4230), .Y(new_n14442));
  nor_5  g12094(.A(new_n14442), .B(new_n14440_1), .Y(new_n14443));
  xnor_4 g12095(.A(new_n14443), .B(new_n14439), .Y(new_n14444));
  not_8  g12096(.A(new_n14444), .Y(new_n14445));
  xnor_4 g12097(.A(new_n14445), .B(new_n10979), .Y(new_n14446));
  not_8  g12098(.A(new_n4251), .Y(new_n14447));
  nor_5  g12099(.A(new_n14447), .B(new_n4222), .Y(new_n14448));
  and_5  g12100(.A(new_n4282), .B(new_n4252), .Y(new_n14449));
  nor_5  g12101(.A(new_n14449), .B(new_n14448), .Y(new_n14450));
  xnor_4 g12102(.A(new_n14450), .B(new_n14446), .Y(new_n14451));
  not_8  g12103(.A(new_n14451), .Y(new_n14452));
  xnor_4 g12104(.A(new_n14452), .B(new_n14434), .Y(new_n14453));
  xor_4  g12105(.A(new_n14431), .B(new_n14417), .Y(new_n14454));
  nor_5  g12106(.A(new_n14454), .B(new_n4283), .Y(new_n14455));
  xnor_4 g12107(.A(new_n14429), .B(new_n14419), .Y(new_n14456));
  and_5  g12108(.A(new_n14456), .B(new_n4287), .Y(new_n14457_1));
  xnor_4 g12109(.A(new_n14456), .B(new_n4287), .Y(new_n14458));
  xnor_4 g12110(.A(n25974), .B(n19005), .Y(new_n14459));
  xnor_4 g12111(.A(new_n14459), .B(new_n14427), .Y(new_n14460));
  and_5  g12112(.A(new_n14460), .B(new_n4292), .Y(new_n14461));
  xnor_4 g12113(.A(new_n14460), .B(new_n4291), .Y(new_n14462));
  xnor_4 g12114(.A(n5438), .B(n1451), .Y(new_n14463));
  nor_5  g12115(.A(new_n14463), .B(new_n4303), .Y(new_n14464_1));
  xnor_4 g12116(.A(n4326), .B(n1630), .Y(new_n14465));
  xnor_4 g12117(.A(new_n14465), .B(new_n14425), .Y(new_n14466));
  not_8  g12118(.A(new_n14466), .Y(new_n14467));
  and_5  g12119(.A(new_n14467), .B(new_n14464_1), .Y(new_n14468));
  xnor_4 g12120(.A(new_n14467), .B(new_n14464_1), .Y(new_n14469));
  nor_5  g12121(.A(new_n14469), .B(new_n4296), .Y(new_n14470));
  nor_5  g12122(.A(new_n14470), .B(new_n14468), .Y(new_n14471_1));
  and_5  g12123(.A(new_n14471_1), .B(new_n14462), .Y(new_n14472));
  nor_5  g12124(.A(new_n14472), .B(new_n14461), .Y(new_n14473));
  nor_5  g12125(.A(new_n14473), .B(new_n14458), .Y(new_n14474));
  nor_5  g12126(.A(new_n14474), .B(new_n14457_1), .Y(new_n14475_1));
  xnor_4 g12127(.A(new_n14454), .B(new_n4283), .Y(new_n14476));
  nor_5  g12128(.A(new_n14476), .B(new_n14475_1), .Y(new_n14477));
  nor_5  g12129(.A(new_n14477), .B(new_n14455), .Y(new_n14478));
  xor_4  g12130(.A(new_n14478), .B(new_n14453), .Y(n2860));
  xnor_4 g12131(.A(new_n13586), .B(new_n13568), .Y(n2887));
  not_8  g12132(.A(new_n14437), .Y(new_n14481));
  nor_5  g12133(.A(new_n14481), .B(n3570), .Y(new_n14482));
  not_8  g12134(.A(new_n14482), .Y(new_n14483));
  nor_5  g12135(.A(new_n14483), .B(n4409), .Y(new_n14484));
  not_8  g12136(.A(new_n14484), .Y(new_n14485));
  nor_5  g12137(.A(new_n14485), .B(n20359), .Y(new_n14486));
  and_5  g12138(.A(new_n14486), .B(new_n6025), .Y(new_n14487));
  xnor_4 g12139(.A(new_n14487), .B(n8526), .Y(new_n14488));
  nor_5  g12140(.A(new_n14488), .B(n21784), .Y(new_n14489));
  xnor_4 g12141(.A(new_n14486), .B(n2816), .Y(new_n14490));
  and_5  g12142(.A(new_n14490), .B(n5521), .Y(new_n14491));
  or_5   g12143(.A(new_n14490), .B(n5521), .Y(new_n14492));
  xnor_4 g12144(.A(new_n14484), .B(n20359), .Y(new_n14493));
  nor_5  g12145(.A(new_n14493), .B(n11926), .Y(new_n14494));
  xnor_4 g12146(.A(new_n14493), .B(n11926), .Y(new_n14495));
  xnor_4 g12147(.A(new_n14482), .B(n4409), .Y(new_n14496));
  and_5  g12148(.A(new_n14496), .B(n4325), .Y(new_n14497));
  nor_5  g12149(.A(new_n14496), .B(n4325), .Y(new_n14498));
  and_5  g12150(.A(new_n14438), .B(n5337), .Y(new_n14499));
  nor_5  g12151(.A(new_n14438), .B(n5337), .Y(new_n14500));
  nor_5  g12152(.A(new_n14443), .B(new_n14500), .Y(new_n14501));
  nor_5  g12153(.A(new_n14501), .B(new_n14499), .Y(new_n14502));
  nor_5  g12154(.A(new_n14502), .B(new_n14498), .Y(new_n14503));
  or_5   g12155(.A(new_n14503), .B(new_n14497), .Y(new_n14504));
  nor_5  g12156(.A(new_n14504), .B(new_n14495), .Y(new_n14505));
  nor_5  g12157(.A(new_n14505), .B(new_n14494), .Y(new_n14506));
  and_5  g12158(.A(new_n14506), .B(new_n14492), .Y(new_n14507));
  nor_5  g12159(.A(new_n14507), .B(new_n14491), .Y(new_n14508));
  nor_5  g12160(.A(new_n14508), .B(new_n14489), .Y(new_n14509));
  and_5  g12161(.A(new_n14487), .B(new_n5981), .Y(new_n14510_1));
  and_5  g12162(.A(new_n14488), .B(n21784), .Y(new_n14511));
  or_5   g12163(.A(new_n14511), .B(new_n14510_1), .Y(new_n14512));
  nor_5  g12164(.A(new_n14512), .B(new_n14509), .Y(new_n14513));
  not_8  g12165(.A(new_n14513), .Y(new_n14514));
  xnor_4 g12166(.A(new_n14514), .B(new_n10955), .Y(new_n14515));
  not_8  g12167(.A(n21784), .Y(new_n14516));
  xnor_4 g12168(.A(new_n14488), .B(new_n14516), .Y(new_n14517));
  xnor_4 g12169(.A(new_n14517), .B(new_n14508), .Y(new_n14518));
  and_5  g12170(.A(new_n14518), .B(new_n10961_1), .Y(new_n14519));
  xnor_4 g12171(.A(new_n14518), .B(new_n10960), .Y(new_n14520));
  xnor_4 g12172(.A(new_n14490), .B(n5521), .Y(new_n14521));
  xnor_4 g12173(.A(new_n14521), .B(new_n14506), .Y(new_n14522));
  nor_5  g12174(.A(new_n14522), .B(new_n10965), .Y(new_n14523));
  xnor_4 g12175(.A(new_n14522), .B(new_n10965), .Y(new_n14524));
  nor_5  g12176(.A(new_n14503), .B(new_n14497), .Y(new_n14525));
  xnor_4 g12177(.A(new_n14525), .B(new_n14495), .Y(new_n14526));
  and_5  g12178(.A(new_n14526), .B(new_n10969), .Y(new_n14527));
  xnor_4 g12179(.A(new_n14496), .B(new_n5991), .Y(new_n14528));
  xnor_4 g12180(.A(new_n14528), .B(new_n14502), .Y(new_n14529));
  and_5  g12181(.A(new_n14529), .B(new_n10974), .Y(new_n14530));
  xnor_4 g12182(.A(new_n14529), .B(new_n10974), .Y(new_n14531));
  and_5  g12183(.A(new_n14444), .B(new_n10979), .Y(new_n14532));
  or_5   g12184(.A(new_n14449), .B(new_n14448), .Y(new_n14533));
  and_5  g12185(.A(new_n14533), .B(new_n14446), .Y(new_n14534));
  nor_5  g12186(.A(new_n14534), .B(new_n14532), .Y(new_n14535));
  nor_5  g12187(.A(new_n14535), .B(new_n14531), .Y(new_n14536));
  nor_5  g12188(.A(new_n14536), .B(new_n14530), .Y(new_n14537));
  xnor_4 g12189(.A(new_n14526), .B(new_n10970), .Y(new_n14538));
  and_5  g12190(.A(new_n14538), .B(new_n14537), .Y(new_n14539));
  nor_5  g12191(.A(new_n14539), .B(new_n14527), .Y(new_n14540));
  nor_5  g12192(.A(new_n14540), .B(new_n14524), .Y(new_n14541_1));
  nor_5  g12193(.A(new_n14541_1), .B(new_n14523), .Y(new_n14542));
  and_5  g12194(.A(new_n14542), .B(new_n14520), .Y(new_n14543));
  nor_5  g12195(.A(new_n14543), .B(new_n14519), .Y(new_n14544));
  xnor_4 g12196(.A(new_n14544), .B(new_n14515), .Y(new_n14545));
  not_8  g12197(.A(new_n14545), .Y(new_n14546_1));
  not_8  g12198(.A(n8827), .Y(new_n14547_1));
  not_8  g12199(.A(new_n4170), .Y(new_n14548));
  nor_5  g12200(.A(new_n14548), .B(n19905), .Y(new_n14549));
  not_8  g12201(.A(new_n14549), .Y(new_n14550));
  nor_5  g12202(.A(new_n14550), .B(n26452), .Y(new_n14551));
  not_8  g12203(.A(new_n14551), .Y(new_n14552));
  nor_5  g12204(.A(new_n14552), .B(n15546), .Y(new_n14553));
  not_8  g12205(.A(new_n14553), .Y(new_n14554));
  nor_5  g12206(.A(new_n14554), .B(n5077), .Y(new_n14555));
  and_5  g12207(.A(new_n14555), .B(new_n12683), .Y(new_n14556));
  and_5  g12208(.A(new_n14556), .B(new_n14547_1), .Y(new_n14557));
  xnor_4 g12209(.A(new_n14556), .B(n8827), .Y(new_n14558));
  nor_5  g12210(.A(new_n14558), .B(n11898), .Y(new_n14559));
  xnor_4 g12211(.A(new_n14555), .B(n18035), .Y(new_n14560));
  nor_5  g12212(.A(new_n14560), .B(n19941), .Y(new_n14561));
  xnor_4 g12213(.A(new_n14560), .B(new_n12673), .Y(new_n14562));
  xnor_4 g12214(.A(new_n14553), .B(n5077), .Y(new_n14563));
  nor_5  g12215(.A(new_n14563), .B(n1099), .Y(new_n14564));
  xnor_4 g12216(.A(new_n14563), .B(n1099), .Y(new_n14565));
  xnor_4 g12217(.A(new_n14551), .B(n15546), .Y(new_n14566));
  nor_5  g12218(.A(new_n14566), .B(n2113), .Y(new_n14567));
  xnor_4 g12219(.A(new_n14549), .B(n26452), .Y(new_n14568));
  nor_5  g12220(.A(new_n14568), .B(n21134), .Y(new_n14569));
  xnor_4 g12221(.A(new_n14568), .B(n21134), .Y(new_n14570_1));
  nor_5  g12222(.A(new_n4171), .B(n6369), .Y(new_n14571));
  and_5  g12223(.A(new_n4193), .B(new_n4172_1), .Y(new_n14572));
  nor_5  g12224(.A(new_n14572), .B(new_n14571), .Y(new_n14573));
  nor_5  g12225(.A(new_n14573), .B(new_n14570_1), .Y(new_n14574));
  or_5   g12226(.A(new_n14574), .B(new_n14569), .Y(new_n14575_1));
  xnor_4 g12227(.A(new_n14566), .B(new_n10434), .Y(new_n14576_1));
  and_5  g12228(.A(new_n14576_1), .B(new_n14575_1), .Y(new_n14577));
  nor_5  g12229(.A(new_n14577), .B(new_n14567), .Y(new_n14578));
  nor_5  g12230(.A(new_n14578), .B(new_n14565), .Y(new_n14579));
  or_5   g12231(.A(new_n14579), .B(new_n14564), .Y(new_n14580));
  and_5  g12232(.A(new_n14580), .B(new_n14562), .Y(new_n14581));
  nor_5  g12233(.A(new_n14581), .B(new_n14561), .Y(new_n14582));
  and_5  g12234(.A(new_n14558), .B(n11898), .Y(new_n14583));
  nor_5  g12235(.A(new_n14583), .B(new_n14582), .Y(new_n14584));
  nor_5  g12236(.A(new_n14584), .B(new_n14559), .Y(new_n14585));
  nor_5  g12237(.A(new_n14585), .B(new_n14557), .Y(new_n14586));
  xnor_4 g12238(.A(new_n14586), .B(new_n14546_1), .Y(new_n14587));
  xnor_4 g12239(.A(new_n14542), .B(new_n14520), .Y(new_n14588));
  not_8  g12240(.A(new_n14588), .Y(new_n14589));
  xnor_4 g12241(.A(new_n14558), .B(new_n12671), .Y(new_n14590));
  xnor_4 g12242(.A(new_n14590), .B(new_n14582), .Y(new_n14591));
  not_8  g12243(.A(new_n14591), .Y(new_n14592));
  nor_5  g12244(.A(new_n14592), .B(new_n14589), .Y(new_n14593_1));
  xnor_4 g12245(.A(new_n14592), .B(new_n14589), .Y(new_n14594));
  xor_4  g12246(.A(new_n14580), .B(new_n14562), .Y(new_n14595));
  not_8  g12247(.A(new_n14595), .Y(new_n14596));
  xnor_4 g12248(.A(new_n14540), .B(new_n14524), .Y(new_n14597));
  nor_5  g12249(.A(new_n14597), .B(new_n14596), .Y(new_n14598));
  xnor_4 g12250(.A(new_n14597), .B(new_n14596), .Y(new_n14599));
  xnor_4 g12251(.A(new_n14578), .B(new_n14565), .Y(new_n14600));
  xnor_4 g12252(.A(new_n14538), .B(new_n14537), .Y(new_n14601));
  nor_5  g12253(.A(new_n14601), .B(new_n14600), .Y(new_n14602));
  not_8  g12254(.A(new_n14600), .Y(new_n14603_1));
  not_8  g12255(.A(new_n14601), .Y(new_n14604));
  xnor_4 g12256(.A(new_n14604), .B(new_n14603_1), .Y(new_n14605));
  xnor_4 g12257(.A(new_n14535), .B(new_n14531), .Y(new_n14606));
  xor_4  g12258(.A(new_n14576_1), .B(new_n14575_1), .Y(new_n14607));
  and_5  g12259(.A(new_n14607), .B(new_n14606), .Y(new_n14608));
  xnor_4 g12260(.A(new_n14607), .B(new_n14606), .Y(new_n14609));
  xnor_4 g12261(.A(new_n14573), .B(new_n14570_1), .Y(new_n14610));
  nor_5  g12262(.A(new_n14610), .B(new_n14451), .Y(new_n14611));
  not_8  g12263(.A(new_n14610), .Y(new_n14612));
  xnor_4 g12264(.A(new_n14612), .B(new_n14452), .Y(new_n14613));
  nor_5  g12265(.A(new_n4283), .B(new_n4194), .Y(new_n14614));
  and_5  g12266(.A(new_n4310), .B(new_n4284), .Y(new_n14615));
  nor_5  g12267(.A(new_n14615), .B(new_n14614), .Y(new_n14616));
  nor_5  g12268(.A(new_n14616), .B(new_n14613), .Y(new_n14617));
  nor_5  g12269(.A(new_n14617), .B(new_n14611), .Y(new_n14618));
  nor_5  g12270(.A(new_n14618), .B(new_n14609), .Y(new_n14619));
  nor_5  g12271(.A(new_n14619), .B(new_n14608), .Y(new_n14620));
  nor_5  g12272(.A(new_n14620), .B(new_n14605), .Y(new_n14621));
  nor_5  g12273(.A(new_n14621), .B(new_n14602), .Y(new_n14622));
  nor_5  g12274(.A(new_n14622), .B(new_n14599), .Y(new_n14623));
  nor_5  g12275(.A(new_n14623), .B(new_n14598), .Y(new_n14624));
  nor_5  g12276(.A(new_n14624), .B(new_n14594), .Y(new_n14625));
  nor_5  g12277(.A(new_n14625), .B(new_n14593_1), .Y(new_n14626));
  xor_4  g12278(.A(new_n14626), .B(new_n14587), .Y(n2929));
  not_8  g12279(.A(new_n7269), .Y(new_n14628));
  xnor_4 g12280(.A(n22793), .B(n767), .Y(new_n14629));
  not_8  g12281(.A(n7330), .Y(new_n14630));
  nor_5  g12282(.A(n8439), .B(new_n14630), .Y(new_n14631));
  xnor_4 g12283(.A(n8439), .B(n7330), .Y(new_n14632));
  nor_5  g12284(.A(n25523), .B(new_n2683), .Y(new_n14633_1));
  xnor_4 g12285(.A(n25523), .B(n22492), .Y(new_n14634));
  not_8  g12286(.A(n12821), .Y(new_n14635));
  nor_5  g12287(.A(new_n14635), .B(n5579), .Y(new_n14636_1));
  xnor_4 g12288(.A(n12821), .B(n5579), .Y(new_n14637));
  nor_5  g12289(.A(n23430), .B(new_n2689), .Y(new_n14638));
  xnor_4 g12290(.A(n23430), .B(n3468), .Y(new_n14639));
  not_8  g12291(.A(n10411), .Y(new_n14640));
  nor_5  g12292(.A(n18558), .B(new_n14640), .Y(new_n14641));
  and_5  g12293(.A(new_n13323), .B(new_n13313), .Y(new_n14642));
  nor_5  g12294(.A(new_n14642), .B(new_n14641), .Y(new_n14643));
  and_5  g12295(.A(new_n14643), .B(new_n14639), .Y(new_n14644));
  or_5   g12296(.A(new_n14644), .B(new_n14638), .Y(new_n14645));
  and_5  g12297(.A(new_n14645), .B(new_n14637), .Y(new_n14646));
  or_5   g12298(.A(new_n14646), .B(new_n14636_1), .Y(new_n14647));
  and_5  g12299(.A(new_n14647), .B(new_n14634), .Y(new_n14648));
  or_5   g12300(.A(new_n14648), .B(new_n14633_1), .Y(new_n14649));
  and_5  g12301(.A(new_n14649), .B(new_n14632), .Y(new_n14650));
  nor_5  g12302(.A(new_n14650), .B(new_n14631), .Y(new_n14651));
  xnor_4 g12303(.A(new_n14651), .B(new_n14629), .Y(new_n14652));
  not_8  g12304(.A(new_n14652), .Y(new_n14653));
  xnor_4 g12305(.A(new_n14653), .B(new_n14628), .Y(new_n14654));
  xor_4  g12306(.A(new_n14649), .B(new_n14632), .Y(new_n14655));
  and_5  g12307(.A(new_n14655), .B(new_n7274), .Y(new_n14656));
  not_8  g12308(.A(new_n7274), .Y(new_n14657));
  xnor_4 g12309(.A(new_n14655), .B(new_n14657), .Y(new_n14658));
  xor_4  g12310(.A(new_n14647), .B(new_n14634), .Y(new_n14659));
  nor_5  g12311(.A(new_n14659), .B(new_n7278), .Y(new_n14660));
  xnor_4 g12312(.A(new_n14659), .B(new_n7278), .Y(new_n14661));
  xor_4  g12313(.A(new_n14645), .B(new_n14637), .Y(new_n14662));
  nor_5  g12314(.A(new_n14662), .B(new_n7282), .Y(new_n14663));
  xnor_4 g12315(.A(new_n14662), .B(new_n11953), .Y(new_n14664));
  xnor_4 g12316(.A(new_n14643), .B(new_n14639), .Y(new_n14665));
  not_8  g12317(.A(new_n14665), .Y(new_n14666));
  and_5  g12318(.A(new_n14666), .B(new_n7285), .Y(new_n14667));
  xnor_4 g12319(.A(new_n14665), .B(new_n7285), .Y(new_n14668));
  nor_5  g12320(.A(new_n13324), .B(new_n7290), .Y(new_n14669));
  or_5   g12321(.A(new_n13606), .B(new_n13599), .Y(new_n14670));
  and_5  g12322(.A(new_n14670), .B(new_n13598), .Y(new_n14671));
  or_5   g12323(.A(new_n14671), .B(new_n14669), .Y(new_n14672));
  and_5  g12324(.A(new_n14672), .B(new_n14668), .Y(new_n14673));
  nor_5  g12325(.A(new_n14673), .B(new_n14667), .Y(new_n14674));
  and_5  g12326(.A(new_n14674), .B(new_n14664), .Y(new_n14675));
  nor_5  g12327(.A(new_n14675), .B(new_n14663), .Y(new_n14676));
  nor_5  g12328(.A(new_n14676), .B(new_n14661), .Y(new_n14677));
  nor_5  g12329(.A(new_n14677), .B(new_n14660), .Y(new_n14678));
  and_5  g12330(.A(new_n14678), .B(new_n14658), .Y(new_n14679));
  nor_5  g12331(.A(new_n14679), .B(new_n14656), .Y(new_n14680_1));
  xnor_4 g12332(.A(new_n14680_1), .B(new_n14654), .Y(new_n14681));
  not_8  g12333(.A(new_n14681), .Y(new_n14682));
  xnor_4 g12334(.A(n22379), .B(n15077), .Y(new_n14683));
  nor_5  g12335(.A(n3710), .B(new_n2850), .Y(new_n14684_1));
  xnor_4 g12336(.A(n3710), .B(n1662), .Y(new_n14685));
  nor_5  g12337(.A(n26318), .B(new_n2853_1), .Y(new_n14686));
  xnor_4 g12338(.A(n26318), .B(n12875), .Y(new_n14687));
  nor_5  g12339(.A(n26054), .B(new_n2856), .Y(new_n14688));
  xnor_4 g12340(.A(n26054), .B(n2035), .Y(new_n14689));
  nor_5  g12341(.A(n19081), .B(new_n2859), .Y(new_n14690));
  or_5   g12342(.A(new_n8753), .B(n5213), .Y(new_n14691));
  nor_5  g12343(.A(new_n8771), .B(n4665), .Y(new_n14692_1));
  and_5  g12344(.A(new_n13619), .B(new_n13610), .Y(new_n14693));
  nor_5  g12345(.A(new_n14693), .B(new_n14692_1), .Y(new_n14694));
  and_5  g12346(.A(new_n14694), .B(new_n14691), .Y(new_n14695));
  or_5   g12347(.A(new_n14695), .B(new_n14690), .Y(new_n14696));
  and_5  g12348(.A(new_n14696), .B(new_n14689), .Y(new_n14697));
  or_5   g12349(.A(new_n14697), .B(new_n14688), .Y(new_n14698));
  and_5  g12350(.A(new_n14698), .B(new_n14687), .Y(new_n14699));
  or_5   g12351(.A(new_n14699), .B(new_n14686), .Y(new_n14700));
  and_5  g12352(.A(new_n14700), .B(new_n14685), .Y(new_n14701_1));
  or_5   g12353(.A(new_n14701_1), .B(new_n14684_1), .Y(new_n14702_1));
  xor_4  g12354(.A(new_n14702_1), .B(new_n14683), .Y(new_n14703));
  xnor_4 g12355(.A(new_n14703), .B(new_n14682), .Y(new_n14704_1));
  xor_4  g12356(.A(new_n14700), .B(new_n14685), .Y(new_n14705));
  xor_4  g12357(.A(new_n14678), .B(new_n14658), .Y(new_n14706));
  nor_5  g12358(.A(new_n14706), .B(new_n14705), .Y(new_n14707));
  xnor_4 g12359(.A(new_n14706), .B(new_n14705), .Y(new_n14708));
  xor_4  g12360(.A(new_n14698), .B(new_n14687), .Y(new_n14709));
  xnor_4 g12361(.A(new_n14676), .B(new_n14661), .Y(new_n14710));
  nor_5  g12362(.A(new_n14710), .B(new_n14709), .Y(new_n14711));
  xnor_4 g12363(.A(new_n14710), .B(new_n14709), .Y(new_n14712));
  xor_4  g12364(.A(new_n14696), .B(new_n14689), .Y(new_n14713));
  xnor_4 g12365(.A(new_n14674), .B(new_n14664), .Y(new_n14714));
  nor_5  g12366(.A(new_n14714), .B(new_n14713), .Y(new_n14715));
  nor_5  g12367(.A(new_n14671), .B(new_n14669), .Y(new_n14716));
  xnor_4 g12368(.A(new_n14716), .B(new_n14668), .Y(new_n14717));
  not_8  g12369(.A(new_n14717), .Y(new_n14718));
  xnor_4 g12370(.A(n19081), .B(n5213), .Y(new_n14719));
  xnor_4 g12371(.A(new_n14719), .B(new_n14694), .Y(new_n14720));
  and_5  g12372(.A(new_n14720), .B(new_n14718), .Y(new_n14721));
  xnor_4 g12373(.A(new_n14720), .B(new_n14718), .Y(new_n14722));
  and_5  g12374(.A(new_n13620), .B(new_n13609), .Y(new_n14723));
  nor_5  g12375(.A(new_n13640), .B(new_n13621), .Y(new_n14724));
  nor_5  g12376(.A(new_n14724), .B(new_n14723), .Y(new_n14725));
  nor_5  g12377(.A(new_n14725), .B(new_n14722), .Y(new_n14726));
  nor_5  g12378(.A(new_n14726), .B(new_n14721), .Y(new_n14727));
  xnor_4 g12379(.A(new_n14714), .B(new_n14713), .Y(new_n14728));
  nor_5  g12380(.A(new_n14728), .B(new_n14727), .Y(new_n14729));
  nor_5  g12381(.A(new_n14729), .B(new_n14715), .Y(new_n14730));
  nor_5  g12382(.A(new_n14730), .B(new_n14712), .Y(new_n14731));
  nor_5  g12383(.A(new_n14731), .B(new_n14711), .Y(new_n14732));
  nor_5  g12384(.A(new_n14732), .B(new_n14708), .Y(new_n14733));
  nor_5  g12385(.A(new_n14733), .B(new_n14707), .Y(new_n14734_1));
  xnor_4 g12386(.A(new_n14734_1), .B(new_n14704_1), .Y(n2948));
  xor_4  g12387(.A(new_n14151), .B(new_n14132), .Y(n2961));
  xnor_4 g12388(.A(new_n11261_1), .B(new_n11239), .Y(n2971));
  xnor_4 g12389(.A(new_n2534), .B(new_n2515_1), .Y(n3010));
  xor_4  g12390(.A(new_n6737), .B(new_n6727), .Y(n3017));
  xnor_4 g12391(.A(new_n11592), .B(new_n8996), .Y(new_n14740));
  xnor_4 g12392(.A(new_n14740), .B(new_n11597), .Y(n3020));
  xnor_4 g12393(.A(new_n6139), .B(new_n6114), .Y(n3067));
  xnor_4 g12394(.A(n23541), .B(new_n2582_1), .Y(new_n14743));
  xnor_4 g12395(.A(n27134), .B(n4588), .Y(new_n14744));
  xnor_4 g12396(.A(new_n14744), .B(new_n14743), .Y(new_n14745));
  xnor_4 g12397(.A(new_n14745), .B(new_n9885), .Y(n3076));
  nor_5  g12398(.A(n15490), .B(n18), .Y(new_n14747));
  not_8  g12399(.A(new_n14747), .Y(new_n14748));
  nor_5  g12400(.A(new_n14748), .B(n2783), .Y(new_n14749));
  xnor_4 g12401(.A(new_n14749), .B(n10611), .Y(new_n14750));
  xnor_4 g12402(.A(new_n14750), .B(new_n6589), .Y(new_n14751));
  xnor_4 g12403(.A(new_n14747), .B(n2783), .Y(new_n14752));
  not_8  g12404(.A(new_n14752), .Y(new_n14753));
  nor_5  g12405(.A(new_n14753), .B(new_n6606), .Y(new_n14754));
  xnor_4 g12406(.A(new_n14753), .B(n19680), .Y(new_n14755));
  xnor_4 g12407(.A(n15490), .B(n18), .Y(new_n14756));
  and_5  g12408(.A(new_n14756), .B(new_n6616), .Y(new_n14757));
  or_5   g12409(.A(new_n4818), .B(new_n6596_1), .Y(new_n14758));
  xnor_4 g12410(.A(new_n14756), .B(n2809), .Y(new_n14759));
  and_5  g12411(.A(new_n14759), .B(new_n14758), .Y(new_n14760));
  nor_5  g12412(.A(new_n14760), .B(new_n14757), .Y(new_n14761));
  and_5  g12413(.A(new_n14761), .B(new_n14755), .Y(new_n14762));
  or_5   g12414(.A(new_n14762), .B(new_n14754), .Y(new_n14763_1));
  xor_4  g12415(.A(new_n14763_1), .B(new_n14751), .Y(new_n14764));
  xnor_4 g12416(.A(new_n14764), .B(new_n10584), .Y(new_n14765));
  xnor_4 g12417(.A(new_n14761), .B(new_n14755), .Y(new_n14766));
  nor_5  g12418(.A(new_n14766), .B(new_n10589), .Y(new_n14767));
  xnor_4 g12419(.A(new_n14766), .B(new_n10588_1), .Y(new_n14768));
  nor_5  g12420(.A(new_n14759), .B(new_n5790), .Y(new_n14769));
  xor_4  g12421(.A(new_n14759), .B(new_n14758), .Y(new_n14770));
  nor_5  g12422(.A(new_n14770), .B(new_n10592), .Y(new_n14771));
  xnor_4 g12423(.A(n15508), .B(n18), .Y(new_n14772_1));
  nor_5  g12424(.A(new_n14772_1), .B(new_n5772), .Y(new_n14773));
  nor_5  g12425(.A(new_n14773), .B(new_n14771), .Y(new_n14774));
  nor_5  g12426(.A(new_n14774), .B(new_n14769), .Y(new_n14775));
  and_5  g12427(.A(new_n14775), .B(new_n14768), .Y(new_n14776));
  nor_5  g12428(.A(new_n14776), .B(new_n14767), .Y(new_n14777));
  xor_4  g12429(.A(new_n14777), .B(new_n14765), .Y(n3089));
  xnor_4 g12430(.A(new_n5201), .B(new_n5200), .Y(n3125));
  xnor_4 g12431(.A(n21839), .B(new_n10958), .Y(new_n14780));
  nor_5  g12432(.A(n27089), .B(n12657), .Y(new_n14781));
  or_5   g12433(.A(new_n2967), .B(new_n2928), .Y(new_n14782));
  and_5  g12434(.A(new_n14782), .B(new_n2927), .Y(new_n14783));
  nor_5  g12435(.A(new_n14783), .B(new_n14781), .Y(new_n14784));
  xnor_4 g12436(.A(new_n14784), .B(new_n14780), .Y(new_n14785));
  nor_5  g12437(.A(new_n14785), .B(new_n10923), .Y(new_n14786));
  xnor_4 g12438(.A(new_n14785), .B(new_n10923), .Y(new_n14787));
  nor_5  g12439(.A(new_n10926), .B(new_n2969), .Y(new_n14788));
  nor_5  g12440(.A(new_n10929), .B(new_n2973), .Y(new_n14789));
  xnor_4 g12441(.A(new_n10929), .B(new_n2974), .Y(new_n14790_1));
  not_8  g12442(.A(new_n2981), .Y(new_n14791));
  nor_5  g12443(.A(new_n10933), .B(new_n14791), .Y(new_n14792));
  xnor_4 g12444(.A(new_n10932), .B(new_n14791), .Y(new_n14793));
  nor_5  g12445(.A(new_n10937), .B(new_n13097), .Y(new_n14794));
  and_5  g12446(.A(new_n13115), .B(new_n13098), .Y(new_n14795));
  or_5   g12447(.A(new_n14795), .B(new_n14794), .Y(new_n14796));
  and_5  g12448(.A(new_n14796), .B(new_n14793), .Y(new_n14797));
  nor_5  g12449(.A(new_n14797), .B(new_n14792), .Y(new_n14798));
  and_5  g12450(.A(new_n14798), .B(new_n14790_1), .Y(new_n14799));
  or_5   g12451(.A(new_n14799), .B(new_n14789), .Y(new_n14800));
  not_8  g12452(.A(new_n2969), .Y(new_n14801_1));
  xnor_4 g12453(.A(new_n10926), .B(new_n14801_1), .Y(new_n14802));
  and_5  g12454(.A(new_n14802), .B(new_n14800), .Y(new_n14803));
  nor_5  g12455(.A(new_n14803), .B(new_n14788), .Y(new_n14804));
  nor_5  g12456(.A(new_n14804), .B(new_n14787), .Y(new_n14805));
  nor_5  g12457(.A(new_n14805), .B(new_n14786), .Y(new_n14806));
  nor_5  g12458(.A(n21839), .B(n19282), .Y(new_n14807));
  or_5   g12459(.A(new_n14783), .B(new_n14781), .Y(new_n14808));
  and_5  g12460(.A(new_n14808), .B(new_n14780), .Y(new_n14809));
  nor_5  g12461(.A(new_n14809), .B(new_n14807), .Y(new_n14810));
  not_8  g12462(.A(new_n14810), .Y(new_n14811));
  and_5  g12463(.A(new_n14811), .B(new_n10925), .Y(new_n14812));
  and_5  g12464(.A(new_n14812), .B(new_n14806), .Y(new_n14813));
  or_5   g12465(.A(new_n14811), .B(new_n10925), .Y(new_n14814));
  nor_5  g12466(.A(new_n14814), .B(new_n14806), .Y(new_n14815));
  nor_5  g12467(.A(new_n14815), .B(new_n14813), .Y(new_n14816));
  xnor_4 g12468(.A(new_n14816), .B(new_n11794), .Y(new_n14817));
  xnor_4 g12469(.A(new_n14810), .B(new_n10925), .Y(new_n14818));
  xnor_4 g12470(.A(new_n14818), .B(new_n14806), .Y(new_n14819_1));
  nor_5  g12471(.A(new_n14819_1), .B(new_n11324), .Y(new_n14820));
  xnor_4 g12472(.A(new_n14819_1), .B(new_n11324), .Y(new_n14821));
  xnor_4 g12473(.A(new_n14804), .B(new_n14787), .Y(new_n14822));
  nor_5  g12474(.A(new_n14822), .B(new_n11339), .Y(new_n14823));
  xnor_4 g12475(.A(new_n14822), .B(new_n11339), .Y(new_n14824));
  xor_4  g12476(.A(new_n14802), .B(new_n14800), .Y(new_n14825));
  and_5  g12477(.A(new_n14825), .B(new_n11858), .Y(new_n14826_1));
  xnor_4 g12478(.A(new_n14825), .B(new_n11858), .Y(new_n14827_1));
  xnor_4 g12479(.A(new_n14798), .B(new_n14790_1), .Y(new_n14828));
  nor_5  g12480(.A(new_n14828), .B(new_n11348_1), .Y(new_n14829));
  xnor_4 g12481(.A(new_n14828), .B(new_n11348_1), .Y(new_n14830));
  xor_4  g12482(.A(new_n14796), .B(new_n14793), .Y(new_n14831));
  nor_5  g12483(.A(new_n14831), .B(new_n11352_1), .Y(new_n14832));
  xnor_4 g12484(.A(new_n14831), .B(new_n11352_1), .Y(new_n14833));
  nor_5  g12485(.A(new_n13116_1), .B(new_n11357), .Y(new_n14834));
  nor_5  g12486(.A(new_n13139), .B(new_n13117), .Y(new_n14835));
  nor_5  g12487(.A(new_n14835), .B(new_n14834), .Y(new_n14836));
  nor_5  g12488(.A(new_n14836), .B(new_n14833), .Y(new_n14837));
  nor_5  g12489(.A(new_n14837), .B(new_n14832), .Y(new_n14838));
  nor_5  g12490(.A(new_n14838), .B(new_n14830), .Y(new_n14839_1));
  nor_5  g12491(.A(new_n14839_1), .B(new_n14829), .Y(new_n14840));
  nor_5  g12492(.A(new_n14840), .B(new_n14827_1), .Y(new_n14841));
  nor_5  g12493(.A(new_n14841), .B(new_n14826_1), .Y(new_n14842));
  nor_5  g12494(.A(new_n14842), .B(new_n14824), .Y(new_n14843));
  nor_5  g12495(.A(new_n14843), .B(new_n14823), .Y(new_n14844));
  nor_5  g12496(.A(new_n14844), .B(new_n14821), .Y(new_n14845));
  nor_5  g12497(.A(new_n14845), .B(new_n14820), .Y(new_n14846));
  not_8  g12498(.A(new_n14846), .Y(new_n14847));
  xnor_4 g12499(.A(new_n14847), .B(new_n14817), .Y(n3126));
  xnor_4 g12500(.A(new_n11898_1), .B(new_n11865), .Y(n3208));
  xnor_4 g12501(.A(new_n13972), .B(new_n13971), .Y(n3219));
  xnor_4 g12502(.A(new_n14395), .B(new_n14388), .Y(n3235));
  xnor_4 g12503(.A(new_n11139), .B(new_n11126), .Y(n3244));
  nor_5  g12504(.A(new_n7926), .B(n5532), .Y(new_n14853));
  not_8  g12505(.A(n11579), .Y(new_n14854));
  nor_5  g12506(.A(new_n14854), .B(n3962), .Y(new_n14855));
  nor_5  g12507(.A(n23513), .B(new_n7931), .Y(new_n14856));
  and_5  g12508(.A(new_n13333_1), .B(new_n9875), .Y(new_n14857));
  nor_5  g12509(.A(n6427), .B(new_n7934), .Y(new_n14858));
  or_5   g12510(.A(new_n14858), .B(new_n14857), .Y(new_n14859));
  and_5  g12511(.A(new_n14859), .B(new_n9823), .Y(new_n14860));
  or_5   g12512(.A(new_n14860), .B(new_n14856), .Y(new_n14861));
  and_5  g12513(.A(new_n14861), .B(new_n9843), .Y(new_n14862));
  or_5   g12514(.A(new_n14862), .B(new_n14855), .Y(new_n14863));
  and_5  g12515(.A(new_n14863), .B(new_n9846), .Y(new_n14864));
  or_5   g12516(.A(new_n14864), .B(new_n14853), .Y(new_n14865));
  xor_4  g12517(.A(new_n14865), .B(new_n9849), .Y(new_n14866));
  xnor_4 g12518(.A(new_n14866), .B(new_n14655), .Y(new_n14867));
  xor_4  g12519(.A(new_n14863), .B(new_n9846), .Y(new_n14868));
  nor_5  g12520(.A(new_n14868), .B(new_n14659), .Y(new_n14869));
  xnor_4 g12521(.A(new_n14868), .B(new_n14659), .Y(new_n14870));
  xor_4  g12522(.A(new_n14861), .B(new_n9843), .Y(new_n14871));
  nor_5  g12523(.A(new_n14871), .B(new_n14662), .Y(new_n14872));
  xnor_4 g12524(.A(new_n14871), .B(new_n14662), .Y(new_n14873));
  xor_4  g12525(.A(new_n14859), .B(new_n9823), .Y(new_n14874));
  nor_5  g12526(.A(new_n14874), .B(new_n14666), .Y(new_n14875));
  xnor_4 g12527(.A(new_n14874), .B(new_n14665), .Y(new_n14876));
  nor_5  g12528(.A(new_n13335), .B(new_n13324), .Y(new_n14877));
  nor_5  g12529(.A(new_n13354), .B(new_n13336), .Y(new_n14878));
  nor_5  g12530(.A(new_n14878), .B(new_n14877), .Y(new_n14879));
  and_5  g12531(.A(new_n14879), .B(new_n14876), .Y(new_n14880));
  nor_5  g12532(.A(new_n14880), .B(new_n14875), .Y(new_n14881));
  nor_5  g12533(.A(new_n14881), .B(new_n14873), .Y(new_n14882));
  nor_5  g12534(.A(new_n14882), .B(new_n14872), .Y(new_n14883));
  nor_5  g12535(.A(new_n14883), .B(new_n14870), .Y(new_n14884));
  nor_5  g12536(.A(new_n14884), .B(new_n14869), .Y(new_n14885));
  xnor_4 g12537(.A(new_n14885), .B(new_n14867), .Y(new_n14886));
  not_8  g12538(.A(new_n14886), .Y(new_n14887));
  nor_5  g12539(.A(n23541), .B(n16247), .Y(new_n14888));
  not_8  g12540(.A(new_n14888), .Y(new_n14889));
  nor_5  g12541(.A(new_n14889), .B(n8638), .Y(new_n14890));
  not_8  g12542(.A(new_n14890), .Y(new_n14891_1));
  nor_5  g12543(.A(new_n14891_1), .B(n15979), .Y(new_n14892));
  not_8  g12544(.A(new_n14892), .Y(new_n14893));
  nor_5  g12545(.A(new_n14893), .B(n26483), .Y(new_n14894));
  not_8  g12546(.A(new_n14894), .Y(new_n14895));
  nor_5  g12547(.A(new_n14895), .B(n24768), .Y(new_n14896));
  not_8  g12548(.A(new_n14896), .Y(new_n14897));
  nor_5  g12549(.A(new_n14897), .B(n8687), .Y(new_n14898));
  xnor_4 g12550(.A(new_n14898), .B(n19270), .Y(new_n14899_1));
  xnor_4 g12551(.A(new_n14899_1), .B(new_n2562), .Y(new_n14900));
  xnor_4 g12552(.A(new_n14896), .B(n8687), .Y(new_n14901));
  nor_5  g12553(.A(new_n14901), .B(n13190), .Y(new_n14902));
  xnor_4 g12554(.A(new_n14901), .B(new_n2566), .Y(new_n14903));
  xnor_4 g12555(.A(new_n14894), .B(n24768), .Y(new_n14904));
  nor_5  g12556(.A(new_n14904), .B(n3460), .Y(new_n14905));
  xnor_4 g12557(.A(new_n14904), .B(new_n11305), .Y(new_n14906));
  xnor_4 g12558(.A(new_n14892), .B(n26483), .Y(new_n14907));
  nor_5  g12559(.A(new_n14907), .B(n5226), .Y(new_n14908));
  xnor_4 g12560(.A(new_n14907), .B(new_n9502), .Y(new_n14909));
  xnor_4 g12561(.A(new_n14890), .B(n15979), .Y(new_n14910));
  nor_5  g12562(.A(new_n14910), .B(n17664), .Y(new_n14911));
  xnor_4 g12563(.A(new_n14888), .B(n8638), .Y(new_n14912));
  nor_5  g12564(.A(new_n14912), .B(n23369), .Y(new_n14913));
  xnor_4 g12565(.A(new_n14912), .B(new_n2578_1), .Y(new_n14914));
  xnor_4 g12566(.A(n23541), .B(n16247), .Y(new_n14915));
  and_5  g12567(.A(new_n14915), .B(new_n8697), .Y(new_n14916));
  or_5   g12568(.A(new_n2629), .B(new_n2582_1), .Y(new_n14917));
  xnor_4 g12569(.A(new_n14915), .B(n1136), .Y(new_n14918));
  and_5  g12570(.A(new_n14918), .B(new_n14917), .Y(new_n14919));
  or_5   g12571(.A(new_n14919), .B(new_n14916), .Y(new_n14920));
  and_5  g12572(.A(new_n14920), .B(new_n14914), .Y(new_n14921));
  or_5   g12573(.A(new_n14921), .B(new_n14913), .Y(new_n14922));
  xnor_4 g12574(.A(new_n14910), .B(new_n2574), .Y(new_n14923));
  and_5  g12575(.A(new_n14923), .B(new_n14922), .Y(new_n14924));
  or_5   g12576(.A(new_n14924), .B(new_n14911), .Y(new_n14925));
  and_5  g12577(.A(new_n14925), .B(new_n14909), .Y(new_n14926));
  or_5   g12578(.A(new_n14926), .B(new_n14908), .Y(new_n14927));
  and_5  g12579(.A(new_n14927), .B(new_n14906), .Y(new_n14928));
  or_5   g12580(.A(new_n14928), .B(new_n14905), .Y(new_n14929));
  and_5  g12581(.A(new_n14929), .B(new_n14903), .Y(new_n14930));
  nor_5  g12582(.A(new_n14930), .B(new_n14902), .Y(new_n14931_1));
  xnor_4 g12583(.A(new_n14931_1), .B(new_n14900), .Y(new_n14932));
  xnor_4 g12584(.A(new_n14932), .B(new_n14887), .Y(new_n14933));
  nor_5  g12585(.A(new_n14928), .B(new_n14905), .Y(new_n14934));
  xnor_4 g12586(.A(new_n14934), .B(new_n14903), .Y(new_n14935));
  not_8  g12587(.A(new_n14935), .Y(new_n14936));
  xnor_4 g12588(.A(new_n14883), .B(new_n14870), .Y(new_n14937));
  nor_5  g12589(.A(new_n14937), .B(new_n14936), .Y(new_n14938));
  nor_5  g12590(.A(new_n14926), .B(new_n14908), .Y(new_n14939));
  xnor_4 g12591(.A(new_n14939), .B(new_n14906), .Y(new_n14940));
  not_8  g12592(.A(new_n14940), .Y(new_n14941));
  xnor_4 g12593(.A(new_n14881), .B(new_n14873), .Y(new_n14942));
  nor_5  g12594(.A(new_n14942), .B(new_n14941), .Y(new_n14943));
  not_8  g12595(.A(new_n14942), .Y(new_n14944_1));
  xnor_4 g12596(.A(new_n14944_1), .B(new_n14940), .Y(new_n14945));
  nor_5  g12597(.A(new_n14924), .B(new_n14911), .Y(new_n14946));
  xnor_4 g12598(.A(new_n14946), .B(new_n14909), .Y(new_n14947));
  not_8  g12599(.A(new_n14947), .Y(new_n14948));
  xnor_4 g12600(.A(new_n14879), .B(new_n14876), .Y(new_n14949));
  nor_5  g12601(.A(new_n14949), .B(new_n14948), .Y(new_n14950));
  nor_5  g12602(.A(new_n14921), .B(new_n14913), .Y(new_n14951));
  xnor_4 g12603(.A(new_n14923), .B(new_n14951), .Y(new_n14952));
  not_8  g12604(.A(new_n14952), .Y(new_n14953));
  nor_5  g12605(.A(new_n14953), .B(new_n13356), .Y(new_n14954_1));
  xnor_4 g12606(.A(new_n14952), .B(new_n13356), .Y(new_n14955));
  xor_4  g12607(.A(new_n14920), .B(new_n14914), .Y(new_n14956));
  nor_5  g12608(.A(new_n14956), .B(new_n13372), .Y(new_n14957));
  xor_4  g12609(.A(new_n14956), .B(new_n13372), .Y(new_n14958));
  nor_5  g12610(.A(new_n2629), .B(new_n2582_1), .Y(new_n14959));
  xnor_4 g12611(.A(new_n14918), .B(new_n14959), .Y(new_n14960));
  and_5  g12612(.A(new_n14960), .B(new_n13385), .Y(new_n14961));
  not_8  g12613(.A(new_n14743), .Y(new_n14962));
  nor_5  g12614(.A(new_n14962), .B(new_n13377), .Y(new_n14963));
  xnor_4 g12615(.A(new_n14960), .B(new_n13385), .Y(new_n14964));
  nor_5  g12616(.A(new_n14964), .B(new_n14963), .Y(new_n14965));
  nor_5  g12617(.A(new_n14965), .B(new_n14961), .Y(new_n14966));
  and_5  g12618(.A(new_n14966), .B(new_n14958), .Y(new_n14967));
  nor_5  g12619(.A(new_n14967), .B(new_n14957), .Y(new_n14968));
  and_5  g12620(.A(new_n14968), .B(new_n14955), .Y(new_n14969));
  nor_5  g12621(.A(new_n14969), .B(new_n14954_1), .Y(new_n14970));
  not_8  g12622(.A(new_n14949), .Y(new_n14971));
  xnor_4 g12623(.A(new_n14971), .B(new_n14947), .Y(new_n14972));
  nor_5  g12624(.A(new_n14972), .B(new_n14970), .Y(new_n14973));
  nor_5  g12625(.A(new_n14973), .B(new_n14950), .Y(new_n14974));
  nor_5  g12626(.A(new_n14974), .B(new_n14945), .Y(new_n14975));
  nor_5  g12627(.A(new_n14975), .B(new_n14943), .Y(new_n14976));
  xnor_4 g12628(.A(new_n14937), .B(new_n14936), .Y(new_n14977_1));
  nor_5  g12629(.A(new_n14977_1), .B(new_n14976), .Y(new_n14978));
  nor_5  g12630(.A(new_n14978), .B(new_n14938), .Y(new_n14979));
  xnor_4 g12631(.A(new_n14979), .B(new_n14933), .Y(n3263));
  xnor_4 g12632(.A(new_n12091), .B(new_n12078), .Y(n3289));
  xnor_4 g12633(.A(n21832), .B(new_n8968), .Y(new_n14982));
  nor_5  g12634(.A(new_n2356), .B(new_n8971_1), .Y(new_n14983));
  or_5   g12635(.A(n26913), .B(n12956), .Y(new_n14984));
  nor_5  g12636(.A(n18295), .B(n16223), .Y(new_n14985));
  or_5   g12637(.A(new_n5035), .B(new_n5031_1), .Y(new_n14986));
  and_5  g12638(.A(new_n14986), .B(new_n5030), .Y(new_n14987));
  nor_5  g12639(.A(new_n14987), .B(new_n14985), .Y(new_n14988));
  and_5  g12640(.A(new_n14988), .B(new_n14984), .Y(new_n14989_1));
  nor_5  g12641(.A(new_n14989_1), .B(new_n14983), .Y(new_n14990));
  xor_4  g12642(.A(new_n14990), .B(new_n14982), .Y(new_n14991));
  xnor_4 g12643(.A(new_n14991), .B(new_n8506), .Y(new_n14992));
  xnor_4 g12644(.A(n26913), .B(new_n8971_1), .Y(new_n14993));
  xnor_4 g12645(.A(new_n14993), .B(new_n14988), .Y(new_n14994));
  nor_5  g12646(.A(new_n14994), .B(n7057), .Y(new_n14995));
  not_8  g12647(.A(new_n14994), .Y(new_n14996));
  xnor_4 g12648(.A(new_n14996), .B(n7057), .Y(new_n14997));
  nor_5  g12649(.A(new_n5037), .B(n8381), .Y(new_n14998));
  or_5   g12650(.A(new_n5049), .B(new_n5044), .Y(new_n14999));
  and_5  g12651(.A(new_n14999), .B(new_n5039), .Y(new_n15000));
  or_5   g12652(.A(new_n15000), .B(new_n14998), .Y(new_n15001));
  and_5  g12653(.A(new_n15001), .B(new_n14997), .Y(new_n15002_1));
  nor_5  g12654(.A(new_n15002_1), .B(new_n14995), .Y(new_n15003));
  xnor_4 g12655(.A(new_n15003), .B(new_n14992), .Y(new_n15004_1));
  not_8  g12656(.A(new_n15004_1), .Y(new_n15005));
  xnor_4 g12657(.A(new_n14048), .B(n21649), .Y(new_n15006));
  nor_5  g12658(.A(new_n9409), .B(n18274), .Y(new_n15007));
  xnor_4 g12659(.A(new_n14050), .B(n18274), .Y(new_n15008));
  nor_5  g12660(.A(new_n9427), .B(n3828), .Y(new_n15009));
  nor_5  g12661(.A(new_n14057), .B(n23842), .Y(new_n15010));
  not_8  g12662(.A(n21654), .Y(new_n15011_1));
  or_5   g12663(.A(new_n9434), .B(new_n15011_1), .Y(new_n15012));
  xnor_4 g12664(.A(new_n14057), .B(new_n5172), .Y(new_n15013));
  and_5  g12665(.A(new_n15013), .B(new_n15012), .Y(new_n15014));
  or_5   g12666(.A(new_n15014), .B(new_n15010), .Y(new_n15015));
  xnor_4 g12667(.A(new_n9428), .B(n3828), .Y(new_n15016));
  and_5  g12668(.A(new_n15016), .B(new_n15015), .Y(new_n15017));
  or_5   g12669(.A(new_n15017), .B(new_n15009), .Y(new_n15018));
  and_5  g12670(.A(new_n15018), .B(new_n15008), .Y(new_n15019_1));
  nor_5  g12671(.A(new_n15019_1), .B(new_n15007), .Y(new_n15020));
  xor_4  g12672(.A(new_n15020), .B(new_n15006), .Y(new_n15021));
  xnor_4 g12673(.A(new_n15021), .B(new_n15005), .Y(new_n15022));
  nor_5  g12674(.A(new_n15000), .B(new_n14998), .Y(new_n15023));
  xnor_4 g12675(.A(new_n15023), .B(new_n14997), .Y(new_n15024));
  xor_4  g12676(.A(new_n15018), .B(new_n15008), .Y(new_n15025));
  and_5  g12677(.A(new_n15025), .B(new_n15024), .Y(new_n15026));
  xnor_4 g12678(.A(new_n15025), .B(new_n15024), .Y(new_n15027));
  xor_4  g12679(.A(new_n15016), .B(new_n15015), .Y(new_n15028));
  and_5  g12680(.A(new_n15028), .B(new_n5051), .Y(new_n15029));
  xor_4  g12681(.A(new_n15013), .B(new_n15012), .Y(new_n15030));
  and_5  g12682(.A(new_n15030), .B(new_n5077_1), .Y(new_n15031_1));
  xnor_4 g12683(.A(new_n9434), .B(n21654), .Y(new_n15032));
  not_8  g12684(.A(new_n15032), .Y(new_n15033_1));
  nor_5  g12685(.A(new_n15033_1), .B(new_n5081), .Y(new_n15034));
  xnor_4 g12686(.A(new_n15030), .B(new_n5077_1), .Y(new_n15035));
  nor_5  g12687(.A(new_n15035), .B(new_n15034), .Y(new_n15036));
  nor_5  g12688(.A(new_n15036), .B(new_n15031_1), .Y(new_n15037));
  xnor_4 g12689(.A(new_n15028), .B(new_n5051), .Y(new_n15038));
  nor_5  g12690(.A(new_n15038), .B(new_n15037), .Y(new_n15039));
  nor_5  g12691(.A(new_n15039), .B(new_n15029), .Y(new_n15040));
  nor_5  g12692(.A(new_n15040), .B(new_n15027), .Y(new_n15041));
  nor_5  g12693(.A(new_n15041), .B(new_n15026), .Y(new_n15042));
  xnor_4 g12694(.A(new_n15042), .B(new_n15022), .Y(n3301));
  xnor_4 g12695(.A(new_n10639), .B(n3030), .Y(new_n15044));
  not_8  g12696(.A(n19515), .Y(new_n15045));
  nor_5  g12697(.A(new_n10629), .B(new_n15045), .Y(new_n15046));
  xnor_4 g12698(.A(new_n10630), .B(new_n15045), .Y(new_n15047));
  nor_5  g12699(.A(new_n10619), .B(new_n13358), .Y(new_n15048));
  xnor_4 g12700(.A(new_n10620), .B(new_n13358), .Y(new_n15049));
  nor_5  g12701(.A(new_n10611_1), .B(n12209), .Y(new_n15050));
  or_5   g12702(.A(new_n10607), .B(new_n13145), .Y(new_n15051));
  and_5  g12703(.A(new_n13148), .B(new_n15051), .Y(new_n15052_1));
  nor_5  g12704(.A(new_n15052_1), .B(new_n15050), .Y(new_n15053_1));
  and_5  g12705(.A(new_n15053_1), .B(new_n15049), .Y(new_n15054));
  or_5   g12706(.A(new_n15054), .B(new_n15048), .Y(new_n15055));
  and_5  g12707(.A(new_n15055), .B(new_n15047), .Y(new_n15056));
  nor_5  g12708(.A(new_n15056), .B(new_n15046), .Y(new_n15057));
  xnor_4 g12709(.A(new_n15057), .B(new_n15044), .Y(new_n15058));
  not_8  g12710(.A(new_n15058), .Y(new_n15059));
  xnor_4 g12711(.A(new_n15059), .B(new_n9943), .Y(new_n15060));
  nor_5  g12712(.A(new_n15054), .B(new_n15048), .Y(new_n15061));
  xnor_4 g12713(.A(new_n15061), .B(new_n15047), .Y(new_n15062));
  not_8  g12714(.A(new_n15062), .Y(new_n15063));
  nor_5  g12715(.A(new_n15063), .B(new_n9947), .Y(new_n15064));
  xnor_4 g12716(.A(new_n15062), .B(new_n9948), .Y(new_n15065));
  xnor_4 g12717(.A(new_n15053_1), .B(new_n15049), .Y(new_n15066));
  nor_5  g12718(.A(new_n15066), .B(new_n9952), .Y(new_n15067));
  not_8  g12719(.A(new_n15066), .Y(new_n15068));
  xnor_4 g12720(.A(new_n15068), .B(new_n9953), .Y(new_n15069));
  nor_5  g12721(.A(new_n13149), .B(new_n9965), .Y(new_n15070));
  and_5  g12722(.A(new_n13151), .B(new_n13144_1), .Y(new_n15071));
  nor_5  g12723(.A(new_n15071), .B(new_n15070), .Y(new_n15072));
  nor_5  g12724(.A(new_n15072), .B(new_n15069), .Y(new_n15073));
  nor_5  g12725(.A(new_n15073), .B(new_n15067), .Y(new_n15074));
  nor_5  g12726(.A(new_n15074), .B(new_n15065), .Y(new_n15075));
  nor_5  g12727(.A(new_n15075), .B(new_n15064), .Y(new_n15076));
  xor_4  g12728(.A(new_n15076), .B(new_n15060), .Y(n3316));
  xnor_4 g12729(.A(new_n13135), .B(new_n13123), .Y(n3332));
  nor_5  g12730(.A(new_n7961), .B(n17458), .Y(new_n15079));
  xnor_4 g12731(.A(new_n7961), .B(new_n10870), .Y(new_n15080));
  nor_5  g12732(.A(new_n7966), .B(n1222), .Y(new_n15081));
  xnor_4 g12733(.A(new_n7966), .B(new_n10873), .Y(new_n15082_1));
  nor_5  g12734(.A(new_n7971), .B(n25240), .Y(new_n15083));
  nor_5  g12735(.A(new_n10429), .B(new_n10412), .Y(new_n15084));
  or_5   g12736(.A(new_n15084), .B(new_n15083), .Y(new_n15085));
  and_5  g12737(.A(new_n15085), .B(new_n15082_1), .Y(new_n15086));
  or_5   g12738(.A(new_n15086), .B(new_n15081), .Y(new_n15087));
  and_5  g12739(.A(new_n15087), .B(new_n15080), .Y(new_n15088));
  nor_5  g12740(.A(new_n15088), .B(new_n15079), .Y(new_n15089));
  and_5  g12741(.A(new_n15089), .B(new_n8026), .Y(new_n15090));
  nor_5  g12742(.A(new_n12681), .B(new_n14547_1), .Y(new_n15091));
  and_5  g12743(.A(new_n12693), .B(new_n12682), .Y(new_n15092));
  nor_5  g12744(.A(new_n15092), .B(new_n15091), .Y(new_n15093));
  nor_5  g12745(.A(n23166), .B(n11898), .Y(new_n15094_1));
  and_5  g12746(.A(new_n12680), .B(new_n12672), .Y(new_n15095));
  or_5   g12747(.A(new_n15095), .B(new_n15094_1), .Y(new_n15096));
  nor_5  g12748(.A(new_n15096), .B(new_n15093), .Y(new_n15097));
  not_8  g12749(.A(new_n15097), .Y(new_n15098));
  xnor_4 g12750(.A(new_n15098), .B(new_n15090), .Y(new_n15099));
  xnor_4 g12751(.A(new_n15089), .B(new_n8027_1), .Y(new_n15100));
  xnor_4 g12752(.A(new_n15096), .B(new_n15093), .Y(new_n15101));
  nor_5  g12753(.A(new_n15101), .B(new_n15100), .Y(new_n15102));
  xnor_4 g12754(.A(new_n15101), .B(new_n15100), .Y(new_n15103));
  not_8  g12755(.A(new_n15103), .Y(new_n15104));
  xor_4  g12756(.A(new_n15087), .B(new_n15080), .Y(new_n15105));
  nor_5  g12757(.A(new_n15105), .B(new_n12694), .Y(new_n15106));
  xor_4  g12758(.A(new_n15105), .B(new_n12694), .Y(new_n15107));
  xor_4  g12759(.A(new_n15085), .B(new_n15082_1), .Y(new_n15108));
  and_5  g12760(.A(new_n15108), .B(new_n12699), .Y(new_n15109));
  nor_5  g12761(.A(new_n10477), .B(new_n10430), .Y(new_n15110));
  nor_5  g12762(.A(new_n10503), .B(new_n10478), .Y(new_n15111));
  nor_5  g12763(.A(new_n15111), .B(new_n15110), .Y(new_n15112));
  xnor_4 g12764(.A(new_n15108), .B(new_n12699), .Y(new_n15113));
  nor_5  g12765(.A(new_n15113), .B(new_n15112), .Y(new_n15114));
  nor_5  g12766(.A(new_n15114), .B(new_n15109), .Y(new_n15115));
  and_5  g12767(.A(new_n15115), .B(new_n15107), .Y(new_n15116));
  nor_5  g12768(.A(new_n15116), .B(new_n15106), .Y(new_n15117));
  and_5  g12769(.A(new_n15117), .B(new_n15104), .Y(new_n15118_1));
  nor_5  g12770(.A(new_n15118_1), .B(new_n15102), .Y(new_n15119));
  xnor_4 g12771(.A(new_n15119), .B(new_n15099), .Y(n3340));
  xnor_4 g12772(.A(n13851), .B(n5077), .Y(new_n15121));
  nor_5  g12773(.A(n24937), .B(new_n10452), .Y(new_n15122));
  xnor_4 g12774(.A(n24937), .B(n15546), .Y(new_n15123));
  not_8  g12775(.A(n5098), .Y(new_n15124));
  and_5  g12776(.A(n26452), .B(new_n15124), .Y(new_n15125));
  xnor_4 g12777(.A(n26452), .B(n5098), .Y(new_n15126));
  nor_5  g12778(.A(new_n10460), .B(n3030), .Y(new_n15127));
  xnor_4 g12779(.A(n19905), .B(n3030), .Y(new_n15128_1));
  nor_5  g12780(.A(new_n15045), .B(n17035), .Y(new_n15129));
  or_5   g12781(.A(new_n13367_1), .B(new_n13359), .Y(new_n15130));
  and_5  g12782(.A(new_n15130), .B(new_n13357), .Y(new_n15131));
  nor_5  g12783(.A(new_n15131), .B(new_n15129), .Y(new_n15132));
  and_5  g12784(.A(new_n15132), .B(new_n15128_1), .Y(new_n15133));
  or_5   g12785(.A(new_n15133), .B(new_n15127), .Y(new_n15134));
  and_5  g12786(.A(new_n15134), .B(new_n15126), .Y(new_n15135));
  or_5   g12787(.A(new_n15135), .B(new_n15125), .Y(new_n15136));
  and_5  g12788(.A(new_n15136), .B(new_n15123), .Y(new_n15137));
  or_5   g12789(.A(new_n15137), .B(new_n15122), .Y(new_n15138));
  xor_4  g12790(.A(new_n15138), .B(new_n15121), .Y(new_n15139_1));
  xnor_4 g12791(.A(new_n15139_1), .B(new_n14887), .Y(new_n15140));
  xor_4  g12792(.A(new_n15136), .B(new_n15123), .Y(new_n15141));
  nor_5  g12793(.A(new_n15141), .B(new_n14937), .Y(new_n15142));
  xnor_4 g12794(.A(new_n15141), .B(new_n14937), .Y(new_n15143));
  xor_4  g12795(.A(new_n15134), .B(new_n15126), .Y(new_n15144));
  nor_5  g12796(.A(new_n15144), .B(new_n14942), .Y(new_n15145_1));
  xnor_4 g12797(.A(new_n15144), .B(new_n14944_1), .Y(new_n15146_1));
  xnor_4 g12798(.A(new_n15132), .B(new_n15128_1), .Y(new_n15147));
  nor_5  g12799(.A(new_n15147), .B(new_n14971), .Y(new_n15148));
  not_8  g12800(.A(new_n15147), .Y(new_n15149));
  xnor_4 g12801(.A(new_n15149), .B(new_n14971), .Y(new_n15150));
  nor_5  g12802(.A(new_n13370), .B(new_n13356), .Y(new_n15151));
  nor_5  g12803(.A(new_n13390), .B(new_n13371), .Y(new_n15152));
  nor_5  g12804(.A(new_n15152), .B(new_n15151), .Y(new_n15153));
  and_5  g12805(.A(new_n15153), .B(new_n15150), .Y(new_n15154));
  nor_5  g12806(.A(new_n15154), .B(new_n15148), .Y(new_n15155));
  and_5  g12807(.A(new_n15155), .B(new_n15146_1), .Y(new_n15156));
  nor_5  g12808(.A(new_n15156), .B(new_n15145_1), .Y(new_n15157));
  nor_5  g12809(.A(new_n15157), .B(new_n15143), .Y(new_n15158));
  nor_5  g12810(.A(new_n15158), .B(new_n15142), .Y(new_n15159));
  xor_4  g12811(.A(new_n15159), .B(new_n15140), .Y(n3343));
  not_8  g12812(.A(new_n14898), .Y(new_n15161));
  nor_5  g12813(.A(new_n15161), .B(n19270), .Y(new_n15162));
  not_8  g12814(.A(new_n15162), .Y(new_n15163));
  nor_5  g12815(.A(new_n15163), .B(n14704), .Y(new_n15164));
  and_5  g12816(.A(new_n15164), .B(new_n14347), .Y(new_n15165_1));
  xnor_4 g12817(.A(new_n15164), .B(n25365), .Y(new_n15166));
  nor_5  g12818(.A(new_n15166), .B(n20040), .Y(new_n15167_1));
  xnor_4 g12819(.A(new_n15162), .B(n14704), .Y(new_n15168));
  nor_5  g12820(.A(new_n15168), .B(n19531), .Y(new_n15169));
  xnor_4 g12821(.A(new_n15168), .B(new_n2558), .Y(new_n15170));
  nor_5  g12822(.A(new_n14899_1), .B(n18345), .Y(new_n15171));
  or_5   g12823(.A(new_n14930), .B(new_n14902), .Y(new_n15172));
  and_5  g12824(.A(new_n15172), .B(new_n14900), .Y(new_n15173));
  or_5   g12825(.A(new_n15173), .B(new_n15171), .Y(new_n15174));
  and_5  g12826(.A(new_n15174), .B(new_n15170), .Y(new_n15175));
  nor_5  g12827(.A(new_n15175), .B(new_n15169), .Y(new_n15176_1));
  and_5  g12828(.A(new_n15166), .B(n20040), .Y(new_n15177));
  nor_5  g12829(.A(new_n15177), .B(new_n15176_1), .Y(new_n15178));
  nor_5  g12830(.A(new_n15178), .B(new_n15167_1), .Y(new_n15179));
  nor_5  g12831(.A(new_n15179), .B(new_n15165_1), .Y(new_n15180_1));
  xnor_4 g12832(.A(new_n15166), .B(new_n11289), .Y(new_n15181));
  xnor_4 g12833(.A(new_n15181), .B(new_n15176_1), .Y(new_n15182_1));
  nor_5  g12834(.A(new_n15182_1), .B(new_n13702), .Y(new_n15183));
  not_8  g12835(.A(new_n15182_1), .Y(new_n15184));
  nor_5  g12836(.A(new_n15184), .B(new_n13701), .Y(new_n15185));
  nor_5  g12837(.A(new_n15173), .B(new_n15171), .Y(new_n15186));
  xnor_4 g12838(.A(new_n15186), .B(new_n15170), .Y(new_n15187));
  nor_5  g12839(.A(new_n15187), .B(new_n13685), .Y(new_n15188));
  not_8  g12840(.A(new_n15187), .Y(new_n15189));
  xnor_4 g12841(.A(new_n15189), .B(new_n13685), .Y(new_n15190));
  nor_5  g12842(.A(new_n14932), .B(new_n13688), .Y(new_n15191));
  not_8  g12843(.A(new_n14932), .Y(new_n15192));
  xnor_4 g12844(.A(new_n15192), .B(new_n13688), .Y(new_n15193));
  nor_5  g12845(.A(new_n14935), .B(new_n6472), .Y(new_n15194));
  xnor_4 g12846(.A(new_n14936), .B(new_n6472), .Y(new_n15195));
  nor_5  g12847(.A(new_n14940), .B(new_n6476_1), .Y(new_n15196));
  nor_5  g12848(.A(new_n14947), .B(new_n6480), .Y(new_n15197));
  xnor_4 g12849(.A(new_n14948), .B(new_n6480), .Y(new_n15198));
  nor_5  g12850(.A(new_n14953), .B(new_n6482), .Y(new_n15199));
  xnor_4 g12851(.A(new_n14953), .B(new_n6499), .Y(new_n15200));
  nor_5  g12852(.A(new_n14956), .B(new_n6486), .Y(new_n15201));
  xnor_4 g12853(.A(new_n14956), .B(new_n6484), .Y(new_n15202));
  not_8  g12854(.A(new_n14960), .Y(new_n15203));
  nor_5  g12855(.A(new_n15203), .B(new_n6489), .Y(new_n15204));
  or_5   g12856(.A(new_n14962), .B(new_n6491), .Y(new_n15205_1));
  xnor_4 g12857(.A(new_n15203), .B(new_n6488), .Y(new_n15206));
  and_5  g12858(.A(new_n15206), .B(new_n15205_1), .Y(new_n15207));
  nor_5  g12859(.A(new_n15207), .B(new_n15204), .Y(new_n15208));
  and_5  g12860(.A(new_n15208), .B(new_n15202), .Y(new_n15209));
  nor_5  g12861(.A(new_n15209), .B(new_n15201), .Y(new_n15210));
  and_5  g12862(.A(new_n15210), .B(new_n15200), .Y(new_n15211));
  nor_5  g12863(.A(new_n15211), .B(new_n15199), .Y(new_n15212));
  and_5  g12864(.A(new_n15212), .B(new_n15198), .Y(new_n15213));
  or_5   g12865(.A(new_n15213), .B(new_n15197), .Y(new_n15214));
  xnor_4 g12866(.A(new_n14941), .B(new_n6476_1), .Y(new_n15215));
  and_5  g12867(.A(new_n15215), .B(new_n15214), .Y(new_n15216));
  or_5   g12868(.A(new_n15216), .B(new_n15196), .Y(new_n15217));
  and_5  g12869(.A(new_n15217), .B(new_n15195), .Y(new_n15218));
  or_5   g12870(.A(new_n15218), .B(new_n15194), .Y(new_n15219));
  and_5  g12871(.A(new_n15219), .B(new_n15193), .Y(new_n15220));
  or_5   g12872(.A(new_n15220), .B(new_n15191), .Y(new_n15221));
  and_5  g12873(.A(new_n15221), .B(new_n15190), .Y(new_n15222));
  nor_5  g12874(.A(new_n15222), .B(new_n15188), .Y(new_n15223));
  nor_5  g12875(.A(new_n15223), .B(new_n15185), .Y(new_n15224));
  or_5   g12876(.A(new_n15224), .B(new_n13724), .Y(new_n15225));
  or_5   g12877(.A(new_n15225), .B(new_n15183), .Y(new_n15226));
  xnor_4 g12878(.A(new_n15226), .B(new_n15180_1), .Y(new_n15227));
  and_5  g12879(.A(new_n12251), .B(new_n11795), .Y(new_n15228));
  xnor_4 g12880(.A(new_n12251), .B(new_n11795), .Y(new_n15229));
  and_5  g12881(.A(new_n12255), .B(new_n6155), .Y(new_n15230_1));
  xnor_4 g12882(.A(new_n12255), .B(new_n6155), .Y(new_n15231));
  and_5  g12883(.A(new_n12259), .B(new_n6158), .Y(new_n15232));
  xnor_4 g12884(.A(new_n12259), .B(new_n6158), .Y(new_n15233));
  and_5  g12885(.A(new_n12263), .B(new_n6161), .Y(new_n15234));
  xnor_4 g12886(.A(new_n12263), .B(new_n6161), .Y(new_n15235));
  and_5  g12887(.A(new_n12267), .B(new_n11812), .Y(new_n15236));
  xnor_4 g12888(.A(new_n12267), .B(new_n11812), .Y(new_n15237));
  not_8  g12889(.A(n21226), .Y(new_n15238));
  and_5  g12890(.A(new_n12271), .B(new_n15238), .Y(new_n15239));
  xnor_4 g12891(.A(new_n12271), .B(new_n15238), .Y(new_n15240));
  nor_5  g12892(.A(new_n12275), .B(n4426), .Y(new_n15241_1));
  xnor_4 g12893(.A(new_n12275), .B(new_n6170), .Y(new_n15242));
  nor_5  g12894(.A(new_n12282), .B(n20036), .Y(new_n15243));
  xnor_4 g12895(.A(new_n12282), .B(new_n8659), .Y(new_n15244));
  nor_5  g12896(.A(new_n12291), .B(new_n4120), .Y(new_n15245));
  or_5   g12897(.A(new_n12287), .B(n9380), .Y(new_n15246));
  xnor_4 g12898(.A(new_n12290), .B(new_n4120), .Y(new_n15247));
  and_5  g12899(.A(new_n15247), .B(new_n15246), .Y(new_n15248));
  nor_5  g12900(.A(new_n15248), .B(new_n15245), .Y(new_n15249));
  and_5  g12901(.A(new_n15249), .B(new_n15244), .Y(new_n15250));
  or_5   g12902(.A(new_n15250), .B(new_n15243), .Y(new_n15251));
  and_5  g12903(.A(new_n15251), .B(new_n15242), .Y(new_n15252));
  nor_5  g12904(.A(new_n15252), .B(new_n15241_1), .Y(new_n15253));
  nor_5  g12905(.A(new_n15253), .B(new_n15240), .Y(new_n15254));
  nor_5  g12906(.A(new_n15254), .B(new_n15239), .Y(new_n15255_1));
  nor_5  g12907(.A(new_n15255_1), .B(new_n15237), .Y(new_n15256));
  nor_5  g12908(.A(new_n15256), .B(new_n15236), .Y(new_n15257));
  nor_5  g12909(.A(new_n15257), .B(new_n15235), .Y(new_n15258_1));
  nor_5  g12910(.A(new_n15258_1), .B(new_n15234), .Y(new_n15259));
  nor_5  g12911(.A(new_n15259), .B(new_n15233), .Y(new_n15260));
  nor_5  g12912(.A(new_n15260), .B(new_n15232), .Y(new_n15261));
  nor_5  g12913(.A(new_n15261), .B(new_n15231), .Y(new_n15262));
  nor_5  g12914(.A(new_n15262), .B(new_n15230_1), .Y(new_n15263));
  nor_5  g12915(.A(new_n15263), .B(new_n15229), .Y(new_n15264));
  nor_5  g12916(.A(new_n15264), .B(new_n15228), .Y(new_n15265));
  xnor_4 g12917(.A(new_n15265), .B(new_n12156), .Y(new_n15266));
  nor_5  g12918(.A(new_n15266), .B(new_n15227), .Y(new_n15267));
  xnor_4 g12919(.A(new_n15263), .B(new_n15229), .Y(new_n15268));
  xnor_4 g12920(.A(new_n15184), .B(new_n13702), .Y(new_n15269));
  xnor_4 g12921(.A(new_n15269), .B(new_n15223), .Y(new_n15270));
  nor_5  g12922(.A(new_n15270), .B(new_n15268), .Y(new_n15271_1));
  xnor_4 g12923(.A(new_n15270), .B(new_n15268), .Y(new_n15272));
  xnor_4 g12924(.A(new_n15261), .B(new_n15231), .Y(new_n15273));
  xor_4  g12925(.A(new_n15221), .B(new_n15190), .Y(new_n15274));
  nor_5  g12926(.A(new_n15274), .B(new_n15273), .Y(new_n15275_1));
  xnor_4 g12927(.A(new_n15274), .B(new_n15273), .Y(new_n15276));
  xnor_4 g12928(.A(new_n15259), .B(new_n15233), .Y(new_n15277));
  xor_4  g12929(.A(new_n15219), .B(new_n15193), .Y(new_n15278));
  nor_5  g12930(.A(new_n15278), .B(new_n15277), .Y(new_n15279));
  xnor_4 g12931(.A(new_n15278), .B(new_n15277), .Y(new_n15280));
  xnor_4 g12932(.A(new_n15257), .B(new_n15235), .Y(new_n15281));
  xor_4  g12933(.A(new_n15217), .B(new_n15195), .Y(new_n15282));
  nor_5  g12934(.A(new_n15282), .B(new_n15281), .Y(new_n15283));
  xnor_4 g12935(.A(new_n15282), .B(new_n15281), .Y(new_n15284));
  xnor_4 g12936(.A(new_n15255_1), .B(new_n15237), .Y(new_n15285));
  xor_4  g12937(.A(new_n15215), .B(new_n15214), .Y(new_n15286));
  nor_5  g12938(.A(new_n15286), .B(new_n15285), .Y(new_n15287));
  xnor_4 g12939(.A(new_n15286), .B(new_n15285), .Y(new_n15288));
  xnor_4 g12940(.A(new_n15253), .B(new_n15240), .Y(new_n15289_1));
  xnor_4 g12941(.A(new_n15212), .B(new_n15198), .Y(new_n15290));
  not_8  g12942(.A(new_n15290), .Y(new_n15291));
  nor_5  g12943(.A(new_n15291), .B(new_n15289_1), .Y(new_n15292));
  xnor_4 g12944(.A(new_n15291), .B(new_n15289_1), .Y(new_n15293));
  xor_4  g12945(.A(new_n15251), .B(new_n15242), .Y(new_n15294));
  xnor_4 g12946(.A(new_n15210), .B(new_n15200), .Y(new_n15295));
  not_8  g12947(.A(new_n15295), .Y(new_n15296));
  and_5  g12948(.A(new_n15296), .B(new_n15294), .Y(new_n15297));
  xnor_4 g12949(.A(new_n15296), .B(new_n15294), .Y(new_n15298));
  xnor_4 g12950(.A(new_n15249), .B(new_n15244), .Y(new_n15299));
  xnor_4 g12951(.A(new_n15208), .B(new_n15202), .Y(new_n15300_1));
  not_8  g12952(.A(new_n15300_1), .Y(new_n15301));
  nor_5  g12953(.A(new_n15301), .B(new_n15299), .Y(new_n15302));
  nor_5  g12954(.A(new_n14962), .B(new_n6491), .Y(new_n15303));
  xnor_4 g12955(.A(new_n15206), .B(new_n15303), .Y(new_n15304));
  not_8  g12956(.A(new_n15304), .Y(new_n15305));
  xor_4  g12957(.A(new_n15247), .B(new_n15246), .Y(new_n15306));
  and_5  g12958(.A(new_n15306), .B(new_n15305), .Y(new_n15307_1));
  xnor_4 g12959(.A(new_n14962), .B(n4939), .Y(new_n15308));
  not_8  g12960(.A(new_n15308), .Y(new_n15309));
  xnor_4 g12961(.A(new_n12287), .B(new_n6176), .Y(new_n15310));
  nor_5  g12962(.A(new_n15310), .B(new_n15309), .Y(new_n15311));
  xnor_4 g12963(.A(new_n15306), .B(new_n15304), .Y(new_n15312));
  and_5  g12964(.A(new_n15312), .B(new_n15311), .Y(new_n15313));
  nor_5  g12965(.A(new_n15313), .B(new_n15307_1), .Y(new_n15314));
  xnor_4 g12966(.A(new_n15300_1), .B(new_n15299), .Y(new_n15315));
  and_5  g12967(.A(new_n15315), .B(new_n15314), .Y(new_n15316));
  nor_5  g12968(.A(new_n15316), .B(new_n15302), .Y(new_n15317));
  nor_5  g12969(.A(new_n15317), .B(new_n15298), .Y(new_n15318));
  nor_5  g12970(.A(new_n15318), .B(new_n15297), .Y(new_n15319));
  nor_5  g12971(.A(new_n15319), .B(new_n15293), .Y(new_n15320));
  nor_5  g12972(.A(new_n15320), .B(new_n15292), .Y(new_n15321));
  nor_5  g12973(.A(new_n15321), .B(new_n15288), .Y(new_n15322));
  nor_5  g12974(.A(new_n15322), .B(new_n15287), .Y(new_n15323));
  nor_5  g12975(.A(new_n15323), .B(new_n15284), .Y(new_n15324));
  nor_5  g12976(.A(new_n15324), .B(new_n15283), .Y(new_n15325));
  nor_5  g12977(.A(new_n15325), .B(new_n15280), .Y(new_n15326));
  nor_5  g12978(.A(new_n15326), .B(new_n15279), .Y(new_n15327_1));
  nor_5  g12979(.A(new_n15327_1), .B(new_n15276), .Y(new_n15328));
  nor_5  g12980(.A(new_n15328), .B(new_n15275_1), .Y(new_n15329));
  nor_5  g12981(.A(new_n15329), .B(new_n15272), .Y(new_n15330));
  nor_5  g12982(.A(new_n15330), .B(new_n15271_1), .Y(new_n15331));
  xnor_4 g12983(.A(new_n15266), .B(new_n15227), .Y(new_n15332_1));
  nor_5  g12984(.A(new_n15332_1), .B(new_n15331), .Y(new_n15333));
  nor_5  g12985(.A(new_n15333), .B(new_n15267), .Y(new_n15334));
  nor_5  g12986(.A(new_n15226), .B(new_n15180_1), .Y(new_n15335));
  or_5   g12987(.A(new_n12155), .B(new_n12111), .Y(new_n15336));
  and_5  g12988(.A(new_n15265), .B(new_n15336), .Y(new_n15337));
  xor_4  g12989(.A(new_n15337), .B(new_n15335), .Y(new_n15338));
  xnor_4 g12990(.A(new_n15338), .B(new_n15334), .Y(n3390));
  xnor_4 g12991(.A(new_n6573), .B(new_n6572), .Y(n3426));
  not_8  g12992(.A(new_n4740), .Y(new_n15341));
  xnor_4 g12993(.A(new_n15341), .B(new_n4739), .Y(n3451));
  xnor_4 g12994(.A(new_n12008), .B(new_n11991), .Y(n3459));
  xnor_4 g12995(.A(n6773), .B(new_n5587), .Y(new_n15344));
  xnor_4 g12996(.A(new_n15344), .B(n21687), .Y(new_n15345_1));
  nor_5  g12997(.A(new_n15345_1), .B(new_n13471), .Y(new_n15346));
  nor_5  g12998(.A(new_n15344), .B(new_n2548), .Y(new_n15347));
  nor_5  g12999(.A(new_n15347), .B(n6729), .Y(new_n15348));
  or_5   g13000(.A(new_n2548), .B(new_n6178), .Y(new_n15349));
  nor_5  g13001(.A(new_n15344), .B(new_n15349), .Y(new_n15350));
  nor_5  g13002(.A(new_n15350), .B(new_n15348), .Y(new_n15351));
  nor_5  g13003(.A(new_n4030), .B(new_n5587), .Y(new_n15352));
  xnor_4 g13004(.A(n22173), .B(n17090), .Y(new_n15353_1));
  xor_4  g13005(.A(new_n15353_1), .B(new_n15352), .Y(new_n15354));
  xnor_4 g13006(.A(new_n15354), .B(new_n15351), .Y(new_n15355));
  not_8  g13007(.A(new_n15355), .Y(new_n15356));
  xnor_4 g13008(.A(new_n15356), .B(new_n13466), .Y(new_n15357));
  xnor_4 g13009(.A(new_n15357), .B(new_n15346), .Y(n3502));
  xnor_4 g13010(.A(new_n10771), .B(new_n10738), .Y(n3516));
  nor_5  g13011(.A(n24129), .B(n22274), .Y(new_n15360));
  not_8  g13012(.A(new_n15360), .Y(new_n15361));
  nor_5  g13013(.A(new_n15361), .B(n1689), .Y(new_n15362));
  not_8  g13014(.A(new_n15362), .Y(new_n15363));
  nor_5  g13015(.A(new_n15363), .B(n19608), .Y(new_n15364));
  not_8  g13016(.A(new_n15364), .Y(new_n15365));
  nor_5  g13017(.A(new_n15365), .B(n25126), .Y(new_n15366_1));
  not_8  g13018(.A(new_n15366_1), .Y(new_n15367));
  nor_5  g13019(.A(new_n15367), .B(n10712), .Y(new_n15368));
  xnor_4 g13020(.A(new_n15368), .B(n18145), .Y(new_n15369));
  xnor_4 g13021(.A(new_n15369), .B(n15761), .Y(new_n15370));
  xnor_4 g13022(.A(new_n15366_1), .B(n10712), .Y(new_n15371));
  nor_5  g13023(.A(new_n15371), .B(new_n10179), .Y(new_n15372));
  xnor_4 g13024(.A(new_n15371), .B(n11201), .Y(new_n15373));
  xnor_4 g13025(.A(new_n15364), .B(n25126), .Y(new_n15374));
  nor_5  g13026(.A(new_n15374), .B(new_n10182), .Y(new_n15375));
  xnor_4 g13027(.A(new_n15374), .B(n18690), .Y(new_n15376));
  xnor_4 g13028(.A(new_n15363), .B(n19608), .Y(new_n15377));
  and_5  g13029(.A(new_n15377), .B(n12153), .Y(new_n15378_1));
  xnor_4 g13030(.A(new_n15362), .B(n19608), .Y(new_n15379));
  xnor_4 g13031(.A(new_n15379), .B(n12153), .Y(new_n15380));
  xnor_4 g13032(.A(new_n15360), .B(n1689), .Y(new_n15381));
  nor_5  g13033(.A(new_n15381), .B(new_n10186), .Y(new_n15382_1));
  xnor_4 g13034(.A(new_n15381), .B(n13044), .Y(new_n15383));
  xnor_4 g13035(.A(n24129), .B(new_n4118), .Y(new_n15384));
  nor_5  g13036(.A(new_n15384), .B(new_n5807), .Y(new_n15385));
  nor_5  g13037(.A(n24129), .B(new_n5805), .Y(new_n15386));
  xnor_4 g13038(.A(new_n15384), .B(n18745), .Y(new_n15387));
  and_5  g13039(.A(new_n15387), .B(new_n15386), .Y(new_n15388));
  or_5   g13040(.A(new_n15388), .B(new_n15385), .Y(new_n15389));
  and_5  g13041(.A(new_n15389), .B(new_n15383), .Y(new_n15390));
  or_5   g13042(.A(new_n15390), .B(new_n15382_1), .Y(new_n15391));
  and_5  g13043(.A(new_n15391), .B(new_n15380), .Y(new_n15392));
  or_5   g13044(.A(new_n15392), .B(new_n15378_1), .Y(new_n15393));
  and_5  g13045(.A(new_n15393), .B(new_n15376), .Y(new_n15394));
  or_5   g13046(.A(new_n15394), .B(new_n15375), .Y(new_n15395));
  and_5  g13047(.A(new_n15395), .B(new_n15373), .Y(new_n15396));
  or_5   g13048(.A(new_n15396), .B(new_n15372), .Y(new_n15397));
  xor_4  g13049(.A(new_n15397), .B(new_n15370), .Y(new_n15398));
  xnor_4 g13050(.A(new_n15398), .B(new_n6874), .Y(new_n15399));
  xor_4  g13051(.A(new_n15395), .B(new_n15373), .Y(new_n15400));
  and_5  g13052(.A(new_n15400), .B(new_n6877), .Y(new_n15401));
  xnor_4 g13053(.A(new_n15400), .B(new_n6877), .Y(new_n15402));
  xor_4  g13054(.A(new_n15393), .B(new_n15376), .Y(new_n15403));
  and_5  g13055(.A(new_n15403), .B(new_n6882), .Y(new_n15404));
  xnor_4 g13056(.A(new_n15403), .B(new_n6882), .Y(new_n15405));
  xor_4  g13057(.A(new_n15391), .B(new_n15380), .Y(new_n15406));
  and_5  g13058(.A(new_n15406), .B(new_n6886), .Y(new_n15407_1));
  xnor_4 g13059(.A(new_n15406), .B(new_n6888), .Y(new_n15408));
  xor_4  g13060(.A(new_n15389), .B(new_n15383), .Y(new_n15409));
  nor_5  g13061(.A(new_n15409), .B(new_n4115), .Y(new_n15410));
  xnor_4 g13062(.A(new_n15409), .B(new_n4116), .Y(new_n15411));
  xor_4  g13063(.A(new_n15387), .B(new_n15386), .Y(new_n15412));
  nor_5  g13064(.A(new_n15412), .B(new_n4130), .Y(new_n15413));
  xnor_4 g13065(.A(n24129), .B(n16167), .Y(new_n15414));
  nor_5  g13066(.A(new_n15414), .B(new_n4135), .Y(new_n15415));
  xnor_4 g13067(.A(new_n15412), .B(new_n4138), .Y(new_n15416));
  and_5  g13068(.A(new_n15416), .B(new_n15415), .Y(new_n15417));
  or_5   g13069(.A(new_n15417), .B(new_n15413), .Y(new_n15418));
  and_5  g13070(.A(new_n15418), .B(new_n15411), .Y(new_n15419));
  nor_5  g13071(.A(new_n15419), .B(new_n15410), .Y(new_n15420));
  and_5  g13072(.A(new_n15420), .B(new_n15408), .Y(new_n15421));
  nor_5  g13073(.A(new_n15421), .B(new_n15407_1), .Y(new_n15422));
  nor_5  g13074(.A(new_n15422), .B(new_n15405), .Y(new_n15423));
  nor_5  g13075(.A(new_n15423), .B(new_n15404), .Y(new_n15424_1));
  nor_5  g13076(.A(new_n15424_1), .B(new_n15402), .Y(new_n15425));
  or_5   g13077(.A(new_n15425), .B(new_n15401), .Y(new_n15426));
  xor_4  g13078(.A(new_n15426), .B(new_n15399), .Y(new_n15427));
  xnor_4 g13079(.A(new_n15427), .B(new_n10305), .Y(new_n15428_1));
  xnor_4 g13080(.A(new_n15424_1), .B(new_n15402), .Y(new_n15429));
  nor_5  g13081(.A(new_n15429), .B(new_n10310), .Y(new_n15430));
  xnor_4 g13082(.A(new_n15429), .B(new_n10310), .Y(new_n15431));
  xnor_4 g13083(.A(new_n15422), .B(new_n15405), .Y(new_n15432));
  nor_5  g13084(.A(new_n15432), .B(new_n10314), .Y(new_n15433));
  xnor_4 g13085(.A(new_n15432), .B(new_n10314), .Y(new_n15434));
  xnor_4 g13086(.A(new_n15420), .B(new_n15408), .Y(new_n15435_1));
  nor_5  g13087(.A(new_n15435_1), .B(new_n10319), .Y(new_n15436));
  xor_4  g13088(.A(new_n15418), .B(new_n15411), .Y(new_n15437));
  nor_5  g13089(.A(new_n15437), .B(new_n10322), .Y(new_n15438_1));
  xnor_4 g13090(.A(new_n15437), .B(new_n10322), .Y(new_n15439));
  xor_4  g13091(.A(new_n15416), .B(new_n15415), .Y(new_n15440));
  nor_5  g13092(.A(new_n15440), .B(new_n5814), .Y(new_n15441));
  xnor_4 g13093(.A(new_n15414), .B(new_n4134_1), .Y(new_n15442));
  and_5  g13094(.A(new_n15442), .B(new_n5799), .Y(new_n15443));
  xnor_4 g13095(.A(new_n15440), .B(new_n5814), .Y(new_n15444));
  nor_5  g13096(.A(new_n15444), .B(new_n15443), .Y(new_n15445));
  nor_5  g13097(.A(new_n15445), .B(new_n15441), .Y(new_n15446));
  nor_5  g13098(.A(new_n15446), .B(new_n15439), .Y(new_n15447));
  nor_5  g13099(.A(new_n15447), .B(new_n15438_1), .Y(new_n15448));
  xnor_4 g13100(.A(new_n15435_1), .B(new_n10319), .Y(new_n15449));
  nor_5  g13101(.A(new_n15449), .B(new_n15448), .Y(new_n15450));
  nor_5  g13102(.A(new_n15450), .B(new_n15436), .Y(new_n15451));
  nor_5  g13103(.A(new_n15451), .B(new_n15434), .Y(new_n15452));
  nor_5  g13104(.A(new_n15452), .B(new_n15433), .Y(new_n15453));
  nor_5  g13105(.A(new_n15453), .B(new_n15431), .Y(new_n15454));
  nor_5  g13106(.A(new_n15454), .B(new_n15430), .Y(new_n15455));
  xor_4  g13107(.A(new_n15455), .B(new_n15428_1), .Y(n3528));
  xnor_4 g13108(.A(new_n9057), .B(new_n9001), .Y(n3555));
  nor_5  g13109(.A(new_n10052), .B(new_n2673), .Y(new_n15458));
  and_5  g13110(.A(new_n2782), .B(new_n2720), .Y(new_n15459));
  nor_5  g13111(.A(new_n15459), .B(new_n15458), .Y(new_n15460));
  not_8  g13112(.A(new_n15460), .Y(new_n15461));
  nor_5  g13113(.A(new_n2672), .B(n13951), .Y(new_n15462));
  and_5  g13114(.A(new_n10050), .B(new_n15462), .Y(new_n15463));
  and_5  g13115(.A(new_n15463), .B(new_n15461), .Y(new_n15464));
  or_5   g13116(.A(new_n10050), .B(new_n15462), .Y(new_n15465_1));
  nor_5  g13117(.A(new_n15465_1), .B(new_n15461), .Y(new_n15466));
  nor_5  g13118(.A(new_n15466), .B(new_n15464), .Y(new_n15467_1));
  nor_5  g13119(.A(new_n15467_1), .B(new_n14356), .Y(new_n15468));
  xnor_4 g13120(.A(new_n15467_1), .B(new_n14356), .Y(new_n15469));
  xnor_4 g13121(.A(new_n10049), .B(new_n15462), .Y(new_n15470_1));
  xnor_4 g13122(.A(new_n15470_1), .B(new_n15461), .Y(new_n15471));
  nor_5  g13123(.A(new_n15471), .B(new_n14361), .Y(new_n15472));
  xnor_4 g13124(.A(new_n15471), .B(new_n14361), .Y(new_n15473));
  nor_5  g13125(.A(new_n2783_1), .B(new_n2655), .Y(new_n15474));
  and_5  g13126(.A(new_n2847), .B(new_n2784), .Y(new_n15475));
  nor_5  g13127(.A(new_n15475), .B(new_n15474), .Y(new_n15476));
  nor_5  g13128(.A(new_n15476), .B(new_n15473), .Y(new_n15477_1));
  nor_5  g13129(.A(new_n15477_1), .B(new_n15472), .Y(new_n15478));
  nor_5  g13130(.A(new_n15478), .B(new_n15469), .Y(new_n15479));
  nor_5  g13131(.A(new_n15479), .B(new_n15468), .Y(new_n15480));
  nor_5  g13132(.A(new_n15480), .B(new_n15464), .Y(n3561));
  xnor_4 g13133(.A(n16439), .B(n14680), .Y(new_n15482));
  and_5  g13134(.A(n17250), .B(new_n4369), .Y(new_n15483));
  and_5  g13135(.A(new_n10525_1), .B(new_n10505), .Y(new_n15484));
  or_5   g13136(.A(new_n15484), .B(new_n15483), .Y(new_n15485));
  xor_4  g13137(.A(new_n15485), .B(new_n15482), .Y(new_n15486));
  xnor_4 g13138(.A(new_n9613), .B(new_n7613), .Y(new_n15487));
  not_8  g13139(.A(new_n15487), .Y(new_n15488));
  nor_5  g13140(.A(new_n9617), .B(n13783), .Y(new_n15489));
  nor_5  g13141(.A(new_n10540_1), .B(new_n10528), .Y(new_n15490_1));
  nor_5  g13142(.A(new_n15490_1), .B(new_n15489), .Y(new_n15491));
  xnor_4 g13143(.A(new_n15491), .B(new_n15488), .Y(new_n15492));
  xnor_4 g13144(.A(new_n15492), .B(new_n15486), .Y(new_n15493));
  and_5  g13145(.A(new_n10541), .B(new_n10526), .Y(new_n15494));
  nor_5  g13146(.A(new_n10574), .B(new_n10542), .Y(new_n15495));
  nor_5  g13147(.A(new_n15495), .B(new_n15494), .Y(new_n15496_1));
  xnor_4 g13148(.A(new_n15496_1), .B(new_n15493), .Y(new_n15497));
  not_8  g13149(.A(new_n15497), .Y(new_n15498));
  xnor_4 g13150(.A(new_n15498), .B(new_n5625), .Y(new_n15499));
  nor_5  g13151(.A(new_n10575), .B(new_n5632), .Y(new_n15500));
  and_5  g13152(.A(new_n10605), .B(new_n10577_1), .Y(new_n15501_1));
  nor_5  g13153(.A(new_n15501_1), .B(new_n15500), .Y(new_n15502));
  xor_4  g13154(.A(new_n15502), .B(new_n15499), .Y(n3563));
  xor_4  g13155(.A(new_n6133), .B(new_n6131), .Y(n3617));
  xnor_4 g13156(.A(n22253), .B(n8305), .Y(new_n15505));
  and_5  g13157(.A(new_n7043), .B(n1255), .Y(new_n15506_1));
  xnor_4 g13158(.A(n12861), .B(n1255), .Y(new_n15507));
  and_5  g13159(.A(new_n7046), .B(n9512), .Y(new_n15508_1));
  xnor_4 g13160(.A(n13333), .B(n9512), .Y(new_n15509));
  and_5  g13161(.A(n16608), .B(new_n7049), .Y(new_n15510));
  and_5  g13162(.A(n21735), .B(new_n5125), .Y(new_n15511));
  and_5  g13163(.A(new_n4635), .B(new_n4613), .Y(new_n15512));
  or_5   g13164(.A(new_n15512), .B(new_n15511), .Y(new_n15513));
  xnor_4 g13165(.A(n16608), .B(n2210), .Y(new_n15514));
  and_5  g13166(.A(new_n15514), .B(new_n15513), .Y(new_n15515));
  or_5   g13167(.A(new_n15515), .B(new_n15510), .Y(new_n15516));
  and_5  g13168(.A(new_n15516), .B(new_n15509), .Y(new_n15517));
  or_5   g13169(.A(new_n15517), .B(new_n15508_1), .Y(new_n15518));
  and_5  g13170(.A(new_n15518), .B(new_n15507), .Y(new_n15519));
  or_5   g13171(.A(new_n15519), .B(new_n15506_1), .Y(new_n15520));
  xor_4  g13172(.A(new_n15520), .B(new_n15505), .Y(new_n15521));
  xnor_4 g13173(.A(new_n15521), .B(new_n11226), .Y(new_n15522));
  xor_4  g13174(.A(new_n15518), .B(new_n15507), .Y(new_n15523));
  nor_5  g13175(.A(new_n15523), .B(new_n11229), .Y(new_n15524));
  xnor_4 g13176(.A(new_n15523), .B(new_n11229), .Y(new_n15525));
  xor_4  g13177(.A(new_n15516), .B(new_n15509), .Y(new_n15526));
  nor_5  g13178(.A(new_n15526), .B(new_n11233), .Y(new_n15527));
  xor_4  g13179(.A(new_n15514), .B(new_n15513), .Y(new_n15528));
  and_5  g13180(.A(new_n15528), .B(new_n11237), .Y(new_n15529));
  xnor_4 g13181(.A(new_n15528), .B(new_n11236), .Y(new_n15530));
  and_5  g13182(.A(new_n11240), .B(new_n4636), .Y(new_n15531));
  and_5  g13183(.A(new_n4756), .B(new_n4724), .Y(new_n15532));
  or_5   g13184(.A(new_n15532), .B(new_n15531), .Y(new_n15533));
  and_5  g13185(.A(new_n15533), .B(new_n15530), .Y(new_n15534));
  nor_5  g13186(.A(new_n15534), .B(new_n15529), .Y(new_n15535));
  xnor_4 g13187(.A(new_n15526), .B(new_n11233), .Y(new_n15536));
  not_8  g13188(.A(new_n15536), .Y(new_n15537));
  and_5  g13189(.A(new_n15537), .B(new_n15535), .Y(new_n15538));
  nor_5  g13190(.A(new_n15538), .B(new_n15527), .Y(new_n15539_1));
  nor_5  g13191(.A(new_n15539_1), .B(new_n15525), .Y(new_n15540));
  nor_5  g13192(.A(new_n15540), .B(new_n15524), .Y(new_n15541));
  xor_4  g13193(.A(new_n15541), .B(new_n15522), .Y(n3642));
  xnor_4 g13194(.A(n16544), .B(new_n3087), .Y(new_n15543));
  nor_5  g13195(.A(n23463), .B(n6814), .Y(new_n15544));
  xnor_4 g13196(.A(n23463), .B(new_n2887_1), .Y(new_n15545));
  nor_5  g13197(.A(n19701), .B(n13074), .Y(new_n15546_1));
  xnor_4 g13198(.A(n19701), .B(new_n3095), .Y(new_n15547));
  nor_5  g13199(.A(n23529), .B(n10739), .Y(new_n15548));
  xnor_4 g13200(.A(n23529), .B(new_n3099), .Y(new_n15549));
  nor_5  g13201(.A(n24620), .B(n21753), .Y(new_n15550));
  xnor_4 g13202(.A(n24620), .B(new_n2350), .Y(new_n15551));
  nor_5  g13203(.A(n21832), .B(n5211), .Y(new_n15552));
  and_5  g13204(.A(new_n14990), .B(new_n14982), .Y(new_n15553));
  or_5   g13205(.A(new_n15553), .B(new_n15552), .Y(new_n15554));
  and_5  g13206(.A(new_n15554), .B(new_n15551), .Y(new_n15555_1));
  or_5   g13207(.A(new_n15555_1), .B(new_n15550), .Y(new_n15556));
  and_5  g13208(.A(new_n15556), .B(new_n15549), .Y(new_n15557));
  or_5   g13209(.A(new_n15557), .B(new_n15548), .Y(new_n15558_1));
  and_5  g13210(.A(new_n15558_1), .B(new_n15547), .Y(new_n15559_1));
  or_5   g13211(.A(new_n15559_1), .B(new_n15546_1), .Y(new_n15560));
  and_5  g13212(.A(new_n15560), .B(new_n15545), .Y(new_n15561));
  nor_5  g13213(.A(new_n15561), .B(new_n15544), .Y(new_n15562));
  xnor_4 g13214(.A(new_n15562), .B(new_n15543), .Y(new_n15563));
  not_8  g13215(.A(new_n15563), .Y(new_n15564));
  xnor_4 g13216(.A(new_n15564), .B(n3324), .Y(new_n15565));
  nor_5  g13217(.A(new_n15559_1), .B(new_n15546_1), .Y(new_n15566));
  xnor_4 g13218(.A(new_n15566), .B(new_n15545), .Y(new_n15567));
  nor_5  g13219(.A(new_n15567), .B(n17911), .Y(new_n15568));
  not_8  g13220(.A(new_n15567), .Y(new_n15569));
  xnor_4 g13221(.A(new_n15569), .B(n17911), .Y(new_n15570_1));
  nor_5  g13222(.A(new_n15557), .B(new_n15548), .Y(new_n15571));
  xnor_4 g13223(.A(new_n15571), .B(new_n15547), .Y(new_n15572));
  nor_5  g13224(.A(new_n15572), .B(n21997), .Y(new_n15573_1));
  not_8  g13225(.A(new_n15572), .Y(new_n15574));
  xnor_4 g13226(.A(new_n15574), .B(n21997), .Y(new_n15575));
  nor_5  g13227(.A(new_n15555_1), .B(new_n15550), .Y(new_n15576));
  xnor_4 g13228(.A(new_n15576), .B(new_n15549), .Y(new_n15577));
  nor_5  g13229(.A(new_n15577), .B(n25119), .Y(new_n15578));
  xnor_4 g13230(.A(new_n15577), .B(new_n8501), .Y(new_n15579));
  nor_5  g13231(.A(new_n15553), .B(new_n15552), .Y(new_n15580));
  xnor_4 g13232(.A(new_n15580), .B(new_n15551), .Y(new_n15581));
  not_8  g13233(.A(new_n15581), .Y(new_n15582));
  nor_5  g13234(.A(new_n15582), .B(new_n8503), .Y(new_n15583));
  nor_5  g13235(.A(new_n14991), .B(n18537), .Y(new_n15584));
  or_5   g13236(.A(new_n15002_1), .B(new_n14995), .Y(new_n15585));
  and_5  g13237(.A(new_n15585), .B(new_n14992), .Y(new_n15586));
  nor_5  g13238(.A(new_n15586), .B(new_n15584), .Y(new_n15587));
  xnor_4 g13239(.A(new_n15582), .B(n1163), .Y(new_n15588_1));
  and_5  g13240(.A(new_n15588_1), .B(new_n15587), .Y(new_n15589));
  nor_5  g13241(.A(new_n15589), .B(new_n15583), .Y(new_n15590_1));
  and_5  g13242(.A(new_n15590_1), .B(new_n15579), .Y(new_n15591));
  or_5   g13243(.A(new_n15591), .B(new_n15578), .Y(new_n15592));
  and_5  g13244(.A(new_n15592), .B(new_n15575), .Y(new_n15593));
  or_5   g13245(.A(new_n15593), .B(new_n15573_1), .Y(new_n15594));
  and_5  g13246(.A(new_n15594), .B(new_n15570_1), .Y(new_n15595));
  nor_5  g13247(.A(new_n15595), .B(new_n15568), .Y(new_n15596));
  xnor_4 g13248(.A(new_n15596), .B(new_n15565), .Y(new_n15597));
  xnor_4 g13249(.A(n23250), .B(n16507), .Y(new_n15598_1));
  not_8  g13250(.A(n11455), .Y(new_n15599));
  nor_5  g13251(.A(n22470), .B(new_n15599), .Y(new_n15600));
  xnor_4 g13252(.A(n22470), .B(n11455), .Y(new_n15601));
  not_8  g13253(.A(n3945), .Y(new_n15602_1));
  nor_5  g13254(.A(n19116), .B(new_n15602_1), .Y(new_n15603));
  xnor_4 g13255(.A(n19116), .B(n3945), .Y(new_n15604));
  not_8  g13256(.A(n5255), .Y(new_n15605));
  nor_5  g13257(.A(n6861), .B(new_n15605), .Y(new_n15606));
  xnor_4 g13258(.A(n6861), .B(n5255), .Y(new_n15607));
  nor_5  g13259(.A(new_n5163), .B(n19357), .Y(new_n15608));
  xnor_4 g13260(.A(n21649), .B(n19357), .Y(new_n15609));
  nor_5  g13261(.A(new_n5166), .B(n2328), .Y(new_n15610));
  not_8  g13262(.A(n15053), .Y(new_n15611));
  nor_5  g13263(.A(new_n15611), .B(n3828), .Y(new_n15612));
  nor_5  g13264(.A(new_n5069), .B(new_n5065), .Y(new_n15613));
  nor_5  g13265(.A(new_n15613), .B(new_n15612), .Y(new_n15614_1));
  xnor_4 g13266(.A(n18274), .B(n2328), .Y(new_n15615));
  and_5  g13267(.A(new_n15615), .B(new_n15614_1), .Y(new_n15616));
  or_5   g13268(.A(new_n15616), .B(new_n15610), .Y(new_n15617));
  and_5  g13269(.A(new_n15617), .B(new_n15609), .Y(new_n15618));
  or_5   g13270(.A(new_n15618), .B(new_n15608), .Y(new_n15619));
  and_5  g13271(.A(new_n15619), .B(new_n15607), .Y(new_n15620));
  or_5   g13272(.A(new_n15620), .B(new_n15606), .Y(new_n15621));
  and_5  g13273(.A(new_n15621), .B(new_n15604), .Y(new_n15622));
  or_5   g13274(.A(new_n15622), .B(new_n15603), .Y(new_n15623));
  and_5  g13275(.A(new_n15623), .B(new_n15601), .Y(new_n15624));
  or_5   g13276(.A(new_n15624), .B(new_n15600), .Y(new_n15625));
  xor_4  g13277(.A(new_n15625), .B(new_n15598_1), .Y(new_n15626));
  nor_5  g13278(.A(new_n15626), .B(n4967), .Y(new_n15627));
  xnor_4 g13279(.A(new_n15626), .B(n4967), .Y(new_n15628));
  xor_4  g13280(.A(new_n15623), .B(new_n15601), .Y(new_n15629));
  nor_5  g13281(.A(new_n15629), .B(n15602), .Y(new_n15630));
  xor_4  g13282(.A(new_n15621), .B(new_n15604), .Y(new_n15631));
  and_5  g13283(.A(new_n15631), .B(n8694), .Y(new_n15632));
  xor_4  g13284(.A(new_n15619), .B(new_n15607), .Y(new_n15633));
  nor_5  g13285(.A(new_n15633), .B(n12380), .Y(new_n15634));
  xnor_4 g13286(.A(new_n15633), .B(n12380), .Y(new_n15635));
  xor_4  g13287(.A(new_n15617), .B(new_n15609), .Y(new_n15636_1));
  nor_5  g13288(.A(new_n15636_1), .B(n8943), .Y(new_n15637));
  xnor_4 g13289(.A(new_n15636_1), .B(n8943), .Y(new_n15638));
  not_8  g13290(.A(new_n15638), .Y(new_n15639));
  not_8  g13291(.A(n8255), .Y(new_n15640));
  xnor_4 g13292(.A(new_n15615), .B(new_n15614_1), .Y(new_n15641));
  nor_5  g13293(.A(new_n15641), .B(new_n15640), .Y(new_n15642));
  xnor_4 g13294(.A(new_n5069), .B(new_n5065), .Y(new_n15643));
  and_5  g13295(.A(new_n15643), .B(n11184), .Y(new_n15644));
  not_8  g13296(.A(new_n5071), .Y(new_n15645));
  nor_5  g13297(.A(new_n15645), .B(new_n5063), .Y(new_n15646));
  nor_5  g13298(.A(new_n15646), .B(new_n15644), .Y(new_n15647));
  xnor_4 g13299(.A(new_n15641), .B(n8255), .Y(new_n15648));
  not_8  g13300(.A(new_n15648), .Y(new_n15649));
  nor_5  g13301(.A(new_n15649), .B(new_n15647), .Y(new_n15650));
  nor_5  g13302(.A(new_n15650), .B(new_n15642), .Y(new_n15651));
  and_5  g13303(.A(new_n15651), .B(new_n15639), .Y(new_n15652_1));
  nor_5  g13304(.A(new_n15652_1), .B(new_n15637), .Y(new_n15653));
  nor_5  g13305(.A(new_n15653), .B(new_n15635), .Y(new_n15654));
  nor_5  g13306(.A(new_n15654), .B(new_n15634), .Y(new_n15655));
  xnor_4 g13307(.A(new_n15631), .B(n8694), .Y(new_n15656));
  not_8  g13308(.A(new_n15656), .Y(new_n15657));
  and_5  g13309(.A(new_n15657), .B(new_n15655), .Y(new_n15658));
  nor_5  g13310(.A(new_n15658), .B(new_n15632), .Y(new_n15659));
  not_8  g13311(.A(n15602), .Y(new_n15660));
  xnor_4 g13312(.A(new_n15629), .B(new_n15660), .Y(new_n15661));
  and_5  g13313(.A(new_n15661), .B(new_n15659), .Y(new_n15662_1));
  nor_5  g13314(.A(new_n15662_1), .B(new_n15630), .Y(new_n15663));
  nor_5  g13315(.A(new_n15663), .B(new_n15628), .Y(new_n15664));
  nor_5  g13316(.A(new_n15664), .B(new_n15627), .Y(new_n15665));
  xnor_4 g13317(.A(n6659), .B(n5101), .Y(new_n15666));
  not_8  g13318(.A(n23250), .Y(new_n15667));
  nor_5  g13319(.A(new_n15667), .B(n16507), .Y(new_n15668));
  and_5  g13320(.A(new_n15625), .B(new_n15598_1), .Y(new_n15669));
  or_5   g13321(.A(new_n15669), .B(new_n15668), .Y(new_n15670));
  xor_4  g13322(.A(new_n15670), .B(new_n15666), .Y(new_n15671));
  xnor_4 g13323(.A(new_n15671), .B(n13419), .Y(new_n15672));
  xor_4  g13324(.A(new_n15672), .B(new_n15665), .Y(new_n15673));
  xor_4  g13325(.A(new_n15673), .B(new_n15597), .Y(new_n15674));
  nor_5  g13326(.A(new_n15593), .B(new_n15573_1), .Y(new_n15675));
  xnor_4 g13327(.A(new_n15675), .B(new_n15570_1), .Y(new_n15676));
  not_8  g13328(.A(new_n15676), .Y(new_n15677));
  xnor_4 g13329(.A(new_n15663), .B(new_n15628), .Y(new_n15678));
  nor_5  g13330(.A(new_n15678), .B(new_n15677), .Y(new_n15679));
  xnor_4 g13331(.A(new_n15678), .B(new_n15677), .Y(new_n15680));
  xor_4  g13332(.A(new_n15592), .B(new_n15575), .Y(new_n15681));
  not_8  g13333(.A(new_n15661), .Y(new_n15682));
  xnor_4 g13334(.A(new_n15682), .B(new_n15659), .Y(new_n15683));
  and_5  g13335(.A(new_n15683), .B(new_n15681), .Y(new_n15684));
  xnor_4 g13336(.A(new_n15683), .B(new_n15681), .Y(new_n15685));
  xnor_4 g13337(.A(new_n15590_1), .B(new_n15579), .Y(new_n15686));
  xnor_4 g13338(.A(new_n15656), .B(new_n15655), .Y(new_n15687));
  nor_5  g13339(.A(new_n15687), .B(new_n15686), .Y(new_n15688));
  xnor_4 g13340(.A(new_n15687), .B(new_n15686), .Y(new_n15689));
  xnor_4 g13341(.A(new_n15653), .B(new_n15635), .Y(new_n15690));
  xor_4  g13342(.A(new_n15588_1), .B(new_n15587), .Y(new_n15691));
  nor_5  g13343(.A(new_n15691), .B(new_n15690), .Y(new_n15692));
  xnor_4 g13344(.A(new_n15691), .B(new_n15690), .Y(new_n15693));
  xnor_4 g13345(.A(new_n15651), .B(new_n15638), .Y(new_n15694));
  and_5  g13346(.A(new_n15694), .B(new_n15004_1), .Y(new_n15695));
  xnor_4 g13347(.A(new_n15694), .B(new_n15004_1), .Y(new_n15696));
  not_8  g13348(.A(new_n15024), .Y(new_n15697));
  xnor_4 g13349(.A(new_n15648), .B(new_n15647), .Y(new_n15698));
  nor_5  g13350(.A(new_n15698), .B(new_n15697), .Y(new_n15699));
  xnor_4 g13351(.A(new_n15698), .B(new_n15697), .Y(new_n15700));
  nor_5  g13352(.A(new_n5072), .B(new_n5052), .Y(new_n15701));
  nor_5  g13353(.A(new_n5088), .B(new_n5073), .Y(new_n15702));
  nor_5  g13354(.A(new_n15702), .B(new_n15701), .Y(new_n15703));
  nor_5  g13355(.A(new_n15703), .B(new_n15700), .Y(new_n15704));
  nor_5  g13356(.A(new_n15704), .B(new_n15699), .Y(new_n15705));
  nor_5  g13357(.A(new_n15705), .B(new_n15696), .Y(new_n15706));
  nor_5  g13358(.A(new_n15706), .B(new_n15695), .Y(new_n15707));
  nor_5  g13359(.A(new_n15707), .B(new_n15693), .Y(new_n15708));
  nor_5  g13360(.A(new_n15708), .B(new_n15692), .Y(new_n15709));
  nor_5  g13361(.A(new_n15709), .B(new_n15689), .Y(new_n15710));
  nor_5  g13362(.A(new_n15710), .B(new_n15688), .Y(new_n15711));
  nor_5  g13363(.A(new_n15711), .B(new_n15685), .Y(new_n15712));
  nor_5  g13364(.A(new_n15712), .B(new_n15684), .Y(new_n15713));
  nor_5  g13365(.A(new_n15713), .B(new_n15680), .Y(new_n15714));
  nor_5  g13366(.A(new_n15714), .B(new_n15679), .Y(new_n15715));
  xor_4  g13367(.A(new_n15715), .B(new_n15674), .Y(n3649));
  nor_5  g13368(.A(n26625), .B(n14230), .Y(new_n15717));
  not_8  g13369(.A(new_n15717), .Y(new_n15718));
  nor_5  g13370(.A(new_n15718), .B(n26744), .Y(new_n15719));
  not_8  g13371(.A(new_n15719), .Y(new_n15720));
  nor_5  g13372(.A(new_n15720), .B(n11566), .Y(new_n15721));
  not_8  g13373(.A(new_n15721), .Y(new_n15722));
  nor_5  g13374(.A(new_n15722), .B(n3959), .Y(new_n15723));
  not_8  g13375(.A(new_n15723), .Y(new_n15724));
  nor_5  g13376(.A(new_n15724), .B(n26565), .Y(new_n15725));
  xnor_4 g13377(.A(new_n15725), .B(n3366), .Y(new_n15726));
  xnor_4 g13378(.A(new_n15726), .B(n26191), .Y(new_n15727));
  xnor_4 g13379(.A(new_n15723), .B(n26565), .Y(new_n15728));
  not_8  g13380(.A(new_n15728), .Y(new_n15729));
  nor_5  g13381(.A(new_n15729), .B(n26512), .Y(new_n15730));
  xnor_4 g13382(.A(new_n15728), .B(n26512), .Y(new_n15731));
  not_8  g13383(.A(n19575), .Y(new_n15732));
  xnor_4 g13384(.A(new_n15721), .B(n3959), .Y(new_n15733));
  and_5  g13385(.A(new_n15733), .B(new_n15732), .Y(new_n15734));
  xnor_4 g13386(.A(new_n15733), .B(n19575), .Y(new_n15735));
  not_8  g13387(.A(n15378), .Y(new_n15736));
  xnor_4 g13388(.A(new_n15719), .B(n11566), .Y(new_n15737));
  and_5  g13389(.A(new_n15737), .B(new_n15736), .Y(new_n15738));
  xnor_4 g13390(.A(new_n15737), .B(n15378), .Y(new_n15739));
  xnor_4 g13391(.A(new_n15717), .B(n26744), .Y(new_n15740));
  not_8  g13392(.A(new_n15740), .Y(new_n15741));
  nor_5  g13393(.A(new_n15741), .B(n17095), .Y(new_n15742));
  xnor_4 g13394(.A(n26625), .B(new_n9484), .Y(new_n15743_1));
  nor_5  g13395(.A(new_n15743_1), .B(new_n9531), .Y(new_n15744));
  nor_5  g13396(.A(new_n9532), .B(n14230), .Y(new_n15745));
  xnor_4 g13397(.A(new_n15743_1), .B(n22591), .Y(new_n15746));
  and_5  g13398(.A(new_n15746), .B(new_n15745), .Y(new_n15747));
  nor_5  g13399(.A(new_n15747), .B(new_n15744), .Y(new_n15748));
  xnor_4 g13400(.A(new_n15740), .B(n17095), .Y(new_n15749_1));
  and_5  g13401(.A(new_n15749_1), .B(new_n15748), .Y(new_n15750));
  or_5   g13402(.A(new_n15750), .B(new_n15742), .Y(new_n15751));
  and_5  g13403(.A(new_n15751), .B(new_n15739), .Y(new_n15752));
  or_5   g13404(.A(new_n15752), .B(new_n15738), .Y(new_n15753));
  and_5  g13405(.A(new_n15753), .B(new_n15735), .Y(new_n15754));
  or_5   g13406(.A(new_n15754), .B(new_n15734), .Y(new_n15755));
  and_5  g13407(.A(new_n15755), .B(new_n15731), .Y(new_n15756));
  or_5   g13408(.A(new_n15756), .B(new_n15730), .Y(new_n15757));
  xor_4  g13409(.A(new_n15757), .B(new_n15727), .Y(new_n15758));
  xnor_4 g13410(.A(new_n15758), .B(n7917), .Y(new_n15759));
  xor_4  g13411(.A(new_n15755), .B(new_n15731), .Y(new_n15760));
  and_5  g13412(.A(new_n15760), .B(new_n14174_1), .Y(new_n15761_1));
  xnor_4 g13413(.A(new_n15760), .B(n17302), .Y(new_n15762_1));
  xor_4  g13414(.A(new_n15753), .B(new_n15735), .Y(new_n15763));
  nor_5  g13415(.A(new_n15763), .B(new_n14177), .Y(new_n15764));
  xnor_4 g13416(.A(new_n15763), .B(new_n14177), .Y(new_n15765));
  xor_4  g13417(.A(new_n15751), .B(new_n15739), .Y(new_n15766_1));
  nor_5  g13418(.A(new_n15766_1), .B(new_n14191), .Y(new_n15767));
  xnor_4 g13419(.A(new_n15766_1), .B(new_n14191), .Y(new_n15768));
  xor_4  g13420(.A(new_n15749_1), .B(new_n15748), .Y(new_n15769));
  nor_5  g13421(.A(new_n15769), .B(new_n14181), .Y(new_n15770));
  xnor_4 g13422(.A(new_n15769), .B(new_n14181), .Y(new_n15771));
  xnor_4 g13423(.A(new_n15746), .B(new_n15745), .Y(new_n15772));
  nor_5  g13424(.A(new_n15772), .B(new_n14183), .Y(new_n15773));
  not_8  g13425(.A(new_n15772), .Y(new_n15774));
  or_5   g13426(.A(new_n15774), .B(n22358), .Y(new_n15775));
  xnor_4 g13427(.A(n26167), .B(n14230), .Y(new_n15776));
  and_5  g13428(.A(new_n15776), .B(n9646), .Y(new_n15777));
  and_5  g13429(.A(new_n15777), .B(new_n15775), .Y(new_n15778));
  nor_5  g13430(.A(new_n15778), .B(new_n15773), .Y(new_n15779));
  nor_5  g13431(.A(new_n15779), .B(new_n15771), .Y(new_n15780_1));
  nor_5  g13432(.A(new_n15780_1), .B(new_n15770), .Y(new_n15781));
  nor_5  g13433(.A(new_n15781), .B(new_n15768), .Y(new_n15782));
  nor_5  g13434(.A(new_n15782), .B(new_n15767), .Y(new_n15783));
  nor_5  g13435(.A(new_n15783), .B(new_n15765), .Y(new_n15784));
  nor_5  g13436(.A(new_n15784), .B(new_n15764), .Y(new_n15785));
  and_5  g13437(.A(new_n15785), .B(new_n15762_1), .Y(new_n15786));
  or_5   g13438(.A(new_n15786), .B(new_n15761_1), .Y(new_n15787));
  xor_4  g13439(.A(new_n15787), .B(new_n15759), .Y(new_n15788));
  xnor_4 g13440(.A(new_n15788), .B(new_n6918), .Y(new_n15789));
  xor_4  g13441(.A(new_n15785), .B(new_n15762_1), .Y(new_n15790));
  nor_5  g13442(.A(new_n15790), .B(new_n6923), .Y(new_n15791));
  xnor_4 g13443(.A(new_n15790), .B(new_n6923), .Y(new_n15792));
  xnor_4 g13444(.A(new_n15783), .B(new_n15765), .Y(new_n15793_1));
  nor_5  g13445(.A(new_n15793_1), .B(new_n6926), .Y(new_n15794));
  xnor_4 g13446(.A(new_n15793_1), .B(new_n6926), .Y(new_n15795));
  not_8  g13447(.A(new_n6931), .Y(new_n15796));
  xnor_4 g13448(.A(new_n15781), .B(new_n15768), .Y(new_n15797));
  nor_5  g13449(.A(new_n15797), .B(new_n15796), .Y(new_n15798));
  xnor_4 g13450(.A(new_n15797), .B(new_n15796), .Y(new_n15799));
  xnor_4 g13451(.A(new_n15779), .B(new_n15771), .Y(new_n15800));
  nor_5  g13452(.A(new_n15800), .B(new_n6937), .Y(new_n15801));
  xnor_4 g13453(.A(new_n15800), .B(new_n6936), .Y(new_n15802));
  xnor_4 g13454(.A(new_n15774), .B(n22358), .Y(new_n15803));
  xnor_4 g13455(.A(new_n15803), .B(new_n15777), .Y(new_n15804));
  nor_5  g13456(.A(new_n15804), .B(new_n6943), .Y(new_n15805));
  xnor_4 g13457(.A(new_n15776), .B(new_n6585), .Y(new_n15806));
  nor_5  g13458(.A(new_n15806), .B(new_n6947), .Y(new_n15807));
  xnor_4 g13459(.A(new_n15804), .B(new_n6944), .Y(new_n15808));
  and_5  g13460(.A(new_n15808), .B(new_n15807), .Y(new_n15809));
  nor_5  g13461(.A(new_n15809), .B(new_n15805), .Y(new_n15810));
  and_5  g13462(.A(new_n15810), .B(new_n15802), .Y(new_n15811));
  nor_5  g13463(.A(new_n15811), .B(new_n15801), .Y(new_n15812_1));
  nor_5  g13464(.A(new_n15812_1), .B(new_n15799), .Y(new_n15813));
  nor_5  g13465(.A(new_n15813), .B(new_n15798), .Y(new_n15814));
  nor_5  g13466(.A(new_n15814), .B(new_n15795), .Y(new_n15815_1));
  nor_5  g13467(.A(new_n15815_1), .B(new_n15794), .Y(new_n15816_1));
  nor_5  g13468(.A(new_n15816_1), .B(new_n15792), .Y(new_n15817));
  nor_5  g13469(.A(new_n15817), .B(new_n15791), .Y(new_n15818));
  xnor_4 g13470(.A(new_n15818), .B(new_n15789), .Y(n3665));
  xnor_4 g13471(.A(new_n5802), .B(new_n5801), .Y(n3679));
  nor_5  g13472(.A(n16521), .B(n7139), .Y(new_n15821));
  not_8  g13473(.A(new_n15821), .Y(new_n15822));
  nor_5  g13474(.A(new_n15822), .B(n16824), .Y(new_n15823));
  not_8  g13475(.A(new_n15823), .Y(new_n15824));
  nor_5  g13476(.A(new_n15824), .B(n604), .Y(new_n15825));
  not_8  g13477(.A(new_n15825), .Y(new_n15826));
  nor_5  g13478(.A(new_n15826), .B(n4913), .Y(new_n15827));
  not_8  g13479(.A(new_n15827), .Y(new_n15828));
  nor_5  g13480(.A(new_n15828), .B(n9172), .Y(new_n15829));
  not_8  g13481(.A(new_n15829), .Y(new_n15830));
  nor_5  g13482(.A(new_n15830), .B(n442), .Y(new_n15831_1));
  not_8  g13483(.A(new_n15831_1), .Y(new_n15832));
  nor_5  g13484(.A(new_n15832), .B(n13719), .Y(new_n15833));
  xnor_4 g13485(.A(new_n15833), .B(n7026), .Y(new_n15834));
  xnor_4 g13486(.A(new_n15834), .B(new_n5921), .Y(new_n15835));
  xnor_4 g13487(.A(new_n15831_1), .B(n13719), .Y(new_n15836));
  and_5  g13488(.A(new_n15836), .B(new_n5925), .Y(new_n15837));
  not_8  g13489(.A(new_n5925), .Y(new_n15838));
  xnor_4 g13490(.A(new_n15836), .B(new_n15838), .Y(new_n15839));
  xnor_4 g13491(.A(new_n15829), .B(n442), .Y(new_n15840));
  nor_5  g13492(.A(new_n15840), .B(new_n5930), .Y(new_n15841));
  not_8  g13493(.A(new_n5930), .Y(new_n15842));
  xnor_4 g13494(.A(new_n15840), .B(new_n15842), .Y(new_n15843));
  xnor_4 g13495(.A(new_n15827), .B(n9172), .Y(new_n15844));
  nor_5  g13496(.A(new_n15844), .B(new_n5935), .Y(new_n15845));
  xnor_4 g13497(.A(new_n15844), .B(new_n13211), .Y(new_n15846_1));
  xnor_4 g13498(.A(new_n15825), .B(n4913), .Y(new_n15847));
  nor_5  g13499(.A(new_n15847), .B(new_n5940), .Y(new_n15848));
  xnor_4 g13500(.A(new_n15847), .B(new_n13213), .Y(new_n15849));
  xnor_4 g13501(.A(new_n15823), .B(n604), .Y(new_n15850));
  nor_5  g13502(.A(new_n15850), .B(new_n5945), .Y(new_n15851));
  xnor_4 g13503(.A(new_n15850), .B(new_n5947), .Y(new_n15852));
  xnor_4 g13504(.A(new_n15821), .B(n16824), .Y(new_n15853));
  nor_5  g13505(.A(new_n15853), .B(new_n5952), .Y(new_n15854));
  xnor_4 g13506(.A(new_n15853), .B(new_n5953), .Y(new_n15855));
  nor_5  g13507(.A(new_n15822), .B(new_n5956), .Y(new_n15856));
  nor_5  g13508(.A(new_n10777), .B(n7139), .Y(new_n15857));
  xnor_4 g13509(.A(new_n15857), .B(new_n3560), .Y(new_n15858));
  and_5  g13510(.A(new_n15858), .B(new_n5959), .Y(new_n15859_1));
  or_5   g13511(.A(new_n15859_1), .B(new_n15856), .Y(new_n15860));
  and_5  g13512(.A(new_n15860), .B(new_n15855), .Y(new_n15861));
  or_5   g13513(.A(new_n15861), .B(new_n15854), .Y(new_n15862));
  and_5  g13514(.A(new_n15862), .B(new_n15852), .Y(new_n15863));
  or_5   g13515(.A(new_n15863), .B(new_n15851), .Y(new_n15864));
  and_5  g13516(.A(new_n15864), .B(new_n15849), .Y(new_n15865));
  or_5   g13517(.A(new_n15865), .B(new_n15848), .Y(new_n15866));
  and_5  g13518(.A(new_n15866), .B(new_n15846_1), .Y(new_n15867));
  or_5   g13519(.A(new_n15867), .B(new_n15845), .Y(new_n15868));
  and_5  g13520(.A(new_n15868), .B(new_n15843), .Y(new_n15869_1));
  nor_5  g13521(.A(new_n15869_1), .B(new_n15841), .Y(new_n15870));
  and_5  g13522(.A(new_n15870), .B(new_n15839), .Y(new_n15871));
  or_5   g13523(.A(new_n15871), .B(new_n15837), .Y(new_n15872));
  xor_4  g13524(.A(new_n15872), .B(new_n15835), .Y(new_n15873));
  xnor_4 g13525(.A(new_n6029), .B(new_n4909), .Y(new_n15874));
  nor_5  g13526(.A(new_n6033), .B(new_n4913_1), .Y(new_n15875));
  xnor_4 g13527(.A(new_n6035), .B(new_n4913_1), .Y(new_n15876));
  nor_5  g13528(.A(new_n6039), .B(new_n4917), .Y(new_n15877));
  or_5   g13529(.A(new_n8497), .B(new_n8477), .Y(new_n15878));
  and_5  g13530(.A(new_n15878), .B(new_n8476), .Y(new_n15879));
  or_5   g13531(.A(new_n15879), .B(new_n15877), .Y(new_n15880));
  and_5  g13532(.A(new_n15880), .B(new_n15876), .Y(new_n15881));
  nor_5  g13533(.A(new_n15881), .B(new_n15875), .Y(new_n15882));
  xnor_4 g13534(.A(new_n15882), .B(new_n15874), .Y(new_n15883));
  xnor_4 g13535(.A(new_n15883), .B(new_n15873), .Y(new_n15884_1));
  xor_4  g13536(.A(new_n15880), .B(new_n15876), .Y(new_n15885_1));
  xor_4  g13537(.A(new_n15870), .B(new_n15839), .Y(new_n15886));
  nor_5  g13538(.A(new_n15886), .B(new_n15885_1), .Y(new_n15887));
  xnor_4 g13539(.A(new_n15886), .B(new_n15885_1), .Y(new_n15888));
  xor_4  g13540(.A(new_n15868), .B(new_n15843), .Y(new_n15889_1));
  and_5  g13541(.A(new_n15889_1), .B(new_n8500), .Y(new_n15890));
  xnor_4 g13542(.A(new_n15889_1), .B(new_n8500), .Y(new_n15891));
  xor_4  g13543(.A(new_n15866), .B(new_n15846_1), .Y(new_n15892));
  and_5  g13544(.A(new_n15892), .B(new_n8531), .Y(new_n15893));
  xnor_4 g13545(.A(new_n15892), .B(new_n8531), .Y(new_n15894));
  not_8  g13546(.A(new_n8537), .Y(new_n15895));
  xor_4  g13547(.A(new_n15864), .B(new_n15849), .Y(new_n15896));
  and_5  g13548(.A(new_n15896), .B(new_n15895), .Y(new_n15897));
  xnor_4 g13549(.A(new_n15896), .B(new_n15895), .Y(new_n15898));
  xor_4  g13550(.A(new_n15862), .B(new_n15852), .Y(new_n15899));
  and_5  g13551(.A(new_n15899), .B(new_n8543), .Y(new_n15900));
  xnor_4 g13552(.A(new_n15899), .B(new_n8542), .Y(new_n15901));
  xor_4  g13553(.A(new_n15860), .B(new_n15855), .Y(new_n15902));
  nor_5  g13554(.A(new_n15902), .B(new_n8547), .Y(new_n15903));
  xnor_4 g13555(.A(new_n15902), .B(new_n8548), .Y(new_n15904));
  xnor_4 g13556(.A(new_n15858), .B(new_n6127), .Y(new_n15905));
  and_5  g13557(.A(new_n15905), .B(new_n8552), .Y(new_n15906));
  xnor_4 g13558(.A(new_n5956), .B(n7139), .Y(new_n15907));
  and_5  g13559(.A(new_n15907), .B(new_n8556), .Y(new_n15908));
  xnor_4 g13560(.A(new_n15905), .B(new_n8552), .Y(new_n15909));
  nor_5  g13561(.A(new_n15909), .B(new_n15908), .Y(new_n15910));
  nor_5  g13562(.A(new_n15910), .B(new_n15906), .Y(new_n15911));
  and_5  g13563(.A(new_n15911), .B(new_n15904), .Y(new_n15912));
  nor_5  g13564(.A(new_n15912), .B(new_n15903), .Y(new_n15913));
  and_5  g13565(.A(new_n15913), .B(new_n15901), .Y(new_n15914));
  nor_5  g13566(.A(new_n15914), .B(new_n15900), .Y(new_n15915));
  nor_5  g13567(.A(new_n15915), .B(new_n15898), .Y(new_n15916));
  nor_5  g13568(.A(new_n15916), .B(new_n15897), .Y(new_n15917_1));
  nor_5  g13569(.A(new_n15917_1), .B(new_n15894), .Y(new_n15918_1));
  nor_5  g13570(.A(new_n15918_1), .B(new_n15893), .Y(new_n15919));
  nor_5  g13571(.A(new_n15919), .B(new_n15891), .Y(new_n15920));
  nor_5  g13572(.A(new_n15920), .B(new_n15890), .Y(new_n15921));
  nor_5  g13573(.A(new_n15921), .B(new_n15888), .Y(new_n15922_1));
  nor_5  g13574(.A(new_n15922_1), .B(new_n15887), .Y(new_n15923));
  xnor_4 g13575(.A(new_n15923), .B(new_n15884_1), .Y(n3725));
  nor_5  g13576(.A(n11220), .B(n3425), .Y(new_n15925));
  nor_5  g13577(.A(new_n12817), .B(new_n12814), .Y(new_n15926));
  nor_5  g13578(.A(new_n15926), .B(new_n15925), .Y(new_n15927));
  nor_5  g13579(.A(n7335), .B(n2160), .Y(new_n15928));
  and_5  g13580(.A(new_n12812_1), .B(new_n12809), .Y(new_n15929));
  nor_5  g13581(.A(new_n15929), .B(new_n15928), .Y(new_n15930));
  xnor_4 g13582(.A(new_n15930), .B(new_n15927), .Y(new_n15931));
  nor_5  g13583(.A(new_n12818), .B(new_n12813), .Y(new_n15932));
  nor_5  g13584(.A(new_n12822), .B(new_n12819), .Y(new_n15933));
  nor_5  g13585(.A(new_n15933), .B(new_n15932), .Y(new_n15934));
  not_8  g13586(.A(new_n15934), .Y(new_n15935));
  xnor_4 g13587(.A(new_n15935), .B(new_n15931), .Y(new_n15936_1));
  xnor_4 g13588(.A(new_n15936_1), .B(new_n14514), .Y(new_n15937));
  nor_5  g13589(.A(new_n14518), .B(new_n12824), .Y(new_n15938));
  xnor_4 g13590(.A(new_n14518), .B(new_n12823), .Y(new_n15939));
  and_5  g13591(.A(new_n14522), .B(new_n5400_1), .Y(new_n15940));
  xnor_4 g13592(.A(new_n14522), .B(new_n5399_1), .Y(new_n15941));
  nor_5  g13593(.A(new_n14526), .B(new_n5403_1), .Y(new_n15942));
  not_8  g13594(.A(new_n5409), .Y(new_n15943));
  nor_5  g13595(.A(new_n14529), .B(new_n15943), .Y(new_n15944));
  xnor_4 g13596(.A(new_n14529), .B(new_n15943), .Y(new_n15945));
  nor_5  g13597(.A(new_n14444), .B(new_n5413), .Y(new_n15946));
  xnor_4 g13598(.A(new_n14445), .B(new_n5414), .Y(new_n15947_1));
  nor_5  g13599(.A(new_n5418), .B(new_n4251), .Y(new_n15948));
  nor_5  g13600(.A(new_n5421), .B(new_n4258), .Y(new_n15949));
  xnor_4 g13601(.A(new_n5421), .B(new_n4257), .Y(new_n15950));
  nor_5  g13602(.A(new_n5427), .B(new_n4261), .Y(new_n15951));
  xnor_4 g13603(.A(new_n5427), .B(new_n4277), .Y(new_n15952));
  nor_5  g13604(.A(new_n5432), .B(new_n4264), .Y(new_n15953));
  or_5   g13605(.A(new_n5430_1), .B(new_n4244), .Y(new_n15954));
  nor_5  g13606(.A(new_n5436), .B(new_n4266_1), .Y(new_n15955));
  and_5  g13607(.A(new_n15955), .B(new_n15954), .Y(new_n15956_1));
  or_5   g13608(.A(new_n15956_1), .B(new_n15953), .Y(new_n15957));
  and_5  g13609(.A(new_n15957), .B(new_n15952), .Y(new_n15958_1));
  or_5   g13610(.A(new_n15958_1), .B(new_n15951), .Y(new_n15959));
  and_5  g13611(.A(new_n15959), .B(new_n15950), .Y(new_n15960));
  nor_5  g13612(.A(new_n15960), .B(new_n15949), .Y(new_n15961));
  xnor_4 g13613(.A(new_n5418), .B(new_n14447), .Y(new_n15962));
  and_5  g13614(.A(new_n15962), .B(new_n15961), .Y(new_n15963));
  nor_5  g13615(.A(new_n15963), .B(new_n15948), .Y(new_n15964));
  nor_5  g13616(.A(new_n15964), .B(new_n15947_1), .Y(new_n15965));
  nor_5  g13617(.A(new_n15965), .B(new_n15946), .Y(new_n15966));
  nor_5  g13618(.A(new_n15966), .B(new_n15945), .Y(new_n15967_1));
  nor_5  g13619(.A(new_n15967_1), .B(new_n15944), .Y(new_n15968));
  xnor_4 g13620(.A(new_n14526), .B(new_n5404), .Y(new_n15969));
  and_5  g13621(.A(new_n15969), .B(new_n15968), .Y(new_n15970));
  or_5   g13622(.A(new_n15970), .B(new_n15942), .Y(new_n15971));
  and_5  g13623(.A(new_n15971), .B(new_n15941), .Y(new_n15972));
  nor_5  g13624(.A(new_n15972), .B(new_n15940), .Y(new_n15973));
  and_5  g13625(.A(new_n15973), .B(new_n15939), .Y(new_n15974));
  nor_5  g13626(.A(new_n15974), .B(new_n15938), .Y(new_n15975));
  xnor_4 g13627(.A(new_n15975), .B(new_n15937), .Y(n3733));
  xnor_4 g13628(.A(new_n10658), .B(n24937), .Y(new_n15977));
  nor_5  g13629(.A(new_n10649), .B(new_n15124), .Y(new_n15978));
  xnor_4 g13630(.A(new_n10650_1), .B(new_n15124), .Y(new_n15979_1));
  and_5  g13631(.A(new_n10640), .B(n3030), .Y(new_n15980));
  or_5   g13632(.A(new_n15056), .B(new_n15046), .Y(new_n15981));
  and_5  g13633(.A(new_n15981), .B(new_n15044), .Y(new_n15982));
  or_5   g13634(.A(new_n15982), .B(new_n15980), .Y(new_n15983));
  and_5  g13635(.A(new_n15983), .B(new_n15979_1), .Y(new_n15984));
  nor_5  g13636(.A(new_n15984), .B(new_n15978), .Y(new_n15985));
  xnor_4 g13637(.A(new_n15985), .B(new_n15977), .Y(new_n15986_1));
  not_8  g13638(.A(new_n15986_1), .Y(new_n15987));
  xnor_4 g13639(.A(new_n15987), .B(new_n9934_1), .Y(new_n15988));
  nor_5  g13640(.A(new_n15982), .B(new_n15980), .Y(new_n15989));
  xnor_4 g13641(.A(new_n15989), .B(new_n15979_1), .Y(new_n15990));
  nor_5  g13642(.A(new_n15990), .B(new_n9939), .Y(new_n15991));
  not_8  g13643(.A(new_n15990), .Y(new_n15992));
  xnor_4 g13644(.A(new_n15992), .B(new_n9939), .Y(new_n15993));
  nor_5  g13645(.A(new_n15058), .B(new_n9943), .Y(new_n15994));
  and_5  g13646(.A(new_n15076), .B(new_n15060), .Y(new_n15995));
  or_5   g13647(.A(new_n15995), .B(new_n15994), .Y(new_n15996));
  and_5  g13648(.A(new_n15996), .B(new_n15993), .Y(new_n15997));
  or_5   g13649(.A(new_n15997), .B(new_n15991), .Y(new_n15998));
  xor_4  g13650(.A(new_n15998), .B(new_n15988), .Y(n3755));
  xnor_4 g13651(.A(new_n9049), .B(new_n9017), .Y(n3758));
  not_8  g13652(.A(new_n15368), .Y(new_n16001));
  nor_5  g13653(.A(new_n16001), .B(n18145), .Y(new_n16002));
  not_8  g13654(.A(new_n16002), .Y(new_n16003));
  nor_5  g13655(.A(new_n16003), .B(n655), .Y(new_n16004));
  not_8  g13656(.A(new_n16004), .Y(new_n16005));
  nor_5  g13657(.A(new_n16005), .B(n19033), .Y(new_n16006));
  xnor_4 g13658(.A(new_n16006), .B(n2570), .Y(new_n16007));
  xnor_4 g13659(.A(new_n16007), .B(n14692), .Y(new_n16008));
  xnor_4 g13660(.A(new_n16004), .B(n19033), .Y(new_n16009));
  nor_5  g13661(.A(new_n16009), .B(new_n10170), .Y(new_n16010));
  xnor_4 g13662(.A(new_n16009), .B(n4100), .Y(new_n16011));
  xnor_4 g13663(.A(new_n16002), .B(n655), .Y(new_n16012));
  nor_5  g13664(.A(new_n16012), .B(new_n10173), .Y(new_n16013_1));
  xnor_4 g13665(.A(new_n16012), .B(n21957), .Y(new_n16014));
  nor_5  g13666(.A(new_n15369), .B(new_n10176), .Y(new_n16015));
  and_5  g13667(.A(new_n15397), .B(new_n15370), .Y(new_n16016));
  or_5   g13668(.A(new_n16016), .B(new_n16015), .Y(new_n16017));
  and_5  g13669(.A(new_n16017), .B(new_n16014), .Y(new_n16018));
  or_5   g13670(.A(new_n16018), .B(new_n16013_1), .Y(new_n16019));
  and_5  g13671(.A(new_n16019), .B(new_n16011), .Y(new_n16020));
  or_5   g13672(.A(new_n16020), .B(new_n16010), .Y(new_n16021));
  xor_4  g13673(.A(new_n16021), .B(new_n16008), .Y(new_n16022));
  and_5  g13674(.A(new_n16022), .B(new_n11803), .Y(new_n16023));
  xnor_4 g13675(.A(new_n16022), .B(new_n11803), .Y(new_n16024));
  xor_4  g13676(.A(new_n16019), .B(new_n16011), .Y(new_n16025));
  and_5  g13677(.A(new_n16025), .B(new_n6863_1), .Y(new_n16026));
  xnor_4 g13678(.A(new_n16025), .B(new_n6863_1), .Y(new_n16027));
  xor_4  g13679(.A(new_n16017), .B(new_n16014), .Y(new_n16028));
  and_5  g13680(.A(new_n16028), .B(new_n6867_1), .Y(new_n16029_1));
  xnor_4 g13681(.A(new_n16028), .B(new_n6867_1), .Y(new_n16030));
  and_5  g13682(.A(new_n15398), .B(new_n6872), .Y(new_n16031));
  and_5  g13683(.A(new_n15426), .B(new_n15399), .Y(new_n16032));
  nor_5  g13684(.A(new_n16032), .B(new_n16031), .Y(new_n16033));
  nor_5  g13685(.A(new_n16033), .B(new_n16030), .Y(new_n16034));
  nor_5  g13686(.A(new_n16034), .B(new_n16029_1), .Y(new_n16035));
  nor_5  g13687(.A(new_n16035), .B(new_n16027), .Y(new_n16036));
  nor_5  g13688(.A(new_n16036), .B(new_n16026), .Y(new_n16037));
  nor_5  g13689(.A(new_n16037), .B(new_n16024), .Y(new_n16038));
  nor_5  g13690(.A(new_n16038), .B(new_n16023), .Y(new_n16039));
  not_8  g13691(.A(new_n16006), .Y(new_n16040));
  nor_5  g13692(.A(new_n16040), .B(n2570), .Y(new_n16041));
  xnor_4 g13693(.A(new_n16040), .B(n2570), .Y(new_n16042));
  and_5  g13694(.A(new_n16042), .B(n14692), .Y(new_n16043));
  and_5  g13695(.A(new_n16021), .B(new_n16008), .Y(new_n16044));
  nor_5  g13696(.A(new_n16044), .B(new_n16043), .Y(new_n16045));
  xnor_4 g13697(.A(new_n16045), .B(new_n16041), .Y(new_n16046));
  xnor_4 g13698(.A(new_n16046), .B(new_n11846), .Y(new_n16047));
  xnor_4 g13699(.A(new_n16047), .B(new_n16039), .Y(new_n16048));
  nor_5  g13700(.A(new_n16048), .B(new_n10285), .Y(new_n16049));
  xnor_4 g13701(.A(new_n16048), .B(new_n10285), .Y(new_n16050));
  xnor_4 g13702(.A(new_n16037), .B(new_n16024), .Y(new_n16051));
  nor_5  g13703(.A(new_n16051), .B(new_n10342), .Y(new_n16052));
  xnor_4 g13704(.A(new_n16051), .B(new_n10342), .Y(new_n16053));
  xnor_4 g13705(.A(new_n16035), .B(new_n16027), .Y(new_n16054));
  nor_5  g13706(.A(new_n16054), .B(new_n10295_1), .Y(new_n16055));
  xnor_4 g13707(.A(new_n16054), .B(new_n10295_1), .Y(new_n16056));
  xnor_4 g13708(.A(new_n16033), .B(new_n16030), .Y(new_n16057));
  nor_5  g13709(.A(new_n16057), .B(new_n10300), .Y(new_n16058));
  xnor_4 g13710(.A(new_n16057), .B(new_n10299), .Y(new_n16059));
  nor_5  g13711(.A(new_n15427), .B(new_n10304), .Y(new_n16060_1));
  and_5  g13712(.A(new_n15455), .B(new_n15428_1), .Y(new_n16061));
  nor_5  g13713(.A(new_n16061), .B(new_n16060_1), .Y(new_n16062_1));
  and_5  g13714(.A(new_n16062_1), .B(new_n16059), .Y(new_n16063));
  nor_5  g13715(.A(new_n16063), .B(new_n16058), .Y(new_n16064));
  nor_5  g13716(.A(new_n16064), .B(new_n16056), .Y(new_n16065));
  nor_5  g13717(.A(new_n16065), .B(new_n16055), .Y(new_n16066));
  nor_5  g13718(.A(new_n16066), .B(new_n16053), .Y(new_n16067));
  nor_5  g13719(.A(new_n16067), .B(new_n16052), .Y(new_n16068_1));
  nor_5  g13720(.A(new_n16068_1), .B(new_n16050), .Y(new_n16069));
  nor_5  g13721(.A(new_n16069), .B(new_n16049), .Y(new_n16070));
  not_8  g13722(.A(new_n16070), .Y(new_n16071));
  nor_5  g13723(.A(new_n16046), .B(new_n11846), .Y(new_n16072));
  and_5  g13724(.A(new_n16045), .B(new_n16041), .Y(new_n16073));
  nand_5 g13725(.A(new_n16046), .B(new_n11846), .Y(new_n16074));
  and_5  g13726(.A(new_n16074), .B(new_n16039), .Y(new_n16075));
  or_5   g13727(.A(new_n16075), .B(new_n16073), .Y(new_n16076));
  nor_5  g13728(.A(new_n16076), .B(new_n16072), .Y(new_n16077));
  xnor_4 g13729(.A(new_n16077), .B(new_n16071), .Y(n3760));
  xnor_4 g13730(.A(new_n3922), .B(new_n3898), .Y(n3781));
  xnor_4 g13731(.A(new_n13298), .B(new_n13276), .Y(n3794));
  xnor_4 g13732(.A(n9246), .B(new_n3755_1), .Y(new_n16081));
  and_5  g13733(.A(new_n10779), .B(new_n16081), .Y(new_n16082));
  nor_5  g13734(.A(new_n16082), .B(new_n5008), .Y(new_n16083));
  and_5  g13735(.A(new_n16082), .B(new_n4777_1), .Y(new_n16084));
  nor_5  g13736(.A(new_n16084), .B(new_n16083), .Y(new_n16085));
  nor_5  g13737(.A(new_n10778), .B(new_n5956), .Y(new_n16086));
  nor_5  g13738(.A(new_n5956), .B(new_n5897), .Y(new_n16087));
  nor_5  g13739(.A(new_n5959), .B(new_n10777), .Y(new_n16088));
  nor_5  g13740(.A(new_n16088), .B(new_n16087), .Y(new_n16089));
  xnor_4 g13741(.A(new_n16089), .B(new_n12869), .Y(new_n16090));
  xnor_4 g13742(.A(new_n16090), .B(new_n16086), .Y(new_n16091));
  xor_4  g13743(.A(new_n16091), .B(new_n16085), .Y(n3842));
  xnor_4 g13744(.A(new_n12085), .B(new_n8891), .Y(n3850));
  xnor_4 g13745(.A(new_n14469), .B(new_n4297), .Y(n3869));
  xnor_4 g13746(.A(n21749), .B(n919), .Y(new_n16095));
  nor_5  g13747(.A(n25316), .B(n7769), .Y(new_n16096));
  or_5   g13748(.A(new_n9485), .B(new_n4146_1), .Y(new_n16097));
  xnor_4 g13749(.A(n25316), .B(new_n9487), .Y(new_n16098_1));
  and_5  g13750(.A(new_n16098_1), .B(new_n16097), .Y(new_n16099));
  nor_5  g13751(.A(new_n16099), .B(new_n16096), .Y(new_n16100));
  xnor_4 g13752(.A(new_n16100), .B(new_n16095), .Y(new_n16101));
  xnor_4 g13753(.A(new_n16101), .B(n19584), .Y(new_n16102));
  not_8  g13754(.A(n15332), .Y(new_n16103));
  xnor_4 g13755(.A(n21138), .B(new_n4146_1), .Y(new_n16104));
  nor_5  g13756(.A(new_n16104), .B(new_n16103), .Y(new_n16105));
  nor_5  g13757(.A(new_n16105), .B(n5060), .Y(new_n16106));
  xor_4  g13758(.A(new_n16098_1), .B(new_n16097), .Y(new_n16107));
  xnor_4 g13759(.A(new_n16105), .B(n5060), .Y(new_n16108));
  nor_5  g13760(.A(new_n16108), .B(new_n16107), .Y(new_n16109));
  nor_5  g13761(.A(new_n16109), .B(new_n16106), .Y(new_n16110_1));
  xnor_4 g13762(.A(new_n16110_1), .B(new_n16102), .Y(new_n16111));
  xnor_4 g13763(.A(new_n16111), .B(new_n15301), .Y(new_n16112));
  xor_4  g13764(.A(new_n16108), .B(new_n16107), .Y(new_n16113));
  nor_5  g13765(.A(new_n16113), .B(new_n15305), .Y(new_n16114));
  xnor_4 g13766(.A(new_n16104), .B(n15332), .Y(new_n16115));
  nor_5  g13767(.A(new_n16115), .B(new_n15309), .Y(new_n16116));
  xnor_4 g13768(.A(new_n16113), .B(new_n15305), .Y(new_n16117));
  nor_5  g13769(.A(new_n16117), .B(new_n16116), .Y(new_n16118));
  nor_5  g13770(.A(new_n16118), .B(new_n16114), .Y(new_n16119));
  xnor_4 g13771(.A(new_n16119), .B(new_n16112), .Y(n3871));
  xor_4  g13772(.A(new_n15911), .B(new_n15904), .Y(n3891));
  xnor_4 g13773(.A(n10250), .B(n2570), .Y(new_n16122));
  nor_5  g13774(.A(n19033), .B(new_n6155), .Y(new_n16123));
  xnor_4 g13775(.A(n19033), .B(n7674), .Y(new_n16124));
  nor_5  g13776(.A(new_n6158), .B(n655), .Y(new_n16125));
  xnor_4 g13777(.A(n6397), .B(n655), .Y(new_n16126));
  nor_5  g13778(.A(new_n6161), .B(n18145), .Y(new_n16127));
  xnor_4 g13779(.A(n19196), .B(n18145), .Y(new_n16128));
  nor_5  g13780(.A(new_n11812), .B(n10712), .Y(new_n16129));
  xnor_4 g13781(.A(n23586), .B(n10712), .Y(new_n16130));
  nor_5  g13782(.A(n25126), .B(new_n15238), .Y(new_n16131));
  xnor_4 g13783(.A(n25126), .B(n21226), .Y(new_n16132));
  nor_5  g13784(.A(n19608), .B(new_n6170), .Y(new_n16133));
  not_8  g13785(.A(n1689), .Y(new_n16134));
  nor_5  g13786(.A(n20036), .B(new_n16134), .Y(new_n16135));
  or_5   g13787(.A(new_n4125), .B(new_n4119_1), .Y(new_n16136));
  and_5  g13788(.A(new_n16136), .B(new_n4117), .Y(new_n16137));
  nor_5  g13789(.A(new_n16137), .B(new_n16135), .Y(new_n16138));
  xnor_4 g13790(.A(n19608), .B(n4426), .Y(new_n16139));
  and_5  g13791(.A(new_n16139), .B(new_n16138), .Y(new_n16140));
  or_5   g13792(.A(new_n16140), .B(new_n16133), .Y(new_n16141));
  and_5  g13793(.A(new_n16141), .B(new_n16132), .Y(new_n16142_1));
  or_5   g13794(.A(new_n16142_1), .B(new_n16131), .Y(new_n16143));
  and_5  g13795(.A(new_n16143), .B(new_n16130), .Y(new_n16144));
  or_5   g13796(.A(new_n16144), .B(new_n16129), .Y(new_n16145));
  and_5  g13797(.A(new_n16145), .B(new_n16128), .Y(new_n16146));
  or_5   g13798(.A(new_n16146), .B(new_n16127), .Y(new_n16147));
  and_5  g13799(.A(new_n16147), .B(new_n16126), .Y(new_n16148));
  or_5   g13800(.A(new_n16148), .B(new_n16125), .Y(new_n16149));
  and_5  g13801(.A(new_n16149), .B(new_n16124), .Y(new_n16150));
  or_5   g13802(.A(new_n16150), .B(new_n16123), .Y(new_n16151));
  xor_4  g13803(.A(new_n16151), .B(new_n16122), .Y(new_n16152));
  xnor_4 g13804(.A(new_n16152), .B(new_n11802), .Y(new_n16153));
  xor_4  g13805(.A(new_n16149), .B(new_n16124), .Y(new_n16154));
  nor_5  g13806(.A(new_n16154), .B(new_n6864), .Y(new_n16155));
  xnor_4 g13807(.A(new_n16154), .B(new_n6863_1), .Y(new_n16156));
  xor_4  g13808(.A(new_n16147), .B(new_n16126), .Y(new_n16157));
  nor_5  g13809(.A(new_n16157), .B(new_n6869), .Y(new_n16158_1));
  xnor_4 g13810(.A(new_n16157), .B(new_n6867_1), .Y(new_n16159));
  xor_4  g13811(.A(new_n16145), .B(new_n16128), .Y(new_n16160));
  nor_5  g13812(.A(new_n16160), .B(new_n6874), .Y(new_n16161));
  xnor_4 g13813(.A(new_n16160), .B(new_n6872), .Y(new_n16162));
  xor_4  g13814(.A(new_n16143), .B(new_n16130), .Y(new_n16163));
  nor_5  g13815(.A(new_n16163), .B(new_n6879), .Y(new_n16164));
  xnor_4 g13816(.A(new_n16163), .B(new_n6877), .Y(new_n16165));
  xor_4  g13817(.A(new_n16141), .B(new_n16132), .Y(new_n16166));
  nor_5  g13818(.A(new_n16166), .B(new_n6881), .Y(new_n16167_1));
  xnor_4 g13819(.A(new_n16166), .B(new_n6881), .Y(new_n16168));
  xnor_4 g13820(.A(new_n16139), .B(new_n16138), .Y(new_n16169));
  not_8  g13821(.A(new_n16169), .Y(new_n16170));
  nor_5  g13822(.A(new_n16170), .B(new_n6888), .Y(new_n16171));
  xnor_4 g13823(.A(new_n16169), .B(new_n6888), .Y(new_n16172));
  not_8  g13824(.A(new_n4127), .Y(new_n16173));
  nor_5  g13825(.A(new_n16173), .B(new_n4116), .Y(new_n16174));
  and_5  g13826(.A(new_n4141), .B(new_n4128), .Y(new_n16175));
  or_5   g13827(.A(new_n16175), .B(new_n16174), .Y(new_n16176));
  and_5  g13828(.A(new_n16176), .B(new_n16172), .Y(new_n16177));
  nor_5  g13829(.A(new_n16177), .B(new_n16171), .Y(new_n16178));
  nor_5  g13830(.A(new_n16178), .B(new_n16168), .Y(new_n16179));
  or_5   g13831(.A(new_n16179), .B(new_n16167_1), .Y(new_n16180));
  and_5  g13832(.A(new_n16180), .B(new_n16165), .Y(new_n16181));
  or_5   g13833(.A(new_n16181), .B(new_n16164), .Y(new_n16182));
  and_5  g13834(.A(new_n16182), .B(new_n16162), .Y(new_n16183));
  or_5   g13835(.A(new_n16183), .B(new_n16161), .Y(new_n16184));
  and_5  g13836(.A(new_n16184), .B(new_n16159), .Y(new_n16185_1));
  or_5   g13837(.A(new_n16185_1), .B(new_n16158_1), .Y(new_n16186));
  and_5  g13838(.A(new_n16186), .B(new_n16156), .Y(new_n16187));
  nor_5  g13839(.A(new_n16187), .B(new_n16155), .Y(new_n16188));
  xnor_4 g13840(.A(new_n16188), .B(new_n16153), .Y(new_n16189));
  xnor_4 g13841(.A(new_n16189), .B(new_n6361), .Y(new_n16190));
  xor_4  g13842(.A(new_n16186), .B(new_n16156), .Y(new_n16191));
  and_5  g13843(.A(new_n16191), .B(new_n6368), .Y(new_n16192));
  xnor_4 g13844(.A(new_n16191), .B(new_n6368), .Y(new_n16193));
  not_8  g13845(.A(new_n6373), .Y(new_n16194));
  xor_4  g13846(.A(new_n16184), .B(new_n16159), .Y(new_n16195));
  and_5  g13847(.A(new_n16195), .B(new_n16194), .Y(new_n16196_1));
  xnor_4 g13848(.A(new_n16195), .B(new_n16194), .Y(new_n16197));
  xor_4  g13849(.A(new_n16182), .B(new_n16162), .Y(new_n16198));
  and_5  g13850(.A(new_n16198), .B(new_n6377), .Y(new_n16199));
  xnor_4 g13851(.A(new_n16198), .B(new_n6377), .Y(new_n16200));
  xor_4  g13852(.A(new_n16180), .B(new_n16165), .Y(new_n16201));
  and_5  g13853(.A(new_n16201), .B(new_n6382), .Y(new_n16202));
  xnor_4 g13854(.A(new_n16201), .B(new_n6382), .Y(new_n16203));
  xnor_4 g13855(.A(new_n16178), .B(new_n16168), .Y(new_n16204));
  nor_5  g13856(.A(new_n16204), .B(new_n6386), .Y(new_n16205));
  xnor_4 g13857(.A(new_n16204), .B(new_n6386), .Y(new_n16206_1));
  not_8  g13858(.A(new_n6391), .Y(new_n16207));
  xor_4  g13859(.A(new_n16176), .B(new_n16172), .Y(new_n16208));
  and_5  g13860(.A(new_n16208), .B(new_n16207), .Y(new_n16209));
  xnor_4 g13861(.A(new_n16208), .B(new_n16207), .Y(new_n16210));
  nor_5  g13862(.A(new_n4151_1), .B(new_n4142), .Y(new_n16211));
  nor_5  g13863(.A(new_n4163), .B(new_n4152_1), .Y(new_n16212));
  nor_5  g13864(.A(new_n16212), .B(new_n16211), .Y(new_n16213));
  nor_5  g13865(.A(new_n16213), .B(new_n16210), .Y(new_n16214));
  nor_5  g13866(.A(new_n16214), .B(new_n16209), .Y(new_n16215_1));
  nor_5  g13867(.A(new_n16215_1), .B(new_n16206_1), .Y(new_n16216));
  nor_5  g13868(.A(new_n16216), .B(new_n16205), .Y(new_n16217_1));
  nor_5  g13869(.A(new_n16217_1), .B(new_n16203), .Y(new_n16218_1));
  nor_5  g13870(.A(new_n16218_1), .B(new_n16202), .Y(new_n16219_1));
  nor_5  g13871(.A(new_n16219_1), .B(new_n16200), .Y(new_n16220));
  nor_5  g13872(.A(new_n16220), .B(new_n16199), .Y(new_n16221));
  nor_5  g13873(.A(new_n16221), .B(new_n16197), .Y(new_n16222));
  nor_5  g13874(.A(new_n16222), .B(new_n16196_1), .Y(new_n16223_1));
  nor_5  g13875(.A(new_n16223_1), .B(new_n16193), .Y(new_n16224));
  nor_5  g13876(.A(new_n16224), .B(new_n16192), .Y(new_n16225));
  xnor_4 g13877(.A(new_n16225), .B(new_n16190), .Y(n3932));
  xnor_4 g13878(.A(new_n3916), .B(new_n3915), .Y(n3934));
  xnor_4 g13879(.A(new_n4096), .B(new_n4095), .Y(n3971));
  nor_5  g13880(.A(n8581), .B(n5026), .Y(new_n16229));
  not_8  g13881(.A(new_n16229), .Y(new_n16230_1));
  nor_5  g13882(.A(new_n16230_1), .B(n12161), .Y(new_n16231));
  not_8  g13883(.A(new_n16231), .Y(new_n16232));
  nor_5  g13884(.A(new_n16232), .B(n18157), .Y(new_n16233));
  not_8  g13885(.A(new_n16233), .Y(new_n16234));
  nor_5  g13886(.A(new_n16234), .B(n20923), .Y(new_n16235));
  not_8  g13887(.A(new_n16235), .Y(new_n16236));
  nor_5  g13888(.A(new_n16236), .B(n8067), .Y(new_n16237));
  not_8  g13889(.A(new_n16237), .Y(new_n16238));
  nor_5  g13890(.A(new_n16238), .B(n10125), .Y(new_n16239));
  not_8  g13891(.A(new_n16239), .Y(new_n16240));
  nor_5  g13892(.A(new_n16240), .B(n25240), .Y(new_n16241));
  xnor_4 g13893(.A(new_n16241), .B(n1222), .Y(new_n16242));
  xnor_4 g13894(.A(new_n16242), .B(new_n8789), .Y(new_n16243_1));
  xnor_4 g13895(.A(new_n16239), .B(n25240), .Y(new_n16244));
  nor_5  g13896(.A(new_n16244), .B(n3710), .Y(new_n16245));
  xnor_4 g13897(.A(new_n16244), .B(new_n9992), .Y(new_n16246));
  xnor_4 g13898(.A(new_n16237), .B(n10125), .Y(new_n16247_1));
  and_5  g13899(.A(new_n16247_1), .B(n26318), .Y(new_n16248));
  or_5   g13900(.A(new_n16247_1), .B(n26318), .Y(new_n16249));
  xnor_4 g13901(.A(new_n16235), .B(n8067), .Y(new_n16250));
  nor_5  g13902(.A(new_n16250), .B(n26054), .Y(new_n16251));
  xnor_4 g13903(.A(new_n16250), .B(new_n8749), .Y(new_n16252));
  xnor_4 g13904(.A(new_n16233), .B(n20923), .Y(new_n16253));
  nor_5  g13905(.A(new_n16253), .B(n19081), .Y(new_n16254));
  xnor_4 g13906(.A(new_n16253), .B(new_n8753), .Y(new_n16255));
  xnor_4 g13907(.A(new_n16231), .B(n18157), .Y(new_n16256));
  nor_5  g13908(.A(new_n16256), .B(n8309), .Y(new_n16257));
  xnor_4 g13909(.A(new_n16229), .B(n12161), .Y(new_n16258));
  nor_5  g13910(.A(new_n16258), .B(n19144), .Y(new_n16259));
  xnor_4 g13911(.A(new_n16258), .B(new_n8759), .Y(new_n16260));
  xnor_4 g13912(.A(n8581), .B(new_n7220), .Y(new_n16261));
  nor_5  g13913(.A(new_n16261), .B(n12593), .Y(new_n16262));
  or_5   g13914(.A(new_n8763), .B(new_n6628_1), .Y(new_n16263));
  xnor_4 g13915(.A(new_n16261), .B(new_n10007), .Y(new_n16264));
  and_5  g13916(.A(new_n16264), .B(new_n16263), .Y(new_n16265));
  or_5   g13917(.A(new_n16265), .B(new_n16262), .Y(new_n16266));
  and_5  g13918(.A(new_n16266), .B(new_n16260), .Y(new_n16267));
  or_5   g13919(.A(new_n16267), .B(new_n16259), .Y(new_n16268));
  xnor_4 g13920(.A(new_n16256), .B(new_n8771), .Y(new_n16269));
  and_5  g13921(.A(new_n16269), .B(new_n16268), .Y(new_n16270));
  or_5   g13922(.A(new_n16270), .B(new_n16257), .Y(new_n16271));
  and_5  g13923(.A(new_n16271), .B(new_n16255), .Y(new_n16272));
  or_5   g13924(.A(new_n16272), .B(new_n16254), .Y(new_n16273));
  and_5  g13925(.A(new_n16273), .B(new_n16252), .Y(new_n16274));
  nor_5  g13926(.A(new_n16274), .B(new_n16251), .Y(new_n16275_1));
  and_5  g13927(.A(new_n16275_1), .B(new_n16249), .Y(new_n16276));
  nor_5  g13928(.A(new_n16276), .B(new_n16248), .Y(new_n16277));
  and_5  g13929(.A(new_n16277), .B(new_n16246), .Y(new_n16278));
  or_5   g13930(.A(new_n16278), .B(new_n16245), .Y(new_n16279_1));
  xor_4  g13931(.A(new_n16279_1), .B(new_n16243_1), .Y(new_n16280));
  xnor_4 g13932(.A(new_n16280), .B(n26797), .Y(new_n16281));
  xnor_4 g13933(.A(new_n16277), .B(new_n16246), .Y(new_n16282));
  not_8  g13934(.A(new_n16282), .Y(new_n16283));
  nor_5  g13935(.A(new_n16283), .B(new_n8033), .Y(new_n16284));
  xnor_4 g13936(.A(new_n16283), .B(n23913), .Y(new_n16285));
  xnor_4 g13937(.A(new_n16247_1), .B(new_n8745_1), .Y(new_n16286));
  xnor_4 g13938(.A(new_n16286), .B(new_n16275_1), .Y(new_n16287));
  nor_5  g13939(.A(new_n16287), .B(new_n8036), .Y(new_n16288));
  not_8  g13940(.A(new_n16287), .Y(new_n16289));
  xnor_4 g13941(.A(new_n16289), .B(new_n8036), .Y(new_n16290));
  nor_5  g13942(.A(new_n16272), .B(new_n16254), .Y(new_n16291));
  xnor_4 g13943(.A(new_n16291), .B(new_n16252), .Y(new_n16292));
  nor_5  g13944(.A(new_n16292), .B(new_n8039), .Y(new_n16293));
  not_8  g13945(.A(new_n16292), .Y(new_n16294));
  xnor_4 g13946(.A(new_n16294), .B(new_n8039), .Y(new_n16295));
  xor_4  g13947(.A(new_n16271), .B(new_n16255), .Y(new_n16296));
  nor_5  g13948(.A(new_n16296), .B(new_n8042_1), .Y(new_n16297));
  xnor_4 g13949(.A(new_n16296), .B(n3909), .Y(new_n16298));
  xor_4  g13950(.A(new_n16269), .B(new_n16268), .Y(new_n16299));
  nor_5  g13951(.A(new_n16299), .B(new_n8045), .Y(new_n16300));
  xnor_4 g13952(.A(new_n16299), .B(n23974), .Y(new_n16301));
  xor_4  g13953(.A(new_n16266), .B(new_n16260), .Y(new_n16302));
  nor_5  g13954(.A(new_n16302), .B(new_n8050), .Y(new_n16303));
  xnor_4 g13955(.A(new_n16302), .B(n2146), .Y(new_n16304));
  xor_4  g13956(.A(new_n16264), .B(new_n16263), .Y(new_n16305));
  nor_5  g13957(.A(new_n16305), .B(new_n8055), .Y(new_n16306));
  xnor_4 g13958(.A(n13714), .B(n8581), .Y(new_n16307));
  nor_5  g13959(.A(new_n16307), .B(new_n5587), .Y(new_n16308));
  xnor_4 g13960(.A(new_n16305), .B(n22173), .Y(new_n16309));
  and_5  g13961(.A(new_n16309), .B(new_n16308), .Y(new_n16310));
  or_5   g13962(.A(new_n16310), .B(new_n16306), .Y(new_n16311));
  and_5  g13963(.A(new_n16311), .B(new_n16304), .Y(new_n16312));
  or_5   g13964(.A(new_n16312), .B(new_n16303), .Y(new_n16313));
  and_5  g13965(.A(new_n16313), .B(new_n16301), .Y(new_n16314));
  or_5   g13966(.A(new_n16314), .B(new_n16300), .Y(new_n16315));
  and_5  g13967(.A(new_n16315), .B(new_n16298), .Y(new_n16316));
  or_5   g13968(.A(new_n16316), .B(new_n16297), .Y(new_n16317));
  and_5  g13969(.A(new_n16317), .B(new_n16295), .Y(new_n16318));
  or_5   g13970(.A(new_n16318), .B(new_n16293), .Y(new_n16319));
  and_5  g13971(.A(new_n16319), .B(new_n16290), .Y(new_n16320));
  or_5   g13972(.A(new_n16320), .B(new_n16288), .Y(new_n16321));
  and_5  g13973(.A(new_n16321), .B(new_n16285), .Y(new_n16322_1));
  nor_5  g13974(.A(new_n16322_1), .B(new_n16284), .Y(new_n16323));
  xnor_4 g13975(.A(new_n16323), .B(new_n16281), .Y(new_n16324));
  xnor_4 g13976(.A(new_n16324), .B(new_n8144), .Y(new_n16325));
  xor_4  g13977(.A(new_n16321), .B(new_n16285), .Y(new_n16326));
  nor_5  g13978(.A(new_n16326), .B(new_n8149_1), .Y(new_n16327_1));
  xnor_4 g13979(.A(new_n16326), .B(new_n8149_1), .Y(new_n16328));
  xor_4  g13980(.A(new_n16319), .B(new_n16290), .Y(new_n16329));
  nor_5  g13981(.A(new_n16329), .B(new_n8154), .Y(new_n16330));
  xnor_4 g13982(.A(new_n16329), .B(new_n8154), .Y(new_n16331));
  not_8  g13983(.A(new_n8159_1), .Y(new_n16332));
  xor_4  g13984(.A(new_n16317), .B(new_n16295), .Y(new_n16333));
  nor_5  g13985(.A(new_n16333), .B(new_n16332), .Y(new_n16334));
  xnor_4 g13986(.A(new_n16333), .B(new_n16332), .Y(new_n16335));
  xor_4  g13987(.A(new_n16315), .B(new_n16298), .Y(new_n16336));
  nor_5  g13988(.A(new_n16336), .B(new_n8164), .Y(new_n16337));
  xnor_4 g13989(.A(new_n16336), .B(new_n8164), .Y(new_n16338));
  xor_4  g13990(.A(new_n16313), .B(new_n16301), .Y(new_n16339));
  nor_5  g13991(.A(new_n16339), .B(new_n8168), .Y(new_n16340));
  xnor_4 g13992(.A(new_n16339), .B(new_n8168), .Y(new_n16341));
  xor_4  g13993(.A(new_n16311), .B(new_n16304), .Y(new_n16342));
  nor_5  g13994(.A(new_n16342), .B(new_n8173), .Y(new_n16343));
  xor_4  g13995(.A(new_n16309), .B(new_n16308), .Y(new_n16344));
  nor_5  g13996(.A(new_n16344), .B(new_n8183), .Y(new_n16345));
  xnor_4 g13997(.A(new_n16307), .B(n583), .Y(new_n16346));
  and_5  g13998(.A(new_n16346), .B(new_n8181), .Y(new_n16347));
  xnor_4 g13999(.A(new_n16344), .B(new_n8183), .Y(new_n16348));
  nor_5  g14000(.A(new_n16348), .B(new_n16347), .Y(new_n16349));
  nor_5  g14001(.A(new_n16349), .B(new_n16345), .Y(new_n16350_1));
  xnor_4 g14002(.A(new_n16342), .B(new_n8173), .Y(new_n16351));
  nor_5  g14003(.A(new_n16351), .B(new_n16350_1), .Y(new_n16352));
  nor_5  g14004(.A(new_n16352), .B(new_n16343), .Y(new_n16353));
  nor_5  g14005(.A(new_n16353), .B(new_n16341), .Y(new_n16354));
  nor_5  g14006(.A(new_n16354), .B(new_n16340), .Y(new_n16355));
  nor_5  g14007(.A(new_n16355), .B(new_n16338), .Y(new_n16356));
  nor_5  g14008(.A(new_n16356), .B(new_n16337), .Y(new_n16357));
  nor_5  g14009(.A(new_n16357), .B(new_n16335), .Y(new_n16358));
  nor_5  g14010(.A(new_n16358), .B(new_n16334), .Y(new_n16359));
  nor_5  g14011(.A(new_n16359), .B(new_n16331), .Y(new_n16360));
  nor_5  g14012(.A(new_n16360), .B(new_n16330), .Y(new_n16361));
  nor_5  g14013(.A(new_n16361), .B(new_n16328), .Y(new_n16362));
  nor_5  g14014(.A(new_n16362), .B(new_n16327_1), .Y(new_n16363));
  xnor_4 g14015(.A(new_n16363), .B(new_n16325), .Y(n3983));
  not_8  g14016(.A(new_n6666), .Y(new_n16365));
  xnor_4 g14017(.A(n13714), .B(n583), .Y(new_n16366));
  xnor_4 g14018(.A(new_n16366), .B(n6611), .Y(new_n16367_1));
  nor_5  g14019(.A(new_n16367_1), .B(new_n16365), .Y(new_n16368));
  or_5   g14020(.A(new_n16366), .B(new_n5588), .Y(new_n16369));
  nor_5  g14021(.A(new_n8763), .B(new_n5587), .Y(new_n16370));
  xnor_4 g14022(.A(n22173), .B(n12593), .Y(new_n16371));
  xnor_4 g14023(.A(new_n16371), .B(new_n16370), .Y(new_n16372));
  xnor_4 g14024(.A(new_n16372), .B(new_n5584), .Y(new_n16373));
  xor_4  g14025(.A(new_n16373), .B(new_n16369), .Y(new_n16374));
  xnor_4 g14026(.A(new_n16374), .B(new_n16368), .Y(new_n16375));
  xnor_4 g14027(.A(new_n16375), .B(new_n6662), .Y(n4000));
  xnor_4 g14028(.A(n26823), .B(n20179), .Y(new_n16377));
  nor_5  g14029(.A(n19228), .B(new_n5280), .Y(new_n16378));
  xnor_4 g14030(.A(n19228), .B(n4812), .Y(new_n16379_1));
  nor_5  g14031(.A(new_n8394), .B(n15539), .Y(new_n16380));
  xnor_4 g14032(.A(n24278), .B(n15539), .Y(new_n16381));
  nor_5  g14033(.A(new_n8398), .B(n8052), .Y(new_n16382));
  or_5   g14034(.A(n24618), .B(new_n6767), .Y(new_n16383));
  nor_5  g14035(.A(new_n7448), .B(n3952), .Y(new_n16384));
  and_5  g14036(.A(new_n11150), .B(new_n11149), .Y(new_n16385));
  nor_5  g14037(.A(new_n16385), .B(new_n16384), .Y(new_n16386));
  and_5  g14038(.A(new_n16386), .B(new_n16383), .Y(new_n16387));
  or_5   g14039(.A(new_n16387), .B(new_n16382), .Y(new_n16388));
  and_5  g14040(.A(new_n16388), .B(new_n16381), .Y(new_n16389));
  or_5   g14041(.A(new_n16389), .B(new_n16380), .Y(new_n16390));
  and_5  g14042(.A(new_n16390), .B(new_n16379_1), .Y(new_n16391));
  or_5   g14043(.A(new_n16391), .B(new_n16378), .Y(new_n16392));
  xor_4  g14044(.A(new_n16392), .B(new_n16377), .Y(new_n16393));
  xnor_4 g14045(.A(new_n16393), .B(new_n7381), .Y(new_n16394));
  xor_4  g14046(.A(new_n16390), .B(new_n16379_1), .Y(new_n16395));
  nor_5  g14047(.A(new_n16395), .B(new_n7385), .Y(new_n16396_1));
  xnor_4 g14048(.A(new_n16395), .B(new_n7385), .Y(new_n16397));
  not_8  g14049(.A(new_n7389), .Y(new_n16398_1));
  xor_4  g14050(.A(new_n16388), .B(new_n16381), .Y(new_n16399));
  nor_5  g14051(.A(new_n16399), .B(new_n16398_1), .Y(new_n16400));
  xnor_4 g14052(.A(n24618), .B(n8052), .Y(new_n16401));
  xnor_4 g14053(.A(new_n16401), .B(new_n16386), .Y(new_n16402));
  and_5  g14054(.A(new_n16402), .B(new_n7393), .Y(new_n16403));
  xnor_4 g14055(.A(new_n16402), .B(new_n7392), .Y(new_n16404));
  and_5  g14056(.A(new_n11151), .B(new_n11148), .Y(new_n16405));
  nor_5  g14057(.A(new_n11152), .B(new_n7406), .Y(new_n16406_1));
  nor_5  g14058(.A(new_n16406_1), .B(new_n16405), .Y(new_n16407_1));
  and_5  g14059(.A(new_n16407_1), .B(new_n16404), .Y(new_n16408));
  nor_5  g14060(.A(new_n16408), .B(new_n16403), .Y(new_n16409));
  xnor_4 g14061(.A(new_n16399), .B(new_n16398_1), .Y(new_n16410));
  nor_5  g14062(.A(new_n16410), .B(new_n16409), .Y(new_n16411));
  nor_5  g14063(.A(new_n16411), .B(new_n16400), .Y(new_n16412));
  nor_5  g14064(.A(new_n16412), .B(new_n16397), .Y(new_n16413));
  nor_5  g14065(.A(new_n16413), .B(new_n16396_1), .Y(new_n16414));
  xnor_4 g14066(.A(new_n16414), .B(new_n16394), .Y(n4010));
  xnor_4 g14067(.A(n11220), .B(n2160), .Y(new_n16416));
  nor_5  g14068(.A(n22379), .B(new_n11674_1), .Y(new_n16417));
  xnor_4 g14069(.A(n22379), .B(n10763), .Y(new_n16418));
  nor_5  g14070(.A(new_n2890), .B(n1662), .Y(new_n16419_1));
  xnor_4 g14071(.A(n7437), .B(n1662), .Y(new_n16420));
  nor_5  g14072(.A(new_n2893), .B(n12875), .Y(new_n16421));
  nor_5  g14073(.A(new_n2896), .B(n2035), .Y(new_n16422));
  and_5  g14074(.A(new_n14433), .B(new_n14415), .Y(new_n16423));
  or_5   g14075(.A(new_n16423), .B(new_n16422), .Y(new_n16424_1));
  xnor_4 g14076(.A(n20700), .B(n12875), .Y(new_n16425));
  and_5  g14077(.A(new_n16425), .B(new_n16424_1), .Y(new_n16426));
  or_5   g14078(.A(new_n16426), .B(new_n16421), .Y(new_n16427));
  and_5  g14079(.A(new_n16427), .B(new_n16420), .Y(new_n16428_1));
  or_5   g14080(.A(new_n16428_1), .B(new_n16419_1), .Y(new_n16429));
  and_5  g14081(.A(new_n16429), .B(new_n16418), .Y(new_n16430));
  or_5   g14082(.A(new_n16430), .B(new_n16417), .Y(new_n16431));
  xor_4  g14083(.A(new_n16431), .B(new_n16416), .Y(new_n16432));
  xnor_4 g14084(.A(new_n16432), .B(new_n14588), .Y(new_n16433_1));
  xor_4  g14085(.A(new_n16429), .B(new_n16418), .Y(new_n16434));
  nor_5  g14086(.A(new_n16434), .B(new_n14597), .Y(new_n16435));
  xnor_4 g14087(.A(new_n16434), .B(new_n14597), .Y(new_n16436));
  xor_4  g14088(.A(new_n16427), .B(new_n16420), .Y(new_n16437));
  nor_5  g14089(.A(new_n16437), .B(new_n14601), .Y(new_n16438));
  xor_4  g14090(.A(new_n16425), .B(new_n16424_1), .Y(new_n16439_1));
  not_8  g14091(.A(new_n16439_1), .Y(new_n16440_1));
  nor_5  g14092(.A(new_n16440_1), .B(new_n14606), .Y(new_n16441));
  xnor_4 g14093(.A(new_n16439_1), .B(new_n14606), .Y(new_n16442));
  and_5  g14094(.A(new_n14451), .B(new_n14434), .Y(new_n16443));
  and_5  g14095(.A(new_n14478), .B(new_n14453), .Y(new_n16444));
  or_5   g14096(.A(new_n16444), .B(new_n16443), .Y(new_n16445_1));
  and_5  g14097(.A(new_n16445_1), .B(new_n16442), .Y(new_n16446));
  nor_5  g14098(.A(new_n16446), .B(new_n16441), .Y(new_n16447));
  xnor_4 g14099(.A(new_n16437), .B(new_n14604), .Y(new_n16448));
  and_5  g14100(.A(new_n16448), .B(new_n16447), .Y(new_n16449));
  nor_5  g14101(.A(new_n16449), .B(new_n16438), .Y(new_n16450));
  nor_5  g14102(.A(new_n16450), .B(new_n16436), .Y(new_n16451));
  nor_5  g14103(.A(new_n16451), .B(new_n16435), .Y(new_n16452));
  xor_4  g14104(.A(new_n16452), .B(new_n16433_1), .Y(n4014));
  xnor_4 g14105(.A(new_n13881), .B(new_n11636), .Y(new_n16454));
  nor_5  g14106(.A(new_n13884), .B(n26224), .Y(new_n16455));
  xnor_4 g14107(.A(new_n13884), .B(new_n12526), .Y(new_n16456));
  nor_5  g14108(.A(new_n3736), .B(n19327), .Y(new_n16457));
  or_5   g14109(.A(new_n3769), .B(new_n3739), .Y(new_n16458));
  and_5  g14110(.A(new_n16458), .B(new_n3737), .Y(new_n16459));
  or_5   g14111(.A(new_n16459), .B(new_n16457), .Y(new_n16460_1));
  and_5  g14112(.A(new_n16460_1), .B(new_n16456), .Y(new_n16461));
  nor_5  g14113(.A(new_n16461), .B(new_n16455), .Y(new_n16462));
  xnor_4 g14114(.A(new_n16462), .B(new_n16454), .Y(new_n16463));
  not_8  g14115(.A(new_n16463), .Y(new_n16464));
  xnor_4 g14116(.A(new_n16464), .B(new_n4801), .Y(new_n16465));
  nor_5  g14117(.A(new_n16459), .B(new_n16457), .Y(new_n16466));
  xnor_4 g14118(.A(new_n16466), .B(new_n16456), .Y(new_n16467));
  nor_5  g14119(.A(new_n16467), .B(new_n7328), .Y(new_n16468));
  not_8  g14120(.A(new_n16467), .Y(new_n16469));
  xnor_4 g14121(.A(new_n16469), .B(new_n7328), .Y(new_n16470));
  nor_5  g14122(.A(new_n3771), .B(new_n3725_1), .Y(new_n16471));
  and_5  g14123(.A(new_n3812), .B(new_n3773), .Y(new_n16472));
  or_5   g14124(.A(new_n16472), .B(new_n16471), .Y(new_n16473));
  and_5  g14125(.A(new_n16473), .B(new_n16470), .Y(new_n16474));
  or_5   g14126(.A(new_n16474), .B(new_n16468), .Y(new_n16475));
  xor_4  g14127(.A(new_n16475), .B(new_n16465), .Y(new_n16476_1));
  xnor_4 g14128(.A(new_n16476_1), .B(new_n11745), .Y(new_n16477));
  xor_4  g14129(.A(new_n16473), .B(new_n16470), .Y(new_n16478));
  nor_5  g14130(.A(new_n16478), .B(new_n11750), .Y(new_n16479));
  xnor_4 g14131(.A(new_n16478), .B(new_n11750), .Y(new_n16480));
  nor_5  g14132(.A(new_n3889), .B(new_n3813), .Y(new_n16481_1));
  nor_5  g14133(.A(new_n3926), .B(new_n3890), .Y(new_n16482_1));
  nor_5  g14134(.A(new_n16482_1), .B(new_n16481_1), .Y(new_n16483));
  nor_5  g14135(.A(new_n16483), .B(new_n16480), .Y(new_n16484));
  nor_5  g14136(.A(new_n16484), .B(new_n16479), .Y(new_n16485));
  xnor_4 g14137(.A(new_n16485), .B(new_n16477), .Y(n4071));
  xnor_4 g14138(.A(new_n12718), .B(new_n12713), .Y(n4088));
  not_8  g14139(.A(n7593), .Y(new_n16488));
  and_5  g14140(.A(new_n12826), .B(new_n16488), .Y(new_n16489));
  nor_5  g14141(.A(new_n12827), .B(n5025), .Y(new_n16490));
  and_5  g14142(.A(new_n12827), .B(n5025), .Y(new_n16491));
  nor_5  g14143(.A(new_n12831), .B(new_n16491), .Y(new_n16492));
  nor_5  g14144(.A(new_n16492), .B(new_n16490), .Y(new_n16493_1));
  nor_5  g14145(.A(new_n16493_1), .B(new_n16489), .Y(new_n16494));
  not_8  g14146(.A(new_n16494), .Y(new_n16495));
  not_8  g14147(.A(new_n15927), .Y(new_n16496));
  nor_5  g14148(.A(new_n15930), .B(new_n16496), .Y(new_n16497));
  and_5  g14149(.A(new_n15930), .B(new_n16496), .Y(new_n16498));
  nor_5  g14150(.A(new_n15935), .B(new_n16498), .Y(new_n16499));
  nor_5  g14151(.A(new_n16499), .B(new_n16497), .Y(new_n16500));
  not_8  g14152(.A(new_n16500), .Y(new_n16501));
  nor_5  g14153(.A(new_n16501), .B(new_n16495), .Y(new_n16502_1));
  not_8  g14154(.A(new_n15936_1), .Y(new_n16503));
  nor_5  g14155(.A(new_n16494), .B(new_n16503), .Y(new_n16504));
  or_5   g14156(.A(new_n16495), .B(new_n15936_1), .Y(new_n16505));
  nor_5  g14157(.A(new_n12832), .B(new_n12823), .Y(new_n16506_1));
  and_5  g14158(.A(new_n12836), .B(new_n12833), .Y(new_n16507_1));
  nor_5  g14159(.A(new_n16507_1), .B(new_n16506_1), .Y(new_n16508));
  and_5  g14160(.A(new_n16508), .B(new_n16505), .Y(new_n16509));
  nor_5  g14161(.A(new_n16509), .B(new_n16504), .Y(new_n16510));
  nor_5  g14162(.A(new_n16510), .B(new_n16502_1), .Y(new_n16511));
  nor_5  g14163(.A(new_n16500), .B(new_n16494), .Y(new_n16512));
  nor_5  g14164(.A(new_n16512), .B(new_n16509), .Y(new_n16513));
  nor_5  g14165(.A(new_n16513), .B(new_n16511), .Y(n4089));
  not_8  g14166(.A(new_n11950), .Y(new_n16515));
  nor_5  g14167(.A(new_n16515), .B(n1112), .Y(new_n16516_1));
  xnor_4 g14168(.A(new_n16516_1), .B(n2289), .Y(new_n16517_1));
  not_8  g14169(.A(new_n16517_1), .Y(new_n16518));
  xnor_4 g14170(.A(new_n16518), .B(n3228), .Y(new_n16519));
  nor_5  g14171(.A(new_n11951), .B(n5302), .Y(new_n16520));
  xnor_4 g14172(.A(new_n11951), .B(n5302), .Y(new_n16521_1));
  and_5  g14173(.A(new_n11954), .B(n25738), .Y(new_n16522));
  or_5   g14174(.A(new_n11954), .B(n25738), .Y(new_n16523));
  nor_5  g14175(.A(new_n8578), .B(n21471), .Y(new_n16524_1));
  not_8  g14176(.A(new_n8598), .Y(new_n16525));
  nor_5  g14177(.A(new_n16525), .B(new_n8579), .Y(new_n16526));
  nor_5  g14178(.A(new_n16526), .B(new_n16524_1), .Y(new_n16527_1));
  and_5  g14179(.A(new_n16527_1), .B(new_n16523), .Y(new_n16528));
  nor_5  g14180(.A(new_n16528), .B(new_n16522), .Y(new_n16529));
  not_8  g14181(.A(new_n16529), .Y(new_n16530));
  nor_5  g14182(.A(new_n16530), .B(new_n16521_1), .Y(new_n16531));
  nor_5  g14183(.A(new_n16531), .B(new_n16520), .Y(new_n16532));
  xnor_4 g14184(.A(new_n16532), .B(new_n16519), .Y(new_n16533));
  not_8  g14185(.A(new_n16533), .Y(new_n16534));
  xnor_4 g14186(.A(new_n16534), .B(n13775), .Y(new_n16535));
  xnor_4 g14187(.A(new_n16529), .B(new_n16521_1), .Y(new_n16536));
  not_8  g14188(.A(new_n16536), .Y(new_n16537));
  nor_5  g14189(.A(new_n16537), .B(n1293), .Y(new_n16538));
  xnor_4 g14190(.A(new_n16537), .B(new_n6839), .Y(new_n16539));
  xnor_4 g14191(.A(new_n11955), .B(n25738), .Y(new_n16540));
  xnor_4 g14192(.A(new_n16540), .B(new_n16527_1), .Y(new_n16541));
  nor_5  g14193(.A(new_n16541), .B(new_n6842), .Y(new_n16542));
  nor_5  g14194(.A(new_n8599), .B(new_n8572), .Y(new_n16543));
  and_5  g14195(.A(new_n8622), .B(new_n8601), .Y(new_n16544_1));
  or_5   g14196(.A(new_n16544_1), .B(new_n16543), .Y(new_n16545));
  xnor_4 g14197(.A(new_n16541), .B(n19042), .Y(new_n16546));
  and_5  g14198(.A(new_n16546), .B(new_n16545), .Y(new_n16547));
  nor_5  g14199(.A(new_n16547), .B(new_n16542), .Y(new_n16548));
  and_5  g14200(.A(new_n16548), .B(new_n16539), .Y(new_n16549));
  nor_5  g14201(.A(new_n16549), .B(new_n16538), .Y(new_n16550));
  xnor_4 g14202(.A(new_n16550), .B(new_n16535), .Y(new_n16551));
  xnor_4 g14203(.A(new_n7533), .B(new_n5459), .Y(new_n16552));
  nor_5  g14204(.A(new_n2460), .B(new_n5462), .Y(new_n16553));
  xnor_4 g14205(.A(new_n2460), .B(new_n5462), .Y(new_n16554_1));
  nor_5  g14206(.A(new_n2463), .B(new_n5465), .Y(new_n16555));
  xnor_4 g14207(.A(new_n2463), .B(new_n5465), .Y(new_n16556));
  nor_5  g14208(.A(new_n2466), .B(new_n5468), .Y(new_n16557));
  nor_5  g14209(.A(new_n6695), .B(new_n6681), .Y(new_n16558));
  nor_5  g14210(.A(new_n16558), .B(new_n16557), .Y(new_n16559));
  nor_5  g14211(.A(new_n16559), .B(new_n16556), .Y(new_n16560));
  nor_5  g14212(.A(new_n16560), .B(new_n16555), .Y(new_n16561));
  nor_5  g14213(.A(new_n16561), .B(new_n16554_1), .Y(new_n16562));
  nor_5  g14214(.A(new_n16562), .B(new_n16553), .Y(new_n16563));
  xor_4  g14215(.A(new_n16563), .B(new_n16552), .Y(new_n16564));
  xnor_4 g14216(.A(new_n16564), .B(new_n16551), .Y(new_n16565));
  xnor_4 g14217(.A(new_n16548), .B(new_n16539), .Y(new_n16566));
  xor_4  g14218(.A(new_n16561), .B(new_n16554_1), .Y(new_n16567));
  nor_5  g14219(.A(new_n16567), .B(new_n16566), .Y(new_n16568));
  xnor_4 g14220(.A(new_n16567), .B(new_n16566), .Y(new_n16569));
  xnor_4 g14221(.A(new_n16559), .B(new_n16556), .Y(new_n16570));
  not_8  g14222(.A(new_n16570), .Y(new_n16571));
  xor_4  g14223(.A(new_n16546), .B(new_n16545), .Y(new_n16572));
  nor_5  g14224(.A(new_n16572), .B(new_n16571), .Y(new_n16573));
  nor_5  g14225(.A(new_n8623), .B(new_n6696), .Y(new_n16574));
  nor_5  g14226(.A(new_n8643), .B(new_n8624), .Y(new_n16575));
  nor_5  g14227(.A(new_n16575), .B(new_n16574), .Y(new_n16576));
  xnor_4 g14228(.A(new_n16572), .B(new_n16571), .Y(new_n16577));
  nor_5  g14229(.A(new_n16577), .B(new_n16576), .Y(new_n16578));
  nor_5  g14230(.A(new_n16578), .B(new_n16573), .Y(new_n16579));
  nor_5  g14231(.A(new_n16579), .B(new_n16569), .Y(new_n16580));
  nor_5  g14232(.A(new_n16580), .B(new_n16568), .Y(new_n16581));
  xnor_4 g14233(.A(new_n16581), .B(new_n16565), .Y(n4103));
  nor_5  g14234(.A(new_n14513), .B(new_n12595), .Y(new_n16583_1));
  xnor_4 g14235(.A(new_n14514), .B(new_n12595), .Y(new_n16584_1));
  not_8  g14236(.A(new_n12518), .Y(new_n16585));
  nor_5  g14237(.A(new_n14518), .B(new_n16585), .Y(new_n16586));
  not_8  g14238(.A(new_n12523), .Y(new_n16587));
  nor_5  g14239(.A(new_n14522), .B(new_n16587), .Y(new_n16588));
  xnor_4 g14240(.A(new_n14522), .B(new_n12523), .Y(new_n16589_1));
  and_5  g14241(.A(new_n14526), .B(new_n12528), .Y(new_n16590));
  xnor_4 g14242(.A(new_n14526), .B(new_n12528), .Y(new_n16591));
  not_8  g14243(.A(new_n12533), .Y(new_n16592));
  nor_5  g14244(.A(new_n14529), .B(new_n16592), .Y(new_n16593));
  xnor_4 g14245(.A(new_n14529), .B(new_n12533), .Y(new_n16594));
  and_5  g14246(.A(new_n14445), .B(new_n12537), .Y(new_n16595));
  nor_5  g14247(.A(new_n12545_1), .B(new_n4251), .Y(new_n16596_1));
  xnor_4 g14248(.A(new_n12545_1), .B(new_n14447), .Y(new_n16597));
  nor_5  g14249(.A(new_n12550), .B(new_n4258), .Y(new_n16598));
  xnor_4 g14250(.A(new_n12550), .B(new_n4257), .Y(new_n16599));
  nor_5  g14251(.A(new_n12554), .B(new_n4277), .Y(new_n16600));
  xnor_4 g14252(.A(new_n12553), .B(new_n4277), .Y(new_n16601));
  not_8  g14253(.A(new_n4264), .Y(new_n16602));
  nor_5  g14254(.A(new_n12565), .B(new_n16602), .Y(new_n16603));
  or_5   g14255(.A(new_n12563), .B(new_n4266_1), .Y(new_n16604));
  xnor_4 g14256(.A(new_n12560), .B(new_n16602), .Y(new_n16605));
  and_5  g14257(.A(new_n16605), .B(new_n16604), .Y(new_n16606));
  or_5   g14258(.A(new_n16606), .B(new_n16603), .Y(new_n16607));
  and_5  g14259(.A(new_n16607), .B(new_n16601), .Y(new_n16608_1));
  nor_5  g14260(.A(new_n16608_1), .B(new_n16600), .Y(new_n16609));
  and_5  g14261(.A(new_n16609), .B(new_n16599), .Y(new_n16610));
  nor_5  g14262(.A(new_n16610), .B(new_n16598), .Y(new_n16611));
  and_5  g14263(.A(new_n16611), .B(new_n16597), .Y(new_n16612));
  nor_5  g14264(.A(new_n16612), .B(new_n16596_1), .Y(new_n16613));
  xnor_4 g14265(.A(new_n14445), .B(new_n12537), .Y(new_n16614));
  nor_5  g14266(.A(new_n16614), .B(new_n16613), .Y(new_n16615));
  or_5   g14267(.A(new_n16615), .B(new_n16595), .Y(new_n16616));
  and_5  g14268(.A(new_n16616), .B(new_n16594), .Y(new_n16617_1));
  nor_5  g14269(.A(new_n16617_1), .B(new_n16593), .Y(new_n16618));
  nor_5  g14270(.A(new_n16618), .B(new_n16591), .Y(new_n16619));
  or_5   g14271(.A(new_n16619), .B(new_n16590), .Y(new_n16620));
  and_5  g14272(.A(new_n16620), .B(new_n16589_1), .Y(new_n16621));
  or_5   g14273(.A(new_n16621), .B(new_n16588), .Y(new_n16622));
  xnor_4 g14274(.A(new_n14518), .B(new_n12518), .Y(new_n16623));
  and_5  g14275(.A(new_n16623), .B(new_n16622), .Y(new_n16624));
  nor_5  g14276(.A(new_n16624), .B(new_n16586), .Y(new_n16625));
  and_5  g14277(.A(new_n16625), .B(new_n16584_1), .Y(new_n16626));
  nor_5  g14278(.A(new_n16626), .B(new_n16583_1), .Y(new_n16627));
  not_8  g14279(.A(new_n16627), .Y(new_n16628));
  nor_5  g14280(.A(new_n13508), .B(new_n5872), .Y(new_n16629));
  or_5   g14281(.A(new_n5871), .B(n6456), .Y(new_n16630_1));
  nor_5  g14282(.A(new_n5917), .B(n4085), .Y(new_n16631));
  xnor_4 g14283(.A(new_n5917), .B(new_n5875), .Y(new_n16632));
  nor_5  g14284(.A(new_n5923), .B(n26725), .Y(new_n16633));
  xnor_4 g14285(.A(new_n5923), .B(n26725), .Y(new_n16634));
  nor_5  g14286(.A(new_n5928), .B(n11980), .Y(new_n16635));
  xnor_4 g14287(.A(new_n5928), .B(new_n5880), .Y(new_n16636));
  nor_5  g14288(.A(new_n5933), .B(n3253), .Y(new_n16637));
  xnor_4 g14289(.A(new_n5933), .B(new_n5883), .Y(new_n16638));
  nor_5  g14290(.A(new_n5938), .B(n7759), .Y(new_n16639));
  xnor_4 g14291(.A(new_n5938), .B(new_n5886), .Y(new_n16640_1));
  nor_5  g14292(.A(new_n5943_1), .B(n12562), .Y(new_n16641));
  nor_5  g14293(.A(new_n5949), .B(n7949), .Y(new_n16642));
  xnor_4 g14294(.A(new_n5950), .B(n7949), .Y(new_n16643));
  nor_5  g14295(.A(new_n5960), .B(n24374), .Y(new_n16644));
  or_5   g14296(.A(new_n3798), .B(new_n5895), .Y(new_n16645));
  xnor_4 g14297(.A(new_n5961), .B(n24374), .Y(new_n16646));
  and_5  g14298(.A(new_n16646), .B(new_n16645), .Y(new_n16647));
  or_5   g14299(.A(new_n16647), .B(new_n16644), .Y(new_n16648));
  and_5  g14300(.A(new_n16648), .B(new_n16643), .Y(new_n16649));
  or_5   g14301(.A(new_n16649), .B(new_n16642), .Y(new_n16650));
  xnor_4 g14302(.A(new_n5943_1), .B(new_n5889), .Y(new_n16651));
  and_5  g14303(.A(new_n16651), .B(new_n16650), .Y(new_n16652));
  or_5   g14304(.A(new_n16652), .B(new_n16641), .Y(new_n16653));
  and_5  g14305(.A(new_n16653), .B(new_n16640_1), .Y(new_n16654));
  or_5   g14306(.A(new_n16654), .B(new_n16639), .Y(new_n16655));
  and_5  g14307(.A(new_n16655), .B(new_n16638), .Y(new_n16656_1));
  or_5   g14308(.A(new_n16656_1), .B(new_n16637), .Y(new_n16657));
  and_5  g14309(.A(new_n16657), .B(new_n16636), .Y(new_n16658));
  nor_5  g14310(.A(new_n16658), .B(new_n16635), .Y(new_n16659));
  nor_5  g14311(.A(new_n16659), .B(new_n16634), .Y(new_n16660));
  or_5   g14312(.A(new_n16660), .B(new_n16633), .Y(new_n16661));
  and_5  g14313(.A(new_n16661), .B(new_n16632), .Y(new_n16662));
  nor_5  g14314(.A(new_n16662), .B(new_n16631), .Y(new_n16663));
  and_5  g14315(.A(new_n16663), .B(new_n16630_1), .Y(new_n16664));
  or_5   g14316(.A(new_n16664), .B(new_n13550), .Y(new_n16665));
  nor_5  g14317(.A(new_n16665), .B(new_n16629), .Y(new_n16666));
  and_5  g14318(.A(new_n16666), .B(new_n16628), .Y(new_n16667));
  xor_4  g14319(.A(new_n16625), .B(new_n16584_1), .Y(new_n16668));
  nor_5  g14320(.A(new_n16668), .B(new_n16666), .Y(new_n16669));
  xnor_4 g14321(.A(new_n16668), .B(new_n16666), .Y(new_n16670));
  xor_4  g14322(.A(new_n16623), .B(new_n16622), .Y(new_n16671));
  xnor_4 g14323(.A(new_n13508), .B(n6456), .Y(new_n16672));
  xnor_4 g14324(.A(new_n16672), .B(new_n16663), .Y(new_n16673));
  and_5  g14325(.A(new_n16673), .B(new_n16671), .Y(new_n16674_1));
  xnor_4 g14326(.A(new_n16673), .B(new_n16671), .Y(new_n16675));
  xor_4  g14327(.A(new_n16661), .B(new_n16632), .Y(new_n16676));
  xor_4  g14328(.A(new_n16620), .B(new_n16589_1), .Y(new_n16677));
  and_5  g14329(.A(new_n16677), .B(new_n16676), .Y(new_n16678));
  xnor_4 g14330(.A(new_n16677), .B(new_n16676), .Y(new_n16679));
  xnor_4 g14331(.A(new_n16659), .B(new_n16634), .Y(new_n16680));
  xnor_4 g14332(.A(new_n16618), .B(new_n16591), .Y(new_n16681));
  nor_5  g14333(.A(new_n16681), .B(new_n16680), .Y(new_n16682_1));
  xnor_4 g14334(.A(new_n16681), .B(new_n16680), .Y(new_n16683));
  xor_4  g14335(.A(new_n16657), .B(new_n16636), .Y(new_n16684_1));
  xor_4  g14336(.A(new_n16616), .B(new_n16594), .Y(new_n16685));
  and_5  g14337(.A(new_n16685), .B(new_n16684_1), .Y(new_n16686));
  xnor_4 g14338(.A(new_n16685), .B(new_n16684_1), .Y(new_n16687));
  xor_4  g14339(.A(new_n16655), .B(new_n16638), .Y(new_n16688_1));
  xnor_4 g14340(.A(new_n16614), .B(new_n16613), .Y(new_n16689));
  not_8  g14341(.A(new_n16689), .Y(new_n16690));
  and_5  g14342(.A(new_n16690), .B(new_n16688_1), .Y(new_n16691));
  xnor_4 g14343(.A(new_n16690), .B(new_n16688_1), .Y(new_n16692));
  xor_4  g14344(.A(new_n16653), .B(new_n16640_1), .Y(new_n16693));
  xnor_4 g14345(.A(new_n16611), .B(new_n16597), .Y(new_n16694));
  not_8  g14346(.A(new_n16694), .Y(new_n16695));
  and_5  g14347(.A(new_n16695), .B(new_n16693), .Y(new_n16696));
  xnor_4 g14348(.A(new_n16695), .B(new_n16693), .Y(new_n16697));
  xnor_4 g14349(.A(new_n16609), .B(new_n16599), .Y(new_n16698));
  xor_4  g14350(.A(new_n16651), .B(new_n16650), .Y(new_n16699));
  and_5  g14351(.A(new_n16699), .B(new_n16698), .Y(new_n16700));
  not_8  g14352(.A(new_n16698), .Y(new_n16701));
  xnor_4 g14353(.A(new_n16699), .B(new_n16701), .Y(new_n16702));
  xor_4  g14354(.A(new_n16648), .B(new_n16643), .Y(new_n16703));
  xor_4  g14355(.A(new_n16607), .B(new_n16601), .Y(new_n16704));
  nor_5  g14356(.A(new_n16704), .B(new_n16703), .Y(new_n16705));
  xor_4  g14357(.A(new_n16704), .B(new_n16703), .Y(new_n16706));
  nor_5  g14358(.A(new_n12563), .B(new_n4266_1), .Y(new_n16707));
  xnor_4 g14359(.A(new_n16605), .B(new_n16707), .Y(new_n16708));
  not_8  g14360(.A(new_n16708), .Y(new_n16709));
  nor_5  g14361(.A(new_n16709), .B(new_n16646), .Y(new_n16710));
  xor_4  g14362(.A(new_n16646), .B(new_n16645), .Y(new_n16711));
  nor_5  g14363(.A(new_n16711), .B(new_n16708), .Y(new_n16712));
  xnor_4 g14364(.A(n20658), .B(n14575), .Y(new_n16713));
  xnor_4 g14365(.A(new_n12562_1), .B(new_n4266_1), .Y(new_n16714));
  not_8  g14366(.A(new_n16714), .Y(new_n16715));
  nor_5  g14367(.A(new_n16715), .B(new_n16713), .Y(new_n16716));
  nor_5  g14368(.A(new_n16716), .B(new_n16712), .Y(new_n16717));
  nor_5  g14369(.A(new_n16717), .B(new_n16710), .Y(new_n16718));
  and_5  g14370(.A(new_n16718), .B(new_n16706), .Y(new_n16719));
  nor_5  g14371(.A(new_n16719), .B(new_n16705), .Y(new_n16720));
  and_5  g14372(.A(new_n16720), .B(new_n16702), .Y(new_n16721));
  nor_5  g14373(.A(new_n16721), .B(new_n16700), .Y(new_n16722_1));
  nor_5  g14374(.A(new_n16722_1), .B(new_n16697), .Y(new_n16723));
  nor_5  g14375(.A(new_n16723), .B(new_n16696), .Y(new_n16724));
  nor_5  g14376(.A(new_n16724), .B(new_n16692), .Y(new_n16725));
  nor_5  g14377(.A(new_n16725), .B(new_n16691), .Y(new_n16726));
  nor_5  g14378(.A(new_n16726), .B(new_n16687), .Y(new_n16727));
  nor_5  g14379(.A(new_n16727), .B(new_n16686), .Y(new_n16728));
  nor_5  g14380(.A(new_n16728), .B(new_n16683), .Y(new_n16729));
  nor_5  g14381(.A(new_n16729), .B(new_n16682_1), .Y(new_n16730));
  nor_5  g14382(.A(new_n16730), .B(new_n16679), .Y(new_n16731));
  nor_5  g14383(.A(new_n16731), .B(new_n16678), .Y(new_n16732));
  nor_5  g14384(.A(new_n16732), .B(new_n16675), .Y(new_n16733_1));
  nor_5  g14385(.A(new_n16733_1), .B(new_n16674_1), .Y(new_n16734));
  nor_5  g14386(.A(new_n16734), .B(new_n16670), .Y(new_n16735));
  nor_5  g14387(.A(new_n16735), .B(new_n16669), .Y(new_n16736));
  nor_5  g14388(.A(new_n16736), .B(new_n16667), .Y(new_n16737));
  nor_5  g14389(.A(new_n16666), .B(new_n16628), .Y(new_n16738));
  nor_5  g14390(.A(new_n16738), .B(new_n16735), .Y(new_n16739));
  nor_5  g14391(.A(new_n16739), .B(new_n16737), .Y(n4123));
  xnor_4 g14392(.A(new_n13068), .B(new_n7870), .Y(new_n16741));
  nor_5  g14393(.A(new_n13071), .B(new_n7877), .Y(new_n16742));
  xnor_4 g14394(.A(new_n13072), .B(new_n7876_1), .Y(new_n16743_1));
  not_8  g14395(.A(new_n13076), .Y(new_n16744));
  nor_5  g14396(.A(new_n16744), .B(new_n7899), .Y(new_n16745));
  xnor_4 g14397(.A(new_n16744), .B(new_n7898), .Y(new_n16746));
  and_5  g14398(.A(new_n13086), .B(new_n7885), .Y(new_n16747));
  nor_5  g14399(.A(new_n9708), .B(new_n7887), .Y(new_n16748));
  xnor_4 g14400(.A(new_n13085), .B(new_n7885), .Y(new_n16749));
  and_5  g14401(.A(new_n16749), .B(new_n16748), .Y(new_n16750));
  nor_5  g14402(.A(new_n16750), .B(new_n16747), .Y(new_n16751));
  and_5  g14403(.A(new_n16751), .B(new_n16746), .Y(new_n16752));
  nor_5  g14404(.A(new_n16752), .B(new_n16745), .Y(new_n16753));
  nor_5  g14405(.A(new_n16753), .B(new_n16743_1), .Y(new_n16754));
  nor_5  g14406(.A(new_n16754), .B(new_n16742), .Y(new_n16755));
  xnor_4 g14407(.A(new_n16755), .B(new_n16741), .Y(n4134));
  xnor_4 g14408(.A(new_n9055), .B(new_n9005), .Y(n4146));
  xnor_4 g14409(.A(new_n15062), .B(new_n13958), .Y(new_n16758));
  nor_5  g14410(.A(new_n15068), .B(new_n13963), .Y(new_n16759));
  xnor_4 g14411(.A(new_n15066), .B(new_n13963), .Y(new_n16760));
  and_5  g14412(.A(new_n13966), .B(new_n13150), .Y(new_n16761));
  nor_5  g14413(.A(new_n13969), .B(new_n13143), .Y(new_n16762));
  xnor_4 g14414(.A(new_n13966), .B(new_n13149), .Y(new_n16763));
  and_5  g14415(.A(new_n16763), .B(new_n16762), .Y(new_n16764));
  nor_5  g14416(.A(new_n16764), .B(new_n16761), .Y(new_n16765));
  and_5  g14417(.A(new_n16765), .B(new_n16760), .Y(new_n16766));
  nor_5  g14418(.A(new_n16766), .B(new_n16759), .Y(new_n16767));
  xnor_4 g14419(.A(new_n16767), .B(new_n16758), .Y(n4150));
  xnor_4 g14420(.A(new_n12342), .B(new_n12341_1), .Y(n4151));
  xnor_4 g14421(.A(new_n12663), .B(new_n12604), .Y(n4152));
  xnor_4 g14422(.A(new_n6143), .B(new_n6104_1), .Y(n4153));
  nor_5  g14423(.A(new_n11842_1), .B(n10250), .Y(new_n16772));
  and_5  g14424(.A(new_n8680), .B(new_n8645), .Y(new_n16773));
  nor_5  g14425(.A(new_n16773), .B(new_n16772), .Y(new_n16774));
  xnor_4 g14426(.A(new_n16774), .B(new_n12059), .Y(new_n16775));
  not_8  g14427(.A(new_n16774), .Y(new_n16776));
  nor_5  g14428(.A(new_n16776), .B(new_n12063), .Y(new_n16777));
  nor_5  g14429(.A(new_n16774), .B(new_n12064), .Y(new_n16778));
  and_5  g14430(.A(new_n12067), .B(new_n8681), .Y(new_n16779));
  and_5  g14431(.A(new_n8909_1), .B(new_n8854), .Y(new_n16780));
  nor_5  g14432(.A(new_n16780), .B(new_n16779), .Y(new_n16781));
  nor_5  g14433(.A(new_n16781), .B(new_n16778), .Y(new_n16782));
  nor_5  g14434(.A(new_n16782), .B(new_n16777), .Y(new_n16783));
  xnor_4 g14435(.A(new_n16783), .B(new_n16775), .Y(n4165));
  xnor_4 g14436(.A(new_n11411), .B(new_n11382), .Y(n4172));
  xnor_4 g14437(.A(new_n11249), .B(new_n4745_1), .Y(n4173));
  xnor_4 g14438(.A(new_n6579), .B(new_n6559), .Y(n4176));
  xnor_4 g14439(.A(new_n9040), .B(new_n9039), .Y(n4186));
  xnor_4 g14440(.A(new_n16357), .B(new_n16335), .Y(n4204));
  nor_5  g14441(.A(new_n11296), .B(new_n5500), .Y(new_n16790));
  xnor_4 g14442(.A(new_n11296), .B(new_n5500), .Y(new_n16791));
  nor_5  g14443(.A(new_n6789), .B(new_n5503), .Y(new_n16792));
  nor_5  g14444(.A(new_n6832), .B(new_n6790_1), .Y(new_n16793));
  nor_5  g14445(.A(new_n16793), .B(new_n16792), .Y(new_n16794));
  nor_5  g14446(.A(new_n16794), .B(new_n16791), .Y(new_n16795));
  nor_5  g14447(.A(new_n16795), .B(new_n16790), .Y(new_n16796));
  nor_5  g14448(.A(new_n16796), .B(new_n11792), .Y(new_n16797));
  not_8  g14449(.A(new_n15725), .Y(new_n16798_1));
  nor_5  g14450(.A(new_n16798_1), .B(n3366), .Y(new_n16799));
  not_8  g14451(.A(new_n16799), .Y(new_n16800));
  nor_5  g14452(.A(new_n16800), .B(n19652), .Y(new_n16801));
  xnor_4 g14453(.A(new_n16801), .B(n3984), .Y(new_n16802));
  and_5  g14454(.A(new_n16802), .B(new_n11326_1), .Y(new_n16803));
  xnor_4 g14455(.A(new_n16802), .B(n17037), .Y(new_n16804));
  xnor_4 g14456(.A(new_n16800), .B(n19652), .Y(new_n16805));
  and_5  g14457(.A(new_n16805), .B(n5386), .Y(new_n16806));
  not_8  g14458(.A(new_n15726), .Y(new_n16807));
  nor_5  g14459(.A(new_n16807), .B(n26191), .Y(new_n16808));
  and_5  g14460(.A(new_n15757), .B(new_n15727), .Y(new_n16809));
  nor_5  g14461(.A(new_n16809), .B(new_n16808), .Y(new_n16810));
  xor_4  g14462(.A(new_n16805), .B(n5386), .Y(new_n16811));
  and_5  g14463(.A(new_n16811), .B(new_n16810), .Y(new_n16812_1));
  nor_5  g14464(.A(new_n16812_1), .B(new_n16806), .Y(new_n16813));
  and_5  g14465(.A(new_n16813), .B(new_n16804), .Y(new_n16814));
  nor_5  g14466(.A(new_n16814), .B(new_n16803), .Y(new_n16815));
  not_8  g14467(.A(new_n16801), .Y(new_n16816));
  nor_5  g14468(.A(new_n16816), .B(n3984), .Y(new_n16817));
  xnor_4 g14469(.A(new_n16817), .B(n4514), .Y(new_n16818_1));
  xnor_4 g14470(.A(new_n16818_1), .B(n7569), .Y(new_n16819));
  xnor_4 g14471(.A(new_n16819), .B(new_n16815), .Y(new_n16820));
  nor_5  g14472(.A(new_n16820), .B(new_n14303), .Y(new_n16821));
  xnor_4 g14473(.A(new_n16820), .B(new_n14303), .Y(new_n16822));
  xor_4  g14474(.A(new_n16813), .B(new_n16804), .Y(new_n16823));
  nor_5  g14475(.A(new_n16823), .B(new_n14165), .Y(new_n16824_1));
  xnor_4 g14476(.A(new_n16823), .B(n25751), .Y(new_n16825));
  xor_4  g14477(.A(new_n16811), .B(new_n16810), .Y(new_n16826));
  nor_5  g14478(.A(new_n16826), .B(n26053), .Y(new_n16827));
  xnor_4 g14479(.A(new_n16826), .B(new_n14168), .Y(new_n16828));
  and_5  g14480(.A(new_n15758), .B(new_n14171), .Y(new_n16829));
  and_5  g14481(.A(new_n15787), .B(new_n15759), .Y(new_n16830));
  or_5   g14482(.A(new_n16830), .B(new_n16829), .Y(new_n16831));
  and_5  g14483(.A(new_n16831), .B(new_n16828), .Y(new_n16832));
  nor_5  g14484(.A(new_n16832), .B(new_n16827), .Y(new_n16833));
  and_5  g14485(.A(new_n16833), .B(new_n16825), .Y(new_n16834_1));
  nor_5  g14486(.A(new_n16834_1), .B(new_n16824_1), .Y(new_n16835));
  nor_5  g14487(.A(new_n16835), .B(new_n16822), .Y(new_n16836));
  nor_5  g14488(.A(new_n16836), .B(new_n16821), .Y(new_n16837_1));
  and_5  g14489(.A(new_n16817), .B(new_n11273_1), .Y(new_n16838));
  nor_5  g14490(.A(new_n16818_1), .B(new_n11325_1), .Y(new_n16839));
  nor_5  g14491(.A(new_n16839), .B(new_n16815), .Y(new_n16840));
  and_5  g14492(.A(new_n16840), .B(new_n16838), .Y(new_n16841_1));
  and_5  g14493(.A(new_n16841_1), .B(new_n16837_1), .Y(new_n16842));
  and_5  g14494(.A(new_n16818_1), .B(new_n11325_1), .Y(new_n16843));
  xor_4  g14495(.A(new_n16840), .B(new_n16838), .Y(new_n16844));
  nor_5  g14496(.A(new_n16844), .B(new_n16843), .Y(new_n16845));
  not_8  g14497(.A(new_n16845), .Y(new_n16846));
  or_5   g14498(.A(new_n16846), .B(new_n16837_1), .Y(new_n16847));
  nor_5  g14499(.A(new_n16847), .B(new_n16841_1), .Y(new_n16848));
  nor_5  g14500(.A(new_n16848), .B(new_n16842), .Y(new_n16849));
  or_5   g14501(.A(new_n16849), .B(new_n16797), .Y(new_n16850));
  xnor_4 g14502(.A(new_n16845), .B(new_n16837_1), .Y(new_n16851));
  xnor_4 g14503(.A(new_n16796), .B(new_n11323), .Y(new_n16852));
  not_8  g14504(.A(new_n16852), .Y(new_n16853));
  and_5  g14505(.A(new_n16853), .B(new_n16851), .Y(new_n16854));
  xnor_4 g14506(.A(new_n16853), .B(new_n16851), .Y(new_n16855));
  xnor_4 g14507(.A(new_n16835), .B(new_n16822), .Y(new_n16856));
  xnor_4 g14508(.A(new_n16794), .B(new_n16791), .Y(new_n16857));
  not_8  g14509(.A(new_n16857), .Y(new_n16858));
  nor_5  g14510(.A(new_n16858), .B(new_n16856), .Y(new_n16859));
  xnor_4 g14511(.A(new_n16858), .B(new_n16856), .Y(new_n16860));
  not_8  g14512(.A(new_n6833), .Y(new_n16861));
  xnor_4 g14513(.A(new_n16833), .B(new_n16825), .Y(new_n16862));
  nor_5  g14514(.A(new_n16862), .B(new_n16861), .Y(new_n16863));
  xnor_4 g14515(.A(new_n16862), .B(new_n16861), .Y(new_n16864));
  xor_4  g14516(.A(new_n16831), .B(new_n16828), .Y(new_n16865));
  nor_5  g14517(.A(new_n16865), .B(new_n6913), .Y(new_n16866));
  nor_5  g14518(.A(new_n15788), .B(new_n6918), .Y(new_n16867));
  nor_5  g14519(.A(new_n15818), .B(new_n15789), .Y(new_n16868));
  nor_5  g14520(.A(new_n16868), .B(new_n16867), .Y(new_n16869));
  xnor_4 g14521(.A(new_n16865), .B(new_n6913), .Y(new_n16870));
  nor_5  g14522(.A(new_n16870), .B(new_n16869), .Y(new_n16871));
  nor_5  g14523(.A(new_n16871), .B(new_n16866), .Y(new_n16872));
  nor_5  g14524(.A(new_n16872), .B(new_n16864), .Y(new_n16873));
  nor_5  g14525(.A(new_n16873), .B(new_n16863), .Y(new_n16874));
  nor_5  g14526(.A(new_n16874), .B(new_n16860), .Y(new_n16875));
  nor_5  g14527(.A(new_n16875), .B(new_n16859), .Y(new_n16876));
  nor_5  g14528(.A(new_n16876), .B(new_n16855), .Y(new_n16877));
  nor_5  g14529(.A(new_n16877), .B(new_n16854), .Y(new_n16878));
  and_5  g14530(.A(new_n16878), .B(new_n16850), .Y(new_n16879));
  and_5  g14531(.A(new_n16849), .B(new_n16797), .Y(new_n16880));
  or_5   g14532(.A(new_n16880), .B(new_n16842), .Y(new_n16881));
  nor_5  g14533(.A(new_n16881), .B(new_n16879), .Y(n4205));
  not_8  g14534(.A(new_n12997), .Y(new_n16883));
  nor_5  g14535(.A(new_n16883), .B(n22198), .Y(new_n16884));
  not_8  g14536(.A(new_n16884), .Y(new_n16885_1));
  nor_5  g14537(.A(new_n16885_1), .B(n24327), .Y(new_n16886));
  xnor_4 g14538(.A(new_n16886), .B(n2659), .Y(new_n16887));
  xnor_4 g14539(.A(new_n16887), .B(n18444), .Y(new_n16888));
  xnor_4 g14540(.A(new_n16884), .B(n24327), .Y(new_n16889));
  nor_5  g14541(.A(new_n16889), .B(n24638), .Y(new_n16890));
  xnor_4 g14542(.A(new_n16889), .B(n24638), .Y(new_n16891));
  nor_5  g14543(.A(new_n12998), .B(n21674), .Y(new_n16892));
  nor_5  g14544(.A(new_n13020), .B(new_n12999), .Y(new_n16893));
  nor_5  g14545(.A(new_n16893), .B(new_n16892), .Y(new_n16894));
  nor_5  g14546(.A(new_n16894), .B(new_n16891), .Y(new_n16895));
  nor_5  g14547(.A(new_n16895), .B(new_n16890), .Y(new_n16896));
  xor_4  g14548(.A(new_n16896), .B(new_n16888), .Y(new_n16897));
  xnor_4 g14549(.A(new_n16897), .B(new_n7715), .Y(new_n16898));
  xnor_4 g14550(.A(new_n16894), .B(new_n16891), .Y(new_n16899));
  and_5  g14551(.A(new_n16899), .B(new_n7718), .Y(new_n16900));
  xor_4  g14552(.A(new_n16899), .B(new_n7718), .Y(new_n16901));
  nor_5  g14553(.A(new_n13021), .B(new_n7722), .Y(new_n16902));
  nor_5  g14554(.A(new_n13043_1), .B(new_n13022), .Y(new_n16903));
  nor_5  g14555(.A(new_n16903), .B(new_n16902), .Y(new_n16904));
  and_5  g14556(.A(new_n16904), .B(new_n16901), .Y(new_n16905_1));
  nor_5  g14557(.A(new_n16905_1), .B(new_n16900), .Y(new_n16906));
  xnor_4 g14558(.A(new_n16906), .B(new_n16898), .Y(new_n16907));
  xnor_4 g14559(.A(n21997), .B(n5400), .Y(new_n16908));
  nor_5  g14560(.A(n25119), .B(new_n8284), .Y(new_n16909));
  xnor_4 g14561(.A(n25119), .B(n23923), .Y(new_n16910));
  nor_5  g14562(.A(n1163), .B(new_n8353), .Y(new_n16911_1));
  and_5  g14563(.A(new_n13064), .B(new_n13045), .Y(new_n16912));
  or_5   g14564(.A(new_n16912), .B(new_n16911_1), .Y(new_n16913));
  and_5  g14565(.A(new_n16913), .B(new_n16910), .Y(new_n16914));
  or_5   g14566(.A(new_n16914), .B(new_n16909), .Y(new_n16915));
  xor_4  g14567(.A(new_n16915), .B(new_n16908), .Y(new_n16916));
  xnor_4 g14568(.A(new_n16916), .B(new_n16907), .Y(new_n16917));
  xor_4  g14569(.A(new_n16913), .B(new_n16910), .Y(new_n16918));
  xnor_4 g14570(.A(new_n16904), .B(new_n16901), .Y(new_n16919));
  not_8  g14571(.A(new_n16919), .Y(new_n16920));
  and_5  g14572(.A(new_n16920), .B(new_n16918), .Y(new_n16921));
  xnor_4 g14573(.A(new_n16919), .B(new_n16918), .Y(new_n16922));
  nor_5  g14574(.A(new_n13065), .B(new_n13044_1), .Y(new_n16923));
  nor_5  g14575(.A(new_n13095), .B(new_n13066), .Y(new_n16924));
  nor_5  g14576(.A(new_n16924), .B(new_n16923), .Y(new_n16925));
  and_5  g14577(.A(new_n16925), .B(new_n16922), .Y(new_n16926));
  or_5   g14578(.A(new_n16926), .B(new_n16921), .Y(new_n16927));
  xor_4  g14579(.A(new_n16927), .B(new_n16917), .Y(n4215));
  and_5  g14580(.A(new_n14005), .B(new_n5985), .Y(new_n16929));
  xnor_4 g14581(.A(new_n16929), .B(n3582), .Y(new_n16930));
  xnor_4 g14582(.A(new_n16930), .B(new_n4907), .Y(new_n16931));
  and_5  g14583(.A(new_n14006), .B(n2858), .Y(new_n16932));
  or_5   g14584(.A(new_n14006), .B(n2858), .Y(new_n16933));
  and_5  g14585(.A(new_n14031), .B(new_n16933), .Y(new_n16934));
  nor_5  g14586(.A(new_n16934), .B(new_n16932), .Y(new_n16935));
  xnor_4 g14587(.A(new_n16935), .B(new_n16931), .Y(new_n16936));
  not_8  g14588(.A(new_n9610), .Y(new_n16937));
  nor_5  g14589(.A(new_n16937), .B(n27089), .Y(new_n16938));
  xnor_4 g14590(.A(new_n16938), .B(n21839), .Y(new_n16939));
  not_8  g14591(.A(new_n16939), .Y(new_n16940));
  xnor_4 g14592(.A(new_n16940), .B(n22626), .Y(new_n16941));
  nor_5  g14593(.A(new_n9611), .B(n14440), .Y(new_n16942));
  xnor_4 g14594(.A(new_n9611), .B(new_n7482), .Y(new_n16943));
  not_8  g14595(.A(new_n16943), .Y(new_n16944));
  nor_5  g14596(.A(new_n9613), .B(n1654), .Y(new_n16945));
  nor_5  g14597(.A(new_n15491), .B(new_n15488), .Y(new_n16946));
  nor_5  g14598(.A(new_n16946), .B(new_n16945), .Y(new_n16947));
  nor_5  g14599(.A(new_n16947), .B(new_n16944), .Y(new_n16948));
  or_5   g14600(.A(new_n16948), .B(new_n16942), .Y(new_n16949));
  xnor_4 g14601(.A(new_n16949), .B(new_n16941), .Y(new_n16950));
  xnor_4 g14602(.A(new_n16950), .B(new_n16936), .Y(new_n16951_1));
  xnor_4 g14603(.A(new_n16947), .B(new_n16943), .Y(new_n16952));
  nor_5  g14604(.A(new_n16952), .B(new_n14032), .Y(new_n16953));
  not_8  g14605(.A(new_n14035), .Y(new_n16954_1));
  nor_5  g14606(.A(new_n15492), .B(new_n16954_1), .Y(new_n16955));
  xnor_4 g14607(.A(new_n15492), .B(new_n16954_1), .Y(new_n16956));
  nor_5  g14608(.A(new_n14038), .B(new_n10541), .Y(new_n16957));
  xnor_4 g14609(.A(new_n14038), .B(new_n10541), .Y(new_n16958));
  nor_5  g14610(.A(new_n14041), .B(new_n10543), .Y(new_n16959));
  xnor_4 g14611(.A(new_n14043), .B(new_n10546), .Y(new_n16960));
  nor_5  g14612(.A(new_n14048), .B(new_n10554), .Y(new_n16961));
  xnor_4 g14613(.A(new_n14048), .B(new_n10554), .Y(new_n16962));
  and_5  g14614(.A(new_n9423_1), .B(new_n9409), .Y(new_n16963));
  nor_5  g14615(.A(new_n9440), .B(new_n9424), .Y(new_n16964));
  nor_5  g14616(.A(new_n16964), .B(new_n16963), .Y(new_n16965));
  nor_5  g14617(.A(new_n16965), .B(new_n16962), .Y(new_n16966));
  or_5   g14618(.A(new_n16966), .B(new_n16961), .Y(new_n16967));
  nor_5  g14619(.A(new_n16967), .B(new_n16960), .Y(new_n16968_1));
  nor_5  g14620(.A(new_n16968_1), .B(new_n16959), .Y(new_n16969));
  nor_5  g14621(.A(new_n16969), .B(new_n16958), .Y(new_n16970));
  nor_5  g14622(.A(new_n16970), .B(new_n16957), .Y(new_n16971_1));
  nor_5  g14623(.A(new_n16971_1), .B(new_n16956), .Y(new_n16972));
  nor_5  g14624(.A(new_n16972), .B(new_n16955), .Y(new_n16973));
  not_8  g14625(.A(new_n16952), .Y(new_n16974));
  xnor_4 g14626(.A(new_n16974), .B(new_n14032), .Y(new_n16975));
  and_5  g14627(.A(new_n16975), .B(new_n16973), .Y(new_n16976));
  nor_5  g14628(.A(new_n16976), .B(new_n16953), .Y(new_n16977));
  xnor_4 g14629(.A(new_n16977), .B(new_n16951_1), .Y(new_n16978));
  not_8  g14630(.A(new_n16978), .Y(new_n16979));
  not_8  g14631(.A(new_n14749), .Y(new_n16980));
  nor_5  g14632(.A(new_n16980), .B(n10611), .Y(new_n16981));
  not_8  g14633(.A(new_n16981), .Y(new_n16982));
  nor_5  g14634(.A(new_n16982), .B(n3164), .Y(new_n16983));
  not_8  g14635(.A(new_n16983), .Y(new_n16984));
  nor_5  g14636(.A(new_n16984), .B(n11356), .Y(new_n16985));
  not_8  g14637(.A(new_n16985), .Y(new_n16986));
  nor_5  g14638(.A(new_n16986), .B(n14345), .Y(new_n16987));
  not_8  g14639(.A(new_n16987), .Y(new_n16988_1));
  nor_5  g14640(.A(new_n16988_1), .B(n6381), .Y(new_n16989_1));
  not_8  g14641(.A(new_n16989_1), .Y(new_n16990));
  nor_5  g14642(.A(new_n16990), .B(n10577), .Y(new_n16991));
  xnor_4 g14643(.A(new_n16991), .B(n23166), .Y(new_n16992));
  xnor_4 g14644(.A(new_n16992), .B(new_n7772), .Y(new_n16993));
  xnor_4 g14645(.A(new_n16989_1), .B(n10577), .Y(new_n16994_1));
  nor_5  g14646(.A(new_n16994_1), .B(n26408), .Y(new_n16995));
  xnor_4 g14647(.A(new_n16994_1), .B(n26408), .Y(new_n16996));
  xnor_4 g14648(.A(new_n16987), .B(n6381), .Y(new_n16997));
  nor_5  g14649(.A(new_n16997), .B(n18227), .Y(new_n16998));
  xnor_4 g14650(.A(new_n16997), .B(new_n4804_1), .Y(new_n16999));
  xnor_4 g14651(.A(new_n16985), .B(n14345), .Y(new_n17000));
  nor_5  g14652(.A(new_n17000), .B(n7377), .Y(new_n17001));
  xnor_4 g14653(.A(new_n17000), .B(new_n4807), .Y(new_n17002));
  xnor_4 g14654(.A(new_n16983), .B(n11356), .Y(new_n17003));
  nor_5  g14655(.A(new_n17003), .B(n11630), .Y(new_n17004));
  xnor_4 g14656(.A(new_n16981), .B(n3164), .Y(new_n17005));
  nor_5  g14657(.A(new_n17005), .B(n13453), .Y(new_n17006_1));
  xnor_4 g14658(.A(new_n17005), .B(new_n12754), .Y(new_n17007));
  and_5  g14659(.A(new_n14750), .B(n7421), .Y(new_n17008));
  and_5  g14660(.A(new_n14763_1), .B(new_n14751), .Y(new_n17009));
  nor_5  g14661(.A(new_n17009), .B(new_n17008), .Y(new_n17010));
  and_5  g14662(.A(new_n17010), .B(new_n17007), .Y(new_n17011));
  or_5   g14663(.A(new_n17011), .B(new_n17006_1), .Y(new_n17012));
  not_8  g14664(.A(n11630), .Y(new_n17013));
  xnor_4 g14665(.A(new_n17003), .B(new_n17013), .Y(new_n17014));
  and_5  g14666(.A(new_n17014), .B(new_n17012), .Y(new_n17015));
  or_5   g14667(.A(new_n17015), .B(new_n17004), .Y(new_n17016));
  and_5  g14668(.A(new_n17016), .B(new_n17002), .Y(new_n17017));
  or_5   g14669(.A(new_n17017), .B(new_n17001), .Y(new_n17018));
  and_5  g14670(.A(new_n17018), .B(new_n16999), .Y(new_n17019));
  nor_5  g14671(.A(new_n17019), .B(new_n16998), .Y(new_n17020));
  nor_5  g14672(.A(new_n17020), .B(new_n16996), .Y(new_n17021));
  nor_5  g14673(.A(new_n17021), .B(new_n16995), .Y(new_n17022));
  xnor_4 g14674(.A(new_n17022), .B(new_n16993), .Y(new_n17023));
  not_8  g14675(.A(new_n17023), .Y(new_n17024));
  xnor_4 g14676(.A(new_n17024), .B(new_n16979), .Y(new_n17025));
  xnor_4 g14677(.A(new_n17020), .B(new_n16996), .Y(new_n17026));
  xor_4  g14678(.A(new_n16975), .B(new_n16973), .Y(new_n17027));
  nor_5  g14679(.A(new_n17027), .B(new_n17026), .Y(new_n17028));
  xnor_4 g14680(.A(new_n17027), .B(new_n17026), .Y(new_n17029));
  nor_5  g14681(.A(new_n17017), .B(new_n17001), .Y(new_n17030));
  xnor_4 g14682(.A(new_n17030), .B(new_n16999), .Y(new_n17031));
  not_8  g14683(.A(new_n17031), .Y(new_n17032));
  xor_4  g14684(.A(new_n16971_1), .B(new_n16956), .Y(new_n17033));
  not_8  g14685(.A(new_n17033), .Y(new_n17034));
  nor_5  g14686(.A(new_n17034), .B(new_n17032), .Y(new_n17035_1));
  xnor_4 g14687(.A(new_n17034), .B(new_n17032), .Y(new_n17036));
  nor_5  g14688(.A(new_n17015), .B(new_n17004), .Y(new_n17037_1));
  xnor_4 g14689(.A(new_n17037_1), .B(new_n17002), .Y(new_n17038));
  not_8  g14690(.A(new_n17038), .Y(new_n17039));
  xor_4  g14691(.A(new_n16969), .B(new_n16958), .Y(new_n17040));
  not_8  g14692(.A(new_n17040), .Y(new_n17041));
  nor_5  g14693(.A(new_n17041), .B(new_n17039), .Y(new_n17042));
  xnor_4 g14694(.A(new_n17041), .B(new_n17039), .Y(new_n17043));
  nor_5  g14695(.A(new_n16966), .B(new_n16961), .Y(new_n17044));
  xnor_4 g14696(.A(new_n17044), .B(new_n16960), .Y(new_n17045));
  not_8  g14697(.A(new_n17045), .Y(new_n17046));
  xor_4  g14698(.A(new_n17014), .B(new_n17012), .Y(new_n17047));
  not_8  g14699(.A(new_n17047), .Y(new_n17048));
  nor_5  g14700(.A(new_n17048), .B(new_n17046), .Y(new_n17049));
  xnor_4 g14701(.A(new_n17048), .B(new_n17046), .Y(new_n17050));
  xnor_4 g14702(.A(new_n17010), .B(new_n17007), .Y(new_n17051));
  xor_4  g14703(.A(new_n16965), .B(new_n16962), .Y(new_n17052));
  nor_5  g14704(.A(new_n17052), .B(new_n17051), .Y(new_n17053));
  not_8  g14705(.A(new_n17051), .Y(new_n17054));
  not_8  g14706(.A(new_n17052), .Y(new_n17055));
  xnor_4 g14707(.A(new_n17055), .B(new_n17054), .Y(new_n17056));
  nor_5  g14708(.A(new_n14764), .B(new_n9441), .Y(new_n17057));
  xnor_4 g14709(.A(new_n14764), .B(new_n9441), .Y(new_n17058));
  not_8  g14710(.A(new_n17058), .Y(new_n17059));
  nor_5  g14711(.A(new_n14766), .B(new_n9455), .Y(new_n17060));
  xnor_4 g14712(.A(new_n14766), .B(new_n9455), .Y(new_n17061));
  nor_5  g14713(.A(new_n14770), .B(new_n9467), .Y(new_n17062));
  nor_5  g14714(.A(new_n14772_1), .B(new_n9462), .Y(new_n17063));
  xnor_4 g14715(.A(new_n14770), .B(new_n9468), .Y(new_n17064));
  and_5  g14716(.A(new_n17064), .B(new_n17063), .Y(new_n17065));
  nor_5  g14717(.A(new_n17065), .B(new_n17062), .Y(new_n17066));
  nor_5  g14718(.A(new_n17066), .B(new_n17061), .Y(new_n17067));
  nor_5  g14719(.A(new_n17067), .B(new_n17060), .Y(new_n17068_1));
  and_5  g14720(.A(new_n17068_1), .B(new_n17059), .Y(new_n17069_1));
  nor_5  g14721(.A(new_n17069_1), .B(new_n17057), .Y(new_n17070_1));
  nor_5  g14722(.A(new_n17070_1), .B(new_n17056), .Y(new_n17071));
  nor_5  g14723(.A(new_n17071), .B(new_n17053), .Y(new_n17072));
  nor_5  g14724(.A(new_n17072), .B(new_n17050), .Y(new_n17073));
  nor_5  g14725(.A(new_n17073), .B(new_n17049), .Y(new_n17074));
  nor_5  g14726(.A(new_n17074), .B(new_n17043), .Y(new_n17075_1));
  nor_5  g14727(.A(new_n17075_1), .B(new_n17042), .Y(new_n17076));
  nor_5  g14728(.A(new_n17076), .B(new_n17036), .Y(new_n17077_1));
  nor_5  g14729(.A(new_n17077_1), .B(new_n17035_1), .Y(new_n17078));
  nor_5  g14730(.A(new_n17078), .B(new_n17029), .Y(new_n17079));
  or_5   g14731(.A(new_n17079), .B(new_n17028), .Y(new_n17080));
  xor_4  g14732(.A(new_n17080), .B(new_n17025), .Y(n4221));
  xnor_4 g14733(.A(new_n10450), .B(new_n4804_1), .Y(new_n17082));
  nor_5  g14734(.A(new_n10454), .B(new_n4807), .Y(new_n17083));
  xnor_4 g14735(.A(new_n10456), .B(new_n4807), .Y(new_n17084_1));
  nor_5  g14736(.A(new_n10471), .B(new_n17013), .Y(new_n17085));
  nor_5  g14737(.A(new_n10462), .B(new_n12754), .Y(new_n17086));
  or_5   g14738(.A(new_n12757), .B(new_n12756_1), .Y(new_n17087));
  and_5  g14739(.A(new_n17087), .B(new_n12755), .Y(new_n17088));
  or_5   g14740(.A(new_n17088), .B(new_n17086), .Y(new_n17089));
  xnor_4 g14741(.A(new_n10471), .B(n11630), .Y(new_n17090_1));
  and_5  g14742(.A(new_n17090_1), .B(new_n17089), .Y(new_n17091));
  or_5   g14743(.A(new_n17091), .B(new_n17085), .Y(new_n17092));
  and_5  g14744(.A(new_n17092), .B(new_n17084_1), .Y(new_n17093));
  nor_5  g14745(.A(new_n17093), .B(new_n17083), .Y(new_n17094));
  xnor_4 g14746(.A(new_n17094), .B(new_n17082), .Y(new_n17095_1));
  not_8  g14747(.A(new_n17095_1), .Y(new_n17096));
  xnor_4 g14748(.A(new_n17096), .B(new_n15885_1), .Y(new_n17097));
  nor_5  g14749(.A(new_n17091), .B(new_n17085), .Y(new_n17098));
  xnor_4 g14750(.A(new_n17098), .B(new_n17084_1), .Y(new_n17099));
  not_8  g14751(.A(new_n17099), .Y(new_n17100));
  nor_5  g14752(.A(new_n17100), .B(new_n8499), .Y(new_n17101));
  xnor_4 g14753(.A(new_n17099), .B(new_n8500), .Y(new_n17102));
  nor_5  g14754(.A(new_n17088), .B(new_n17086), .Y(new_n17103));
  xnor_4 g14755(.A(new_n17090_1), .B(new_n17103), .Y(new_n17104_1));
  and_5  g14756(.A(new_n17104_1), .B(new_n8531), .Y(new_n17105));
  xnor_4 g14757(.A(new_n17104_1), .B(new_n8531), .Y(new_n17106_1));
  not_8  g14758(.A(new_n12759), .Y(new_n17107));
  nor_5  g14759(.A(new_n17107), .B(new_n8537), .Y(new_n17108));
  xnor_4 g14760(.A(new_n12759), .B(new_n15895), .Y(new_n17109));
  nor_5  g14761(.A(new_n8542), .B(new_n6623), .Y(new_n17110));
  xnor_4 g14762(.A(new_n8542), .B(new_n6623), .Y(new_n17111));
  nor_5  g14763(.A(new_n8548), .B(new_n6654), .Y(new_n17112));
  xnor_4 g14764(.A(new_n8548), .B(new_n6654), .Y(new_n17113));
  nor_5  g14765(.A(new_n8553), .B(new_n6660), .Y(new_n17114));
  nor_5  g14766(.A(new_n8556), .B(new_n6665), .Y(new_n17115));
  xnor_4 g14767(.A(new_n8553), .B(new_n6668), .Y(new_n17116));
  and_5  g14768(.A(new_n17116), .B(new_n17115), .Y(new_n17117));
  nor_5  g14769(.A(new_n17117), .B(new_n17114), .Y(new_n17118));
  nor_5  g14770(.A(new_n17118), .B(new_n17113), .Y(new_n17119_1));
  nor_5  g14771(.A(new_n17119_1), .B(new_n17112), .Y(new_n17120));
  nor_5  g14772(.A(new_n17120), .B(new_n17111), .Y(new_n17121));
  nor_5  g14773(.A(new_n17121), .B(new_n17110), .Y(new_n17122));
  nor_5  g14774(.A(new_n17122), .B(new_n17109), .Y(new_n17123));
  nor_5  g14775(.A(new_n17123), .B(new_n17108), .Y(new_n17124));
  nor_5  g14776(.A(new_n17124), .B(new_n17106_1), .Y(new_n17125));
  nor_5  g14777(.A(new_n17125), .B(new_n17105), .Y(new_n17126));
  nor_5  g14778(.A(new_n17126), .B(new_n17102), .Y(new_n17127));
  nor_5  g14779(.A(new_n17127), .B(new_n17101), .Y(new_n17128));
  xnor_4 g14780(.A(new_n17128), .B(new_n17097), .Y(n4224));
  xor_4  g14781(.A(new_n10595_1), .B(new_n10594), .Y(n4231));
  xnor_4 g14782(.A(new_n13879), .B(n9934), .Y(new_n17131));
  nor_5  g14783(.A(new_n13881), .B(n18496), .Y(new_n17132));
  or_5   g14784(.A(new_n16461), .B(new_n16455), .Y(new_n17133));
  and_5  g14785(.A(new_n17133), .B(new_n16454), .Y(new_n17134));
  nor_5  g14786(.A(new_n17134), .B(new_n17132), .Y(new_n17135));
  xnor_4 g14787(.A(new_n17135), .B(new_n17131), .Y(new_n17136));
  not_8  g14788(.A(new_n17136), .Y(new_n17137));
  xnor_4 g14789(.A(new_n17137), .B(new_n4798), .Y(new_n17138_1));
  nor_5  g14790(.A(new_n16463), .B(new_n4801), .Y(new_n17139));
  and_5  g14791(.A(new_n16475), .B(new_n16465), .Y(new_n17140));
  or_5   g14792(.A(new_n17140), .B(new_n17139), .Y(new_n17141));
  xor_4  g14793(.A(new_n17141), .B(new_n17138_1), .Y(new_n17142));
  xnor_4 g14794(.A(new_n17142), .B(new_n11741_1), .Y(new_n17143));
  nor_5  g14795(.A(new_n16476_1), .B(new_n11745), .Y(new_n17144));
  nor_5  g14796(.A(new_n16485), .B(new_n16477), .Y(new_n17145));
  nor_5  g14797(.A(new_n17145), .B(new_n17144), .Y(new_n17146));
  xnor_4 g14798(.A(new_n17146), .B(new_n17143), .Y(n4266));
  xnor_4 g14799(.A(new_n6956), .B(new_n6930), .Y(n4340));
  xnor_4 g14800(.A(new_n16088), .B(new_n5953), .Y(new_n17149));
  xnor_4 g14801(.A(new_n17149), .B(new_n12853), .Y(new_n17150));
  nor_5  g14802(.A(new_n16089), .B(new_n12869), .Y(new_n17151));
  nor_5  g14803(.A(new_n16090), .B(new_n16086), .Y(new_n17152));
  nor_5  g14804(.A(new_n17152), .B(new_n17151), .Y(new_n17153));
  xor_4  g14805(.A(new_n17153), .B(new_n17150), .Y(new_n17154));
  xnor_4 g14806(.A(new_n17154), .B(new_n4999), .Y(new_n17155));
  and_5  g14807(.A(new_n16091), .B(new_n16085), .Y(new_n17156));
  or_5   g14808(.A(new_n17156), .B(new_n16084), .Y(new_n17157));
  xor_4  g14809(.A(new_n17157), .B(new_n17155), .Y(n4374));
  xnor_4 g14810(.A(new_n11085), .B(new_n11034), .Y(n4401));
  xor_4  g14811(.A(new_n12804), .B(new_n12803), .Y(n4424));
  not_8  g14812(.A(n1881), .Y(new_n17161));
  nor_5  g14813(.A(new_n10685), .B(new_n17161), .Y(new_n17162));
  xnor_4 g14814(.A(new_n10685), .B(n1881), .Y(new_n17163_1));
  nor_5  g14815(.A(new_n10677), .B(n5834), .Y(new_n17164));
  xnor_4 g14816(.A(new_n10676), .B(n5834), .Y(new_n17165));
  and_5  g14817(.A(new_n10668), .B(n13851), .Y(new_n17166));
  xnor_4 g14818(.A(new_n10667), .B(n13851), .Y(new_n17167));
  and_5  g14819(.A(new_n10659), .B(n24937), .Y(new_n17168_1));
  or_5   g14820(.A(new_n15984), .B(new_n15978), .Y(new_n17169));
  and_5  g14821(.A(new_n17169), .B(new_n15977), .Y(new_n17170));
  or_5   g14822(.A(new_n17170), .B(new_n17168_1), .Y(new_n17171));
  and_5  g14823(.A(new_n17171), .B(new_n17167), .Y(new_n17172));
  nor_5  g14824(.A(new_n17172), .B(new_n17166), .Y(new_n17173));
  and_5  g14825(.A(new_n17173), .B(new_n17165), .Y(new_n17174));
  nor_5  g14826(.A(new_n17174), .B(new_n17164), .Y(new_n17175));
  and_5  g14827(.A(new_n17175), .B(new_n17163_1), .Y(new_n17176));
  nor_5  g14828(.A(new_n17176), .B(new_n17162), .Y(new_n17177));
  nor_5  g14829(.A(n8827), .B(n4306), .Y(new_n17178));
  not_8  g14830(.A(new_n10680), .Y(new_n17179));
  nor_5  g14831(.A(new_n10684), .B(new_n17179), .Y(new_n17180));
  nor_5  g14832(.A(new_n17180), .B(new_n17178), .Y(new_n17181));
  xnor_4 g14833(.A(new_n17181), .B(new_n17177), .Y(new_n17182));
  not_8  g14834(.A(new_n17182), .Y(new_n17183));
  xnor_4 g14835(.A(new_n17183), .B(new_n9914), .Y(new_n17184));
  xnor_4 g14836(.A(new_n17175), .B(new_n17163_1), .Y(new_n17185));
  nor_5  g14837(.A(new_n17185), .B(new_n9918), .Y(new_n17186));
  xnor_4 g14838(.A(new_n17185), .B(new_n9918), .Y(new_n17187));
  xor_4  g14839(.A(new_n17173), .B(new_n17165), .Y(new_n17188));
  nor_5  g14840(.A(new_n17188), .B(new_n9923), .Y(new_n17189));
  nor_5  g14841(.A(new_n17170), .B(new_n17168_1), .Y(new_n17190));
  xnor_4 g14842(.A(new_n17190), .B(new_n17167), .Y(new_n17191));
  nor_5  g14843(.A(new_n17191), .B(new_n9929), .Y(new_n17192));
  not_8  g14844(.A(new_n17191), .Y(new_n17193));
  xnor_4 g14845(.A(new_n17193), .B(new_n9929), .Y(new_n17194));
  nor_5  g14846(.A(new_n15986_1), .B(new_n9934_1), .Y(new_n17195));
  and_5  g14847(.A(new_n15998), .B(new_n15988), .Y(new_n17196));
  or_5   g14848(.A(new_n17196), .B(new_n17195), .Y(new_n17197));
  and_5  g14849(.A(new_n17197), .B(new_n17194), .Y(new_n17198));
  nor_5  g14850(.A(new_n17198), .B(new_n17192), .Y(new_n17199));
  xnor_4 g14851(.A(new_n17188), .B(new_n9924), .Y(new_n17200));
  and_5  g14852(.A(new_n17200), .B(new_n17199), .Y(new_n17201));
  nor_5  g14853(.A(new_n17201), .B(new_n17189), .Y(new_n17202_1));
  nor_5  g14854(.A(new_n17202_1), .B(new_n17187), .Y(new_n17203));
  nor_5  g14855(.A(new_n17203), .B(new_n17186), .Y(new_n17204));
  xnor_4 g14856(.A(new_n17204), .B(new_n17184), .Y(n4432));
  xnor_4 g14857(.A(new_n14476), .B(new_n14475_1), .Y(n4441));
  nor_5  g14858(.A(n27120), .B(n23065), .Y(new_n17207));
  not_8  g14859(.A(new_n17207), .Y(new_n17208));
  nor_5  g14860(.A(new_n17208), .B(n24786), .Y(new_n17209));
  not_8  g14861(.A(new_n17209), .Y(new_n17210));
  nor_5  g14862(.A(new_n17210), .B(n25370), .Y(new_n17211));
  not_8  g14863(.A(new_n17211), .Y(new_n17212));
  nor_5  g14864(.A(new_n17212), .B(n19472), .Y(new_n17213));
  not_8  g14865(.A(new_n17213), .Y(new_n17214));
  nor_5  g14866(.A(new_n17214), .B(n19042), .Y(new_n17215));
  not_8  g14867(.A(new_n17215), .Y(new_n17216));
  nor_5  g14868(.A(new_n17216), .B(n1293), .Y(new_n17217));
  xnor_4 g14869(.A(new_n17217), .B(n13775), .Y(new_n17218));
  xnor_4 g14870(.A(new_n17218), .B(new_n16533), .Y(new_n17219_1));
  xnor_4 g14871(.A(new_n17215), .B(n1293), .Y(new_n17220));
  nor_5  g14872(.A(new_n17220), .B(new_n16537), .Y(new_n17221));
  xnor_4 g14873(.A(new_n17220), .B(new_n16537), .Y(new_n17222));
  not_8  g14874(.A(new_n16541), .Y(new_n17223));
  xnor_4 g14875(.A(new_n17213), .B(n19042), .Y(new_n17224));
  nor_5  g14876(.A(new_n17224), .B(new_n17223), .Y(new_n17225));
  xnor_4 g14877(.A(new_n17211), .B(n19472), .Y(new_n17226));
  nor_5  g14878(.A(new_n17226), .B(new_n8600), .Y(new_n17227));
  xnor_4 g14879(.A(new_n17226), .B(new_n8599), .Y(new_n17228));
  xnor_4 g14880(.A(new_n17209), .B(n25370), .Y(new_n17229));
  and_5  g14881(.A(new_n17229), .B(new_n8603), .Y(new_n17230));
  xnor_4 g14882(.A(new_n17229), .B(new_n8602), .Y(new_n17231));
  xnor_4 g14883(.A(new_n17207), .B(n24786), .Y(new_n17232_1));
  nor_5  g14884(.A(new_n17232_1), .B(new_n8608_1), .Y(new_n17233));
  xnor_4 g14885(.A(new_n17232_1), .B(new_n8608_1), .Y(new_n17234));
  xnor_4 g14886(.A(n27120), .B(new_n4109), .Y(new_n17235));
  nor_5  g14887(.A(new_n17235), .B(new_n8612), .Y(new_n17236_1));
  nor_5  g14888(.A(new_n17236_1), .B(new_n8614_1), .Y(new_n17237));
  nor_5  g14889(.A(new_n17237), .B(new_n17234), .Y(new_n17238));
  nor_5  g14890(.A(new_n17238), .B(new_n17233), .Y(new_n17239));
  and_5  g14891(.A(new_n17239), .B(new_n17231), .Y(new_n17240));
  nor_5  g14892(.A(new_n17240), .B(new_n17230), .Y(new_n17241));
  and_5  g14893(.A(new_n17241), .B(new_n17228), .Y(new_n17242));
  nor_5  g14894(.A(new_n17242), .B(new_n17227), .Y(new_n17243_1));
  xnor_4 g14895(.A(new_n17224), .B(new_n17223), .Y(new_n17244));
  nor_5  g14896(.A(new_n17244), .B(new_n17243_1), .Y(new_n17245));
  nor_5  g14897(.A(new_n17245), .B(new_n17225), .Y(new_n17246));
  nor_5  g14898(.A(new_n17246), .B(new_n17222), .Y(new_n17247));
  nor_5  g14899(.A(new_n17247), .B(new_n17221), .Y(new_n17248));
  xor_4  g14900(.A(new_n17248), .B(new_n17219_1), .Y(new_n17249));
  not_8  g14901(.A(new_n11917), .Y(new_n17250_1));
  nor_5  g14902(.A(new_n17250_1), .B(n26318), .Y(new_n17251_1));
  xnor_4 g14903(.A(new_n17251_1), .B(n3710), .Y(new_n17252));
  xnor_4 g14904(.A(new_n17252), .B(new_n5340), .Y(new_n17253));
  nor_5  g14905(.A(new_n11918), .B(new_n5348), .Y(new_n17254));
  nor_5  g14906(.A(new_n11945), .B(new_n11919), .Y(new_n17255));
  nor_5  g14907(.A(new_n17255), .B(new_n17254), .Y(new_n17256));
  xor_4  g14908(.A(new_n17256), .B(new_n17253), .Y(new_n17257));
  xnor_4 g14909(.A(new_n17257), .B(new_n17249), .Y(new_n17258));
  xnor_4 g14910(.A(new_n17246), .B(new_n17222), .Y(new_n17259));
  nor_5  g14911(.A(new_n17259), .B(new_n11946), .Y(new_n17260));
  xnor_4 g14912(.A(new_n17259), .B(new_n11946), .Y(new_n17261));
  xnor_4 g14913(.A(new_n17244), .B(new_n17243_1), .Y(new_n17262));
  nor_5  g14914(.A(new_n17262), .B(new_n11980_1), .Y(new_n17263_1));
  xnor_4 g14915(.A(new_n17262), .B(new_n11981), .Y(new_n17264));
  not_8  g14916(.A(new_n11984), .Y(new_n17265));
  xor_4  g14917(.A(new_n17241), .B(new_n17228), .Y(new_n17266));
  nor_5  g14918(.A(new_n17266), .B(new_n17265), .Y(new_n17267));
  xor_4  g14919(.A(new_n17239), .B(new_n17231), .Y(new_n17268));
  nor_5  g14920(.A(new_n17268), .B(new_n11988), .Y(new_n17269));
  xnor_4 g14921(.A(new_n17268), .B(new_n11988), .Y(new_n17270));
  xnor_4 g14922(.A(new_n17237), .B(new_n17234), .Y(new_n17271));
  and_5  g14923(.A(new_n17271), .B(new_n11992), .Y(new_n17272));
  nor_5  g14924(.A(new_n17271), .B(new_n11992), .Y(new_n17273));
  xor_4  g14925(.A(new_n17235), .B(new_n8615), .Y(new_n17274));
  nor_5  g14926(.A(new_n17274), .B(new_n11998), .Y(new_n17275));
  nor_5  g14927(.A(new_n12002), .B(new_n8632), .Y(new_n17276));
  xnor_4 g14928(.A(new_n17274), .B(new_n11998), .Y(new_n17277));
  nor_5  g14929(.A(new_n17277), .B(new_n17276), .Y(new_n17278));
  or_5   g14930(.A(new_n17278), .B(new_n17275), .Y(new_n17279));
  nor_5  g14931(.A(new_n17279), .B(new_n17273), .Y(new_n17280));
  or_5   g14932(.A(new_n17280), .B(new_n17272), .Y(new_n17281));
  nor_5  g14933(.A(new_n17281), .B(new_n17270), .Y(new_n17282));
  or_5   g14934(.A(new_n17282), .B(new_n17269), .Y(new_n17283));
  xnor_4 g14935(.A(new_n17266), .B(new_n17265), .Y(new_n17284));
  nor_5  g14936(.A(new_n17284), .B(new_n17283), .Y(new_n17285_1));
  or_5   g14937(.A(new_n17285_1), .B(new_n17267), .Y(new_n17286));
  not_8  g14938(.A(new_n17286), .Y(new_n17287));
  and_5  g14939(.A(new_n17287), .B(new_n17264), .Y(new_n17288));
  nor_5  g14940(.A(new_n17288), .B(new_n17263_1), .Y(new_n17289));
  nor_5  g14941(.A(new_n17289), .B(new_n17261), .Y(new_n17290));
  nor_5  g14942(.A(new_n17290), .B(new_n17260), .Y(new_n17291));
  xnor_4 g14943(.A(new_n17291), .B(new_n17258), .Y(n4451));
  xnor_4 g14944(.A(n25494), .B(n6659), .Y(new_n17293));
  nor_5  g14945(.A(new_n15667), .B(n10117), .Y(new_n17294));
  xnor_4 g14946(.A(n23250), .B(n10117), .Y(new_n17295));
  nor_5  g14947(.A(n13460), .B(new_n15599), .Y(new_n17296));
  xnor_4 g14948(.A(n13460), .B(n11455), .Y(new_n17297));
  nor_5  g14949(.A(n6104), .B(new_n15602_1), .Y(new_n17298));
  xnor_4 g14950(.A(n6104), .B(n3945), .Y(new_n17299));
  nor_5  g14951(.A(new_n15605), .B(n4119), .Y(new_n17300));
  and_5  g14952(.A(new_n5183), .B(new_n5162), .Y(new_n17301));
  or_5   g14953(.A(new_n17301), .B(new_n17300), .Y(new_n17302_1));
  and_5  g14954(.A(new_n17302_1), .B(new_n17299), .Y(new_n17303));
  or_5   g14955(.A(new_n17303), .B(new_n17298), .Y(new_n17304));
  and_5  g14956(.A(new_n17304), .B(new_n17297), .Y(new_n17305));
  or_5   g14957(.A(new_n17305), .B(new_n17296), .Y(new_n17306));
  and_5  g14958(.A(new_n17306), .B(new_n17295), .Y(new_n17307));
  or_5   g14959(.A(new_n17307), .B(new_n17294), .Y(new_n17308));
  xor_4  g14960(.A(new_n17308), .B(new_n17293), .Y(new_n17309));
  xor_4  g14961(.A(new_n17309), .B(new_n12956_1), .Y(new_n17310));
  xor_4  g14962(.A(new_n17306), .B(new_n17295), .Y(new_n17311));
  nor_5  g14963(.A(new_n17311), .B(new_n12960), .Y(new_n17312));
  xnor_4 g14964(.A(new_n17311), .B(new_n12960), .Y(new_n17313));
  xor_4  g14965(.A(new_n17304), .B(new_n17297), .Y(new_n17314));
  nor_5  g14966(.A(new_n17314), .B(new_n12964), .Y(new_n17315));
  xnor_4 g14967(.A(new_n17314), .B(new_n12964), .Y(new_n17316));
  not_8  g14968(.A(new_n17316), .Y(new_n17317));
  xor_4  g14969(.A(new_n17302_1), .B(new_n17299), .Y(new_n17318));
  and_5  g14970(.A(new_n17318), .B(new_n12968), .Y(new_n17319));
  xnor_4 g14971(.A(new_n17318), .B(new_n12970), .Y(new_n17320_1));
  and_5  g14972(.A(new_n5184_1), .B(new_n5160), .Y(new_n17321));
  and_5  g14973(.A(new_n5217), .B(new_n5185), .Y(new_n17322));
  or_5   g14974(.A(new_n17322), .B(new_n17321), .Y(new_n17323));
  and_5  g14975(.A(new_n17323), .B(new_n17320_1), .Y(new_n17324));
  nor_5  g14976(.A(new_n17324), .B(new_n17319), .Y(new_n17325));
  and_5  g14977(.A(new_n17325), .B(new_n17317), .Y(new_n17326));
  nor_5  g14978(.A(new_n17326), .B(new_n17315), .Y(new_n17327));
  nor_5  g14979(.A(new_n17327), .B(new_n17313), .Y(new_n17328));
  nor_5  g14980(.A(new_n17328), .B(new_n17312), .Y(new_n17329));
  xor_4  g14981(.A(new_n17329), .B(new_n17310), .Y(n4476));
  not_8  g14982(.A(new_n11525), .Y(new_n17331));
  not_8  g14983(.A(new_n4003), .Y(new_n17332));
  nor_5  g14984(.A(new_n17332), .B(n12398), .Y(new_n17333));
  not_8  g14985(.A(new_n17333), .Y(new_n17334));
  nor_5  g14986(.A(new_n17334), .B(n21317), .Y(new_n17335));
  not_8  g14987(.A(new_n17335), .Y(new_n17336));
  nor_5  g14988(.A(new_n17336), .B(n18452), .Y(new_n17337_1));
  and_5  g14989(.A(new_n17337_1), .B(new_n13645), .Y(new_n17338));
  and_5  g14990(.A(new_n17338), .B(new_n6152), .Y(new_n17339));
  xnor_4 g14991(.A(new_n17339), .B(new_n6240), .Y(new_n17340));
  xnor_4 g14992(.A(new_n17338), .B(n1831), .Y(new_n17341));
  nor_5  g14993(.A(new_n17341), .B(new_n6312), .Y(new_n17342));
  xnor_4 g14994(.A(new_n17337_1), .B(n13137), .Y(new_n17343));
  nor_5  g14995(.A(new_n17343), .B(new_n6248_1), .Y(new_n17344_1));
  xnor_4 g14996(.A(new_n17343), .B(new_n6248_1), .Y(new_n17345));
  xnor_4 g14997(.A(new_n17335), .B(n18452), .Y(new_n17346));
  nor_5  g14998(.A(new_n17346), .B(new_n6254), .Y(new_n17347));
  xnor_4 g14999(.A(new_n17346), .B(new_n6259), .Y(new_n17348));
  xnor_4 g15000(.A(new_n17333), .B(n21317), .Y(new_n17349));
  and_5  g15001(.A(new_n17349), .B(new_n6264), .Y(new_n17350));
  xnor_4 g15002(.A(new_n17349), .B(new_n6265), .Y(new_n17351_1));
  and_5  g15003(.A(new_n4043), .B(new_n4004), .Y(new_n17352));
  and_5  g15004(.A(new_n4076), .B(new_n4045), .Y(new_n17353));
  or_5   g15005(.A(new_n17353), .B(new_n17352), .Y(new_n17354));
  and_5  g15006(.A(new_n17354), .B(new_n17351_1), .Y(new_n17355));
  nor_5  g15007(.A(new_n17355), .B(new_n17350), .Y(new_n17356));
  and_5  g15008(.A(new_n17356), .B(new_n17348), .Y(new_n17357));
  nor_5  g15009(.A(new_n17357), .B(new_n17347), .Y(new_n17358));
  nor_5  g15010(.A(new_n17358), .B(new_n17345), .Y(new_n17359_1));
  nor_5  g15011(.A(new_n17359_1), .B(new_n17344_1), .Y(new_n17360));
  xnor_4 g15012(.A(new_n17341), .B(new_n6312), .Y(new_n17361));
  nor_5  g15013(.A(new_n17361), .B(new_n17360), .Y(new_n17362));
  nor_5  g15014(.A(new_n17362), .B(new_n17342), .Y(new_n17363));
  xnor_4 g15015(.A(new_n17363), .B(new_n17340), .Y(new_n17364));
  xnor_4 g15016(.A(new_n17364), .B(new_n17331), .Y(new_n17365));
  xnor_4 g15017(.A(new_n17361), .B(new_n17360), .Y(new_n17366));
  nor_5  g15018(.A(new_n17366), .B(new_n11530), .Y(new_n17367));
  xnor_4 g15019(.A(new_n17366), .B(new_n11530), .Y(new_n17368));
  xnor_4 g15020(.A(new_n17358), .B(new_n17345), .Y(new_n17369));
  nor_5  g15021(.A(new_n17369), .B(new_n11534), .Y(new_n17370));
  xnor_4 g15022(.A(new_n17369), .B(new_n11534), .Y(new_n17371));
  xnor_4 g15023(.A(new_n17356), .B(new_n17348), .Y(new_n17372));
  nor_5  g15024(.A(new_n17372), .B(new_n11539), .Y(new_n17373));
  xnor_4 g15025(.A(new_n17372), .B(new_n11539), .Y(new_n17374));
  xor_4  g15026(.A(new_n17354), .B(new_n17351_1), .Y(new_n17375));
  nor_5  g15027(.A(new_n17375), .B(new_n11543), .Y(new_n17376));
  xnor_4 g15028(.A(new_n17375), .B(new_n11543), .Y(new_n17377));
  nor_5  g15029(.A(new_n4077), .B(new_n3996), .Y(new_n17378));
  nor_5  g15030(.A(new_n4104), .B(new_n4078), .Y(new_n17379));
  nor_5  g15031(.A(new_n17379), .B(new_n17378), .Y(new_n17380));
  nor_5  g15032(.A(new_n17380), .B(new_n17377), .Y(new_n17381));
  nor_5  g15033(.A(new_n17381), .B(new_n17376), .Y(new_n17382));
  nor_5  g15034(.A(new_n17382), .B(new_n17374), .Y(new_n17383));
  nor_5  g15035(.A(new_n17383), .B(new_n17373), .Y(new_n17384));
  nor_5  g15036(.A(new_n17384), .B(new_n17371), .Y(new_n17385));
  nor_5  g15037(.A(new_n17385), .B(new_n17370), .Y(new_n17386));
  nor_5  g15038(.A(new_n17386), .B(new_n17368), .Y(new_n17387_1));
  nor_5  g15039(.A(new_n17387_1), .B(new_n17367), .Y(new_n17388));
  xnor_4 g15040(.A(new_n17388), .B(new_n17365), .Y(n4478));
  xnor_4 g15041(.A(new_n12302_1), .B(new_n12270), .Y(n4529));
  xnor_4 g15042(.A(new_n6145), .B(new_n6099), .Y(n4552));
  xnor_4 g15043(.A(new_n6141), .B(new_n6109), .Y(n4595));
  xnor_4 g15044(.A(new_n13982), .B(new_n13948), .Y(n4624));
  not_8  g15045(.A(new_n16886), .Y(new_n17394));
  nor_5  g15046(.A(new_n17394), .B(n2659), .Y(new_n17395));
  xnor_4 g15047(.A(new_n17395), .B(n2858), .Y(new_n17396));
  nor_5  g15048(.A(new_n17396), .B(n14899), .Y(new_n17397));
  xnor_4 g15049(.A(new_n17396), .B(n14899), .Y(new_n17398));
  nor_5  g15050(.A(new_n16887), .B(n18444), .Y(new_n17399));
  nor_5  g15051(.A(new_n16896), .B(new_n16888), .Y(new_n17400));
  nor_5  g15052(.A(new_n17400), .B(new_n17399), .Y(new_n17401));
  nor_5  g15053(.A(new_n17401), .B(new_n17398), .Y(new_n17402));
  nor_5  g15054(.A(new_n17402), .B(new_n17397), .Y(new_n17403));
  and_5  g15055(.A(new_n17395), .B(new_n4909), .Y(new_n17404));
  xnor_4 g15056(.A(new_n17404), .B(n3740), .Y(new_n17405));
  xnor_4 g15057(.A(new_n17405), .B(new_n8323), .Y(new_n17406));
  xnor_4 g15058(.A(new_n17406), .B(new_n17403), .Y(new_n17407));
  nor_5  g15059(.A(new_n17407), .B(new_n7703), .Y(new_n17408));
  xnor_4 g15060(.A(new_n17407), .B(new_n7703), .Y(new_n17409));
  xnor_4 g15061(.A(new_n17401), .B(new_n17398), .Y(new_n17410));
  and_5  g15062(.A(new_n17410), .B(new_n7706), .Y(new_n17411));
  xnor_4 g15063(.A(new_n17410), .B(new_n7706), .Y(new_n17412));
  nor_5  g15064(.A(new_n16897), .B(new_n7715), .Y(new_n17413));
  nor_5  g15065(.A(new_n16906), .B(new_n16898), .Y(new_n17414));
  nor_5  g15066(.A(new_n17414), .B(new_n17413), .Y(new_n17415));
  nor_5  g15067(.A(new_n17415), .B(new_n17412), .Y(new_n17416));
  nor_5  g15068(.A(new_n17416), .B(new_n17411), .Y(new_n17417));
  nor_5  g15069(.A(new_n17417), .B(new_n17409), .Y(new_n17418));
  nor_5  g15070(.A(new_n17418), .B(new_n17408), .Y(new_n17419));
  and_5  g15071(.A(new_n17404), .B(new_n4907), .Y(new_n17420));
  and_5  g15072(.A(new_n17405), .B(n3506), .Y(new_n17421_1));
  or_5   g15073(.A(new_n17405), .B(n3506), .Y(new_n17422));
  and_5  g15074(.A(new_n17422), .B(new_n17403), .Y(new_n17423));
  or_5   g15075(.A(new_n17423), .B(new_n17421_1), .Y(new_n17424));
  nor_5  g15076(.A(new_n17424), .B(new_n17420), .Y(new_n17425));
  xnor_4 g15077(.A(new_n17425), .B(new_n17419), .Y(new_n17426));
  xnor_4 g15078(.A(new_n17426), .B(new_n7649), .Y(new_n17427));
  not_8  g15079(.A(new_n17427), .Y(new_n17428));
  xnor_4 g15080(.A(new_n17428), .B(new_n13394), .Y(new_n17429));
  xor_4  g15081(.A(new_n17417), .B(new_n17409), .Y(new_n17430));
  nor_5  g15082(.A(new_n17430), .B(new_n7840), .Y(new_n17431));
  xnor_4 g15083(.A(new_n17415), .B(new_n17412), .Y(new_n17432_1));
  not_8  g15084(.A(new_n17432_1), .Y(new_n17433));
  nor_5  g15085(.A(new_n17433), .B(new_n7849), .Y(new_n17434));
  xnor_4 g15086(.A(new_n17433), .B(new_n7849), .Y(new_n17435));
  not_8  g15087(.A(new_n16907), .Y(new_n17436_1));
  nor_5  g15088(.A(new_n17436_1), .B(new_n7856), .Y(new_n17437));
  xnor_4 g15089(.A(new_n17436_1), .B(new_n7856), .Y(new_n17438));
  nor_5  g15090(.A(new_n16920), .B(new_n7861), .Y(new_n17439));
  xnor_4 g15091(.A(new_n16920), .B(new_n7860), .Y(new_n17440_1));
  not_8  g15092(.A(new_n13044_1), .Y(new_n17441));
  nor_5  g15093(.A(new_n17441), .B(new_n7866), .Y(new_n17442));
  nor_5  g15094(.A(new_n13068), .B(new_n7870), .Y(new_n17443));
  nor_5  g15095(.A(new_n16755), .B(new_n16741), .Y(new_n17444));
  nor_5  g15096(.A(new_n17444), .B(new_n17443), .Y(new_n17445));
  xnor_4 g15097(.A(new_n13044_1), .B(new_n7866), .Y(new_n17446));
  and_5  g15098(.A(new_n17446), .B(new_n17445), .Y(new_n17447));
  nor_5  g15099(.A(new_n17447), .B(new_n17442), .Y(new_n17448));
  and_5  g15100(.A(new_n17448), .B(new_n17440_1), .Y(new_n17449));
  nor_5  g15101(.A(new_n17449), .B(new_n17439), .Y(new_n17450_1));
  nor_5  g15102(.A(new_n17450_1), .B(new_n17438), .Y(new_n17451));
  nor_5  g15103(.A(new_n17451), .B(new_n17437), .Y(new_n17452));
  nor_5  g15104(.A(new_n17452), .B(new_n17435), .Y(new_n17453));
  nor_5  g15105(.A(new_n17453), .B(new_n17434), .Y(new_n17454));
  xnor_4 g15106(.A(new_n17430), .B(new_n7840), .Y(new_n17455));
  nor_5  g15107(.A(new_n17455), .B(new_n17454), .Y(new_n17456));
  nor_5  g15108(.A(new_n17456), .B(new_n17431), .Y(new_n17457));
  xor_4  g15109(.A(new_n17457), .B(new_n17429), .Y(n4646));
  xnor_4 g15110(.A(new_n13990), .B(new_n13932), .Y(n4674));
  xnor_4 g15111(.A(n7057), .B(n3480), .Y(new_n17460));
  nor_5  g15112(.A(new_n7625), .B(n8381), .Y(new_n17461_1));
  nor_5  g15113(.A(n16722), .B(new_n8510_1), .Y(new_n17462));
  nor_5  g15114(.A(n20235), .B(new_n5784), .Y(new_n17463));
  or_5   g15115(.A(new_n5040), .B(n11486), .Y(new_n17464));
  nor_5  g15116(.A(new_n2383), .B(n12495), .Y(new_n17465));
  and_5  g15117(.A(new_n17465), .B(new_n17464), .Y(new_n17466_1));
  nor_5  g15118(.A(new_n17466_1), .B(new_n17463), .Y(new_n17467));
  nor_5  g15119(.A(new_n17467), .B(new_n17462), .Y(new_n17468));
  or_5   g15120(.A(new_n17468), .B(new_n17461_1), .Y(new_n17469));
  xor_4  g15121(.A(new_n17469), .B(new_n17460), .Y(new_n17470));
  xnor_4 g15122(.A(new_n17470), .B(new_n3052), .Y(new_n17471));
  xnor_4 g15123(.A(n16722), .B(n8381), .Y(new_n17472));
  xnor_4 g15124(.A(new_n17472), .B(new_n17467), .Y(new_n17473));
  and_5  g15125(.A(new_n17473), .B(new_n3057), .Y(new_n17474));
  xnor_4 g15126(.A(new_n17473), .B(new_n3057), .Y(new_n17475));
  xnor_4 g15127(.A(n13781), .B(n12495), .Y(new_n17476));
  nor_5  g15128(.A(new_n17476), .B(new_n3064), .Y(new_n17477));
  nor_5  g15129(.A(new_n17477), .B(new_n3069), .Y(new_n17478));
  xnor_4 g15130(.A(new_n17477), .B(new_n3069), .Y(new_n17479));
  xnor_4 g15131(.A(n20235), .B(n11486), .Y(new_n17480));
  xnor_4 g15132(.A(new_n17480), .B(new_n17465), .Y(new_n17481));
  nor_5  g15133(.A(new_n17481), .B(new_n17479), .Y(new_n17482));
  nor_5  g15134(.A(new_n17482), .B(new_n17478), .Y(new_n17483));
  nor_5  g15135(.A(new_n17483), .B(new_n17475), .Y(new_n17484));
  nor_5  g15136(.A(new_n17484), .B(new_n17474), .Y(new_n17485));
  xor_4  g15137(.A(new_n17485), .B(new_n17471), .Y(n4693));
  xnor_4 g15138(.A(new_n10597), .B(new_n10587), .Y(n4731));
  nor_5  g15139(.A(new_n6022_1), .B(new_n5981), .Y(new_n17488));
  or_5   g15140(.A(new_n6086), .B(new_n6028), .Y(new_n17489));
  and_5  g15141(.A(new_n17489), .B(new_n6024), .Y(new_n17490));
  nor_5  g15142(.A(new_n17490), .B(new_n17488), .Y(new_n17491));
  nor_5  g15143(.A(n21784), .B(n3582), .Y(new_n17492));
  or_5   g15144(.A(new_n6020), .B(new_n5984), .Y(new_n17493_1));
  and_5  g15145(.A(new_n17493_1), .B(new_n5983), .Y(new_n17494));
  nor_5  g15146(.A(new_n17494), .B(new_n17492), .Y(new_n17495));
  not_8  g15147(.A(new_n17495), .Y(new_n17496));
  nor_5  g15148(.A(new_n17496), .B(new_n17491), .Y(new_n17497));
  not_8  g15149(.A(new_n17497), .Y(new_n17498));
  xnor_4 g15150(.A(new_n17498), .B(new_n15097), .Y(new_n17499));
  xnor_4 g15151(.A(new_n17495), .B(new_n17491), .Y(new_n17500_1));
  nor_5  g15152(.A(new_n17500_1), .B(new_n15101), .Y(new_n17501));
  xnor_4 g15153(.A(new_n17500_1), .B(new_n15101), .Y(new_n17502));
  and_5  g15154(.A(new_n12694), .B(new_n12670_1), .Y(new_n17503));
  nor_5  g15155(.A(new_n12732), .B(new_n12695), .Y(new_n17504));
  nor_5  g15156(.A(new_n17504), .B(new_n17503), .Y(new_n17505));
  nor_5  g15157(.A(new_n17505), .B(new_n17502), .Y(new_n17506));
  nor_5  g15158(.A(new_n17506), .B(new_n17501), .Y(new_n17507));
  xnor_4 g15159(.A(new_n17507), .B(new_n17499), .Y(n4745));
  xnor_4 g15160(.A(new_n6288), .B(n6773), .Y(new_n17509));
  xnor_4 g15161(.A(new_n17509), .B(new_n9686), .Y(n4747));
  xnor_4 g15162(.A(new_n5747), .B(new_n5746), .Y(n4766));
  xnor_4 g15163(.A(new_n13478), .B(new_n13461), .Y(n4770));
  xnor_4 g15164(.A(new_n16115), .B(new_n15308), .Y(n4777));
  xnor_4 g15165(.A(n17959), .B(n6861), .Y(new_n17514));
  and_5  g15166(.A(n19357), .B(new_n5468), .Y(new_n17515));
  xnor_4 g15167(.A(n19357), .B(n7566), .Y(new_n17516));
  and_5  g15168(.A(new_n5471), .B(n2328), .Y(new_n17517));
  xnor_4 g15169(.A(n7731), .B(n2328), .Y(new_n17518));
  nor_5  g15170(.A(n15053), .B(new_n5475), .Y(new_n17519));
  nor_5  g15171(.A(new_n15611), .B(n12341), .Y(new_n17520));
  nor_5  g15172(.A(n25471), .B(new_n5478), .Y(new_n17521));
  or_5   g15173(.A(new_n5066), .B(n20986), .Y(new_n17522));
  nor_5  g15174(.A(n16502), .B(new_n5798), .Y(new_n17523));
  and_5  g15175(.A(new_n17523), .B(new_n17522), .Y(new_n17524_1));
  nor_5  g15176(.A(new_n17524_1), .B(new_n17521), .Y(new_n17525));
  nor_5  g15177(.A(new_n17525), .B(new_n17520), .Y(new_n17526));
  nor_5  g15178(.A(new_n17526), .B(new_n17519), .Y(new_n17527));
  and_5  g15179(.A(new_n17527), .B(new_n17518), .Y(new_n17528));
  or_5   g15180(.A(new_n17528), .B(new_n17517), .Y(new_n17529_1));
  and_5  g15181(.A(new_n17529_1), .B(new_n17516), .Y(new_n17530));
  or_5   g15182(.A(new_n17530), .B(new_n17515), .Y(new_n17531));
  xor_4  g15183(.A(new_n17531), .B(new_n17514), .Y(new_n17532));
  nor_5  g15184(.A(n20077), .B(n6794), .Y(new_n17533));
  not_8  g15185(.A(new_n17533), .Y(new_n17534));
  nor_5  g15186(.A(new_n17534), .B(n15636), .Y(new_n17535));
  not_8  g15187(.A(new_n17535), .Y(new_n17536));
  nor_5  g15188(.A(new_n17536), .B(n8745), .Y(new_n17537));
  not_8  g15189(.A(new_n17537), .Y(new_n17538));
  nor_5  g15190(.A(new_n17538), .B(n1777), .Y(new_n17539));
  xnor_4 g15191(.A(new_n17539), .B(n22660), .Y(new_n17540));
  xnor_4 g15192(.A(new_n17540), .B(n11580), .Y(new_n17541));
  xnor_4 g15193(.A(new_n17537), .B(n1777), .Y(new_n17542));
  nor_5  g15194(.A(new_n17542), .B(new_n5576), .Y(new_n17543));
  xnor_4 g15195(.A(new_n17542), .B(n15884), .Y(new_n17544));
  xnor_4 g15196(.A(new_n17535), .B(n8745), .Y(new_n17545));
  nor_5  g15197(.A(new_n17545), .B(new_n5595), .Y(new_n17546));
  xnor_4 g15198(.A(new_n17545), .B(new_n5595), .Y(new_n17547));
  xnor_4 g15199(.A(new_n17533), .B(n15636), .Y(new_n17548));
  nor_5  g15200(.A(new_n17548), .B(new_n5582), .Y(new_n17549));
  xnor_4 g15201(.A(new_n17548), .B(n27104), .Y(new_n17550));
  xnor_4 g15202(.A(n20077), .B(new_n2447), .Y(new_n17551));
  nor_5  g15203(.A(new_n17551), .B(new_n5584), .Y(new_n17552));
  nor_5  g15204(.A(n6794), .B(new_n5588), .Y(new_n17553));
  xnor_4 g15205(.A(new_n17551), .B(n27188), .Y(new_n17554));
  and_5  g15206(.A(new_n17554), .B(new_n17553), .Y(new_n17555));
  or_5   g15207(.A(new_n17555), .B(new_n17552), .Y(new_n17556));
  and_5  g15208(.A(new_n17556), .B(new_n17550), .Y(new_n17557_1));
  nor_5  g15209(.A(new_n17557_1), .B(new_n17549), .Y(new_n17558));
  nor_5  g15210(.A(new_n17558), .B(new_n17547), .Y(new_n17559));
  or_5   g15211(.A(new_n17559), .B(new_n17546), .Y(new_n17560));
  and_5  g15212(.A(new_n17560), .B(new_n17544), .Y(new_n17561));
  or_5   g15213(.A(new_n17561), .B(new_n17543), .Y(new_n17562));
  xor_4  g15214(.A(new_n17562), .B(new_n17541), .Y(new_n17563));
  xnor_4 g15215(.A(new_n17563), .B(new_n15581), .Y(new_n17564));
  xor_4  g15216(.A(new_n17560), .B(new_n17544), .Y(new_n17565));
  nor_5  g15217(.A(new_n17565), .B(new_n14991), .Y(new_n17566));
  xnor_4 g15218(.A(new_n17558), .B(new_n17547), .Y(new_n17567));
  nor_5  g15219(.A(new_n17567), .B(new_n14996), .Y(new_n17568));
  xnor_4 g15220(.A(new_n17567), .B(new_n14994), .Y(new_n17569));
  xor_4  g15221(.A(new_n17556), .B(new_n17550), .Y(new_n17570));
  nor_5  g15222(.A(new_n17570), .B(new_n5037), .Y(new_n17571));
  xnor_4 g15223(.A(new_n17570), .B(new_n5037), .Y(new_n17572));
  xnor_4 g15224(.A(new_n17554), .B(new_n17553), .Y(new_n17573));
  not_8  g15225(.A(new_n17573), .Y(new_n17574));
  nor_5  g15226(.A(new_n17574), .B(new_n5048), .Y(new_n17575));
  xnor_4 g15227(.A(n6794), .B(n6611), .Y(new_n17576));
  nor_5  g15228(.A(new_n17576), .B(new_n5042), .Y(new_n17577));
  xnor_4 g15229(.A(new_n17574), .B(new_n5076), .Y(new_n17578));
  and_5  g15230(.A(new_n17578), .B(new_n17577), .Y(new_n17579));
  nor_5  g15231(.A(new_n17579), .B(new_n17575), .Y(new_n17580));
  nor_5  g15232(.A(new_n17580), .B(new_n17572), .Y(new_n17581));
  nor_5  g15233(.A(new_n17581), .B(new_n17571), .Y(new_n17582));
  and_5  g15234(.A(new_n17582), .B(new_n17569), .Y(new_n17583_1));
  nor_5  g15235(.A(new_n17583_1), .B(new_n17568), .Y(new_n17584));
  xor_4  g15236(.A(new_n17565), .B(new_n14991), .Y(new_n17585));
  and_5  g15237(.A(new_n17585), .B(new_n17584), .Y(new_n17586));
  nor_5  g15238(.A(new_n17586), .B(new_n17566), .Y(new_n17587));
  xnor_4 g15239(.A(new_n17587), .B(new_n17564), .Y(new_n17588));
  xnor_4 g15240(.A(new_n17588), .B(new_n17532), .Y(new_n17589));
  xor_4  g15241(.A(new_n17529_1), .B(new_n17516), .Y(new_n17590));
  xor_4  g15242(.A(new_n17585), .B(new_n17584), .Y(new_n17591));
  nor_5  g15243(.A(new_n17591), .B(new_n17590), .Y(new_n17592_1));
  xnor_4 g15244(.A(new_n17591), .B(new_n17590), .Y(new_n17593));
  xnor_4 g15245(.A(new_n17582), .B(new_n17569), .Y(new_n17594));
  not_8  g15246(.A(new_n17594), .Y(new_n17595));
  xnor_4 g15247(.A(new_n17527), .B(new_n17518), .Y(new_n17596));
  and_5  g15248(.A(new_n17596), .B(new_n17595), .Y(new_n17597));
  xnor_4 g15249(.A(new_n17596), .B(new_n17595), .Y(new_n17598));
  xnor_4 g15250(.A(new_n17580), .B(new_n17572), .Y(new_n17599));
  xnor_4 g15251(.A(n15053), .B(n12341), .Y(new_n17600));
  xnor_4 g15252(.A(new_n17600), .B(new_n17525), .Y(new_n17601));
  and_5  g15253(.A(new_n17601), .B(new_n17599), .Y(new_n17602));
  xnor_4 g15254(.A(new_n17601), .B(new_n17599), .Y(new_n17603));
  xnor_4 g15255(.A(new_n17576), .B(new_n5041), .Y(new_n17604));
  not_8  g15256(.A(new_n17604), .Y(new_n17605));
  xnor_4 g15257(.A(n16502), .B(n12384), .Y(new_n17606));
  nor_5  g15258(.A(new_n17606), .B(new_n17605), .Y(new_n17607));
  xnor_4 g15259(.A(n25471), .B(n20986), .Y(new_n17608));
  xnor_4 g15260(.A(new_n17608), .B(new_n17523), .Y(new_n17609));
  nor_5  g15261(.A(new_n17609), .B(new_n17607), .Y(new_n17610));
  xnor_4 g15262(.A(new_n17578), .B(new_n17577), .Y(new_n17611));
  not_8  g15263(.A(new_n17611), .Y(new_n17612));
  xnor_4 g15264(.A(new_n17609), .B(new_n17607), .Y(new_n17613));
  nor_5  g15265(.A(new_n17613), .B(new_n17612), .Y(new_n17614));
  nor_5  g15266(.A(new_n17614), .B(new_n17610), .Y(new_n17615));
  nor_5  g15267(.A(new_n17615), .B(new_n17603), .Y(new_n17616));
  nor_5  g15268(.A(new_n17616), .B(new_n17602), .Y(new_n17617));
  nor_5  g15269(.A(new_n17617), .B(new_n17598), .Y(new_n17618));
  nor_5  g15270(.A(new_n17618), .B(new_n17597), .Y(new_n17619));
  nor_5  g15271(.A(new_n17619), .B(new_n17593), .Y(new_n17620));
  nor_5  g15272(.A(new_n17620), .B(new_n17592_1), .Y(new_n17621));
  xor_4  g15273(.A(new_n17621), .B(new_n17589), .Y(n4785));
  xnor_4 g15274(.A(new_n13777), .B(new_n13745), .Y(n4804));
  xnor_4 g15275(.A(new_n15317), .B(new_n15298), .Y(n4810));
  not_8  g15276(.A(n23166), .Y(new_n17625));
  nor_5  g15277(.A(new_n17625), .B(n18105), .Y(new_n17626));
  or_5   g15278(.A(new_n9117), .B(new_n9080), .Y(new_n17627));
  and_5  g15279(.A(new_n17627), .B(new_n9078), .Y(new_n17628));
  nor_5  g15280(.A(new_n17628), .B(new_n17626), .Y(new_n17629));
  nor_5  g15281(.A(new_n10686), .B(new_n7961), .Y(new_n17630));
  and_5  g15282(.A(new_n10730), .B(new_n10687), .Y(new_n17631));
  nor_5  g15283(.A(new_n17631), .B(new_n17630), .Y(new_n17632));
  and_5  g15284(.A(new_n10685), .B(new_n10678), .Y(new_n17633));
  not_8  g15285(.A(new_n17181), .Y(new_n17634));
  nor_5  g15286(.A(new_n17634), .B(new_n17633), .Y(new_n17635));
  and_5  g15287(.A(new_n17633), .B(new_n17178), .Y(new_n17636));
  nor_5  g15288(.A(new_n17636), .B(new_n17635), .Y(new_n17637));
  xnor_4 g15289(.A(new_n17637), .B(new_n8027_1), .Y(new_n17638_1));
  xnor_4 g15290(.A(new_n17638_1), .B(new_n17632), .Y(new_n17639));
  and_5  g15291(.A(new_n17639), .B(new_n17629), .Y(new_n17640));
  xnor_4 g15292(.A(new_n17639), .B(new_n17629), .Y(new_n17641));
  and_5  g15293(.A(new_n10731), .B(new_n9119), .Y(new_n17642));
  nor_5  g15294(.A(new_n10775_1), .B(new_n10732), .Y(new_n17643));
  nor_5  g15295(.A(new_n17643), .B(new_n17642), .Y(new_n17644));
  nor_5  g15296(.A(new_n17644), .B(new_n17641), .Y(new_n17645));
  nor_5  g15297(.A(new_n17645), .B(new_n17640), .Y(new_n17646));
  or_5   g15298(.A(new_n17637), .B(new_n8026), .Y(new_n17647));
  and_5  g15299(.A(new_n17647), .B(new_n17632), .Y(new_n17648));
  and_5  g15300(.A(new_n17637), .B(new_n8026), .Y(new_n17649));
  or_5   g15301(.A(new_n17649), .B(new_n17636), .Y(new_n17650));
  or_5   g15302(.A(new_n17650), .B(new_n17648), .Y(new_n17651));
  nand_5 g15303(.A(new_n17651), .B(new_n17646), .Y(n4814));
  xnor_4 g15304(.A(new_n15909), .B(new_n15908), .Y(n4850));
  xnor_4 g15305(.A(new_n16726), .B(new_n16687), .Y(n4891));
  xnor_4 g15306(.A(new_n16876), .B(new_n16855), .Y(n4925));
  xnor_4 g15307(.A(new_n15915), .B(new_n15898), .Y(n4947));
  xnor_4 g15308(.A(new_n9378), .B(new_n9377), .Y(n4952));
  xnor_4 g15309(.A(n25068), .B(n6790), .Y(new_n17658));
  not_8  g15310(.A(n2331), .Y(new_n17659));
  nor_5  g15311(.A(n22879), .B(new_n17659), .Y(new_n17660));
  xnor_4 g15312(.A(n22879), .B(n2331), .Y(new_n17661));
  not_8  g15313(.A(n22631), .Y(new_n17662));
  nor_5  g15314(.A(new_n17662), .B(n2117), .Y(new_n17663));
  xnor_4 g15315(.A(n22631), .B(n2117), .Y(new_n17664_1));
  and_5  g15316(.A(new_n7993), .B(n5882), .Y(new_n17665));
  nor_5  g15317(.A(new_n7993), .B(n5882), .Y(new_n17666));
  nor_5  g15318(.A(n15258), .B(new_n9793), .Y(new_n17667));
  nor_5  g15319(.A(new_n9790), .B(n4588), .Y(new_n17668));
  not_8  g15320(.A(new_n17668), .Y(new_n17669));
  nor_5  g15321(.A(new_n7998), .B(n11775), .Y(new_n17670));
  nor_5  g15322(.A(new_n17670), .B(new_n17669), .Y(new_n17671));
  nor_5  g15323(.A(new_n17671), .B(new_n17667), .Y(new_n17672));
  nor_5  g15324(.A(new_n17672), .B(new_n17666), .Y(new_n17673));
  nor_5  g15325(.A(new_n17673), .B(new_n17665), .Y(new_n17674));
  and_5  g15326(.A(new_n17674), .B(new_n17664_1), .Y(new_n17675));
  or_5   g15327(.A(new_n17675), .B(new_n17663), .Y(new_n17676));
  and_5  g15328(.A(new_n17676), .B(new_n17661), .Y(new_n17677));
  or_5   g15329(.A(new_n17677), .B(new_n17660), .Y(new_n17678));
  xor_4  g15330(.A(new_n17678), .B(new_n17658), .Y(new_n17679));
  xnor_4 g15331(.A(new_n17679), .B(new_n14940), .Y(new_n17680));
  xor_4  g15332(.A(new_n17676), .B(new_n17661), .Y(new_n17681));
  nor_5  g15333(.A(new_n17681), .B(new_n14948), .Y(new_n17682));
  xnor_4 g15334(.A(new_n17681), .B(new_n14948), .Y(new_n17683));
  xnor_4 g15335(.A(new_n17674), .B(new_n17664_1), .Y(new_n17684));
  and_5  g15336(.A(new_n17684), .B(new_n14952), .Y(new_n17685));
  xnor_4 g15337(.A(new_n17684), .B(new_n14953), .Y(new_n17686));
  xnor_4 g15338(.A(n16743), .B(n5882), .Y(new_n17687_1));
  xnor_4 g15339(.A(new_n17687_1), .B(new_n17672), .Y(new_n17688));
  nor_5  g15340(.A(new_n17688), .B(new_n14956), .Y(new_n17689));
  xnor_4 g15341(.A(new_n17688), .B(new_n14956), .Y(new_n17690));
  xnor_4 g15342(.A(n15258), .B(n11775), .Y(new_n17691));
  xnor_4 g15343(.A(new_n17691), .B(new_n17669), .Y(new_n17692));
  nor_5  g15344(.A(new_n17692), .B(new_n14960), .Y(new_n17693));
  nor_5  g15345(.A(new_n14744), .B(new_n14962), .Y(new_n17694));
  xnor_4 g15346(.A(new_n17692), .B(new_n15203), .Y(new_n17695));
  and_5  g15347(.A(new_n17695), .B(new_n17694), .Y(new_n17696));
  nor_5  g15348(.A(new_n17696), .B(new_n17693), .Y(new_n17697));
  nor_5  g15349(.A(new_n17697), .B(new_n17690), .Y(new_n17698));
  nor_5  g15350(.A(new_n17698), .B(new_n17689), .Y(new_n17699));
  and_5  g15351(.A(new_n17699), .B(new_n17686), .Y(new_n17700));
  nor_5  g15352(.A(new_n17700), .B(new_n17685), .Y(new_n17701));
  nor_5  g15353(.A(new_n17701), .B(new_n17683), .Y(new_n17702));
  nor_5  g15354(.A(new_n17702), .B(new_n17682), .Y(new_n17703));
  xor_4  g15355(.A(new_n17703), .B(new_n17680), .Y(new_n17704));
  xnor_4 g15356(.A(new_n17704), .B(new_n14871), .Y(new_n17705));
  xnor_4 g15357(.A(new_n17701), .B(new_n17683), .Y(new_n17706));
  nor_5  g15358(.A(new_n17706), .B(new_n14874), .Y(new_n17707));
  xnor_4 g15359(.A(new_n17706), .B(new_n14874), .Y(new_n17708));
  xnor_4 g15360(.A(new_n17699), .B(new_n17686), .Y(new_n17709));
  nor_5  g15361(.A(new_n17709), .B(new_n13334), .Y(new_n17710));
  not_8  g15362(.A(new_n17709), .Y(new_n17711));
  xnor_4 g15363(.A(new_n17711), .B(new_n13335), .Y(new_n17712));
  xnor_4 g15364(.A(new_n17697), .B(new_n17690), .Y(new_n17713));
  not_8  g15365(.A(new_n17713), .Y(new_n17714));
  nor_5  g15366(.A(new_n17714), .B(new_n13341), .Y(new_n17715));
  xnor_4 g15367(.A(new_n17714), .B(new_n13341), .Y(new_n17716));
  not_8  g15368(.A(new_n14745), .Y(new_n17717));
  nor_5  g15369(.A(new_n17717), .B(new_n9885), .Y(new_n17718));
  nor_5  g15370(.A(new_n17718), .B(new_n13384), .Y(new_n17719));
  xnor_4 g15371(.A(new_n17718), .B(new_n13384), .Y(new_n17720));
  xor_4  g15372(.A(new_n17695), .B(new_n17694), .Y(new_n17721_1));
  nor_5  g15373(.A(new_n17721_1), .B(new_n17720), .Y(new_n17722));
  nor_5  g15374(.A(new_n17722), .B(new_n17719), .Y(new_n17723));
  nor_5  g15375(.A(new_n17723), .B(new_n17716), .Y(new_n17724));
  nor_5  g15376(.A(new_n17724), .B(new_n17715), .Y(new_n17725));
  nor_5  g15377(.A(new_n17725), .B(new_n17712), .Y(new_n17726));
  nor_5  g15378(.A(new_n17726), .B(new_n17710), .Y(new_n17727));
  nor_5  g15379(.A(new_n17727), .B(new_n17708), .Y(new_n17728));
  nor_5  g15380(.A(new_n17728), .B(new_n17707), .Y(new_n17729));
  xnor_4 g15381(.A(new_n17729), .B(new_n17705), .Y(n4966));
  xnor_4 g15382(.A(new_n17200), .B(new_n17199), .Y(n4972));
  and_5  g15383(.A(new_n7524_1), .B(new_n5453), .Y(new_n17732));
  xnor_4 g15384(.A(new_n7524_1), .B(n23895), .Y(new_n17733));
  nor_5  g15385(.A(new_n7528), .B(new_n5456), .Y(new_n17734));
  xnor_4 g15386(.A(new_n7528), .B(new_n5456), .Y(new_n17735_1));
  nor_5  g15387(.A(new_n7533), .B(new_n5459), .Y(new_n17736));
  nor_5  g15388(.A(new_n16563), .B(new_n16552), .Y(new_n17737));
  nor_5  g15389(.A(new_n17737), .B(new_n17736), .Y(new_n17738_1));
  nor_5  g15390(.A(new_n17738_1), .B(new_n17735_1), .Y(new_n17739));
  nor_5  g15391(.A(new_n17739), .B(new_n17734), .Y(new_n17740));
  and_5  g15392(.A(new_n17740), .B(new_n17733), .Y(new_n17741));
  nor_5  g15393(.A(new_n17741), .B(new_n17732), .Y(new_n17742));
  not_8  g15394(.A(new_n17742), .Y(new_n17743));
  nor_5  g15395(.A(new_n17743), .B(new_n7519), .Y(new_n17744));
  not_8  g15396(.A(new_n17744), .Y(new_n17745));
  not_8  g15397(.A(new_n16516_1), .Y(new_n17746_1));
  nor_5  g15398(.A(new_n17746_1), .B(n2289), .Y(new_n17747));
  and_5  g15399(.A(new_n17747), .B(new_n6744), .Y(new_n17748));
  xnor_4 g15400(.A(new_n17748), .B(n2978), .Y(new_n17749_1));
  xnor_4 g15401(.A(new_n17749_1), .B(new_n16488), .Y(new_n17750));
  xnor_4 g15402(.A(new_n17747), .B(n23697), .Y(new_n17751));
  and_5  g15403(.A(new_n17751), .B(n337), .Y(new_n17752));
  nor_5  g15404(.A(new_n17751), .B(n337), .Y(new_n17753));
  and_5  g15405(.A(new_n16517_1), .B(n3228), .Y(new_n17754));
  or_5   g15406(.A(new_n16517_1), .B(n3228), .Y(new_n17755));
  and_5  g15407(.A(new_n16532), .B(new_n17755), .Y(new_n17756));
  nor_5  g15408(.A(new_n17756), .B(new_n17754), .Y(new_n17757));
  nor_5  g15409(.A(new_n17757), .B(new_n17753), .Y(new_n17758));
  nor_5  g15410(.A(new_n17758), .B(new_n17752), .Y(new_n17759));
  xnor_4 g15411(.A(new_n17759), .B(new_n17750), .Y(new_n17760));
  nor_5  g15412(.A(new_n17760), .B(n25972), .Y(new_n17761));
  xnor_4 g15413(.A(new_n17760), .B(new_n11842_1), .Y(new_n17762));
  xnor_4 g15414(.A(new_n17751), .B(n337), .Y(new_n17763));
  xnor_4 g15415(.A(new_n17763), .B(new_n17757), .Y(new_n17764));
  not_8  g15416(.A(new_n17764), .Y(new_n17765));
  nor_5  g15417(.A(new_n17765), .B(n21915), .Y(new_n17766));
  nor_5  g15418(.A(new_n16534), .B(n13775), .Y(new_n17767));
  nor_5  g15419(.A(new_n16550), .B(new_n16535), .Y(new_n17768));
  or_5   g15420(.A(new_n17768), .B(new_n17767), .Y(new_n17769));
  xnor_4 g15421(.A(new_n17765), .B(new_n8646), .Y(new_n17770));
  and_5  g15422(.A(new_n17770), .B(new_n17769), .Y(new_n17771));
  or_5   g15423(.A(new_n17771), .B(new_n17766), .Y(new_n17772));
  and_5  g15424(.A(new_n17772), .B(new_n17762), .Y(new_n17773));
  nor_5  g15425(.A(new_n17773), .B(new_n17761), .Y(new_n17774));
  not_8  g15426(.A(new_n17774), .Y(new_n17775));
  and_5  g15427(.A(new_n17748), .B(new_n7429), .Y(new_n17776));
  and_5  g15428(.A(new_n17749_1), .B(n7593), .Y(new_n17777));
  nor_5  g15429(.A(new_n17749_1), .B(n7593), .Y(new_n17778));
  nor_5  g15430(.A(new_n17759), .B(new_n17778), .Y(new_n17779));
  or_5   g15431(.A(new_n17779), .B(new_n17777), .Y(new_n17780));
  nor_5  g15432(.A(new_n17780), .B(new_n17776), .Y(new_n17781));
  not_8  g15433(.A(new_n17781), .Y(new_n17782));
  nor_5  g15434(.A(new_n17782), .B(new_n17775), .Y(new_n17783));
  xnor_4 g15435(.A(new_n17742), .B(new_n7519), .Y(new_n17784_1));
  xnor_4 g15436(.A(new_n17781), .B(new_n17775), .Y(new_n17785));
  nor_5  g15437(.A(new_n17785), .B(new_n17784_1), .Y(new_n17786));
  xnor_4 g15438(.A(new_n17785), .B(new_n17784_1), .Y(new_n17787));
  xnor_4 g15439(.A(new_n17740), .B(new_n17733), .Y(new_n17788));
  not_8  g15440(.A(new_n17788), .Y(new_n17789));
  xor_4  g15441(.A(new_n17772), .B(new_n17762), .Y(new_n17790));
  nor_5  g15442(.A(new_n17790), .B(new_n17789), .Y(new_n17791));
  xnor_4 g15443(.A(new_n17790), .B(new_n17788), .Y(new_n17792));
  xnor_4 g15444(.A(new_n17738_1), .B(new_n17735_1), .Y(new_n17793));
  xor_4  g15445(.A(new_n17770), .B(new_n17769), .Y(new_n17794));
  nor_5  g15446(.A(new_n17794), .B(new_n17793), .Y(new_n17795));
  nor_5  g15447(.A(new_n16564), .B(new_n16551), .Y(new_n17796));
  nor_5  g15448(.A(new_n16581), .B(new_n16565), .Y(new_n17797));
  or_5   g15449(.A(new_n17797), .B(new_n17796), .Y(new_n17798));
  xnor_4 g15450(.A(new_n17794), .B(new_n17793), .Y(new_n17799));
  nor_5  g15451(.A(new_n17799), .B(new_n17798), .Y(new_n17800));
  or_5   g15452(.A(new_n17800), .B(new_n17795), .Y(new_n17801));
  and_5  g15453(.A(new_n17801), .B(new_n17792), .Y(new_n17802));
  or_5   g15454(.A(new_n17802), .B(new_n17791), .Y(new_n17803));
  nor_5  g15455(.A(new_n17803), .B(new_n17787), .Y(new_n17804));
  nor_5  g15456(.A(new_n17804), .B(new_n17786), .Y(new_n17805));
  xnor_4 g15457(.A(new_n17805), .B(new_n17783), .Y(new_n17806));
  xnor_4 g15458(.A(new_n17806), .B(new_n17745), .Y(n5011));
  nor_5  g15459(.A(new_n10030), .B(n2944), .Y(new_n17808));
  xnor_4 g15460(.A(n11220), .B(n2944), .Y(new_n17809));
  not_8  g15461(.A(n22379), .Y(new_n17810));
  nor_5  g15462(.A(new_n17810), .B(n767), .Y(new_n17811));
  and_5  g15463(.A(new_n2885), .B(new_n2849), .Y(new_n17812));
  or_5   g15464(.A(new_n17812), .B(new_n17811), .Y(new_n17813));
  and_5  g15465(.A(new_n17813), .B(new_n17809), .Y(new_n17814));
  nor_5  g15466(.A(new_n17814), .B(new_n17808), .Y(new_n17815));
  not_8  g15467(.A(new_n17815), .Y(new_n17816));
  nor_5  g15468(.A(new_n8954), .B(new_n12808), .Y(new_n17817));
  or_5   g15469(.A(n16544), .B(n2160), .Y(new_n17818));
  nor_5  g15470(.A(n10763), .B(n6814), .Y(new_n17819));
  and_5  g15471(.A(new_n2924), .B(new_n2888), .Y(new_n17820_1));
  nor_5  g15472(.A(new_n17820_1), .B(new_n17819), .Y(new_n17821));
  and_5  g15473(.A(new_n17821), .B(new_n17818), .Y(new_n17822));
  nor_5  g15474(.A(new_n17822), .B(new_n17817), .Y(new_n17823));
  nor_5  g15475(.A(new_n17823), .B(new_n14810), .Y(new_n17824));
  not_8  g15476(.A(new_n17823), .Y(new_n17825));
  xnor_4 g15477(.A(new_n17825), .B(new_n14811), .Y(new_n17826));
  not_8  g15478(.A(new_n14785), .Y(new_n17827));
  xnor_4 g15479(.A(n16544), .B(new_n12808), .Y(new_n17828));
  xnor_4 g15480(.A(new_n17828), .B(new_n17821), .Y(new_n17829));
  nor_5  g15481(.A(new_n17829), .B(new_n17827), .Y(new_n17830));
  not_8  g15482(.A(new_n17829), .Y(new_n17831));
  xnor_4 g15483(.A(new_n17831), .B(new_n17827), .Y(new_n17832));
  nor_5  g15484(.A(new_n14801_1), .B(new_n2925), .Y(new_n17833));
  and_5  g15485(.A(new_n3031), .B(new_n2970), .Y(new_n17834));
  or_5   g15486(.A(new_n17834), .B(new_n17833), .Y(new_n17835));
  and_5  g15487(.A(new_n17835), .B(new_n17832), .Y(new_n17836));
  nor_5  g15488(.A(new_n17836), .B(new_n17830), .Y(new_n17837));
  nor_5  g15489(.A(new_n17837), .B(new_n17826), .Y(new_n17838));
  nor_5  g15490(.A(new_n17838), .B(new_n17824), .Y(new_n17839));
  nor_5  g15491(.A(new_n17839), .B(new_n17816), .Y(new_n17840));
  xnor_4 g15492(.A(new_n17837), .B(new_n17826), .Y(new_n17841));
  not_8  g15493(.A(new_n17841), .Y(new_n17842));
  nor_5  g15494(.A(new_n17842), .B(new_n17815), .Y(new_n17843));
  nor_5  g15495(.A(new_n17841), .B(new_n17816), .Y(new_n17844));
  xor_4  g15496(.A(new_n17813), .B(new_n17809), .Y(new_n17845));
  xor_4  g15497(.A(new_n17835), .B(new_n17832), .Y(new_n17846));
  nor_5  g15498(.A(new_n17846), .B(new_n17845), .Y(new_n17847));
  xnor_4 g15499(.A(new_n17846), .B(new_n17845), .Y(new_n17848));
  nor_5  g15500(.A(new_n3032), .B(new_n2886_1), .Y(new_n17849));
  nor_5  g15501(.A(new_n3084), .B(new_n3033), .Y(new_n17850));
  nor_5  g15502(.A(new_n17850), .B(new_n17849), .Y(new_n17851));
  nor_5  g15503(.A(new_n17851), .B(new_n17848), .Y(new_n17852));
  nor_5  g15504(.A(new_n17852), .B(new_n17847), .Y(new_n17853));
  nor_5  g15505(.A(new_n17853), .B(new_n17844), .Y(new_n17854));
  nor_5  g15506(.A(new_n17854), .B(new_n17843), .Y(new_n17855_1));
  nor_5  g15507(.A(new_n17855_1), .B(new_n17840), .Y(new_n17856));
  not_8  g15508(.A(new_n17839), .Y(new_n17857));
  nor_5  g15509(.A(new_n17857), .B(new_n17815), .Y(new_n17858));
  nor_5  g15510(.A(new_n17858), .B(new_n17854), .Y(new_n17859));
  nor_5  g15511(.A(new_n17859), .B(new_n17856), .Y(n5020));
  nor_5  g15512(.A(n13781), .B(n11486), .Y(new_n17861));
  not_8  g15513(.A(new_n17861), .Y(new_n17862));
  nor_5  g15514(.A(new_n17862), .B(n16722), .Y(new_n17863));
  not_8  g15515(.A(new_n17863), .Y(new_n17864));
  nor_5  g15516(.A(new_n17864), .B(n3480), .Y(new_n17865));
  xnor_4 g15517(.A(new_n17865), .B(n3018), .Y(new_n17866));
  xnor_4 g15518(.A(new_n17866), .B(new_n2994), .Y(new_n17867));
  xnor_4 g15519(.A(new_n17863), .B(n3480), .Y(new_n17868));
  nor_5  g15520(.A(new_n17868), .B(new_n2998), .Y(new_n17869));
  xnor_4 g15521(.A(new_n17868), .B(new_n2998), .Y(new_n17870));
  xnor_4 g15522(.A(new_n17861), .B(n16722), .Y(new_n17871));
  nor_5  g15523(.A(new_n17871), .B(new_n3003), .Y(new_n17872));
  xnor_4 g15524(.A(new_n17871), .B(new_n3003), .Y(new_n17873));
  xnor_4 g15525(.A(n13781), .B(new_n5784), .Y(new_n17874));
  nor_5  g15526(.A(new_n17874), .B(new_n3011), .Y(new_n17875));
  nor_5  g15527(.A(new_n3015), .B(n13781), .Y(new_n17876));
  not_8  g15528(.A(new_n17876), .Y(new_n17877_1));
  xnor_4 g15529(.A(new_n17874), .B(new_n3011), .Y(new_n17878));
  nor_5  g15530(.A(new_n17878), .B(new_n17877_1), .Y(new_n17879));
  nor_5  g15531(.A(new_n17879), .B(new_n17875), .Y(new_n17880));
  nor_5  g15532(.A(new_n17880), .B(new_n17873), .Y(new_n17881));
  nor_5  g15533(.A(new_n17881), .B(new_n17872), .Y(new_n17882));
  nor_5  g15534(.A(new_n17882), .B(new_n17870), .Y(new_n17883));
  nor_5  g15535(.A(new_n17883), .B(new_n17869), .Y(new_n17884));
  xor_4  g15536(.A(new_n17884), .B(new_n17867), .Y(new_n17885));
  xnor_4 g15537(.A(new_n17885), .B(new_n6926), .Y(new_n17886));
  xor_4  g15538(.A(new_n17882), .B(new_n17870), .Y(new_n17887));
  and_5  g15539(.A(new_n17887), .B(new_n6931), .Y(new_n17888));
  xnor_4 g15540(.A(new_n17887), .B(new_n6931), .Y(new_n17889_1));
  xor_4  g15541(.A(new_n17880), .B(new_n17873), .Y(new_n17890));
  and_5  g15542(.A(new_n17890), .B(new_n6936), .Y(new_n17891));
  xnor_4 g15543(.A(new_n17878), .B(new_n17876), .Y(new_n17892));
  and_5  g15544(.A(new_n17892), .B(new_n6943), .Y(new_n17893));
  xnor_4 g15545(.A(new_n3015), .B(new_n2383), .Y(new_n17894));
  nor_5  g15546(.A(new_n17894), .B(new_n6947), .Y(new_n17895));
  xnor_4 g15547(.A(new_n17892), .B(new_n6943), .Y(new_n17896));
  nor_5  g15548(.A(new_n17896), .B(new_n17895), .Y(new_n17897));
  nor_5  g15549(.A(new_n17897), .B(new_n17893), .Y(new_n17898));
  xnor_4 g15550(.A(new_n17890), .B(new_n6936), .Y(new_n17899));
  nor_5  g15551(.A(new_n17899), .B(new_n17898), .Y(new_n17900));
  nor_5  g15552(.A(new_n17900), .B(new_n17891), .Y(new_n17901));
  nor_5  g15553(.A(new_n17901), .B(new_n17889_1), .Y(new_n17902));
  nor_5  g15554(.A(new_n17902), .B(new_n17888), .Y(new_n17903));
  xnor_4 g15555(.A(new_n17903), .B(new_n17886), .Y(n5024));
  xnor_4 g15556(.A(new_n3715), .B(new_n3684), .Y(n5046));
  xnor_4 g15557(.A(new_n5848), .B(new_n3800), .Y(n5062));
  xnor_4 g15558(.A(new_n12351), .B(new_n12326), .Y(n5064));
  xnor_4 g15559(.A(n12495), .B(new_n11651), .Y(new_n17908));
  not_8  g15560(.A(new_n17908), .Y(new_n17909));
  xnor_4 g15561(.A(new_n17909), .B(new_n2477), .Y(new_n17910));
  xnor_4 g15562(.A(n9251), .B(n7428), .Y(new_n17911_1));
  nor_5  g15563(.A(new_n17911_1), .B(new_n17910), .Y(new_n17912_1));
  nor_5  g15564(.A(new_n2367), .B(n7428), .Y(new_n17913));
  xnor_4 g15565(.A(n20138), .B(n10372), .Y(new_n17914));
  xnor_4 g15566(.A(new_n17914), .B(new_n17913), .Y(new_n17915));
  xnor_4 g15567(.A(new_n17915), .B(new_n17912_1), .Y(new_n17916));
  nor_5  g15568(.A(new_n17908), .B(new_n2477), .Y(new_n17917));
  or_5   g15569(.A(new_n5080), .B(new_n11651), .Y(new_n17918));
  xnor_4 g15570(.A(n20235), .B(new_n6989), .Y(new_n17919));
  xor_4  g15571(.A(new_n17919), .B(new_n17918), .Y(new_n17920));
  xnor_4 g15572(.A(new_n17920), .B(new_n2386), .Y(new_n17921));
  xnor_4 g15573(.A(new_n17921), .B(new_n17917), .Y(new_n17922));
  not_8  g15574(.A(new_n17922), .Y(new_n17923));
  xnor_4 g15575(.A(new_n17923), .B(new_n17916), .Y(n5082));
  xnor_4 g15576(.A(new_n13470), .B(new_n13469), .Y(n5120));
  xnor_4 g15577(.A(new_n14618), .B(new_n14609), .Y(n5158));
  xnor_4 g15578(.A(new_n15913), .B(new_n15901), .Y(n5168));
  not_8  g15579(.A(new_n16936), .Y(new_n17928));
  xnor_4 g15580(.A(new_n17928), .B(n6659), .Y(new_n17929));
  not_8  g15581(.A(new_n14032), .Y(new_n17930));
  nor_5  g15582(.A(new_n17930), .B(n23250), .Y(new_n17931_1));
  xnor_4 g15583(.A(new_n17930), .B(new_n15667), .Y(new_n17932));
  nor_5  g15584(.A(new_n16954_1), .B(n11455), .Y(new_n17933));
  xnor_4 g15585(.A(new_n16954_1), .B(new_n15599), .Y(new_n17934));
  nor_5  g15586(.A(new_n14038), .B(n3945), .Y(new_n17935));
  xnor_4 g15587(.A(new_n14038), .B(new_n15602_1), .Y(new_n17936));
  nor_5  g15588(.A(new_n14043), .B(new_n15605), .Y(new_n17937));
  xnor_4 g15589(.A(new_n14043), .B(n5255), .Y(new_n17938));
  nor_5  g15590(.A(new_n14048), .B(new_n5163), .Y(new_n17939));
  and_5  g15591(.A(new_n15020), .B(new_n15006), .Y(new_n17940));
  or_5   g15592(.A(new_n17940), .B(new_n17939), .Y(new_n17941));
  and_5  g15593(.A(new_n17941), .B(new_n17938), .Y(new_n17942));
  nor_5  g15594(.A(new_n17942), .B(new_n17937), .Y(new_n17943));
  and_5  g15595(.A(new_n17943), .B(new_n17936), .Y(new_n17944));
  or_5   g15596(.A(new_n17944), .B(new_n17935), .Y(new_n17945));
  and_5  g15597(.A(new_n17945), .B(new_n17934), .Y(new_n17946));
  or_5   g15598(.A(new_n17946), .B(new_n17933), .Y(new_n17947));
  and_5  g15599(.A(new_n17947), .B(new_n17932), .Y(new_n17948_1));
  or_5   g15600(.A(new_n17948_1), .B(new_n17931_1), .Y(new_n17949));
  xor_4  g15601(.A(new_n17949), .B(new_n17929), .Y(new_n17950));
  xnor_4 g15602(.A(new_n17950), .B(new_n15597), .Y(new_n17951));
  xor_4  g15603(.A(new_n17947), .B(new_n17932), .Y(new_n17952));
  and_5  g15604(.A(new_n17952), .B(new_n15676), .Y(new_n17953));
  xnor_4 g15605(.A(new_n17952), .B(new_n15676), .Y(new_n17954_1));
  xor_4  g15606(.A(new_n17945), .B(new_n17934), .Y(new_n17955));
  and_5  g15607(.A(new_n17955), .B(new_n15681), .Y(new_n17956_1));
  xnor_4 g15608(.A(new_n17955), .B(new_n15681), .Y(new_n17957));
  xnor_4 g15609(.A(new_n17943), .B(new_n17936), .Y(new_n17958));
  nor_5  g15610(.A(new_n17958), .B(new_n15686), .Y(new_n17959_1));
  xnor_4 g15611(.A(new_n17958), .B(new_n15686), .Y(new_n17960));
  xor_4  g15612(.A(new_n17941), .B(new_n17938), .Y(new_n17961));
  nor_5  g15613(.A(new_n17961), .B(new_n15691), .Y(new_n17962));
  xnor_4 g15614(.A(new_n17961), .B(new_n15691), .Y(new_n17963_1));
  nor_5  g15615(.A(new_n15021), .B(new_n15005), .Y(new_n17964));
  nor_5  g15616(.A(new_n15042), .B(new_n15022), .Y(new_n17965));
  nor_5  g15617(.A(new_n17965), .B(new_n17964), .Y(new_n17966));
  nor_5  g15618(.A(new_n17966), .B(new_n17963_1), .Y(new_n17967));
  nor_5  g15619(.A(new_n17967), .B(new_n17962), .Y(new_n17968_1));
  nor_5  g15620(.A(new_n17968_1), .B(new_n17960), .Y(new_n17969));
  nor_5  g15621(.A(new_n17969), .B(new_n17959_1), .Y(new_n17970));
  nor_5  g15622(.A(new_n17970), .B(new_n17957), .Y(new_n17971));
  nor_5  g15623(.A(new_n17971), .B(new_n17956_1), .Y(new_n17972));
  nor_5  g15624(.A(new_n17972), .B(new_n17954_1), .Y(new_n17973));
  nor_5  g15625(.A(new_n17973), .B(new_n17953), .Y(new_n17974));
  xnor_4 g15626(.A(new_n17974), .B(new_n17951), .Y(n5184));
  and_5  g15627(.A(new_n4533), .B(new_n4417), .Y(new_n17976_1));
  and_5  g15628(.A(new_n4611), .B(new_n17976_1), .Y(new_n17977));
  or_5   g15629(.A(new_n4533), .B(new_n4417), .Y(new_n17978));
  nor_5  g15630(.A(new_n4611), .B(new_n17978), .Y(new_n17979));
  or_5   g15631(.A(new_n17979), .B(new_n17977), .Y(n5228));
  not_8  g15632(.A(n1314), .Y(new_n17981));
  nor_5  g15633(.A(n25494), .B(new_n17981), .Y(new_n17982));
  and_5  g15634(.A(new_n11185), .B(new_n11170), .Y(new_n17983));
  nor_5  g15635(.A(new_n17983), .B(new_n17982), .Y(new_n17984));
  xnor_4 g15636(.A(new_n17984), .B(new_n7195), .Y(new_n17985));
  nor_5  g15637(.A(new_n11186), .B(new_n7118), .Y(new_n17986));
  xnor_4 g15638(.A(new_n11186), .B(new_n7118), .Y(new_n17987));
  nor_5  g15639(.A(new_n11205), .B(new_n7122), .Y(new_n17988));
  nor_5  g15640(.A(new_n12353), .B(new_n12324_1), .Y(new_n17989));
  nor_5  g15641(.A(new_n17989), .B(new_n17988), .Y(new_n17990));
  nor_5  g15642(.A(new_n17990), .B(new_n17987), .Y(new_n17991));
  nor_5  g15643(.A(new_n17991), .B(new_n17986), .Y(new_n17992));
  xnor_4 g15644(.A(new_n17992), .B(new_n17985), .Y(n5256));
  xor_4  g15645(.A(new_n6671_1), .B(new_n6658), .Y(n5265));
  xnor_4 g15646(.A(new_n16728), .B(new_n16683), .Y(n5273));
  xnor_4 g15647(.A(n20946), .B(n2289), .Y(new_n17996));
  nor_5  g15648(.A(new_n5275), .B(n1112), .Y(new_n17997));
  xnor_4 g15649(.A(n7751), .B(n1112), .Y(new_n17998_1));
  nor_5  g15650(.A(new_n12889), .B(n20179), .Y(new_n17999));
  and_5  g15651(.A(new_n16392), .B(new_n16377), .Y(new_n18000));
  or_5   g15652(.A(new_n18000), .B(new_n17999), .Y(new_n18001));
  and_5  g15653(.A(new_n18001), .B(new_n17998_1), .Y(new_n18002));
  or_5   g15654(.A(new_n18002), .B(new_n17997), .Y(new_n18003));
  xor_4  g15655(.A(new_n18003), .B(new_n17996), .Y(new_n18004));
  xnor_4 g15656(.A(new_n18004), .B(new_n7373), .Y(new_n18005));
  xor_4  g15657(.A(new_n18001), .B(new_n17998_1), .Y(new_n18006));
  nor_5  g15658(.A(new_n18006), .B(new_n7377_1), .Y(new_n18007));
  xnor_4 g15659(.A(new_n18006), .B(new_n7377_1), .Y(new_n18008));
  nor_5  g15660(.A(new_n16393), .B(new_n7381), .Y(new_n18009));
  nor_5  g15661(.A(new_n16414), .B(new_n16394), .Y(new_n18010));
  nor_5  g15662(.A(new_n18010), .B(new_n18009), .Y(new_n18011));
  nor_5  g15663(.A(new_n18011), .B(new_n18008), .Y(new_n18012));
  nor_5  g15664(.A(new_n18012), .B(new_n18007), .Y(new_n18013));
  xnor_4 g15665(.A(new_n18013), .B(new_n18005), .Y(n5274));
  nor_5  g15666(.A(n25316), .B(n20385), .Y(new_n18015));
  not_8  g15667(.A(new_n18015), .Y(new_n18016));
  nor_5  g15668(.A(new_n18016), .B(n919), .Y(new_n18017));
  not_8  g15669(.A(new_n18017), .Y(new_n18018));
  nor_5  g15670(.A(new_n18018), .B(n3918), .Y(new_n18019));
  xnor_4 g15671(.A(new_n18019), .B(n6513), .Y(new_n18020));
  xnor_4 g15672(.A(new_n18020), .B(new_n8814), .Y(new_n18021));
  xnor_4 g15673(.A(new_n18017), .B(n3918), .Y(new_n18022));
  nor_5  g15674(.A(new_n18022), .B(new_n8821_1), .Y(new_n18023));
  xnor_4 g15675(.A(new_n18015), .B(n919), .Y(new_n18024));
  nor_5  g15676(.A(new_n18024), .B(new_n11057), .Y(new_n18025_1));
  xnor_4 g15677(.A(new_n18024), .B(new_n8825), .Y(new_n18026));
  xnor_4 g15678(.A(n25316), .B(n20385), .Y(new_n18027));
  nor_5  g15679(.A(new_n18027), .B(new_n8830), .Y(new_n18028));
  nor_5  g15680(.A(new_n8832), .B(new_n4146_1), .Y(new_n18029));
  xnor_4 g15681(.A(new_n18027), .B(new_n8835), .Y(new_n18030));
  and_5  g15682(.A(new_n18030), .B(new_n18029), .Y(new_n18031));
  nor_5  g15683(.A(new_n18031), .B(new_n18028), .Y(new_n18032));
  and_5  g15684(.A(new_n18032), .B(new_n18026), .Y(new_n18033));
  nor_5  g15685(.A(new_n18033), .B(new_n18025_1), .Y(new_n18034));
  xnor_4 g15686(.A(new_n18022), .B(new_n8821_1), .Y(new_n18035_1));
  nor_5  g15687(.A(new_n18035_1), .B(new_n18034), .Y(new_n18036));
  or_5   g15688(.A(new_n18036), .B(new_n18023), .Y(new_n18037));
  xor_4  g15689(.A(new_n18037), .B(new_n18021), .Y(new_n18038));
  not_8  g15690(.A(new_n18038), .Y(new_n18039));
  xnor_4 g15691(.A(new_n16166), .B(n19472), .Y(new_n18040));
  nor_5  g15692(.A(new_n16170), .B(new_n6846), .Y(new_n18041));
  xnor_4 g15693(.A(new_n16170), .B(n25370), .Y(new_n18042));
  nor_5  g15694(.A(new_n16173), .B(new_n8605), .Y(new_n18043_1));
  xnor_4 g15695(.A(new_n16173), .B(n24786), .Y(new_n18044));
  and_5  g15696(.A(new_n4132), .B(n27120), .Y(new_n18045_1));
  or_5   g15697(.A(new_n4136), .B(n23065), .Y(new_n18046));
  xnor_4 g15698(.A(new_n4132), .B(new_n8628), .Y(new_n18047));
  and_5  g15699(.A(new_n18047), .B(new_n18046), .Y(new_n18048));
  or_5   g15700(.A(new_n18048), .B(new_n18045_1), .Y(new_n18049));
  and_5  g15701(.A(new_n18049), .B(new_n18044), .Y(new_n18050));
  or_5   g15702(.A(new_n18050), .B(new_n18043_1), .Y(new_n18051));
  and_5  g15703(.A(new_n18051), .B(new_n18042), .Y(new_n18052));
  or_5   g15704(.A(new_n18052), .B(new_n18041), .Y(new_n18053));
  xor_4  g15705(.A(new_n18053), .B(new_n18040), .Y(new_n18054));
  xnor_4 g15706(.A(new_n18054), .B(new_n18039), .Y(new_n18055));
  xor_4  g15707(.A(new_n18051), .B(new_n18042), .Y(new_n18056));
  xnor_4 g15708(.A(new_n18035_1), .B(new_n18034), .Y(new_n18057));
  nor_5  g15709(.A(new_n18057), .B(new_n18056), .Y(new_n18058));
  xnor_4 g15710(.A(new_n18057), .B(new_n18056), .Y(new_n18059_1));
  xor_4  g15711(.A(new_n18049), .B(new_n18044), .Y(new_n18060));
  xnor_4 g15712(.A(new_n18032), .B(new_n18026), .Y(new_n18061_1));
  nor_5  g15713(.A(new_n18061_1), .B(new_n18060), .Y(new_n18062));
  xnor_4 g15714(.A(new_n18061_1), .B(new_n18060), .Y(new_n18063));
  xnor_4 g15715(.A(new_n18030), .B(new_n18029), .Y(new_n18064));
  not_8  g15716(.A(new_n18064), .Y(new_n18065));
  xor_4  g15717(.A(new_n18047), .B(new_n18046), .Y(new_n18066));
  nor_5  g15718(.A(new_n18066), .B(new_n18065), .Y(new_n18067));
  not_8  g15719(.A(new_n8911_1), .Y(new_n18068));
  xnor_4 g15720(.A(new_n4136), .B(new_n4109), .Y(new_n18069));
  nor_5  g15721(.A(new_n18069), .B(new_n18068), .Y(new_n18070));
  xnor_4 g15722(.A(new_n18066), .B(new_n18065), .Y(new_n18071_1));
  nor_5  g15723(.A(new_n18071_1), .B(new_n18070), .Y(new_n18072));
  nor_5  g15724(.A(new_n18072), .B(new_n18067), .Y(new_n18073));
  nor_5  g15725(.A(new_n18073), .B(new_n18063), .Y(new_n18074));
  nor_5  g15726(.A(new_n18074), .B(new_n18062), .Y(new_n18075));
  nor_5  g15727(.A(new_n18075), .B(new_n18059_1), .Y(new_n18076));
  nor_5  g15728(.A(new_n18076), .B(new_n18058), .Y(new_n18077));
  xnor_4 g15729(.A(new_n18077), .B(new_n18055), .Y(n5300));
  and_5  g15730(.A(new_n12918), .B(new_n7185), .Y(new_n18079));
  and_5  g15731(.A(new_n7193), .B(new_n7190_1), .Y(new_n18080));
  nor_5  g15732(.A(new_n18080), .B(new_n18079), .Y(new_n18081));
  nor_5  g15733(.A(new_n18081), .B(new_n17984), .Y(new_n18082));
  not_8  g15734(.A(new_n18081), .Y(new_n18083));
  xnor_4 g15735(.A(new_n18083), .B(new_n17984), .Y(new_n18084));
  nor_5  g15736(.A(new_n17984), .B(new_n7195), .Y(new_n18085));
  nor_5  g15737(.A(new_n17992), .B(new_n17985), .Y(new_n18086));
  nor_5  g15738(.A(new_n18086), .B(new_n18085), .Y(new_n18087));
  and_5  g15739(.A(new_n18087), .B(new_n18084), .Y(new_n18088));
  nor_5  g15740(.A(new_n18088), .B(new_n18082), .Y(n5325));
  xnor_4 g15741(.A(n25120), .B(n17458), .Y(new_n18090));
  nor_5  g15742(.A(n8363), .B(n1222), .Y(new_n18091));
  xnor_4 g15743(.A(n8363), .B(n1222), .Y(new_n18092));
  nor_5  g15744(.A(n25240), .B(n14680), .Y(new_n18093));
  xnor_4 g15745(.A(n25240), .B(n14680), .Y(new_n18094));
  nor_5  g15746(.A(n17250), .B(n10125), .Y(new_n18095));
  xnor_4 g15747(.A(n17250), .B(new_n10414), .Y(new_n18096));
  nor_5  g15748(.A(new_n10506), .B(new_n10881), .Y(new_n18097));
  or_5   g15749(.A(n23160), .B(n8067), .Y(new_n18098));
  nor_5  g15750(.A(n20923), .B(n16524), .Y(new_n18099));
  nor_5  g15751(.A(new_n12763), .B(new_n12760), .Y(new_n18100));
  nor_5  g15752(.A(new_n18100), .B(new_n18099), .Y(new_n18101));
  and_5  g15753(.A(new_n18101), .B(new_n18098), .Y(new_n18102));
  nor_5  g15754(.A(new_n18102), .B(new_n18097), .Y(new_n18103));
  and_5  g15755(.A(new_n18103), .B(new_n18096), .Y(new_n18104));
  nor_5  g15756(.A(new_n18104), .B(new_n18095), .Y(new_n18105_1));
  nor_5  g15757(.A(new_n18105_1), .B(new_n18094), .Y(new_n18106));
  nor_5  g15758(.A(new_n18106), .B(new_n18093), .Y(new_n18107));
  nor_5  g15759(.A(new_n18107), .B(new_n18092), .Y(new_n18108));
  nor_5  g15760(.A(new_n18108), .B(new_n18091), .Y(new_n18109));
  xnor_4 g15761(.A(new_n18109), .B(new_n18090), .Y(new_n18110));
  nor_5  g15762(.A(new_n18110), .B(n23272), .Y(new_n18111));
  xnor_4 g15763(.A(new_n18110), .B(n23272), .Y(new_n18112));
  xnor_4 g15764(.A(new_n18107), .B(new_n18092), .Y(new_n18113));
  nor_5  g15765(.A(new_n18113), .B(n11481), .Y(new_n18114));
  xnor_4 g15766(.A(new_n18113), .B(n11481), .Y(new_n18115));
  xnor_4 g15767(.A(new_n18105_1), .B(new_n18094), .Y(new_n18116));
  nor_5  g15768(.A(new_n18116), .B(n16439), .Y(new_n18117));
  xnor_4 g15769(.A(new_n18116), .B(n16439), .Y(new_n18118));
  xnor_4 g15770(.A(new_n18103), .B(new_n18096), .Y(new_n18119));
  nor_5  g15771(.A(new_n18119), .B(n15241), .Y(new_n18120));
  xnor_4 g15772(.A(new_n18119), .B(n15241), .Y(new_n18121));
  xnor_4 g15773(.A(n23160), .B(n8067), .Y(new_n18122));
  xnor_4 g15774(.A(new_n18122), .B(new_n18101), .Y(new_n18123));
  nor_5  g15775(.A(new_n18123), .B(n7678), .Y(new_n18124));
  xnor_4 g15776(.A(new_n18123), .B(new_n4373), .Y(new_n18125));
  nor_5  g15777(.A(new_n12764), .B(n3785), .Y(new_n18126));
  nor_5  g15778(.A(new_n12768), .B(new_n12765), .Y(new_n18127));
  or_5   g15779(.A(new_n18127), .B(new_n18126), .Y(new_n18128));
  and_5  g15780(.A(new_n18128), .B(new_n18125), .Y(new_n18129));
  nor_5  g15781(.A(new_n18129), .B(new_n18124), .Y(new_n18130));
  nor_5  g15782(.A(new_n18130), .B(new_n18121), .Y(new_n18131));
  nor_5  g15783(.A(new_n18131), .B(new_n18120), .Y(new_n18132));
  nor_5  g15784(.A(new_n18132), .B(new_n18118), .Y(new_n18133));
  nor_5  g15785(.A(new_n18133), .B(new_n18117), .Y(new_n18134));
  nor_5  g15786(.A(new_n18134), .B(new_n18115), .Y(new_n18135));
  nor_5  g15787(.A(new_n18135), .B(new_n18114), .Y(new_n18136));
  nor_5  g15788(.A(new_n18136), .B(new_n18112), .Y(new_n18137));
  or_5   g15789(.A(new_n18137), .B(new_n18111), .Y(new_n18138));
  nor_5  g15790(.A(n25120), .B(n17458), .Y(new_n18139));
  nor_5  g15791(.A(new_n18109), .B(new_n18090), .Y(new_n18140));
  nor_5  g15792(.A(new_n18140), .B(new_n18139), .Y(new_n18141));
  not_8  g15793(.A(new_n18141), .Y(new_n18142));
  nor_5  g15794(.A(new_n18142), .B(new_n18138), .Y(new_n18143_1));
  not_8  g15795(.A(new_n18143_1), .Y(new_n18144));
  xnor_4 g15796(.A(n12702), .B(n12507), .Y(new_n18145_1));
  nor_5  g15797(.A(n26797), .B(n15077), .Y(new_n18146));
  xnor_4 g15798(.A(n26797), .B(n15077), .Y(new_n18147));
  nor_5  g15799(.A(n23913), .B(n3710), .Y(new_n18148));
  xnor_4 g15800(.A(n23913), .B(n3710), .Y(new_n18149));
  nor_5  g15801(.A(n26318), .B(n22554), .Y(new_n18150));
  xnor_4 g15802(.A(n26318), .B(n22554), .Y(new_n18151_1));
  nor_5  g15803(.A(n26054), .B(n20429), .Y(new_n18152_1));
  xnor_4 g15804(.A(n26054), .B(n20429), .Y(new_n18153));
  nor_5  g15805(.A(n19081), .B(n3909), .Y(new_n18154));
  xnor_4 g15806(.A(n19081), .B(n3909), .Y(new_n18155));
  nor_5  g15807(.A(n23974), .B(n8309), .Y(new_n18156));
  xnor_4 g15808(.A(n23974), .B(new_n8771), .Y(new_n18157_1));
  nor_5  g15809(.A(new_n8759), .B(new_n8050), .Y(new_n18158));
  or_5   g15810(.A(n19144), .B(n2146), .Y(new_n18159));
  nor_5  g15811(.A(n22173), .B(n12593), .Y(new_n18160));
  nor_5  g15812(.A(new_n16371), .B(new_n16370), .Y(new_n18161));
  nor_5  g15813(.A(new_n18161), .B(new_n18160), .Y(new_n18162));
  and_5  g15814(.A(new_n18162), .B(new_n18159), .Y(new_n18163));
  nor_5  g15815(.A(new_n18163), .B(new_n18158), .Y(new_n18164));
  and_5  g15816(.A(new_n18164), .B(new_n18157_1), .Y(new_n18165));
  nor_5  g15817(.A(new_n18165), .B(new_n18156), .Y(new_n18166));
  nor_5  g15818(.A(new_n18166), .B(new_n18155), .Y(new_n18167));
  nor_5  g15819(.A(new_n18167), .B(new_n18154), .Y(new_n18168));
  nor_5  g15820(.A(new_n18168), .B(new_n18153), .Y(new_n18169));
  nor_5  g15821(.A(new_n18169), .B(new_n18152_1), .Y(new_n18170));
  nor_5  g15822(.A(new_n18170), .B(new_n18151_1), .Y(new_n18171_1));
  nor_5  g15823(.A(new_n18171_1), .B(new_n18150), .Y(new_n18172));
  nor_5  g15824(.A(new_n18172), .B(new_n18149), .Y(new_n18173));
  nor_5  g15825(.A(new_n18173), .B(new_n18148), .Y(new_n18174));
  nor_5  g15826(.A(new_n18174), .B(new_n18147), .Y(new_n18175));
  nor_5  g15827(.A(new_n18175), .B(new_n18146), .Y(new_n18176));
  xnor_4 g15828(.A(new_n18176), .B(new_n18145_1), .Y(new_n18177));
  nor_5  g15829(.A(new_n18177), .B(n12650), .Y(new_n18178));
  xnor_4 g15830(.A(new_n18177), .B(n12650), .Y(new_n18179));
  xnor_4 g15831(.A(new_n18174), .B(new_n18147), .Y(new_n18180));
  nor_5  g15832(.A(new_n18180), .B(n10201), .Y(new_n18181));
  xnor_4 g15833(.A(new_n18180), .B(n10201), .Y(new_n18182));
  xnor_4 g15834(.A(new_n18172), .B(new_n18149), .Y(new_n18183));
  nor_5  g15835(.A(new_n18183), .B(n10593), .Y(new_n18184));
  xnor_4 g15836(.A(new_n18183), .B(n10593), .Y(new_n18185));
  xnor_4 g15837(.A(new_n18170), .B(new_n18151_1), .Y(new_n18186));
  nor_5  g15838(.A(new_n18186), .B(n18290), .Y(new_n18187));
  xnor_4 g15839(.A(new_n18168), .B(new_n18153), .Y(new_n18188));
  nor_5  g15840(.A(new_n18188), .B(n11580), .Y(new_n18189));
  xnor_4 g15841(.A(new_n18188), .B(n11580), .Y(new_n18190));
  xnor_4 g15842(.A(new_n18166), .B(new_n18155), .Y(new_n18191));
  nor_5  g15843(.A(new_n18191), .B(n15884), .Y(new_n18192));
  xnor_4 g15844(.A(new_n18191), .B(n15884), .Y(new_n18193_1));
  xnor_4 g15845(.A(new_n18164), .B(new_n18157_1), .Y(new_n18194));
  nor_5  g15846(.A(new_n18194), .B(n6356), .Y(new_n18195));
  xnor_4 g15847(.A(n19144), .B(new_n8050), .Y(new_n18196));
  xnor_4 g15848(.A(new_n18196), .B(new_n18162), .Y(new_n18197));
  nor_5  g15849(.A(new_n18197), .B(new_n5582), .Y(new_n18198));
  xnor_4 g15850(.A(new_n18197), .B(n27104), .Y(new_n18199));
  nor_5  g15851(.A(new_n16372), .B(n27188), .Y(new_n18200));
  and_5  g15852(.A(new_n16373), .B(new_n16369), .Y(new_n18201));
  nor_5  g15853(.A(new_n18201), .B(new_n18200), .Y(new_n18202));
  and_5  g15854(.A(new_n18202), .B(new_n18199), .Y(new_n18203));
  nor_5  g15855(.A(new_n18203), .B(new_n18198), .Y(new_n18204));
  xnor_4 g15856(.A(new_n18194), .B(new_n5595), .Y(new_n18205));
  and_5  g15857(.A(new_n18205), .B(new_n18204), .Y(new_n18206));
  nor_5  g15858(.A(new_n18206), .B(new_n18195), .Y(new_n18207));
  nor_5  g15859(.A(new_n18207), .B(new_n18193_1), .Y(new_n18208));
  nor_5  g15860(.A(new_n18208), .B(new_n18192), .Y(new_n18209));
  nor_5  g15861(.A(new_n18209), .B(new_n18190), .Y(new_n18210));
  nor_5  g15862(.A(new_n18210), .B(new_n18189), .Y(new_n18211));
  xnor_4 g15863(.A(new_n18186), .B(n18290), .Y(new_n18212));
  nor_5  g15864(.A(new_n18212), .B(new_n18211), .Y(new_n18213));
  nor_5  g15865(.A(new_n18213), .B(new_n18187), .Y(new_n18214));
  nor_5  g15866(.A(new_n18214), .B(new_n18185), .Y(new_n18215));
  nor_5  g15867(.A(new_n18215), .B(new_n18184), .Y(new_n18216));
  nor_5  g15868(.A(new_n18216), .B(new_n18182), .Y(new_n18217));
  nor_5  g15869(.A(new_n18217), .B(new_n18181), .Y(new_n18218));
  nor_5  g15870(.A(new_n18218), .B(new_n18179), .Y(new_n18219));
  nor_5  g15871(.A(new_n18219), .B(new_n18178), .Y(new_n18220));
  nor_5  g15872(.A(n12702), .B(n12507), .Y(new_n18221));
  nor_5  g15873(.A(new_n18176), .B(new_n18145_1), .Y(new_n18222));
  nor_5  g15874(.A(new_n18222), .B(new_n18221), .Y(new_n18223));
  and_5  g15875(.A(new_n18223), .B(new_n18220), .Y(new_n18224));
  xnor_4 g15876(.A(new_n18224), .B(new_n18144), .Y(new_n18225));
  xnor_4 g15877(.A(new_n18141), .B(new_n18138), .Y(new_n18226));
  xnor_4 g15878(.A(new_n18223), .B(new_n18220), .Y(new_n18227_1));
  and_5  g15879(.A(new_n18227_1), .B(new_n18226), .Y(new_n18228));
  xnor_4 g15880(.A(new_n18227_1), .B(new_n18226), .Y(new_n18229));
  xnor_4 g15881(.A(new_n18136), .B(new_n18112), .Y(new_n18230));
  not_8  g15882(.A(new_n18230), .Y(new_n18231));
  xnor_4 g15883(.A(new_n18218), .B(new_n18179), .Y(new_n18232_1));
  nor_5  g15884(.A(new_n18232_1), .B(new_n18231), .Y(new_n18233));
  xnor_4 g15885(.A(new_n18232_1), .B(new_n18231), .Y(new_n18234));
  xnor_4 g15886(.A(new_n18134), .B(new_n18115), .Y(new_n18235));
  not_8  g15887(.A(new_n18235), .Y(new_n18236));
  xnor_4 g15888(.A(new_n18216), .B(new_n18182), .Y(new_n18237));
  nor_5  g15889(.A(new_n18237), .B(new_n18236), .Y(new_n18238_1));
  xnor_4 g15890(.A(new_n18237), .B(new_n18236), .Y(new_n18239));
  xnor_4 g15891(.A(new_n18132), .B(new_n18118), .Y(new_n18240));
  not_8  g15892(.A(new_n18240), .Y(new_n18241_1));
  xnor_4 g15893(.A(new_n18214), .B(new_n18185), .Y(new_n18242));
  nor_5  g15894(.A(new_n18242), .B(new_n18241_1), .Y(new_n18243));
  xnor_4 g15895(.A(new_n18242), .B(new_n18241_1), .Y(new_n18244));
  xnor_4 g15896(.A(new_n18130), .B(new_n18121), .Y(new_n18245));
  not_8  g15897(.A(new_n18245), .Y(new_n18246));
  xnor_4 g15898(.A(new_n18212), .B(new_n18211), .Y(new_n18247));
  nor_5  g15899(.A(new_n18247), .B(new_n18246), .Y(new_n18248));
  xnor_4 g15900(.A(new_n18247), .B(new_n18246), .Y(new_n18249));
  xnor_4 g15901(.A(new_n18209), .B(new_n18190), .Y(new_n18250));
  xor_4  g15902(.A(new_n18128), .B(new_n18125), .Y(new_n18251));
  nor_5  g15903(.A(new_n18251), .B(new_n18250), .Y(new_n18252));
  xnor_4 g15904(.A(new_n18251), .B(new_n18250), .Y(new_n18253));
  xnor_4 g15905(.A(new_n18207), .B(new_n18193_1), .Y(new_n18254_1));
  nor_5  g15906(.A(new_n18254_1), .B(new_n12770), .Y(new_n18255));
  xnor_4 g15907(.A(new_n18254_1), .B(new_n12770), .Y(new_n18256));
  xnor_4 g15908(.A(new_n18205), .B(new_n18204), .Y(new_n18257));
  nor_5  g15909(.A(new_n18257), .B(new_n6652_1), .Y(new_n18258));
  xor_4  g15910(.A(new_n18202), .B(new_n18199), .Y(new_n18259));
  nor_5  g15911(.A(new_n18259), .B(new_n6657), .Y(new_n18260));
  xnor_4 g15912(.A(new_n18259), .B(new_n6657), .Y(new_n18261));
  not_8  g15913(.A(new_n18261), .Y(new_n18262));
  nor_5  g15914(.A(new_n16374), .B(new_n16368), .Y(new_n18263));
  nor_5  g15915(.A(new_n16375), .B(new_n6663), .Y(new_n18264));
  nor_5  g15916(.A(new_n18264), .B(new_n18263), .Y(new_n18265));
  and_5  g15917(.A(new_n18265), .B(new_n18262), .Y(new_n18266));
  nor_5  g15918(.A(new_n18266), .B(new_n18260), .Y(new_n18267));
  xnor_4 g15919(.A(new_n18257), .B(new_n6652_1), .Y(new_n18268));
  nor_5  g15920(.A(new_n18268), .B(new_n18267), .Y(new_n18269));
  nor_5  g15921(.A(new_n18269), .B(new_n18258), .Y(new_n18270));
  nor_5  g15922(.A(new_n18270), .B(new_n18256), .Y(new_n18271));
  nor_5  g15923(.A(new_n18271), .B(new_n18255), .Y(new_n18272));
  nor_5  g15924(.A(new_n18272), .B(new_n18253), .Y(new_n18273));
  nor_5  g15925(.A(new_n18273), .B(new_n18252), .Y(new_n18274_1));
  nor_5  g15926(.A(new_n18274_1), .B(new_n18249), .Y(new_n18275));
  nor_5  g15927(.A(new_n18275), .B(new_n18248), .Y(new_n18276));
  nor_5  g15928(.A(new_n18276), .B(new_n18244), .Y(new_n18277));
  nor_5  g15929(.A(new_n18277), .B(new_n18243), .Y(new_n18278));
  nor_5  g15930(.A(new_n18278), .B(new_n18239), .Y(new_n18279));
  nor_5  g15931(.A(new_n18279), .B(new_n18238_1), .Y(new_n18280));
  nor_5  g15932(.A(new_n18280), .B(new_n18234), .Y(new_n18281));
  nor_5  g15933(.A(new_n18281), .B(new_n18233), .Y(new_n18282));
  nor_5  g15934(.A(new_n18282), .B(new_n18229), .Y(new_n18283));
  nor_5  g15935(.A(new_n18283), .B(new_n18228), .Y(new_n18284));
  xnor_4 g15936(.A(new_n18284), .B(new_n18225), .Y(n5351));
  and_5  g15937(.A(new_n16077), .B(new_n16071), .Y(n5353));
  nor_5  g15938(.A(new_n11670), .B(n2160), .Y(new_n18287));
  nor_5  g15939(.A(new_n11718), .B(new_n11671), .Y(new_n18288_1));
  nor_5  g15940(.A(new_n18288_1), .B(new_n18287), .Y(new_n18289));
  not_8  g15941(.A(new_n18289), .Y(new_n18290_1));
  nor_5  g15942(.A(n9934), .B(n2272), .Y(new_n18291));
  and_5  g15943(.A(new_n11669), .B(new_n11634), .Y(new_n18292));
  nor_5  g15944(.A(new_n18292), .B(new_n18291), .Y(new_n18293));
  nor_5  g15945(.A(new_n18293), .B(new_n18290_1), .Y(new_n18294));
  and_5  g15946(.A(new_n11725), .B(new_n14516), .Y(new_n18295_1));
  or_5   g15947(.A(new_n18295_1), .B(new_n7260), .Y(new_n18296));
  nor_5  g15948(.A(new_n11726), .B(new_n7264), .Y(new_n18297));
  nor_5  g15949(.A(new_n11740), .B(new_n11727), .Y(new_n18298));
  nor_5  g15950(.A(new_n18298), .B(new_n18297), .Y(new_n18299));
  nor_5  g15951(.A(new_n18299), .B(new_n18296), .Y(new_n18300));
  xnor_4 g15952(.A(new_n18300), .B(new_n18294), .Y(new_n18301_1));
  xnor_4 g15953(.A(new_n18293), .B(new_n18289), .Y(new_n18302));
  not_8  g15954(.A(new_n7260), .Y(new_n18303));
  xnor_4 g15955(.A(new_n18295_1), .B(new_n18303), .Y(new_n18304_1));
  xnor_4 g15956(.A(new_n18304_1), .B(new_n18299), .Y(new_n18305));
  not_8  g15957(.A(new_n18305), .Y(new_n18306));
  and_5  g15958(.A(new_n18306), .B(new_n18302), .Y(new_n18307));
  xnor_4 g15959(.A(new_n18306), .B(new_n18302), .Y(new_n18308));
  and_5  g15960(.A(new_n11742), .B(new_n11719), .Y(new_n18309));
  nor_5  g15961(.A(new_n11789), .B(new_n11743), .Y(new_n18310_1));
  nor_5  g15962(.A(new_n18310_1), .B(new_n18309), .Y(new_n18311_1));
  nor_5  g15963(.A(new_n18311_1), .B(new_n18308), .Y(new_n18312));
  nor_5  g15964(.A(new_n18312), .B(new_n18307), .Y(new_n18313));
  xnor_4 g15965(.A(new_n18313), .B(new_n18301_1), .Y(n5399));
  nor_5  g15966(.A(new_n17136), .B(new_n4798), .Y(new_n18315));
  and_5  g15967(.A(new_n17141), .B(new_n17138_1), .Y(new_n18316));
  nor_5  g15968(.A(new_n18316), .B(new_n18315), .Y(new_n18317));
  nor_5  g15969(.A(new_n13879), .B(new_n12443), .Y(new_n18318));
  or_5   g15970(.A(new_n13877), .B(n9934), .Y(new_n18319));
  and_5  g15971(.A(new_n17135), .B(new_n18319), .Y(new_n18320));
  or_5   g15972(.A(new_n18320), .B(new_n13920), .Y(new_n18321));
  nor_5  g15973(.A(new_n18321), .B(new_n18318), .Y(new_n18322));
  not_8  g15974(.A(new_n18322), .Y(new_n18323_1));
  nor_5  g15975(.A(new_n18323_1), .B(new_n18317), .Y(new_n18324));
  xnor_4 g15976(.A(new_n18324), .B(new_n18300), .Y(new_n18325));
  xnor_4 g15977(.A(new_n18322), .B(new_n18317), .Y(new_n18326));
  nor_5  g15978(.A(new_n18326), .B(new_n18305), .Y(new_n18327));
  nor_5  g15979(.A(new_n17142), .B(new_n11741_1), .Y(new_n18328));
  nor_5  g15980(.A(new_n17146), .B(new_n17143), .Y(new_n18329));
  nor_5  g15981(.A(new_n18329), .B(new_n18328), .Y(new_n18330));
  xnor_4 g15982(.A(new_n18326), .B(new_n18305), .Y(new_n18331));
  nor_5  g15983(.A(new_n18331), .B(new_n18330), .Y(new_n18332_1));
  nor_5  g15984(.A(new_n18332_1), .B(new_n18327), .Y(new_n18333));
  xnor_4 g15985(.A(new_n18333), .B(new_n18325), .Y(n5403));
  xnor_4 g15986(.A(new_n15321), .B(new_n15288), .Y(n5430));
  or_5   g15987(.A(new_n14306), .B(new_n14300), .Y(new_n18336));
  and_5  g15988(.A(new_n14295), .B(new_n10348), .Y(new_n18337));
  nor_5  g15989(.A(new_n14295), .B(new_n10348), .Y(new_n18338));
  nor_5  g15990(.A(new_n14307), .B(new_n18338), .Y(new_n18339));
  or_5   g15991(.A(new_n18339), .B(new_n18337), .Y(new_n18340));
  nor_5  g15992(.A(new_n18340), .B(new_n10209), .Y(new_n18341));
  and_5  g15993(.A(new_n18341), .B(new_n18336), .Y(n5439));
  xnor_4 g15994(.A(new_n12093), .B(new_n12076), .Y(n5472));
  xnor_4 g15995(.A(new_n8385), .B(new_n8350), .Y(n5485));
  xnor_4 g15996(.A(new_n17803), .B(new_n17787), .Y(n5524));
  not_8  g15997(.A(new_n16088), .Y(new_n18346));
  nor_5  g15998(.A(new_n18346), .B(new_n5953), .Y(new_n18347));
  not_8  g15999(.A(new_n18347), .Y(new_n18348));
  nor_5  g16000(.A(new_n18348), .B(new_n5947), .Y(new_n18349));
  not_8  g16001(.A(new_n18349), .Y(new_n18350_1));
  nor_5  g16002(.A(new_n18350_1), .B(new_n13213), .Y(new_n18351));
  not_8  g16003(.A(new_n18351), .Y(new_n18352));
  nor_5  g16004(.A(new_n18352), .B(new_n13211), .Y(new_n18353));
  not_8  g16005(.A(new_n18353), .Y(new_n18354));
  nor_5  g16006(.A(new_n18354), .B(new_n15842), .Y(new_n18355));
  not_8  g16007(.A(new_n18355), .Y(new_n18356));
  nor_5  g16008(.A(new_n18356), .B(new_n15838), .Y(new_n18357));
  not_8  g16009(.A(new_n18357), .Y(new_n18358));
  nor_5  g16010(.A(new_n18358), .B(new_n5921), .Y(new_n18359));
  xnor_4 g16011(.A(new_n18359), .B(new_n5915), .Y(new_n18360));
  nor_5  g16012(.A(new_n18360), .B(new_n13511), .Y(new_n18361));
  xnor_4 g16013(.A(new_n18360), .B(new_n13511), .Y(new_n18362_1));
  xnor_4 g16014(.A(new_n18357), .B(new_n5921), .Y(new_n18363));
  nor_5  g16015(.A(new_n18363), .B(new_n13514), .Y(new_n18364));
  xnor_4 g16016(.A(new_n18363), .B(new_n13514), .Y(new_n18365));
  xnor_4 g16017(.A(new_n18355), .B(new_n15838), .Y(new_n18366));
  nor_5  g16018(.A(new_n18366), .B(new_n13518), .Y(new_n18367));
  xnor_4 g16019(.A(new_n18366), .B(new_n13518), .Y(new_n18368));
  xnor_4 g16020(.A(new_n18353), .B(new_n15842), .Y(new_n18369));
  nor_5  g16021(.A(new_n18369), .B(new_n13522), .Y(new_n18370));
  xnor_4 g16022(.A(new_n18369), .B(new_n13522), .Y(new_n18371));
  xnor_4 g16023(.A(new_n18351), .B(new_n13211), .Y(new_n18372));
  nor_5  g16024(.A(new_n18372), .B(new_n13526), .Y(new_n18373));
  xnor_4 g16025(.A(new_n18372), .B(new_n13526), .Y(new_n18374));
  xnor_4 g16026(.A(new_n18349), .B(new_n13213), .Y(new_n18375));
  nor_5  g16027(.A(new_n18375), .B(new_n13531), .Y(new_n18376));
  xnor_4 g16028(.A(new_n18375), .B(new_n13531), .Y(new_n18377_1));
  xnor_4 g16029(.A(new_n18347), .B(new_n5947), .Y(new_n18378));
  nor_5  g16030(.A(new_n17149), .B(new_n12853), .Y(new_n18379));
  nor_5  g16031(.A(new_n17153), .B(new_n17150), .Y(new_n18380));
  nor_5  g16032(.A(new_n18380), .B(new_n18379), .Y(new_n18381));
  nor_5  g16033(.A(new_n18381), .B(new_n18378), .Y(new_n18382));
  xor_4  g16034(.A(new_n18381), .B(new_n18378), .Y(new_n18383));
  and_5  g16035(.A(new_n18383), .B(new_n12851), .Y(new_n18384));
  nor_5  g16036(.A(new_n18384), .B(new_n18382), .Y(new_n18385));
  nor_5  g16037(.A(new_n18385), .B(new_n18377_1), .Y(new_n18386));
  nor_5  g16038(.A(new_n18386), .B(new_n18376), .Y(new_n18387));
  nor_5  g16039(.A(new_n18387), .B(new_n18374), .Y(new_n18388));
  nor_5  g16040(.A(new_n18388), .B(new_n18373), .Y(new_n18389));
  nor_5  g16041(.A(new_n18389), .B(new_n18371), .Y(new_n18390));
  nor_5  g16042(.A(new_n18390), .B(new_n18370), .Y(new_n18391));
  nor_5  g16043(.A(new_n18391), .B(new_n18368), .Y(new_n18392));
  nor_5  g16044(.A(new_n18392), .B(new_n18367), .Y(new_n18393));
  nor_5  g16045(.A(new_n18393), .B(new_n18365), .Y(new_n18394));
  nor_5  g16046(.A(new_n18394), .B(new_n18364), .Y(new_n18395));
  nor_5  g16047(.A(new_n18395), .B(new_n18362_1), .Y(new_n18396));
  nor_5  g16048(.A(new_n18396), .B(new_n18361), .Y(new_n18397));
  and_5  g16049(.A(new_n18359), .B(new_n5914), .Y(new_n18398));
  nor_5  g16050(.A(new_n18398), .B(new_n13194), .Y(new_n18399));
  and_5  g16051(.A(new_n18398), .B(new_n13190_1), .Y(new_n18400));
  nor_5  g16052(.A(new_n18400), .B(new_n18399), .Y(new_n18401));
  xnor_4 g16053(.A(new_n18401), .B(new_n13553), .Y(new_n18402));
  xnor_4 g16054(.A(new_n18402), .B(new_n18397), .Y(new_n18403));
  nor_5  g16055(.A(new_n18403), .B(new_n4796), .Y(new_n18404));
  xnor_4 g16056(.A(new_n18403), .B(new_n4796), .Y(new_n18405_1));
  xnor_4 g16057(.A(new_n18395), .B(new_n18362_1), .Y(new_n18406));
  nor_5  g16058(.A(new_n18406), .B(new_n4968), .Y(new_n18407));
  xnor_4 g16059(.A(new_n18406), .B(new_n4968), .Y(new_n18408));
  xnor_4 g16060(.A(new_n18393), .B(new_n18365), .Y(new_n18409_1));
  nor_5  g16061(.A(new_n18409_1), .B(new_n4972_1), .Y(new_n18410));
  xnor_4 g16062(.A(new_n18409_1), .B(new_n4972_1), .Y(new_n18411));
  xnor_4 g16063(.A(new_n18391), .B(new_n18368), .Y(new_n18412));
  nor_5  g16064(.A(new_n18412), .B(new_n4976), .Y(new_n18413));
  xnor_4 g16065(.A(new_n18412), .B(new_n4976), .Y(new_n18414_1));
  xnor_4 g16066(.A(new_n18389), .B(new_n18371), .Y(new_n18415));
  nor_5  g16067(.A(new_n18415), .B(new_n4980), .Y(new_n18416));
  xnor_4 g16068(.A(new_n18415), .B(new_n4980), .Y(new_n18417));
  xnor_4 g16069(.A(new_n18387), .B(new_n18374), .Y(new_n18418_1));
  nor_5  g16070(.A(new_n18418_1), .B(new_n4984), .Y(new_n18419));
  xnor_4 g16071(.A(new_n18418_1), .B(new_n4984), .Y(new_n18420));
  xnor_4 g16072(.A(new_n18385), .B(new_n18377_1), .Y(new_n18421));
  nor_5  g16073(.A(new_n18421), .B(new_n4988), .Y(new_n18422));
  xnor_4 g16074(.A(new_n18421), .B(new_n4988), .Y(new_n18423));
  xnor_4 g16075(.A(new_n18383), .B(new_n12851), .Y(new_n18424));
  nor_5  g16076(.A(new_n18424), .B(new_n4992), .Y(new_n18425));
  xnor_4 g16077(.A(new_n18424), .B(new_n4992), .Y(new_n18426));
  not_8  g16078(.A(new_n18426), .Y(new_n18427));
  nor_5  g16079(.A(new_n17154), .B(new_n4998), .Y(new_n18428));
  and_5  g16080(.A(new_n17157), .B(new_n17155), .Y(new_n18429));
  nor_5  g16081(.A(new_n18429), .B(new_n18428), .Y(new_n18430));
  and_5  g16082(.A(new_n18430), .B(new_n18427), .Y(new_n18431));
  nor_5  g16083(.A(new_n18431), .B(new_n18425), .Y(new_n18432));
  nor_5  g16084(.A(new_n18432), .B(new_n18423), .Y(new_n18433));
  nor_5  g16085(.A(new_n18433), .B(new_n18422), .Y(new_n18434));
  nor_5  g16086(.A(new_n18434), .B(new_n18420), .Y(new_n18435));
  nor_5  g16087(.A(new_n18435), .B(new_n18419), .Y(new_n18436));
  nor_5  g16088(.A(new_n18436), .B(new_n18417), .Y(new_n18437_1));
  nor_5  g16089(.A(new_n18437_1), .B(new_n18416), .Y(new_n18438));
  nor_5  g16090(.A(new_n18438), .B(new_n18414_1), .Y(new_n18439_1));
  nor_5  g16091(.A(new_n18439_1), .B(new_n18413), .Y(new_n18440));
  nor_5  g16092(.A(new_n18440), .B(new_n18411), .Y(new_n18441));
  nor_5  g16093(.A(new_n18441), .B(new_n18410), .Y(new_n18442));
  nor_5  g16094(.A(new_n18442), .B(new_n18408), .Y(new_n18443));
  nor_5  g16095(.A(new_n18443), .B(new_n18407), .Y(new_n18444_1));
  nor_5  g16096(.A(new_n18444_1), .B(new_n18405_1), .Y(new_n18445_1));
  or_5   g16097(.A(new_n18445_1), .B(new_n18404), .Y(new_n18446));
  nor_5  g16098(.A(new_n18401), .B(new_n13553), .Y(new_n18447));
  and_5  g16099(.A(new_n18401), .B(new_n13553), .Y(new_n18448));
  nor_5  g16100(.A(new_n18448), .B(new_n18397), .Y(new_n18449));
  nor_5  g16101(.A(new_n18449), .B(new_n18447), .Y(new_n18450));
  nor_5  g16102(.A(new_n18450), .B(new_n18400), .Y(new_n18451));
  xnor_4 g16103(.A(new_n18451), .B(new_n18446), .Y(n5564));
  xnor_4 g16104(.A(new_n6952), .B(new_n6939), .Y(n5593));
  xnor_4 g16105(.A(new_n17193), .B(new_n13941), .Y(new_n18454));
  nor_5  g16106(.A(new_n15987), .B(new_n13946), .Y(new_n18455));
  xnor_4 g16107(.A(new_n15987), .B(new_n13946), .Y(new_n18456));
  nor_5  g16108(.A(new_n15992), .B(new_n13950), .Y(new_n18457));
  xnor_4 g16109(.A(new_n15992), .B(new_n13950), .Y(new_n18458));
  nor_5  g16110(.A(new_n15059), .B(new_n13954), .Y(new_n18459));
  xnor_4 g16111(.A(new_n15059), .B(new_n13954), .Y(new_n18460));
  nor_5  g16112(.A(new_n15063), .B(new_n13958), .Y(new_n18461));
  and_5  g16113(.A(new_n16767), .B(new_n16758), .Y(new_n18462));
  nor_5  g16114(.A(new_n18462), .B(new_n18461), .Y(new_n18463));
  nor_5  g16115(.A(new_n18463), .B(new_n18460), .Y(new_n18464));
  nor_5  g16116(.A(new_n18464), .B(new_n18459), .Y(new_n18465));
  nor_5  g16117(.A(new_n18465), .B(new_n18458), .Y(new_n18466));
  nor_5  g16118(.A(new_n18466), .B(new_n18457), .Y(new_n18467_1));
  nor_5  g16119(.A(new_n18467_1), .B(new_n18456), .Y(new_n18468));
  nor_5  g16120(.A(new_n18468), .B(new_n18455), .Y(new_n18469));
  xnor_4 g16121(.A(new_n18469), .B(new_n18454), .Y(n5603));
  xnor_4 g16122(.A(n17911), .B(n14440), .Y(new_n18471));
  not_8  g16123(.A(n21997), .Y(new_n18472));
  nor_5  g16124(.A(new_n18472), .B(n1654), .Y(new_n18473));
  xnor_4 g16125(.A(n21997), .B(n1654), .Y(new_n18474));
  nor_5  g16126(.A(new_n8501), .B(n13783), .Y(new_n18475));
  xnor_4 g16127(.A(n25119), .B(n13783), .Y(new_n18476));
  nor_5  g16128(.A(n26660), .B(new_n8503), .Y(new_n18477));
  xnor_4 g16129(.A(n26660), .B(n1163), .Y(new_n18478));
  nor_5  g16130(.A(new_n8506), .B(n3018), .Y(new_n18479));
  or_5   g16131(.A(n18537), .B(new_n10550), .Y(new_n18480));
  nor_5  g16132(.A(n7057), .B(new_n2398), .Y(new_n18481));
  and_5  g16133(.A(new_n17469), .B(new_n17460), .Y(new_n18482_1));
  nor_5  g16134(.A(new_n18482_1), .B(new_n18481), .Y(new_n18483_1));
  and_5  g16135(.A(new_n18483_1), .B(new_n18480), .Y(new_n18484));
  or_5   g16136(.A(new_n18484), .B(new_n18479), .Y(new_n18485));
  and_5  g16137(.A(new_n18485), .B(new_n18478), .Y(new_n18486));
  or_5   g16138(.A(new_n18486), .B(new_n18477), .Y(new_n18487));
  and_5  g16139(.A(new_n18487), .B(new_n18476), .Y(new_n18488));
  or_5   g16140(.A(new_n18488), .B(new_n18475), .Y(new_n18489));
  and_5  g16141(.A(new_n18489), .B(new_n18474), .Y(new_n18490));
  or_5   g16142(.A(new_n18490), .B(new_n18473), .Y(new_n18491));
  xor_4  g16143(.A(new_n18491), .B(new_n18471), .Y(new_n18492));
  xor_4  g16144(.A(new_n18492), .B(new_n3032), .Y(new_n18493));
  xor_4  g16145(.A(new_n18489), .B(new_n18474), .Y(new_n18494));
  nor_5  g16146(.A(new_n18494), .B(new_n3035), .Y(new_n18495));
  xnor_4 g16147(.A(new_n18494), .B(new_n3035), .Y(new_n18496_1));
  xor_4  g16148(.A(new_n18487), .B(new_n18476), .Y(new_n18497));
  nor_5  g16149(.A(new_n18497), .B(new_n3039), .Y(new_n18498));
  xnor_4 g16150(.A(new_n18497), .B(new_n3039), .Y(new_n18499));
  xor_4  g16151(.A(new_n18485), .B(new_n18478), .Y(new_n18500));
  nor_5  g16152(.A(new_n18500), .B(new_n3043), .Y(new_n18501));
  xnor_4 g16153(.A(new_n18500), .B(new_n3043), .Y(new_n18502));
  not_8  g16154(.A(new_n18502), .Y(new_n18503));
  xnor_4 g16155(.A(n18537), .B(n3018), .Y(new_n18504));
  xnor_4 g16156(.A(new_n18504), .B(new_n18483_1), .Y(new_n18505));
  nor_5  g16157(.A(new_n18505), .B(new_n3048), .Y(new_n18506));
  nor_5  g16158(.A(new_n17470), .B(new_n3053), .Y(new_n18507));
  and_5  g16159(.A(new_n17485), .B(new_n17471), .Y(new_n18508));
  or_5   g16160(.A(new_n18508), .B(new_n18507), .Y(new_n18509_1));
  xnor_4 g16161(.A(new_n18505), .B(new_n3049), .Y(new_n18510));
  and_5  g16162(.A(new_n18510), .B(new_n18509_1), .Y(new_n18511));
  nor_5  g16163(.A(new_n18511), .B(new_n18506), .Y(new_n18512));
  and_5  g16164(.A(new_n18512), .B(new_n18503), .Y(new_n18513_1));
  nor_5  g16165(.A(new_n18513_1), .B(new_n18501), .Y(new_n18514));
  nor_5  g16166(.A(new_n18514), .B(new_n18499), .Y(new_n18515_1));
  nor_5  g16167(.A(new_n18515_1), .B(new_n18498), .Y(new_n18516));
  nor_5  g16168(.A(new_n18516), .B(new_n18496_1), .Y(new_n18517));
  nor_5  g16169(.A(new_n18517), .B(new_n18495), .Y(new_n18518));
  xor_4  g16170(.A(new_n18518), .B(new_n18493), .Y(n5609));
  xnor_4 g16171(.A(new_n13137_1), .B(new_n13120), .Y(n5634));
  nor_5  g16172(.A(new_n3217), .B(n2978), .Y(new_n18521));
  xnor_4 g16173(.A(n3425), .B(n2978), .Y(new_n18522));
  nor_5  g16174(.A(n23697), .B(new_n3198), .Y(new_n18523));
  xnor_4 g16175(.A(n23697), .B(n9967), .Y(new_n18524));
  nor_5  g16176(.A(new_n7508), .B(n2289), .Y(new_n18525));
  and_5  g16177(.A(new_n18003), .B(new_n17996), .Y(new_n18526));
  or_5   g16178(.A(new_n18526), .B(new_n18525), .Y(new_n18527));
  and_5  g16179(.A(new_n18527), .B(new_n18524), .Y(new_n18528));
  or_5   g16180(.A(new_n18528), .B(new_n18523), .Y(new_n18529));
  and_5  g16181(.A(new_n18529), .B(new_n18522), .Y(new_n18530));
  nor_5  g16182(.A(new_n18530), .B(new_n18521), .Y(new_n18531));
  nor_5  g16183(.A(new_n18531), .B(new_n7322), .Y(new_n18532));
  not_8  g16184(.A(new_n18531), .Y(new_n18533));
  nor_5  g16185(.A(new_n18533), .B(new_n7323), .Y(new_n18534));
  xor_4  g16186(.A(new_n18529), .B(new_n18522), .Y(new_n18535));
  nor_5  g16187(.A(new_n18535), .B(new_n7365), .Y(new_n18536));
  xnor_4 g16188(.A(new_n18535), .B(new_n7365), .Y(new_n18537_1));
  xor_4  g16189(.A(new_n18527), .B(new_n18524), .Y(new_n18538));
  nor_5  g16190(.A(new_n18538), .B(new_n7369), .Y(new_n18539));
  xnor_4 g16191(.A(new_n18538), .B(new_n7369), .Y(new_n18540));
  nor_5  g16192(.A(new_n18004), .B(new_n7373), .Y(new_n18541));
  nor_5  g16193(.A(new_n18013), .B(new_n18005), .Y(new_n18542));
  nor_5  g16194(.A(new_n18542), .B(new_n18541), .Y(new_n18543));
  nor_5  g16195(.A(new_n18543), .B(new_n18540), .Y(new_n18544));
  nor_5  g16196(.A(new_n18544), .B(new_n18539), .Y(new_n18545));
  nor_5  g16197(.A(new_n18545), .B(new_n18537_1), .Y(new_n18546));
  nor_5  g16198(.A(new_n18546), .B(new_n18536), .Y(new_n18547));
  nor_5  g16199(.A(new_n18547), .B(new_n18534), .Y(new_n18548));
  nor_5  g16200(.A(new_n18548), .B(new_n18532), .Y(new_n18549));
  nor_5  g16201(.A(new_n18303), .B(new_n7242), .Y(new_n18550));
  and_5  g16202(.A(new_n7321), .B(new_n7261), .Y(new_n18551));
  nor_5  g16203(.A(new_n18551), .B(new_n18550), .Y(new_n18552));
  not_8  g16204(.A(new_n18552), .Y(new_n18553));
  xnor_4 g16205(.A(new_n18553), .B(new_n18531), .Y(new_n18554));
  xnor_4 g16206(.A(new_n18554), .B(new_n18549), .Y(n5643));
  xnor_4 g16207(.A(n18035), .B(n5834), .Y(new_n18556));
  nor_5  g16208(.A(n13851), .B(new_n10431), .Y(new_n18557));
  and_5  g16209(.A(new_n15138), .B(new_n15121), .Y(new_n18558_1));
  or_5   g16210(.A(new_n18558_1), .B(new_n18557), .Y(new_n18559));
  xor_4  g16211(.A(new_n18559), .B(new_n18556), .Y(new_n18560));
  xnor_4 g16212(.A(new_n18560), .B(new_n14681), .Y(new_n18561));
  nor_5  g16213(.A(new_n15139_1), .B(new_n14706), .Y(new_n18562));
  xnor_4 g16214(.A(new_n15139_1), .B(new_n14706), .Y(new_n18563));
  nor_5  g16215(.A(new_n15141), .B(new_n14710), .Y(new_n18564));
  xnor_4 g16216(.A(new_n15141), .B(new_n14710), .Y(new_n18565));
  nor_5  g16217(.A(new_n15144), .B(new_n14714), .Y(new_n18566));
  xnor_4 g16218(.A(new_n15144), .B(new_n14714), .Y(new_n18567));
  nor_5  g16219(.A(new_n15149), .B(new_n14717), .Y(new_n18568));
  nor_5  g16220(.A(new_n13608), .B(new_n13370), .Y(new_n18569));
  xnor_4 g16221(.A(new_n13609), .B(new_n13369), .Y(new_n18570));
  and_5  g16222(.A(new_n13622), .B(new_n13374), .Y(new_n18571));
  xnor_4 g16223(.A(new_n13622), .B(new_n13374), .Y(new_n18572_1));
  nor_5  g16224(.A(new_n13629), .B(new_n13376), .Y(new_n18573));
  nor_5  g16225(.A(new_n18573), .B(new_n13381), .Y(new_n18574_1));
  xnor_4 g16226(.A(new_n18573), .B(new_n13380), .Y(new_n18575));
  and_5  g16227(.A(new_n18575), .B(new_n13634), .Y(new_n18576_1));
  nor_5  g16228(.A(new_n18576_1), .B(new_n18574_1), .Y(new_n18577));
  nor_5  g16229(.A(new_n18577), .B(new_n18572_1), .Y(new_n18578_1));
  nor_5  g16230(.A(new_n18578_1), .B(new_n18571), .Y(new_n18579));
  nor_5  g16231(.A(new_n18579), .B(new_n18570), .Y(new_n18580));
  nor_5  g16232(.A(new_n18580), .B(new_n18569), .Y(new_n18581));
  xnor_4 g16233(.A(new_n15147), .B(new_n14718), .Y(new_n18582_1));
  nor_5  g16234(.A(new_n18582_1), .B(new_n18581), .Y(new_n18583_1));
  nor_5  g16235(.A(new_n18583_1), .B(new_n18568), .Y(new_n18584_1));
  nor_5  g16236(.A(new_n18584_1), .B(new_n18567), .Y(new_n18585));
  nor_5  g16237(.A(new_n18585), .B(new_n18566), .Y(new_n18586));
  nor_5  g16238(.A(new_n18586), .B(new_n18565), .Y(new_n18587));
  nor_5  g16239(.A(new_n18587), .B(new_n18564), .Y(new_n18588));
  nor_5  g16240(.A(new_n18588), .B(new_n18563), .Y(new_n18589));
  nor_5  g16241(.A(new_n18589), .B(new_n18562), .Y(new_n18590));
  xor_4  g16242(.A(new_n18590), .B(new_n18561), .Y(n5680));
  xnor_4 g16243(.A(new_n14393), .B(new_n14392), .Y(n5687));
  xnor_4 g16244(.A(new_n15446), .B(new_n15439), .Y(n5700));
  xor_4  g16245(.A(new_n10405_1), .B(new_n10357), .Y(n5732));
  xnor_4 g16246(.A(n23775), .B(n8381), .Y(new_n18595));
  nor_5  g16247(.A(n20235), .B(n8259), .Y(new_n18596));
  and_5  g16248(.A(new_n17919), .B(new_n17918), .Y(new_n18597));
  nor_5  g16249(.A(new_n18597), .B(new_n18596), .Y(new_n18598));
  xnor_4 g16250(.A(new_n18598), .B(new_n18595), .Y(new_n18599));
  xnor_4 g16251(.A(new_n18599), .B(new_n2395), .Y(new_n18600));
  nor_5  g16252(.A(new_n17920), .B(new_n2386), .Y(new_n18601));
  nor_5  g16253(.A(new_n17921), .B(new_n17917), .Y(new_n18602));
  nor_5  g16254(.A(new_n18602), .B(new_n18601), .Y(new_n18603));
  xnor_4 g16255(.A(new_n18603), .B(new_n18600), .Y(new_n18604));
  xnor_4 g16256(.A(n8869), .B(n6385), .Y(new_n18605));
  nor_5  g16257(.A(new_n2363_1), .B(n10372), .Y(new_n18606));
  and_5  g16258(.A(new_n17914), .B(new_n17913), .Y(new_n18607));
  or_5   g16259(.A(new_n18607), .B(new_n18606), .Y(new_n18608));
  xor_4  g16260(.A(new_n18608), .B(new_n18605), .Y(new_n18609));
  xnor_4 g16261(.A(new_n18609), .B(new_n18604), .Y(new_n18610_1));
  and_5  g16262(.A(new_n17915), .B(new_n17912_1), .Y(new_n18611));
  nor_5  g16263(.A(new_n17922), .B(new_n17916), .Y(new_n18612));
  nor_5  g16264(.A(new_n18612), .B(new_n18611), .Y(new_n18613));
  xnor_4 g16265(.A(new_n18613), .B(new_n18610_1), .Y(n5742));
  xnor_4 g16266(.A(new_n13388), .B(new_n13387), .Y(n5765));
  xnor_4 g16267(.A(new_n12304_1), .B(new_n12266), .Y(n5776));
  xnor_4 g16268(.A(new_n2841), .B(new_n2800), .Y(n5782));
  xnor_4 g16269(.A(n18901), .B(new_n8503), .Y(new_n18618));
  nor_5  g16270(.A(n18537), .B(n4376), .Y(new_n18619));
  xnor_4 g16271(.A(n18537), .B(n4376), .Y(new_n18620));
  nor_5  g16272(.A(n14570), .B(n7057), .Y(new_n18621));
  xnor_4 g16273(.A(n14570), .B(n7057), .Y(new_n18622));
  nor_5  g16274(.A(n23775), .B(n8381), .Y(new_n18623));
  nor_5  g16275(.A(new_n18598), .B(new_n18595), .Y(new_n18624));
  nor_5  g16276(.A(new_n18624), .B(new_n18623), .Y(new_n18625));
  nor_5  g16277(.A(new_n18625), .B(new_n18622), .Y(new_n18626));
  nor_5  g16278(.A(new_n18626), .B(new_n18621), .Y(new_n18627));
  nor_5  g16279(.A(new_n18627), .B(new_n18620), .Y(new_n18628));
  or_5   g16280(.A(new_n18628), .B(new_n18619), .Y(new_n18629));
  xor_4  g16281(.A(new_n18629), .B(new_n18618), .Y(new_n18630));
  xor_4  g16282(.A(new_n18630), .B(new_n2423), .Y(new_n18631));
  xnor_4 g16283(.A(new_n18627), .B(new_n18620), .Y(new_n18632));
  nor_5  g16284(.A(new_n18632), .B(new_n2414), .Y(new_n18633));
  xnor_4 g16285(.A(new_n18625), .B(new_n18622), .Y(new_n18634));
  nor_5  g16286(.A(new_n18599), .B(new_n2394), .Y(new_n18635_1));
  and_5  g16287(.A(new_n18603), .B(new_n18600), .Y(new_n18636));
  nor_5  g16288(.A(new_n18636), .B(new_n18635_1), .Y(new_n18637));
  nor_5  g16289(.A(new_n18637), .B(new_n18634), .Y(new_n18638));
  xnor_4 g16290(.A(new_n18637), .B(new_n18634), .Y(new_n18639));
  nor_5  g16291(.A(new_n18639), .B(new_n2404), .Y(new_n18640));
  or_5   g16292(.A(new_n18640), .B(new_n18638), .Y(new_n18641));
  xnor_4 g16293(.A(new_n18632), .B(new_n2415), .Y(new_n18642));
  and_5  g16294(.A(new_n18642), .B(new_n18641), .Y(new_n18643));
  nor_5  g16295(.A(new_n18643), .B(new_n18633), .Y(new_n18644));
  xor_4  g16296(.A(new_n18644), .B(new_n18631), .Y(new_n18645));
  xnor_4 g16297(.A(n23068), .B(n7099), .Y(new_n18646));
  nor_5  g16298(.A(n19514), .B(new_n11685), .Y(new_n18647));
  xnor_4 g16299(.A(n19514), .B(n12811), .Y(new_n18648));
  nor_5  g16300(.A(n10053), .B(new_n11689), .Y(new_n18649_1));
  xnor_4 g16301(.A(n10053), .B(n1118), .Y(new_n18650));
  nor_5  g16302(.A(n25974), .B(new_n2947), .Y(new_n18651));
  nor_5  g16303(.A(new_n11693), .B(n8399), .Y(new_n18652));
  nor_5  g16304(.A(new_n3824), .B(n1630), .Y(new_n18653_1));
  or_5   g16305(.A(n9507), .B(new_n2909), .Y(new_n18654));
  nor_5  g16306(.A(new_n2952), .B(n1451), .Y(new_n18655));
  and_5  g16307(.A(new_n18655), .B(new_n18654), .Y(new_n18656));
  nor_5  g16308(.A(new_n18656), .B(new_n18653_1), .Y(new_n18657));
  nor_5  g16309(.A(new_n18657), .B(new_n18652), .Y(new_n18658));
  nor_5  g16310(.A(new_n18658), .B(new_n18651), .Y(new_n18659));
  and_5  g16311(.A(new_n18659), .B(new_n18650), .Y(new_n18660));
  or_5   g16312(.A(new_n18660), .B(new_n18649_1), .Y(new_n18661));
  and_5  g16313(.A(new_n18661), .B(new_n18648), .Y(new_n18662));
  or_5   g16314(.A(new_n18662), .B(new_n18647), .Y(new_n18663));
  xor_4  g16315(.A(new_n18663), .B(new_n18646), .Y(new_n18664));
  xnor_4 g16316(.A(new_n18664), .B(new_n18645), .Y(new_n18665));
  not_8  g16317(.A(new_n18665), .Y(new_n18666));
  xor_4  g16318(.A(new_n18661), .B(new_n18648), .Y(new_n18667));
  not_8  g16319(.A(new_n18667), .Y(new_n18668));
  nor_5  g16320(.A(new_n18640), .B(new_n18638), .Y(new_n18669));
  xnor_4 g16321(.A(new_n18642), .B(new_n18669), .Y(new_n18670));
  nor_5  g16322(.A(new_n18670), .B(new_n18668), .Y(new_n18671));
  xnor_4 g16323(.A(new_n18639), .B(new_n2405), .Y(new_n18672));
  xnor_4 g16324(.A(new_n18659), .B(new_n18650), .Y(new_n18673));
  and_5  g16325(.A(new_n18673), .B(new_n18672), .Y(new_n18674));
  xnor_4 g16326(.A(new_n18673), .B(new_n18672), .Y(new_n18675));
  not_8  g16327(.A(new_n18604), .Y(new_n18676));
  xnor_4 g16328(.A(n25974), .B(n8399), .Y(new_n18677));
  xnor_4 g16329(.A(new_n18677), .B(new_n18657), .Y(new_n18678));
  and_5  g16330(.A(new_n18678), .B(new_n18676), .Y(new_n18679_1));
  xnor_4 g16331(.A(new_n18678), .B(new_n18676), .Y(new_n18680));
  xnor_4 g16332(.A(n26979), .B(n1451), .Y(new_n18681));
  nor_5  g16333(.A(new_n18681), .B(new_n17910), .Y(new_n18682));
  xnor_4 g16334(.A(n9507), .B(n1630), .Y(new_n18683));
  xnor_4 g16335(.A(new_n18683), .B(new_n18655), .Y(new_n18684));
  nor_5  g16336(.A(new_n18684), .B(new_n18682), .Y(new_n18685));
  xnor_4 g16337(.A(new_n18684), .B(new_n18682), .Y(new_n18686));
  nor_5  g16338(.A(new_n18686), .B(new_n17923), .Y(new_n18687));
  nor_5  g16339(.A(new_n18687), .B(new_n18685), .Y(new_n18688));
  nor_5  g16340(.A(new_n18688), .B(new_n18680), .Y(new_n18689));
  nor_5  g16341(.A(new_n18689), .B(new_n18679_1), .Y(new_n18690_1));
  nor_5  g16342(.A(new_n18690_1), .B(new_n18675), .Y(new_n18691));
  nor_5  g16343(.A(new_n18691), .B(new_n18674), .Y(new_n18692));
  xnor_4 g16344(.A(new_n18670), .B(new_n18667), .Y(new_n18693_1));
  and_5  g16345(.A(new_n18693_1), .B(new_n18692), .Y(new_n18694));
  nor_5  g16346(.A(new_n18694), .B(new_n18671), .Y(new_n18695));
  xnor_4 g16347(.A(new_n18695), .B(new_n18666), .Y(n5833));
  xnor_4 g16348(.A(new_n12300), .B(new_n12274), .Y(n5840));
  xor_4  g16349(.A(new_n18510), .B(new_n18509_1), .Y(n5841));
  xnor_4 g16350(.A(new_n12744), .B(new_n12743), .Y(n5850));
  xnor_4 g16351(.A(new_n18579), .B(new_n18570), .Y(n5903));
  xnor_4 g16352(.A(new_n16163), .B(n19042), .Y(new_n18701));
  nor_5  g16353(.A(new_n16166), .B(new_n8572), .Y(new_n18702));
  and_5  g16354(.A(new_n18053), .B(new_n18040), .Y(new_n18703));
  or_5   g16355(.A(new_n18703), .B(new_n18702), .Y(new_n18704));
  xor_4  g16356(.A(new_n18704), .B(new_n18701), .Y(new_n18705));
  not_8  g16357(.A(new_n18019), .Y(new_n18706));
  nor_5  g16358(.A(new_n18706), .B(n6513), .Y(new_n18707));
  xnor_4 g16359(.A(new_n18707), .B(n26752), .Y(new_n18708_1));
  xnor_4 g16360(.A(new_n18708_1), .B(new_n8807), .Y(new_n18709));
  nor_5  g16361(.A(new_n18020), .B(new_n8813), .Y(new_n18710));
  and_5  g16362(.A(new_n18037), .B(new_n18021), .Y(new_n18711));
  nor_5  g16363(.A(new_n18711), .B(new_n18710), .Y(new_n18712));
  xnor_4 g16364(.A(new_n18712), .B(new_n18709), .Y(new_n18713));
  xnor_4 g16365(.A(new_n18713), .B(new_n18705), .Y(new_n18714));
  nor_5  g16366(.A(new_n18054), .B(new_n18039), .Y(new_n18715));
  nor_5  g16367(.A(new_n18077), .B(new_n18055), .Y(new_n18716));
  nor_5  g16368(.A(new_n18716), .B(new_n18715), .Y(new_n18717));
  xnor_4 g16369(.A(new_n18717), .B(new_n18714), .Y(n5904));
  xnor_4 g16370(.A(n27089), .B(n6814), .Y(new_n18719));
  nor_5  g16371(.A(new_n8959), .B(n11841), .Y(new_n18720));
  xnor_4 g16372(.A(n19701), .B(n11841), .Y(new_n18721_1));
  nor_5  g16373(.A(new_n8962), .B(n10710), .Y(new_n18722));
  xnor_4 g16374(.A(n23529), .B(n10710), .Y(new_n18723));
  nor_5  g16375(.A(new_n8965), .B(n20929), .Y(new_n18724));
  xnor_4 g16376(.A(n24620), .B(n20929), .Y(new_n18725_1));
  nor_5  g16377(.A(n8006), .B(new_n8968), .Y(new_n18726));
  xnor_4 g16378(.A(n8006), .B(n5211), .Y(new_n18727));
  nor_5  g16379(.A(n25074), .B(new_n8971_1), .Y(new_n18728));
  xnor_4 g16380(.A(n25074), .B(n12956), .Y(new_n18729));
  nor_5  g16381(.A(n18295), .B(new_n4328), .Y(new_n18730));
  nor_5  g16382(.A(new_n2903), .B(n16396), .Y(new_n18731));
  nor_5  g16383(.A(new_n4331), .B(n6502), .Y(new_n18732));
  nor_5  g16384(.A(n9399), .B(new_n5033), .Y(new_n18733));
  nor_5  g16385(.A(n15780), .B(new_n2951), .Y(new_n18734));
  not_8  g16386(.A(new_n18734), .Y(new_n18735));
  nor_5  g16387(.A(new_n18735), .B(new_n18733), .Y(new_n18736));
  nor_5  g16388(.A(new_n18736), .B(new_n18732), .Y(new_n18737_1));
  nor_5  g16389(.A(new_n18737_1), .B(new_n18731), .Y(new_n18738));
  nor_5  g16390(.A(new_n18738), .B(new_n18730), .Y(new_n18739));
  and_5  g16391(.A(new_n18739), .B(new_n18729), .Y(new_n18740));
  or_5   g16392(.A(new_n18740), .B(new_n18728), .Y(new_n18741));
  and_5  g16393(.A(new_n18741), .B(new_n18727), .Y(new_n18742));
  or_5   g16394(.A(new_n18742), .B(new_n18726), .Y(new_n18743));
  and_5  g16395(.A(new_n18743), .B(new_n18725_1), .Y(new_n18744));
  or_5   g16396(.A(new_n18744), .B(new_n18724), .Y(new_n18745_1));
  and_5  g16397(.A(new_n18745_1), .B(new_n18723), .Y(new_n18746));
  or_5   g16398(.A(new_n18746), .B(new_n18722), .Y(new_n18747));
  and_5  g16399(.A(new_n18747), .B(new_n18721_1), .Y(new_n18748));
  or_5   g16400(.A(new_n18748), .B(new_n18720), .Y(new_n18749));
  xor_4  g16401(.A(new_n18749), .B(new_n18719), .Y(new_n18750));
  xnor_4 g16402(.A(new_n18750), .B(new_n10106), .Y(new_n18751_1));
  xor_4  g16403(.A(new_n18747), .B(new_n18721_1), .Y(new_n18752));
  nor_5  g16404(.A(new_n18752), .B(new_n10110), .Y(new_n18753));
  xnor_4 g16405(.A(new_n18752), .B(new_n10110), .Y(new_n18754));
  xor_4  g16406(.A(new_n18745_1), .B(new_n18723), .Y(new_n18755));
  nor_5  g16407(.A(new_n18755), .B(new_n10114), .Y(new_n18756));
  xnor_4 g16408(.A(new_n18755), .B(new_n10114), .Y(new_n18757));
  xor_4  g16409(.A(new_n18743), .B(new_n18725_1), .Y(new_n18758));
  nor_5  g16410(.A(new_n18758), .B(new_n10118), .Y(new_n18759));
  xor_4  g16411(.A(new_n18741), .B(new_n18727), .Y(new_n18760));
  nor_5  g16412(.A(new_n18760), .B(new_n10121), .Y(new_n18761));
  xnor_4 g16413(.A(new_n18760), .B(new_n10121), .Y(new_n18762));
  xnor_4 g16414(.A(new_n18739), .B(new_n18729), .Y(new_n18763));
  and_5  g16415(.A(new_n18763), .B(new_n10124), .Y(new_n18764));
  xnor_4 g16416(.A(n18295), .B(n16396), .Y(new_n18765));
  xnor_4 g16417(.A(new_n18765), .B(new_n18737_1), .Y(new_n18766));
  and_5  g16418(.A(new_n18766), .B(new_n10128), .Y(new_n18767));
  xnor_4 g16419(.A(new_n18766), .B(new_n10132), .Y(new_n18768));
  xnor_4 g16420(.A(n15780), .B(n2088), .Y(new_n18769));
  nor_5  g16421(.A(new_n18769), .B(new_n10134), .Y(new_n18770));
  xnor_4 g16422(.A(n9399), .B(n6502), .Y(new_n18771));
  xnor_4 g16423(.A(new_n18771), .B(new_n18735), .Y(new_n18772));
  not_8  g16424(.A(new_n18772), .Y(new_n18773));
  and_5  g16425(.A(new_n18773), .B(new_n18770), .Y(new_n18774));
  xnor_4 g16426(.A(new_n18773), .B(new_n18770), .Y(new_n18775));
  nor_5  g16427(.A(new_n18775), .B(new_n10142), .Y(new_n18776));
  nor_5  g16428(.A(new_n18776), .B(new_n18774), .Y(new_n18777));
  and_5  g16429(.A(new_n18777), .B(new_n18768), .Y(new_n18778));
  nor_5  g16430(.A(new_n18778), .B(new_n18767), .Y(new_n18779));
  xnor_4 g16431(.A(new_n18763), .B(new_n10124), .Y(new_n18780_1));
  nor_5  g16432(.A(new_n18780_1), .B(new_n18779), .Y(new_n18781));
  nor_5  g16433(.A(new_n18781), .B(new_n18764), .Y(new_n18782_1));
  nor_5  g16434(.A(new_n18782_1), .B(new_n18762), .Y(new_n18783));
  nor_5  g16435(.A(new_n18783), .B(new_n18761), .Y(new_n18784));
  xnor_4 g16436(.A(new_n18758), .B(new_n10118), .Y(new_n18785));
  nor_5  g16437(.A(new_n18785), .B(new_n18784), .Y(new_n18786));
  nor_5  g16438(.A(new_n18786), .B(new_n18759), .Y(new_n18787));
  nor_5  g16439(.A(new_n18787), .B(new_n18757), .Y(new_n18788));
  nor_5  g16440(.A(new_n18788), .B(new_n18756), .Y(new_n18789));
  nor_5  g16441(.A(new_n18789), .B(new_n18754), .Y(new_n18790));
  nor_5  g16442(.A(new_n18790), .B(new_n18753), .Y(new_n18791));
  xnor_4 g16443(.A(new_n18791), .B(new_n18751_1), .Y(n5911));
  xnor_4 g16444(.A(new_n11769), .B(new_n3913), .Y(n5936));
  xnor_4 g16445(.A(new_n9976), .B(new_n9936), .Y(n5943));
  xnor_4 g16446(.A(new_n13980), .B(new_n13952), .Y(n5964));
  nor_5  g16447(.A(new_n5070), .B(n11184), .Y(new_n18796));
  nor_5  g16448(.A(new_n5057), .B(n23146), .Y(new_n18797));
  or_5   g16449(.A(new_n5082_1), .B(n17968), .Y(new_n18798));
  nor_5  g16450(.A(new_n18798), .B(new_n5061), .Y(new_n18799));
  nor_5  g16451(.A(new_n18799), .B(new_n18797), .Y(new_n18800));
  nor_5  g16452(.A(new_n18800), .B(new_n5071), .Y(new_n18801));
  nor_5  g16453(.A(new_n18801), .B(new_n18796), .Y(new_n18802_1));
  and_5  g16454(.A(new_n18802_1), .B(new_n15641), .Y(new_n18803));
  nor_5  g16455(.A(new_n18802_1), .B(new_n15648), .Y(new_n18804));
  nor_5  g16456(.A(new_n18804), .B(new_n15640), .Y(new_n18805));
  nor_5  g16457(.A(new_n18805), .B(new_n18803), .Y(new_n18806));
  nor_5  g16458(.A(new_n18806), .B(new_n15636_1), .Y(new_n18807));
  nand_5 g16459(.A(new_n18806), .B(new_n15638), .Y(new_n18808));
  and_5  g16460(.A(new_n18808), .B(n8943), .Y(new_n18809));
  nor_5  g16461(.A(new_n18809), .B(new_n18807), .Y(new_n18810));
  nor_5  g16462(.A(new_n18810), .B(new_n15633), .Y(new_n18811));
  nand_5 g16463(.A(new_n18810), .B(new_n15635), .Y(new_n18812));
  and_5  g16464(.A(new_n18812), .B(n12380), .Y(new_n18813));
  nor_5  g16465(.A(new_n18813), .B(new_n18811), .Y(new_n18814));
  nor_5  g16466(.A(new_n18814), .B(new_n15631), .Y(new_n18815));
  nand_5 g16467(.A(new_n18814), .B(new_n15656), .Y(new_n18816));
  and_5  g16468(.A(new_n18816), .B(n8694), .Y(new_n18817));
  nor_5  g16469(.A(new_n18817), .B(new_n18815), .Y(new_n18818));
  nor_5  g16470(.A(new_n18818), .B(new_n15629), .Y(new_n18819));
  and_5  g16471(.A(new_n18818), .B(new_n15682), .Y(new_n18820));
  nor_5  g16472(.A(new_n18820), .B(new_n15660), .Y(new_n18821));
  or_5   g16473(.A(new_n18821), .B(new_n18819), .Y(new_n18822));
  xor_4  g16474(.A(new_n18822), .B(new_n15628), .Y(new_n18823));
  xnor_4 g16475(.A(new_n18823), .B(new_n3224), .Y(new_n18824));
  xnor_4 g16476(.A(new_n18818), .B(new_n15661), .Y(new_n18825));
  and_5  g16477(.A(new_n18825), .B(new_n3228_1), .Y(new_n18826));
  xnor_4 g16478(.A(new_n18825), .B(new_n3228_1), .Y(new_n18827));
  xnor_4 g16479(.A(new_n18814), .B(new_n15657), .Y(new_n18828));
  and_5  g16480(.A(new_n18828), .B(new_n3233), .Y(new_n18829));
  xnor_4 g16481(.A(new_n18828), .B(new_n3233), .Y(new_n18830_1));
  xor_4  g16482(.A(new_n18810), .B(new_n15635), .Y(new_n18831_1));
  and_5  g16483(.A(new_n18831_1), .B(new_n3238), .Y(new_n18832));
  xnor_4 g16484(.A(new_n18831_1), .B(new_n3238), .Y(new_n18833));
  xnor_4 g16485(.A(new_n18806), .B(new_n15639), .Y(new_n18834));
  and_5  g16486(.A(new_n18834), .B(new_n3243), .Y(new_n18835));
  xnor_4 g16487(.A(new_n18834), .B(new_n3243), .Y(new_n18836));
  xnor_4 g16488(.A(new_n18802_1), .B(new_n15649), .Y(new_n18837));
  and_5  g16489(.A(new_n18837), .B(new_n3248), .Y(new_n18838));
  xnor_4 g16490(.A(new_n18837), .B(new_n3248), .Y(new_n18839));
  xnor_4 g16491(.A(new_n18800), .B(new_n15645), .Y(new_n18840));
  and_5  g16492(.A(new_n18840), .B(new_n3253_1), .Y(new_n18841));
  xnor_4 g16493(.A(new_n18840), .B(new_n3253_1), .Y(new_n18842));
  xnor_4 g16494(.A(new_n18798), .B(new_n5074), .Y(new_n18843_1));
  and_5  g16495(.A(new_n18843_1), .B(new_n3261), .Y(new_n18844));
  nor_5  g16496(.A(new_n5084), .B(new_n3257), .Y(new_n18845));
  xnor_4 g16497(.A(new_n18843_1), .B(new_n3261), .Y(new_n18846));
  nor_5  g16498(.A(new_n18846), .B(new_n18845), .Y(new_n18847));
  nor_5  g16499(.A(new_n18847), .B(new_n18844), .Y(new_n18848));
  nor_5  g16500(.A(new_n18848), .B(new_n18842), .Y(new_n18849));
  nor_5  g16501(.A(new_n18849), .B(new_n18841), .Y(new_n18850));
  nor_5  g16502(.A(new_n18850), .B(new_n18839), .Y(new_n18851));
  nor_5  g16503(.A(new_n18851), .B(new_n18838), .Y(new_n18852));
  nor_5  g16504(.A(new_n18852), .B(new_n18836), .Y(new_n18853));
  nor_5  g16505(.A(new_n18853), .B(new_n18835), .Y(new_n18854));
  nor_5  g16506(.A(new_n18854), .B(new_n18833), .Y(new_n18855));
  nor_5  g16507(.A(new_n18855), .B(new_n18832), .Y(new_n18856));
  nor_5  g16508(.A(new_n18856), .B(new_n18830_1), .Y(new_n18857));
  nor_5  g16509(.A(new_n18857), .B(new_n18829), .Y(new_n18858_1));
  nor_5  g16510(.A(new_n18858_1), .B(new_n18827), .Y(new_n18859_1));
  nor_5  g16511(.A(new_n18859_1), .B(new_n18826), .Y(new_n18860));
  xnor_4 g16512(.A(new_n18860), .B(new_n18824), .Y(n5980));
  xnor_4 g16513(.A(new_n11143), .B(new_n11120_1), .Y(n6012));
  nor_5  g16514(.A(new_n10095), .B(n16544), .Y(new_n18863));
  xnor_4 g16515(.A(new_n10095), .B(n16544), .Y(new_n18864_1));
  nor_5  g16516(.A(new_n10058), .B(n6814), .Y(new_n18865_1));
  xnor_4 g16517(.A(new_n10058), .B(n6814), .Y(new_n18866));
  nor_5  g16518(.A(new_n10063), .B(n19701), .Y(new_n18867));
  xnor_4 g16519(.A(new_n10063), .B(n19701), .Y(new_n18868));
  nor_5  g16520(.A(new_n9249), .B(n23529), .Y(new_n18869));
  and_5  g16521(.A(new_n9286), .B(new_n9250), .Y(new_n18870));
  nor_5  g16522(.A(new_n18870), .B(new_n18869), .Y(new_n18871));
  nor_5  g16523(.A(new_n18871), .B(new_n18868), .Y(new_n18872));
  nor_5  g16524(.A(new_n18872), .B(new_n18867), .Y(new_n18873));
  nor_5  g16525(.A(new_n18873), .B(new_n18866), .Y(new_n18874));
  nor_5  g16526(.A(new_n18874), .B(new_n18865_1), .Y(new_n18875));
  nor_5  g16527(.A(new_n18875), .B(new_n18864_1), .Y(new_n18876));
  nor_5  g16528(.A(new_n18876), .B(new_n18863), .Y(new_n18877));
  and_5  g16529(.A(new_n18877), .B(new_n10044), .Y(new_n18878));
  nor_5  g16530(.A(new_n13823), .B(n3582), .Y(new_n18879));
  xnor_4 g16531(.A(new_n13823), .B(n3582), .Y(new_n18880_1));
  nor_5  g16532(.A(new_n13859), .B(n2145), .Y(new_n18881));
  xnor_4 g16533(.A(new_n13859), .B(n2145), .Y(new_n18882));
  nor_5  g16534(.A(new_n13829), .B(n5031), .Y(new_n18883));
  xnor_4 g16535(.A(new_n13829), .B(n5031), .Y(new_n18884));
  nor_5  g16536(.A(new_n9311), .B(new_n7657_1), .Y(new_n18885));
  nor_5  g16537(.A(new_n9349), .B(new_n9313), .Y(new_n18886_1));
  or_5   g16538(.A(new_n18886_1), .B(new_n18885), .Y(new_n18887_1));
  nor_5  g16539(.A(new_n18887_1), .B(new_n18884), .Y(new_n18888));
  nor_5  g16540(.A(new_n18888), .B(new_n18883), .Y(new_n18889));
  nor_5  g16541(.A(new_n18889), .B(new_n18882), .Y(new_n18890));
  nor_5  g16542(.A(new_n18890), .B(new_n18881), .Y(new_n18891));
  nor_5  g16543(.A(new_n18891), .B(new_n18880_1), .Y(new_n18892));
  nor_5  g16544(.A(new_n18892), .B(new_n18879), .Y(new_n18893));
  not_8  g16545(.A(new_n18893), .Y(new_n18894));
  nor_5  g16546(.A(new_n18894), .B(new_n13869), .Y(new_n18895));
  not_8  g16547(.A(new_n18895), .Y(new_n18896));
  xnor_4 g16548(.A(new_n18896), .B(new_n18878), .Y(new_n18897));
  xnor_4 g16549(.A(new_n18877), .B(new_n10045), .Y(new_n18898));
  xnor_4 g16550(.A(new_n18894), .B(new_n13868), .Y(new_n18899));
  not_8  g16551(.A(new_n18899), .Y(new_n18900));
  nor_5  g16552(.A(new_n18900), .B(new_n18898), .Y(new_n18901_1));
  xnor_4 g16553(.A(new_n18900), .B(new_n18898), .Y(new_n18902));
  xnor_4 g16554(.A(new_n18875), .B(new_n18864_1), .Y(new_n18903));
  xor_4  g16555(.A(new_n18891), .B(new_n18880_1), .Y(new_n18904));
  nor_5  g16556(.A(new_n18904), .B(new_n18903), .Y(new_n18905));
  xnor_4 g16557(.A(new_n18904), .B(new_n18903), .Y(new_n18906));
  xnor_4 g16558(.A(new_n18873), .B(new_n18866), .Y(new_n18907_1));
  xor_4  g16559(.A(new_n18889), .B(new_n18882), .Y(new_n18908));
  nor_5  g16560(.A(new_n18908), .B(new_n18907_1), .Y(new_n18909));
  xnor_4 g16561(.A(new_n18908), .B(new_n18907_1), .Y(new_n18910));
  xnor_4 g16562(.A(new_n18871), .B(new_n18868), .Y(new_n18911));
  xor_4  g16563(.A(new_n18887_1), .B(new_n18884), .Y(new_n18912));
  nor_5  g16564(.A(new_n18912), .B(new_n18911), .Y(new_n18913));
  xnor_4 g16565(.A(new_n18912), .B(new_n18911), .Y(new_n18914));
  and_5  g16566(.A(new_n9351), .B(new_n9287_1), .Y(new_n18915));
  nor_5  g16567(.A(new_n9391), .B(new_n9352), .Y(new_n18916));
  nor_5  g16568(.A(new_n18916), .B(new_n18915), .Y(new_n18917));
  nor_5  g16569(.A(new_n18917), .B(new_n18914), .Y(new_n18918));
  nor_5  g16570(.A(new_n18918), .B(new_n18913), .Y(new_n18919_1));
  nor_5  g16571(.A(new_n18919_1), .B(new_n18910), .Y(new_n18920));
  nor_5  g16572(.A(new_n18920), .B(new_n18909), .Y(new_n18921));
  nor_5  g16573(.A(new_n18921), .B(new_n18906), .Y(new_n18922));
  nor_5  g16574(.A(new_n18922), .B(new_n18905), .Y(new_n18923));
  nor_5  g16575(.A(new_n18923), .B(new_n18902), .Y(new_n18924));
  nor_5  g16576(.A(new_n18924), .B(new_n18901_1), .Y(new_n18925));
  xnor_4 g16577(.A(new_n18925), .B(new_n18897), .Y(n6022));
  xnor_4 g16578(.A(new_n18584_1), .B(new_n18567), .Y(n6031));
  not_8  g16579(.A(new_n8139_1), .Y(new_n18928));
  and_5  g16580(.A(new_n16241), .B(new_n10873), .Y(new_n18929));
  xnor_4 g16581(.A(new_n18929), .B(n17458), .Y(new_n18930));
  xnor_4 g16582(.A(new_n18930), .B(new_n8719), .Y(new_n18931));
  nor_5  g16583(.A(new_n16242), .B(n15077), .Y(new_n18932));
  and_5  g16584(.A(new_n16279_1), .B(new_n16243_1), .Y(new_n18933));
  nor_5  g16585(.A(new_n18933), .B(new_n18932), .Y(new_n18934));
  xnor_4 g16586(.A(new_n18934), .B(new_n18931), .Y(new_n18935));
  xnor_4 g16587(.A(new_n18935), .B(n12702), .Y(new_n18936));
  and_5  g16588(.A(new_n16280), .B(new_n5611), .Y(new_n18937));
  and_5  g16589(.A(new_n16323), .B(new_n16281), .Y(new_n18938));
  nor_5  g16590(.A(new_n18938), .B(new_n18937), .Y(new_n18939));
  xor_4  g16591(.A(new_n18939), .B(new_n18936), .Y(new_n18940_1));
  xnor_4 g16592(.A(new_n18940_1), .B(new_n18928), .Y(new_n18941));
  nor_5  g16593(.A(new_n16324), .B(new_n8144), .Y(new_n18942));
  nor_5  g16594(.A(new_n16363), .B(new_n16325), .Y(new_n18943));
  nor_5  g16595(.A(new_n18943), .B(new_n18942), .Y(new_n18944));
  xnor_4 g16596(.A(new_n18944), .B(new_n18941), .Y(n6044));
  and_5  g16597(.A(new_n9119), .B(new_n9077), .Y(new_n18946));
  and_5  g16598(.A(new_n9177), .B(new_n9120), .Y(new_n18947));
  nor_5  g16599(.A(new_n18947), .B(new_n18946), .Y(new_n18948));
  and_5  g16600(.A(new_n9076), .B(new_n10679), .Y(new_n18949));
  xnor_4 g16601(.A(new_n17629), .B(new_n18949), .Y(new_n18950));
  xnor_4 g16602(.A(new_n18950), .B(new_n18948), .Y(new_n18951));
  nor_5  g16603(.A(new_n18951), .B(new_n4536), .Y(new_n18952));
  xnor_4 g16604(.A(new_n18951), .B(new_n4536), .Y(new_n18953));
  nor_5  g16605(.A(new_n9178), .B(new_n9061), .Y(new_n18954));
  nor_5  g16606(.A(new_n9221), .B(new_n9179), .Y(new_n18955));
  nor_5  g16607(.A(new_n18955), .B(new_n18954), .Y(new_n18956));
  nor_5  g16608(.A(new_n18956), .B(new_n18953), .Y(new_n18957));
  nor_5  g16609(.A(new_n18957), .B(new_n18952), .Y(new_n18958));
  not_8  g16610(.A(new_n18958), .Y(new_n18959));
  nor_5  g16611(.A(new_n17629), .B(new_n18949), .Y(new_n18960));
  and_5  g16612(.A(new_n18960), .B(new_n18948), .Y(new_n18961));
  and_5  g16613(.A(new_n18961), .B(new_n4417), .Y(new_n18962_1));
  and_5  g16614(.A(new_n18962_1), .B(new_n18959), .Y(new_n18963));
  or_5   g16615(.A(new_n18961), .B(new_n4417), .Y(new_n18964));
  nor_5  g16616(.A(new_n18964), .B(new_n18959), .Y(new_n18965));
  or_5   g16617(.A(new_n18965), .B(new_n18963), .Y(n6046));
  xnor_4 g16618(.A(n17077), .B(n7437), .Y(new_n18967));
  nor_5  g16619(.A(n26510), .B(new_n2893), .Y(new_n18968));
  xnor_4 g16620(.A(n26510), .B(n20700), .Y(new_n18969));
  nor_5  g16621(.A(n23068), .B(new_n2896), .Y(new_n18970_1));
  and_5  g16622(.A(new_n18663), .B(new_n18646), .Y(new_n18971));
  or_5   g16623(.A(new_n18971), .B(new_n18970_1), .Y(new_n18972));
  and_5  g16624(.A(new_n18972), .B(new_n18969), .Y(new_n18973));
  or_5   g16625(.A(new_n18973), .B(new_n18968), .Y(new_n18974));
  xor_4  g16626(.A(new_n18974), .B(new_n18967), .Y(new_n18975));
  xnor_4 g16627(.A(n21997), .B(new_n6970), .Y(new_n18976));
  nor_5  g16628(.A(new_n8501), .B(new_n6973), .Y(new_n18977_1));
  or_5   g16629(.A(n25119), .B(n21934), .Y(new_n18978));
  nor_5  g16630(.A(n18901), .B(n1163), .Y(new_n18979));
  and_5  g16631(.A(new_n18629), .B(new_n18618), .Y(new_n18980));
  nor_5  g16632(.A(new_n18980), .B(new_n18979), .Y(new_n18981));
  and_5  g16633(.A(new_n18981), .B(new_n18978), .Y(new_n18982_1));
  nor_5  g16634(.A(new_n18982_1), .B(new_n18977_1), .Y(new_n18983));
  xor_4  g16635(.A(new_n18983), .B(new_n18976), .Y(new_n18984));
  xor_4  g16636(.A(new_n18984), .B(new_n7479), .Y(new_n18985));
  xnor_4 g16637(.A(n25119), .B(n21934), .Y(new_n18986));
  xnor_4 g16638(.A(new_n18986), .B(new_n18981), .Y(new_n18987));
  nor_5  g16639(.A(new_n18987), .B(new_n2430), .Y(new_n18988));
  nor_5  g16640(.A(new_n18630), .B(new_n2423), .Y(new_n18989));
  and_5  g16641(.A(new_n18644), .B(new_n18631), .Y(new_n18990));
  nor_5  g16642(.A(new_n18990), .B(new_n18989), .Y(new_n18991));
  xnor_4 g16643(.A(new_n18987), .B(new_n2431), .Y(new_n18992));
  and_5  g16644(.A(new_n18992), .B(new_n18991), .Y(new_n18993));
  nor_5  g16645(.A(new_n18993), .B(new_n18988), .Y(new_n18994));
  xor_4  g16646(.A(new_n18994), .B(new_n18985), .Y(new_n18995));
  xnor_4 g16647(.A(new_n18995), .B(new_n18975), .Y(new_n18996));
  not_8  g16648(.A(new_n18996), .Y(new_n18997));
  xor_4  g16649(.A(new_n18972), .B(new_n18969), .Y(new_n18998));
  xnor_4 g16650(.A(new_n18992), .B(new_n18991), .Y(new_n18999_1));
  and_5  g16651(.A(new_n18999_1), .B(new_n18998), .Y(new_n19000));
  nor_5  g16652(.A(new_n18664), .B(new_n18645), .Y(new_n19001));
  and_5  g16653(.A(new_n18695), .B(new_n18666), .Y(new_n19002));
  nor_5  g16654(.A(new_n19002), .B(new_n19001), .Y(new_n19003));
  not_8  g16655(.A(new_n18999_1), .Y(new_n19004));
  xnor_4 g16656(.A(new_n19004), .B(new_n18998), .Y(new_n19005_1));
  and_5  g16657(.A(new_n19005_1), .B(new_n19003), .Y(new_n19006));
  nor_5  g16658(.A(new_n19006), .B(new_n19000), .Y(new_n19007));
  xnor_4 g16659(.A(new_n19007), .B(new_n18997), .Y(n6084));
  xnor_4 g16660(.A(new_n18775), .B(new_n10141), .Y(n6160));
  xnor_4 g16661(.A(new_n18780_1), .B(new_n18779), .Y(n6171));
  nor_5  g16662(.A(n22359), .B(new_n7923), .Y(new_n19011));
  and_5  g16663(.A(new_n14865), .B(new_n9849), .Y(new_n19012));
  or_5   g16664(.A(new_n19012), .B(new_n19011), .Y(new_n19013));
  xor_4  g16665(.A(new_n19013), .B(new_n9852), .Y(new_n19014));
  xnor_4 g16666(.A(n26264), .B(n21905), .Y(new_n19015));
  not_8  g16667(.A(n7841), .Y(new_n19016));
  nor_5  g16668(.A(n22918), .B(new_n19016), .Y(new_n19017));
  xnor_4 g16669(.A(n22918), .B(n7841), .Y(new_n19018));
  not_8  g16670(.A(n16812), .Y(new_n19019));
  nor_5  g16671(.A(n25923), .B(new_n19019), .Y(new_n19020));
  xnor_4 g16672(.A(n25923), .B(n16812), .Y(new_n19021));
  not_8  g16673(.A(n25068), .Y(new_n19022));
  nor_5  g16674(.A(new_n19022), .B(n6790), .Y(new_n19023));
  and_5  g16675(.A(new_n17678), .B(new_n17658), .Y(new_n19024));
  or_5   g16676(.A(new_n19024), .B(new_n19023), .Y(new_n19025));
  and_5  g16677(.A(new_n19025), .B(new_n19021), .Y(new_n19026));
  or_5   g16678(.A(new_n19026), .B(new_n19020), .Y(new_n19027));
  and_5  g16679(.A(new_n19027), .B(new_n19018), .Y(new_n19028));
  or_5   g16680(.A(new_n19028), .B(new_n19017), .Y(new_n19029));
  xor_4  g16681(.A(new_n19029), .B(new_n19015), .Y(new_n19030));
  xnor_4 g16682(.A(new_n19030), .B(new_n15187), .Y(new_n19031));
  xor_4  g16683(.A(new_n19027), .B(new_n19018), .Y(new_n19032));
  nor_5  g16684(.A(new_n19032), .B(new_n15192), .Y(new_n19033_1));
  xnor_4 g16685(.A(new_n19032), .B(new_n14932), .Y(new_n19034));
  xor_4  g16686(.A(new_n19025), .B(new_n19021), .Y(new_n19035));
  and_5  g16687(.A(new_n19035), .B(new_n14936), .Y(new_n19036));
  xnor_4 g16688(.A(new_n19035), .B(new_n14935), .Y(new_n19037));
  and_5  g16689(.A(new_n17679), .B(new_n14941), .Y(new_n19038));
  and_5  g16690(.A(new_n17703), .B(new_n17680), .Y(new_n19039));
  or_5   g16691(.A(new_n19039), .B(new_n19038), .Y(new_n19040));
  and_5  g16692(.A(new_n19040), .B(new_n19037), .Y(new_n19041));
  nor_5  g16693(.A(new_n19041), .B(new_n19036), .Y(new_n19042_1));
  and_5  g16694(.A(new_n19042_1), .B(new_n19034), .Y(new_n19043));
  nor_5  g16695(.A(new_n19043), .B(new_n19033_1), .Y(new_n19044_1));
  xor_4  g16696(.A(new_n19044_1), .B(new_n19031), .Y(new_n19045));
  xnor_4 g16697(.A(new_n19045), .B(new_n19014), .Y(new_n19046));
  xnor_4 g16698(.A(new_n19042_1), .B(new_n19034), .Y(new_n19047));
  nor_5  g16699(.A(new_n19047), .B(new_n14866), .Y(new_n19048));
  xnor_4 g16700(.A(new_n19047), .B(new_n14866), .Y(new_n19049));
  xor_4  g16701(.A(new_n19040), .B(new_n19037), .Y(new_n19050));
  nor_5  g16702(.A(new_n19050), .B(new_n14868), .Y(new_n19051));
  xnor_4 g16703(.A(new_n19050), .B(new_n14868), .Y(new_n19052));
  nor_5  g16704(.A(new_n17704), .B(new_n14871), .Y(new_n19053));
  nor_5  g16705(.A(new_n17729), .B(new_n17705), .Y(new_n19054));
  nor_5  g16706(.A(new_n19054), .B(new_n19053), .Y(new_n19055));
  nor_5  g16707(.A(new_n19055), .B(new_n19052), .Y(new_n19056));
  nor_5  g16708(.A(new_n19056), .B(new_n19051), .Y(new_n19057));
  nor_5  g16709(.A(new_n19057), .B(new_n19049), .Y(new_n19058));
  nor_5  g16710(.A(new_n19058), .B(new_n19048), .Y(new_n19059));
  xnor_4 g16711(.A(new_n19059), .B(new_n19046), .Y(n6183));
  xnor_4 g16712(.A(n14702), .B(n14345), .Y(new_n19061));
  nor_5  g16713(.A(new_n9088), .B(n2999), .Y(new_n19062));
  xnor_4 g16714(.A(n11356), .B(n2999), .Y(new_n19063));
  nor_5  g16715(.A(new_n9091), .B(n2547), .Y(new_n19064));
  xnor_4 g16716(.A(n3164), .B(n2547), .Y(new_n19065));
  nor_5  g16717(.A(n10611), .B(new_n10623), .Y(new_n19066));
  and_5  g16718(.A(new_n13792), .B(new_n13783_1), .Y(new_n19067));
  nor_5  g16719(.A(new_n19067), .B(new_n19066), .Y(new_n19068));
  and_5  g16720(.A(new_n19068), .B(new_n19065), .Y(new_n19069));
  or_5   g16721(.A(new_n19069), .B(new_n19064), .Y(new_n19070));
  and_5  g16722(.A(new_n19070), .B(new_n19063), .Y(new_n19071));
  or_5   g16723(.A(new_n19071), .B(new_n19062), .Y(new_n19072));
  xor_4  g16724(.A(new_n19072), .B(new_n19061), .Y(new_n19073));
  xor_4  g16725(.A(new_n19073), .B(new_n9011), .Y(new_n19074));
  xor_4  g16726(.A(new_n19070), .B(new_n19063), .Y(new_n19075));
  nor_5  g16727(.A(new_n19075), .B(new_n9015), .Y(new_n19076));
  xnor_4 g16728(.A(new_n19075), .B(new_n9015), .Y(new_n19077));
  not_8  g16729(.A(new_n9019), .Y(new_n19078));
  xnor_4 g16730(.A(new_n19068), .B(new_n19065), .Y(new_n19079));
  and_5  g16731(.A(new_n19079), .B(new_n19078), .Y(new_n19080));
  xnor_4 g16732(.A(new_n19079), .B(new_n19078), .Y(new_n19081_1));
  and_5  g16733(.A(new_n13793), .B(new_n9023), .Y(new_n19082));
  nor_5  g16734(.A(new_n13808), .B(new_n13794), .Y(new_n19083));
  nor_5  g16735(.A(new_n19083), .B(new_n19082), .Y(new_n19084));
  nor_5  g16736(.A(new_n19084), .B(new_n19081_1), .Y(new_n19085));
  nor_5  g16737(.A(new_n19085), .B(new_n19080), .Y(new_n19086));
  nor_5  g16738(.A(new_n19086), .B(new_n19077), .Y(new_n19087));
  nor_5  g16739(.A(new_n19087), .B(new_n19076), .Y(new_n19088));
  xor_4  g16740(.A(new_n19088), .B(new_n19074), .Y(n6189));
  xnor_4 g16741(.A(n20036), .B(n15167), .Y(new_n19090));
  nor_5  g16742(.A(new_n12134), .B(n11192), .Y(new_n19091));
  or_5   g16743(.A(n21095), .B(new_n4120), .Y(new_n19092));
  nor_5  g16744(.A(n9380), .B(new_n6492), .Y(new_n19093));
  and_5  g16745(.A(new_n19093), .B(new_n19092), .Y(new_n19094));
  or_5   g16746(.A(new_n19094), .B(new_n19091), .Y(new_n19095));
  xor_4  g16747(.A(new_n19095), .B(new_n19090), .Y(new_n19096));
  xnor_4 g16748(.A(new_n19096), .B(new_n17713), .Y(new_n19097));
  xnor_4 g16749(.A(n9380), .B(n8656), .Y(new_n19098));
  nor_5  g16750(.A(new_n19098), .B(new_n17717), .Y(new_n19099));
  xnor_4 g16751(.A(n21095), .B(n11192), .Y(new_n19100));
  xnor_4 g16752(.A(new_n19100), .B(new_n19093), .Y(new_n19101));
  nor_5  g16753(.A(new_n19101), .B(new_n19099), .Y(new_n19102));
  xnor_4 g16754(.A(new_n19101), .B(new_n19099), .Y(new_n19103));
  nor_5  g16755(.A(new_n19103), .B(new_n17721_1), .Y(new_n19104));
  nor_5  g16756(.A(new_n19104), .B(new_n19102), .Y(new_n19105));
  xnor_4 g16757(.A(new_n19105), .B(new_n19097), .Y(n6223));
  xnor_4 g16758(.A(new_n13806), .B(new_n13798_1), .Y(n6233));
  xnor_4 g16759(.A(new_n18311_1), .B(new_n18308), .Y(n6245));
  xnor_4 g16760(.A(new_n10145), .B(new_n10133), .Y(n6248));
  xnor_4 g16761(.A(n21839), .B(n16544), .Y(new_n19110));
  nor_5  g16762(.A(n27089), .B(new_n2887_1), .Y(new_n19111));
  and_5  g16763(.A(new_n18749), .B(new_n18719), .Y(new_n19112));
  or_5   g16764(.A(new_n19112), .B(new_n19111), .Y(new_n19113));
  xor_4  g16765(.A(new_n19113), .B(new_n19110), .Y(new_n19114));
  xnor_4 g16766(.A(new_n19114), .B(new_n10102), .Y(new_n19115));
  nor_5  g16767(.A(new_n18750), .B(new_n10106), .Y(new_n19116_1));
  nor_5  g16768(.A(new_n18791), .B(new_n18751_1), .Y(new_n19117));
  nor_5  g16769(.A(new_n19117), .B(new_n19116_1), .Y(new_n19118));
  xnor_4 g16770(.A(new_n19118), .B(new_n19115), .Y(n6256));
  xnor_4 g16771(.A(new_n14620), .B(new_n14605), .Y(n6271));
  nor_5  g16772(.A(new_n7918), .B(n13549), .Y(new_n19121));
  not_8  g16773(.A(n23493), .Y(new_n19122));
  nor_5  g16774(.A(new_n19122), .B(n8405), .Y(new_n19123));
  and_5  g16775(.A(new_n19013), .B(new_n9852), .Y(new_n19124));
  or_5   g16776(.A(new_n19124), .B(new_n19123), .Y(new_n19125_1));
  and_5  g16777(.A(new_n19125_1), .B(new_n9855), .Y(new_n19126));
  nor_5  g16778(.A(new_n19126), .B(new_n19121), .Y(new_n19127));
  nor_5  g16779(.A(n13951), .B(new_n2674), .Y(new_n19128));
  xnor_4 g16780(.A(n13951), .B(n2944), .Y(new_n19129));
  nor_5  g16781(.A(n22793), .B(new_n2677), .Y(new_n19130));
  or_5   g16782(.A(new_n14650), .B(new_n14631), .Y(new_n19131));
  and_5  g16783(.A(new_n19131), .B(new_n14629), .Y(new_n19132));
  or_5   g16784(.A(new_n19132), .B(new_n19130), .Y(new_n19133));
  and_5  g16785(.A(new_n19133), .B(new_n19129), .Y(new_n19134));
  nor_5  g16786(.A(new_n19134), .B(new_n19128), .Y(new_n19135));
  and_5  g16787(.A(new_n19135), .B(new_n19127), .Y(new_n19136));
  nor_5  g16788(.A(new_n19132), .B(new_n19130), .Y(new_n19137));
  xnor_4 g16789(.A(new_n19137), .B(new_n19129), .Y(new_n19138));
  xor_4  g16790(.A(new_n19125_1), .B(new_n9855), .Y(new_n19139));
  nor_5  g16791(.A(new_n19139), .B(new_n19138), .Y(new_n19140));
  not_8  g16792(.A(new_n19138), .Y(new_n19141_1));
  xnor_4 g16793(.A(new_n19139), .B(new_n19141_1), .Y(new_n19142));
  and_5  g16794(.A(new_n19014), .B(new_n14652), .Y(new_n19143));
  xnor_4 g16795(.A(new_n19014), .B(new_n14653), .Y(new_n19144_1));
  nor_5  g16796(.A(new_n14866), .B(new_n14655), .Y(new_n19145));
  nor_5  g16797(.A(new_n14885), .B(new_n14867), .Y(new_n19146));
  nor_5  g16798(.A(new_n19146), .B(new_n19145), .Y(new_n19147));
  and_5  g16799(.A(new_n19147), .B(new_n19144_1), .Y(new_n19148));
  nor_5  g16800(.A(new_n19148), .B(new_n19143), .Y(new_n19149));
  and_5  g16801(.A(new_n19149), .B(new_n19142), .Y(new_n19150));
  nor_5  g16802(.A(new_n19150), .B(new_n19140), .Y(new_n19151));
  xnor_4 g16803(.A(new_n19135), .B(new_n19127), .Y(new_n19152));
  nor_5  g16804(.A(new_n19152), .B(new_n19151), .Y(new_n19153));
  nor_5  g16805(.A(new_n19153), .B(new_n19136), .Y(new_n19154));
  not_8  g16806(.A(new_n19154), .Y(new_n19155));
  nor_5  g16807(.A(new_n14547_1), .B(n1881), .Y(new_n19156));
  xnor_4 g16808(.A(n8827), .B(n1881), .Y(new_n19157));
  nor_5  g16809(.A(new_n12683), .B(n5834), .Y(new_n19158));
  and_5  g16810(.A(new_n18559), .B(new_n18556), .Y(new_n19159));
  or_5   g16811(.A(new_n19159), .B(new_n19158), .Y(new_n19160));
  and_5  g16812(.A(new_n19160), .B(new_n19157), .Y(new_n19161));
  nor_5  g16813(.A(new_n19161), .B(new_n19156), .Y(new_n19162));
  not_8  g16814(.A(new_n19162), .Y(new_n19163_1));
  xnor_4 g16815(.A(new_n19163_1), .B(new_n19155), .Y(new_n19164_1));
  xnor_4 g16816(.A(new_n19152), .B(new_n19151), .Y(new_n19165));
  nor_5  g16817(.A(new_n19165), .B(new_n19162), .Y(new_n19166));
  not_8  g16818(.A(new_n19165), .Y(new_n19167));
  xnor_4 g16819(.A(new_n19167), .B(new_n19162), .Y(new_n19168));
  xor_4  g16820(.A(new_n19160), .B(new_n19157), .Y(new_n19169));
  xnor_4 g16821(.A(new_n19149), .B(new_n19142), .Y(new_n19170));
  and_5  g16822(.A(new_n19170), .B(new_n19169), .Y(new_n19171));
  xnor_4 g16823(.A(new_n19147), .B(new_n19144_1), .Y(new_n19172));
  not_8  g16824(.A(new_n19172), .Y(new_n19173));
  nor_5  g16825(.A(new_n19173), .B(new_n18560), .Y(new_n19174_1));
  xnor_4 g16826(.A(new_n19172), .B(new_n18560), .Y(new_n19175));
  and_5  g16827(.A(new_n15139_1), .B(new_n14886), .Y(new_n19176_1));
  and_5  g16828(.A(new_n15159), .B(new_n15140), .Y(new_n19177));
  nor_5  g16829(.A(new_n19177), .B(new_n19176_1), .Y(new_n19178));
  and_5  g16830(.A(new_n19178), .B(new_n19175), .Y(new_n19179));
  nor_5  g16831(.A(new_n19179), .B(new_n19174_1), .Y(new_n19180));
  not_8  g16832(.A(new_n19170), .Y(new_n19181));
  xnor_4 g16833(.A(new_n19181), .B(new_n19169), .Y(new_n19182));
  and_5  g16834(.A(new_n19182), .B(new_n19180), .Y(new_n19183));
  nor_5  g16835(.A(new_n19183), .B(new_n19171), .Y(new_n19184));
  and_5  g16836(.A(new_n19184), .B(new_n19168), .Y(new_n19185));
  nor_5  g16837(.A(new_n19185), .B(new_n19166), .Y(new_n19186));
  xor_4  g16838(.A(new_n19186), .B(new_n19164_1), .Y(n6276));
  xnor_4 g16839(.A(new_n18268), .B(new_n18267), .Y(n6308));
  xnor_4 g16840(.A(new_n16450), .B(new_n16436), .Y(n6311));
  xnor_4 g16841(.A(new_n16217_1), .B(new_n16203), .Y(n6323));
  nor_5  g16842(.A(new_n5915), .B(new_n13508), .Y(new_n19191));
  and_5  g16843(.A(new_n5979), .B(new_n5916), .Y(new_n19192));
  nor_5  g16844(.A(new_n19192), .B(new_n19191), .Y(new_n19193));
  not_8  g16845(.A(new_n19193), .Y(new_n19194));
  and_5  g16846(.A(new_n13194), .B(new_n13550), .Y(new_n19195));
  and_5  g16847(.A(new_n19195), .B(new_n19194), .Y(new_n19196_1));
  or_5   g16848(.A(new_n13194), .B(new_n13550), .Y(new_n19197));
  nor_5  g16849(.A(new_n19197), .B(new_n19194), .Y(new_n19198));
  nor_5  g16850(.A(new_n19198), .B(new_n19196_1), .Y(new_n19199));
  nor_5  g16851(.A(new_n19199), .B(new_n17497), .Y(new_n19200));
  xnor_4 g16852(.A(new_n19199), .B(new_n17497), .Y(new_n19201));
  xnor_4 g16853(.A(new_n13193), .B(new_n13550), .Y(new_n19202_1));
  xnor_4 g16854(.A(new_n19202_1), .B(new_n19194), .Y(new_n19203));
  nor_5  g16855(.A(new_n19203), .B(new_n17500_1), .Y(new_n19204));
  xnor_4 g16856(.A(new_n19203), .B(new_n17500_1), .Y(new_n19205));
  nor_5  g16857(.A(new_n6088), .B(new_n5980_1), .Y(new_n19206));
  nor_5  g16858(.A(new_n6149), .B(new_n6089), .Y(new_n19207));
  nor_5  g16859(.A(new_n19207), .B(new_n19206), .Y(new_n19208));
  nor_5  g16860(.A(new_n19208), .B(new_n19205), .Y(new_n19209));
  nor_5  g16861(.A(new_n19209), .B(new_n19204), .Y(new_n19210));
  nor_5  g16862(.A(new_n19210), .B(new_n19201), .Y(new_n19211));
  nor_5  g16863(.A(new_n19211), .B(new_n19200), .Y(new_n19212));
  nor_5  g16864(.A(new_n19212), .B(new_n19196_1), .Y(n6330));
  xnor_4 g16865(.A(new_n8568), .B(new_n8534), .Y(n6339));
  xnor_4 g16866(.A(new_n13775_1), .B(new_n13749), .Y(n6354));
  or_5   g16867(.A(new_n3213), .B(n7335), .Y(new_n19216));
  nor_5  g16868(.A(new_n3220), .B(n5696), .Y(new_n19217));
  xnor_4 g16869(.A(new_n3221), .B(n5696), .Y(new_n19218));
  nor_5  g16870(.A(new_n3226), .B(n13367), .Y(new_n19219));
  xnor_4 g16871(.A(new_n3227), .B(n13367), .Y(new_n19220_1));
  nor_5  g16872(.A(new_n3231), .B(n932), .Y(new_n19221_1));
  xnor_4 g16873(.A(new_n3232), .B(n932), .Y(new_n19222));
  nor_5  g16874(.A(new_n3236), .B(n6691), .Y(new_n19223_1));
  xnor_4 g16875(.A(new_n3237), .B(n6691), .Y(new_n19224_1));
  nor_5  g16876(.A(new_n3241), .B(n3260), .Y(new_n19225));
  xnor_4 g16877(.A(new_n3242), .B(n3260), .Y(new_n19226));
  nor_5  g16878(.A(new_n3246), .B(n20489), .Y(new_n19227));
  nor_5  g16879(.A(new_n3251), .B(n2355), .Y(new_n19228_1));
  xnor_4 g16880(.A(new_n3252), .B(n2355), .Y(new_n19229));
  nor_5  g16881(.A(new_n3262), .B(n11121), .Y(new_n19230));
  or_5   g16882(.A(new_n3117), .B(new_n2448), .Y(new_n19231));
  xor_4  g16883(.A(new_n3262), .B(n11121), .Y(new_n19232));
  and_5  g16884(.A(new_n19232), .B(new_n19231), .Y(new_n19233_1));
  or_5   g16885(.A(new_n19233_1), .B(new_n19230), .Y(new_n19234_1));
  and_5  g16886(.A(new_n19234_1), .B(new_n19229), .Y(new_n19235));
  or_5   g16887(.A(new_n19235), .B(new_n19228_1), .Y(new_n19236));
  xnor_4 g16888(.A(new_n3247), .B(n20489), .Y(new_n19237));
  and_5  g16889(.A(new_n19237), .B(new_n19236), .Y(new_n19238));
  or_5   g16890(.A(new_n19238), .B(new_n19227), .Y(new_n19239));
  and_5  g16891(.A(new_n19239), .B(new_n19226), .Y(new_n19240));
  or_5   g16892(.A(new_n19240), .B(new_n19225), .Y(new_n19241));
  and_5  g16893(.A(new_n19241), .B(new_n19224_1), .Y(new_n19242));
  or_5   g16894(.A(new_n19242), .B(new_n19223_1), .Y(new_n19243));
  and_5  g16895(.A(new_n19243), .B(new_n19222), .Y(new_n19244_1));
  or_5   g16896(.A(new_n19244_1), .B(new_n19221_1), .Y(new_n19245));
  and_5  g16897(.A(new_n19245), .B(new_n19220_1), .Y(new_n19246));
  or_5   g16898(.A(new_n19246), .B(new_n19219), .Y(new_n19247));
  and_5  g16899(.A(new_n19247), .B(new_n19218), .Y(new_n19248));
  nor_5  g16900(.A(new_n19248), .B(new_n19217), .Y(new_n19249));
  and_5  g16901(.A(new_n19249), .B(new_n19216), .Y(new_n19250));
  and_5  g16902(.A(new_n3213), .B(n7335), .Y(new_n19251));
  or_5   g16903(.A(new_n19251), .B(new_n3218), .Y(new_n19252));
  nor_5  g16904(.A(new_n19252), .B(new_n19250), .Y(new_n19253));
  and_5  g16905(.A(new_n19253), .B(new_n16628), .Y(new_n19254));
  nor_5  g16906(.A(new_n19253), .B(new_n16668), .Y(new_n19255));
  xnor_4 g16907(.A(new_n19253), .B(new_n16668), .Y(new_n19256));
  xnor_4 g16908(.A(new_n3214), .B(n7335), .Y(new_n19257));
  xnor_4 g16909(.A(new_n19257), .B(new_n19249), .Y(new_n19258));
  and_5  g16910(.A(new_n19258), .B(new_n16671), .Y(new_n19259));
  xnor_4 g16911(.A(new_n19258), .B(new_n16671), .Y(new_n19260));
  xor_4  g16912(.A(new_n19247), .B(new_n19218), .Y(new_n19261));
  and_5  g16913(.A(new_n19261), .B(new_n16677), .Y(new_n19262));
  xnor_4 g16914(.A(new_n19261), .B(new_n16677), .Y(new_n19263));
  not_8  g16915(.A(new_n16681), .Y(new_n19264));
  xor_4  g16916(.A(new_n19245), .B(new_n19220_1), .Y(new_n19265));
  and_5  g16917(.A(new_n19265), .B(new_n19264), .Y(new_n19266));
  xnor_4 g16918(.A(new_n19265), .B(new_n19264), .Y(new_n19267));
  xor_4  g16919(.A(new_n19243), .B(new_n19222), .Y(new_n19268));
  and_5  g16920(.A(new_n19268), .B(new_n16685), .Y(new_n19269));
  xnor_4 g16921(.A(new_n19268), .B(new_n16685), .Y(new_n19270_1));
  xor_4  g16922(.A(new_n19241), .B(new_n19224_1), .Y(new_n19271));
  and_5  g16923(.A(new_n19271), .B(new_n16690), .Y(new_n19272));
  xnor_4 g16924(.A(new_n19271), .B(new_n16690), .Y(new_n19273));
  xor_4  g16925(.A(new_n19239), .B(new_n19226), .Y(new_n19274));
  and_5  g16926(.A(new_n19274), .B(new_n16695), .Y(new_n19275));
  xnor_4 g16927(.A(new_n19274), .B(new_n16695), .Y(new_n19276));
  xor_4  g16928(.A(new_n19237), .B(new_n19236), .Y(new_n19277));
  and_5  g16929(.A(new_n19277), .B(new_n16698), .Y(new_n19278));
  xnor_4 g16930(.A(new_n19277), .B(new_n16701), .Y(new_n19279));
  xor_4  g16931(.A(new_n19234_1), .B(new_n19229), .Y(new_n19280));
  nor_5  g16932(.A(new_n19280), .B(new_n16704), .Y(new_n19281));
  xor_4  g16933(.A(new_n19280), .B(new_n16704), .Y(new_n19282_1));
  nor_5  g16934(.A(new_n19232), .B(new_n16709), .Y(new_n19283));
  xor_4  g16935(.A(new_n19232), .B(new_n19231), .Y(new_n19284));
  nor_5  g16936(.A(new_n19284), .B(new_n16708), .Y(new_n19285));
  xnor_4 g16937(.A(n16217), .B(n12315), .Y(new_n19286));
  nor_5  g16938(.A(new_n19286), .B(new_n16715), .Y(new_n19287));
  nor_5  g16939(.A(new_n19287), .B(new_n19285), .Y(new_n19288));
  nor_5  g16940(.A(new_n19288), .B(new_n19283), .Y(new_n19289));
  and_5  g16941(.A(new_n19289), .B(new_n19282_1), .Y(new_n19290));
  nor_5  g16942(.A(new_n19290), .B(new_n19281), .Y(new_n19291));
  and_5  g16943(.A(new_n19291), .B(new_n19279), .Y(new_n19292));
  nor_5  g16944(.A(new_n19292), .B(new_n19278), .Y(new_n19293));
  nor_5  g16945(.A(new_n19293), .B(new_n19276), .Y(new_n19294));
  nor_5  g16946(.A(new_n19294), .B(new_n19275), .Y(new_n19295));
  nor_5  g16947(.A(new_n19295), .B(new_n19273), .Y(new_n19296));
  nor_5  g16948(.A(new_n19296), .B(new_n19272), .Y(new_n19297));
  nor_5  g16949(.A(new_n19297), .B(new_n19270_1), .Y(new_n19298));
  nor_5  g16950(.A(new_n19298), .B(new_n19269), .Y(new_n19299));
  nor_5  g16951(.A(new_n19299), .B(new_n19267), .Y(new_n19300));
  nor_5  g16952(.A(new_n19300), .B(new_n19266), .Y(new_n19301));
  nor_5  g16953(.A(new_n19301), .B(new_n19263), .Y(new_n19302));
  nor_5  g16954(.A(new_n19302), .B(new_n19262), .Y(new_n19303));
  nor_5  g16955(.A(new_n19303), .B(new_n19260), .Y(new_n19304));
  nor_5  g16956(.A(new_n19304), .B(new_n19259), .Y(new_n19305));
  nor_5  g16957(.A(new_n19305), .B(new_n19256), .Y(new_n19306));
  nor_5  g16958(.A(new_n19306), .B(new_n19255), .Y(new_n19307));
  nor_5  g16959(.A(new_n19307), .B(new_n19254), .Y(new_n19308));
  nor_5  g16960(.A(new_n19253), .B(new_n16628), .Y(new_n19309));
  nor_5  g16961(.A(new_n19309), .B(new_n19306), .Y(new_n19310));
  nor_5  g16962(.A(new_n19310), .B(new_n19308), .Y(n6375));
  xnor_4 g16963(.A(new_n18434), .B(new_n18420), .Y(n6383));
  xnor_4 g16964(.A(new_n14158), .B(new_n14118), .Y(n6407));
  xnor_4 g16965(.A(new_n8560), .B(new_n8559), .Y(n6431));
  xnor_4 g16966(.A(new_n16062_1), .B(new_n16059), .Y(n6437));
  xnor_4 g16967(.A(new_n4161), .B(new_n4159), .Y(n6457));
  xnor_4 g16968(.A(new_n12099), .B(new_n12070), .Y(n6465));
  not_8  g16969(.A(new_n8339_1), .Y(new_n19318));
  and_5  g16970(.A(new_n16930), .B(n3740), .Y(new_n19319));
  and_5  g16971(.A(new_n16929), .B(new_n5982), .Y(new_n19320));
  nor_5  g16972(.A(new_n16930), .B(n3740), .Y(new_n19321));
  nor_5  g16973(.A(new_n16935), .B(new_n19321), .Y(new_n19322));
  or_5   g16974(.A(new_n19322), .B(new_n19320), .Y(new_n19323_1));
  nor_5  g16975(.A(new_n19323_1), .B(new_n19319), .Y(new_n19324));
  not_8  g16976(.A(new_n19324), .Y(new_n19325));
  xnor_4 g16977(.A(new_n19325), .B(new_n19318), .Y(new_n19326));
  not_8  g16978(.A(new_n3472), .Y(new_n19327_1));
  nor_5  g16979(.A(new_n17928), .B(new_n19327_1), .Y(new_n19328));
  xnor_4 g16980(.A(new_n16936), .B(new_n19327_1), .Y(new_n19329));
  nor_5  g16981(.A(new_n17930), .B(new_n3476), .Y(new_n19330));
  and_5  g16982(.A(new_n14073), .B(new_n14033), .Y(new_n19331));
  nor_5  g16983(.A(new_n19331), .B(new_n19330), .Y(new_n19332));
  and_5  g16984(.A(new_n19332), .B(new_n19329), .Y(new_n19333_1));
  nor_5  g16985(.A(new_n19333_1), .B(new_n19328), .Y(new_n19334));
  xnor_4 g16986(.A(new_n19334), .B(new_n19326), .Y(new_n19335));
  not_8  g16987(.A(new_n19335), .Y(new_n19336));
  nor_5  g16988(.A(new_n3598), .B(n2743), .Y(new_n19337));
  nor_5  g16989(.A(new_n3603), .B(new_n3537), .Y(new_n19338));
  nor_5  g16990(.A(new_n3602), .B(n7026), .Y(new_n19339));
  nor_5  g16991(.A(new_n14105), .B(new_n19339), .Y(new_n19340));
  nor_5  g16992(.A(new_n19340), .B(new_n19338), .Y(new_n19341));
  nor_5  g16993(.A(new_n19341), .B(new_n19337), .Y(new_n19342));
  and_5  g16994(.A(new_n3597), .B(new_n4797), .Y(new_n19343));
  not_8  g16995(.A(new_n3598), .Y(new_n19344));
  nor_5  g16996(.A(new_n19344), .B(new_n13254), .Y(new_n19345));
  or_5   g16997(.A(new_n19345), .B(new_n19343), .Y(new_n19346));
  nor_5  g16998(.A(new_n19346), .B(new_n19342), .Y(new_n19347));
  xnor_4 g16999(.A(new_n19347), .B(new_n19336), .Y(new_n19348_1));
  xnor_4 g17000(.A(new_n19332), .B(new_n19329), .Y(new_n19349));
  not_8  g17001(.A(new_n19349), .Y(new_n19350));
  xnor_4 g17002(.A(new_n19344), .B(n2743), .Y(new_n19351));
  xnor_4 g17003(.A(new_n19351), .B(new_n19341), .Y(new_n19352));
  nor_5  g17004(.A(new_n19352), .B(new_n19350), .Y(new_n19353));
  xnor_4 g17005(.A(new_n19352), .B(new_n19350), .Y(new_n19354_1));
  nor_5  g17006(.A(new_n14106), .B(new_n14074), .Y(new_n19355));
  and_5  g17007(.A(new_n14162), .B(new_n14107_1), .Y(new_n19356));
  nor_5  g17008(.A(new_n19356), .B(new_n19355), .Y(new_n19357_1));
  nor_5  g17009(.A(new_n19357_1), .B(new_n19354_1), .Y(new_n19358));
  nor_5  g17010(.A(new_n19358), .B(new_n19353), .Y(new_n19359));
  xnor_4 g17011(.A(new_n19359), .B(new_n19348_1), .Y(n6470));
  xnor_4 g17012(.A(new_n11409), .B(new_n11387), .Y(n6476));
  xnor_4 g17013(.A(new_n17968_1), .B(new_n17960), .Y(n6506));
  nor_5  g17014(.A(new_n9334), .B(new_n9332), .Y(new_n19363));
  not_8  g17015(.A(new_n19363), .Y(new_n19364));
  nor_5  g17016(.A(new_n19364), .B(new_n9340), .Y(new_n19365));
  not_8  g17017(.A(new_n19365), .Y(new_n19366));
  nor_5  g17018(.A(new_n19366), .B(new_n9327), .Y(new_n19367_1));
  not_8  g17019(.A(new_n19367_1), .Y(new_n19368));
  nor_5  g17020(.A(new_n19368), .B(new_n9322), .Y(new_n19369));
  not_8  g17021(.A(new_n19369), .Y(new_n19370));
  nor_5  g17022(.A(new_n19370), .B(new_n9317), .Y(new_n19371));
  not_8  g17023(.A(new_n19371), .Y(new_n19372));
  nor_5  g17024(.A(new_n19372), .B(new_n9312), .Y(new_n19373));
  not_8  g17025(.A(new_n19373), .Y(new_n19374));
  nor_5  g17026(.A(new_n19374), .B(new_n13829), .Y(new_n19375));
  xnor_4 g17027(.A(new_n19375), .B(new_n13859), .Y(new_n19376));
  xnor_4 g17028(.A(new_n19376), .B(new_n10057_1), .Y(new_n19377));
  xnor_4 g17029(.A(new_n19373), .B(new_n13829), .Y(new_n19378));
  nor_5  g17030(.A(new_n19378), .B(new_n10063), .Y(new_n19379));
  xnor_4 g17031(.A(new_n19378), .B(new_n10063), .Y(new_n19380));
  xnor_4 g17032(.A(new_n19371), .B(new_n9312), .Y(new_n19381));
  nor_5  g17033(.A(new_n19381), .B(new_n9249), .Y(new_n19382));
  xnor_4 g17034(.A(new_n19381), .B(new_n9249), .Y(new_n19383));
  xnor_4 g17035(.A(new_n19369), .B(new_n9317), .Y(new_n19384));
  nor_5  g17036(.A(new_n19384), .B(new_n9251_1), .Y(new_n19385_1));
  xnor_4 g17037(.A(new_n19384), .B(new_n9251_1), .Y(new_n19386));
  xnor_4 g17038(.A(new_n19367_1), .B(new_n9322), .Y(new_n19387));
  nor_5  g17039(.A(new_n19387), .B(new_n9256), .Y(new_n19388));
  xnor_4 g17040(.A(new_n19387), .B(new_n9255), .Y(new_n19389_1));
  xnor_4 g17041(.A(new_n19365), .B(new_n9327), .Y(new_n19390));
  nor_5  g17042(.A(new_n19390), .B(new_n9261_1), .Y(new_n19391));
  xnor_4 g17043(.A(new_n19363), .B(new_n9340), .Y(new_n19392));
  nor_5  g17044(.A(new_n19392), .B(new_n9266), .Y(new_n19393));
  xnor_4 g17045(.A(new_n19392), .B(new_n9265), .Y(new_n19394));
  nor_5  g17046(.A(new_n9335), .B(new_n9272), .Y(new_n19395));
  nor_5  g17047(.A(new_n19395), .B(new_n9274), .Y(new_n19396));
  nor_5  g17048(.A(new_n9335), .B(new_n9300), .Y(new_n19397));
  or_5   g17049(.A(new_n19397), .B(new_n19363), .Y(new_n19398));
  and_5  g17050(.A(new_n19395), .B(new_n9237), .Y(new_n19399));
  nor_5  g17051(.A(new_n19399), .B(new_n19396), .Y(new_n19400));
  and_5  g17052(.A(new_n19400), .B(new_n19398), .Y(new_n19401_1));
  or_5   g17053(.A(new_n19401_1), .B(new_n19396), .Y(new_n19402));
  and_5  g17054(.A(new_n19402), .B(new_n19394), .Y(new_n19403));
  or_5   g17055(.A(new_n19403), .B(new_n19393), .Y(new_n19404));
  xnor_4 g17056(.A(new_n19390), .B(new_n9260), .Y(new_n19405));
  and_5  g17057(.A(new_n19405), .B(new_n19404), .Y(new_n19406));
  or_5   g17058(.A(new_n19406), .B(new_n19391), .Y(new_n19407));
  and_5  g17059(.A(new_n19407), .B(new_n19389_1), .Y(new_n19408));
  nor_5  g17060(.A(new_n19408), .B(new_n19388), .Y(new_n19409));
  nor_5  g17061(.A(new_n19409), .B(new_n19386), .Y(new_n19410));
  nor_5  g17062(.A(new_n19410), .B(new_n19385_1), .Y(new_n19411));
  nor_5  g17063(.A(new_n19411), .B(new_n19383), .Y(new_n19412));
  nor_5  g17064(.A(new_n19412), .B(new_n19382), .Y(new_n19413));
  nor_5  g17065(.A(new_n19413), .B(new_n19380), .Y(new_n19414_1));
  or_5   g17066(.A(new_n19414_1), .B(new_n19379), .Y(new_n19415));
  xor_4  g17067(.A(new_n19415), .B(new_n19377), .Y(new_n19416));
  xor_4  g17068(.A(new_n19416), .B(new_n16280), .Y(new_n19417));
  xnor_4 g17069(.A(new_n19413), .B(new_n19380), .Y(new_n19418));
  nor_5  g17070(.A(new_n19418), .B(new_n16282), .Y(new_n19419));
  xnor_4 g17071(.A(new_n19418), .B(new_n16282), .Y(new_n19420));
  xnor_4 g17072(.A(new_n19411), .B(new_n19383), .Y(new_n19421));
  nor_5  g17073(.A(new_n19421), .B(new_n16289), .Y(new_n19422));
  xnor_4 g17074(.A(new_n19421), .B(new_n16289), .Y(new_n19423));
  xnor_4 g17075(.A(new_n19409), .B(new_n19386), .Y(new_n19424_1));
  nor_5  g17076(.A(new_n19424_1), .B(new_n16294), .Y(new_n19425));
  xnor_4 g17077(.A(new_n19424_1), .B(new_n16292), .Y(new_n19426));
  xor_4  g17078(.A(new_n19407), .B(new_n19389_1), .Y(new_n19427));
  nor_5  g17079(.A(new_n19427), .B(new_n16296), .Y(new_n19428));
  xor_4  g17080(.A(new_n19405), .B(new_n19404), .Y(new_n19429));
  nor_5  g17081(.A(new_n19429), .B(new_n16299), .Y(new_n19430));
  xnor_4 g17082(.A(new_n19429), .B(new_n16299), .Y(new_n19431));
  xor_4  g17083(.A(new_n19402), .B(new_n19394), .Y(new_n19432));
  nor_5  g17084(.A(new_n19432), .B(new_n16302), .Y(new_n19433));
  xnor_4 g17085(.A(new_n19432), .B(new_n16302), .Y(new_n19434));
  xor_4  g17086(.A(new_n19400), .B(new_n19398), .Y(new_n19435));
  nor_5  g17087(.A(new_n19435), .B(new_n16305), .Y(new_n19436));
  xnor_4 g17088(.A(n13714), .B(new_n6628_1), .Y(new_n19437));
  xnor_4 g17089(.A(new_n9334), .B(new_n9272), .Y(new_n19438));
  and_5  g17090(.A(new_n19438), .B(new_n19437), .Y(new_n19439));
  xor_4  g17091(.A(new_n19435), .B(new_n16305), .Y(new_n19440));
  and_5  g17092(.A(new_n19440), .B(new_n19439), .Y(new_n19441));
  nor_5  g17093(.A(new_n19441), .B(new_n19436), .Y(new_n19442));
  nor_5  g17094(.A(new_n19442), .B(new_n19434), .Y(new_n19443));
  nor_5  g17095(.A(new_n19443), .B(new_n19433), .Y(new_n19444));
  nor_5  g17096(.A(new_n19444), .B(new_n19431), .Y(new_n19445));
  nor_5  g17097(.A(new_n19445), .B(new_n19430), .Y(new_n19446));
  xnor_4 g17098(.A(new_n19427), .B(new_n16296), .Y(new_n19447));
  nor_5  g17099(.A(new_n19447), .B(new_n19446), .Y(new_n19448));
  nor_5  g17100(.A(new_n19448), .B(new_n19428), .Y(new_n19449));
  and_5  g17101(.A(new_n19449), .B(new_n19426), .Y(new_n19450_1));
  nor_5  g17102(.A(new_n19450_1), .B(new_n19425), .Y(new_n19451));
  nor_5  g17103(.A(new_n19451), .B(new_n19423), .Y(new_n19452));
  nor_5  g17104(.A(new_n19452), .B(new_n19422), .Y(new_n19453));
  nor_5  g17105(.A(new_n19453), .B(new_n19420), .Y(new_n19454_1));
  nor_5  g17106(.A(new_n19454_1), .B(new_n19419), .Y(new_n19455));
  xor_4  g17107(.A(new_n19455), .B(new_n19417), .Y(n6514));
  and_5  g17108(.A(new_n11376), .B(new_n11288), .Y(new_n19457));
  nor_5  g17109(.A(new_n11413), .B(new_n11377), .Y(new_n19458_1));
  nor_5  g17110(.A(new_n19458_1), .B(new_n19457), .Y(new_n19459));
  not_8  g17111(.A(new_n19459), .Y(new_n19460));
  xnor_4 g17112(.A(new_n11336), .B(new_n11794), .Y(new_n19461));
  and_5  g17113(.A(new_n19461), .B(new_n11375_1), .Y(new_n19462));
  nor_5  g17114(.A(new_n11336), .B(new_n11850), .Y(new_n19463));
  or_5   g17115(.A(new_n11375_1), .B(new_n19463), .Y(new_n19464));
  nor_5  g17116(.A(new_n19464), .B(new_n19461), .Y(new_n19465));
  nor_5  g17117(.A(new_n19465), .B(new_n19462), .Y(new_n19466));
  xnor_4 g17118(.A(new_n19466), .B(new_n19460), .Y(n6542));
  xnor_4 g17119(.A(new_n15040), .B(new_n15027), .Y(n6558));
  xnor_4 g17120(.A(new_n17481), .B(new_n17479), .Y(n6560));
  xnor_4 g17121(.A(new_n6277), .B(new_n4021), .Y(new_n19470));
  nor_5  g17122(.A(new_n6280), .B(new_n4106), .Y(new_n19471));
  xnor_4 g17123(.A(new_n6282), .B(new_n4106), .Y(new_n19472_1));
  nor_5  g17124(.A(new_n12226), .B(n17090), .Y(new_n19473));
  or_5   g17125(.A(new_n6288), .B(new_n4030), .Y(new_n19474));
  xnor_4 g17126(.A(new_n12226), .B(new_n4111), .Y(new_n19475));
  and_5  g17127(.A(new_n19475), .B(new_n19474), .Y(new_n19476));
  nor_5  g17128(.A(new_n19476), .B(new_n19473), .Y(new_n19477_1));
  and_5  g17129(.A(new_n19477_1), .B(new_n19472_1), .Y(new_n19478));
  or_5   g17130(.A(new_n19478), .B(new_n19471), .Y(new_n19479));
  xor_4  g17131(.A(new_n19479), .B(new_n19470), .Y(new_n19480));
  xnor_4 g17132(.A(new_n19480), .B(new_n9673), .Y(new_n19481));
  xor_4  g17133(.A(new_n19477_1), .B(new_n19472_1), .Y(new_n19482));
  nor_5  g17134(.A(new_n19482), .B(new_n9678), .Y(new_n19483));
  xnor_4 g17135(.A(new_n19482), .B(new_n9678), .Y(new_n19484));
  xor_4  g17136(.A(new_n19475), .B(new_n19474), .Y(new_n19485));
  and_5  g17137(.A(new_n19485), .B(new_n9683), .Y(new_n19486));
  nor_5  g17138(.A(new_n17509), .B(new_n9686), .Y(new_n19487));
  xnor_4 g17139(.A(new_n19485), .B(new_n10808), .Y(new_n19488));
  and_5  g17140(.A(new_n19488), .B(new_n19487), .Y(new_n19489));
  nor_5  g17141(.A(new_n19489), .B(new_n19486), .Y(new_n19490));
  nor_5  g17142(.A(new_n19490), .B(new_n19484), .Y(new_n19491));
  nor_5  g17143(.A(new_n19491), .B(new_n19483), .Y(new_n19492));
  xnor_4 g17144(.A(new_n19492), .B(new_n19481), .Y(n6567));
  not_8  g17145(.A(new_n13408), .Y(new_n19494_1));
  nor_5  g17146(.A(new_n19494_1), .B(n8324), .Y(new_n19495));
  not_8  g17147(.A(new_n19495), .Y(new_n19496_1));
  nor_5  g17148(.A(new_n19496_1), .B(n1279), .Y(new_n19497));
  not_8  g17149(.A(new_n19497), .Y(new_n19498));
  nor_5  g17150(.A(new_n19498), .B(n9445), .Y(new_n19499));
  not_8  g17151(.A(new_n19499), .Y(new_n19500));
  nor_5  g17152(.A(new_n19500), .B(n19454), .Y(new_n19501));
  xnor_4 g17153(.A(new_n19501), .B(n1536), .Y(new_n19502));
  xnor_4 g17154(.A(new_n19502), .B(new_n4473), .Y(new_n19503));
  xnor_4 g17155(.A(new_n19499), .B(n19454), .Y(new_n19504));
  nor_5  g17156(.A(new_n19504), .B(new_n4482), .Y(new_n19505));
  xnor_4 g17157(.A(new_n19504), .B(new_n4481), .Y(new_n19506));
  xnor_4 g17158(.A(new_n19497), .B(n9445), .Y(new_n19507));
  nor_5  g17159(.A(new_n19507), .B(new_n4488), .Y(new_n19508));
  xnor_4 g17160(.A(new_n19507), .B(new_n4487), .Y(new_n19509));
  xnor_4 g17161(.A(new_n19495), .B(n1279), .Y(new_n19510));
  nor_5  g17162(.A(new_n19510), .B(new_n4493), .Y(new_n19511));
  xnor_4 g17163(.A(new_n19510), .B(new_n4493), .Y(new_n19512));
  nor_5  g17164(.A(new_n13409_1), .B(new_n3963), .Y(new_n19513));
  nor_5  g17165(.A(new_n13431), .B(new_n13410), .Y(new_n19514_1));
  nor_5  g17166(.A(new_n19514_1), .B(new_n19513), .Y(new_n19515_1));
  nor_5  g17167(.A(new_n19515_1), .B(new_n19512), .Y(new_n19516));
  or_5   g17168(.A(new_n19516), .B(new_n19511), .Y(new_n19517));
  and_5  g17169(.A(new_n19517), .B(new_n19509), .Y(new_n19518));
  or_5   g17170(.A(new_n19518), .B(new_n19508), .Y(new_n19519));
  and_5  g17171(.A(new_n19519), .B(new_n19506), .Y(new_n19520));
  nor_5  g17172(.A(new_n19520), .B(new_n19505), .Y(new_n19521));
  xnor_4 g17173(.A(new_n19521), .B(new_n19503), .Y(new_n19522));
  not_8  g17174(.A(new_n19522), .Y(new_n19523_1));
  xnor_4 g17175(.A(new_n8079), .B(n23272), .Y(new_n19524));
  nor_5  g17176(.A(new_n8081), .B(n11481), .Y(new_n19525));
  xnor_4 g17177(.A(new_n8081), .B(new_n4361), .Y(new_n19526));
  nor_5  g17178(.A(new_n8084), .B(n16439), .Y(new_n19527));
  xnor_4 g17179(.A(new_n8084), .B(new_n4365), .Y(new_n19528));
  nor_5  g17180(.A(new_n8087), .B(n15241), .Y(new_n19529));
  nor_5  g17181(.A(new_n8093), .B(new_n4373), .Y(new_n19530));
  and_5  g17182(.A(new_n13450), .B(new_n13433), .Y(new_n19531_1));
  nor_5  g17183(.A(new_n19531_1), .B(new_n19530), .Y(new_n19532));
  xnor_4 g17184(.A(new_n8087), .B(new_n4369), .Y(new_n19533));
  and_5  g17185(.A(new_n19533), .B(new_n19532), .Y(new_n19534));
  or_5   g17186(.A(new_n19534), .B(new_n19529), .Y(new_n19535));
  and_5  g17187(.A(new_n19535), .B(new_n19528), .Y(new_n19536));
  or_5   g17188(.A(new_n19536), .B(new_n19527), .Y(new_n19537));
  and_5  g17189(.A(new_n19537), .B(new_n19526), .Y(new_n19538));
  nor_5  g17190(.A(new_n19538), .B(new_n19525), .Y(new_n19539_1));
  xor_4  g17191(.A(new_n19539_1), .B(new_n19524), .Y(new_n19540));
  xnor_4 g17192(.A(new_n19540), .B(new_n19523_1), .Y(new_n19541));
  xor_4  g17193(.A(new_n19519), .B(new_n19506), .Y(new_n19542));
  xor_4  g17194(.A(new_n19537), .B(new_n19526), .Y(new_n19543));
  and_5  g17195(.A(new_n19543), .B(new_n19542), .Y(new_n19544));
  xnor_4 g17196(.A(new_n19543), .B(new_n19542), .Y(new_n19545));
  xor_4  g17197(.A(new_n19517), .B(new_n19509), .Y(new_n19546));
  xor_4  g17198(.A(new_n19535), .B(new_n19528), .Y(new_n19547));
  and_5  g17199(.A(new_n19547), .B(new_n19546), .Y(new_n19548));
  xnor_4 g17200(.A(new_n19547), .B(new_n19546), .Y(new_n19549));
  xnor_4 g17201(.A(new_n19515_1), .B(new_n19512), .Y(new_n19550));
  xnor_4 g17202(.A(new_n19533), .B(new_n19532), .Y(new_n19551));
  nor_5  g17203(.A(new_n19551), .B(new_n19550), .Y(new_n19552));
  xnor_4 g17204(.A(new_n19551), .B(new_n19550), .Y(new_n19553));
  nor_5  g17205(.A(new_n13451), .B(new_n13432), .Y(new_n19554));
  nor_5  g17206(.A(new_n13482), .B(new_n13452), .Y(new_n19555));
  nor_5  g17207(.A(new_n19555), .B(new_n19554), .Y(new_n19556));
  nor_5  g17208(.A(new_n19556), .B(new_n19553), .Y(new_n19557));
  nor_5  g17209(.A(new_n19557), .B(new_n19552), .Y(new_n19558));
  nor_5  g17210(.A(new_n19558), .B(new_n19549), .Y(new_n19559));
  nor_5  g17211(.A(new_n19559), .B(new_n19548), .Y(new_n19560));
  nor_5  g17212(.A(new_n19560), .B(new_n19545), .Y(new_n19561));
  nor_5  g17213(.A(new_n19561), .B(new_n19544), .Y(new_n19562));
  xnor_4 g17214(.A(new_n19562), .B(new_n19541), .Y(n6576));
  xnor_4 g17215(.A(new_n19284), .B(new_n16708), .Y(new_n19564));
  xnor_4 g17216(.A(new_n19564), .B(new_n19287), .Y(n6587));
  xnor_4 g17217(.A(new_n18280), .B(new_n18234), .Y(n6612));
  nor_5  g17218(.A(new_n16992), .B(new_n10685), .Y(new_n19567));
  xnor_4 g17219(.A(new_n16992), .B(new_n10685), .Y(new_n19568));
  nor_5  g17220(.A(new_n16994_1), .B(new_n10676), .Y(new_n19569));
  xnor_4 g17221(.A(new_n16994_1), .B(new_n10676), .Y(new_n19570_1));
  nor_5  g17222(.A(new_n16997), .B(new_n10667), .Y(new_n19571));
  xnor_4 g17223(.A(new_n16997), .B(new_n10667), .Y(new_n19572));
  nor_5  g17224(.A(new_n17000), .B(new_n10658), .Y(new_n19573));
  xnor_4 g17225(.A(new_n17000), .B(new_n10658), .Y(new_n19574));
  nor_5  g17226(.A(new_n17003), .B(new_n10649), .Y(new_n19575_1));
  xnor_4 g17227(.A(new_n17003), .B(new_n10649), .Y(new_n19576));
  nor_5  g17228(.A(new_n17005), .B(new_n10639), .Y(new_n19577));
  xnor_4 g17229(.A(new_n17005), .B(new_n10639), .Y(new_n19578));
  nor_5  g17230(.A(new_n14750), .B(new_n10629), .Y(new_n19579));
  xnor_4 g17231(.A(new_n14750), .B(new_n10629), .Y(new_n19580));
  nor_5  g17232(.A(new_n14753), .B(new_n10620), .Y(new_n19581));
  nor_5  g17233(.A(new_n10607), .B(n18), .Y(new_n19582));
  and_5  g17234(.A(new_n19582), .B(new_n9099), .Y(new_n19583));
  nor_5  g17235(.A(new_n19582), .B(new_n14756), .Y(new_n19584_1));
  nor_5  g17236(.A(new_n19584_1), .B(new_n19583), .Y(new_n19585));
  and_5  g17237(.A(new_n19585), .B(new_n10611_1), .Y(new_n19586));
  nor_5  g17238(.A(new_n19586), .B(new_n19583), .Y(new_n19587));
  xnor_4 g17239(.A(new_n14752), .B(new_n10620), .Y(new_n19588));
  and_5  g17240(.A(new_n19588), .B(new_n19587), .Y(new_n19589));
  or_5   g17241(.A(new_n19589), .B(new_n19581), .Y(new_n19590));
  nor_5  g17242(.A(new_n19590), .B(new_n19580), .Y(new_n19591));
  nor_5  g17243(.A(new_n19591), .B(new_n19579), .Y(new_n19592));
  nor_5  g17244(.A(new_n19592), .B(new_n19578), .Y(new_n19593));
  nor_5  g17245(.A(new_n19593), .B(new_n19577), .Y(new_n19594));
  nor_5  g17246(.A(new_n19594), .B(new_n19576), .Y(new_n19595));
  nor_5  g17247(.A(new_n19595), .B(new_n19575_1), .Y(new_n19596));
  nor_5  g17248(.A(new_n19596), .B(new_n19574), .Y(new_n19597));
  nor_5  g17249(.A(new_n19597), .B(new_n19573), .Y(new_n19598));
  nor_5  g17250(.A(new_n19598), .B(new_n19572), .Y(new_n19599));
  nor_5  g17251(.A(new_n19599), .B(new_n19571), .Y(new_n19600));
  nor_5  g17252(.A(new_n19600), .B(new_n19570_1), .Y(new_n19601));
  nor_5  g17253(.A(new_n19601), .B(new_n19569), .Y(new_n19602_1));
  nor_5  g17254(.A(new_n19602_1), .B(new_n19568), .Y(new_n19603));
  nor_5  g17255(.A(new_n19603), .B(new_n19567), .Y(new_n19604));
  and_5  g17256(.A(new_n16991), .B(new_n17625), .Y(new_n19605));
  and_5  g17257(.A(new_n17634), .B(new_n19605), .Y(new_n19606));
  and_5  g17258(.A(new_n19606), .B(new_n19604), .Y(new_n19607));
  or_5   g17259(.A(new_n17634), .B(new_n19605), .Y(new_n19608_1));
  nor_5  g17260(.A(new_n19608_1), .B(new_n19604), .Y(new_n19609));
  nor_5  g17261(.A(new_n19609), .B(new_n19607), .Y(new_n19610));
  xnor_4 g17262(.A(new_n17181), .B(new_n19605), .Y(new_n19611));
  xnor_4 g17263(.A(new_n19611), .B(new_n19604), .Y(new_n19612));
  nor_5  g17264(.A(new_n19612), .B(new_n18899), .Y(new_n19613));
  xnor_4 g17265(.A(new_n19612), .B(new_n18899), .Y(new_n19614));
  xor_4  g17266(.A(new_n19602_1), .B(new_n19568), .Y(new_n19615));
  and_5  g17267(.A(new_n19615), .B(new_n18904), .Y(new_n19616));
  xnor_4 g17268(.A(new_n19615), .B(new_n18904), .Y(new_n19617_1));
  xor_4  g17269(.A(new_n19600), .B(new_n19570_1), .Y(new_n19618_1));
  and_5  g17270(.A(new_n19618_1), .B(new_n18908), .Y(new_n19619));
  xnor_4 g17271(.A(new_n19618_1), .B(new_n18908), .Y(new_n19620));
  xor_4  g17272(.A(new_n19598), .B(new_n19572), .Y(new_n19621));
  and_5  g17273(.A(new_n19621), .B(new_n18912), .Y(new_n19622));
  xnor_4 g17274(.A(new_n19621), .B(new_n18912), .Y(new_n19623_1));
  xor_4  g17275(.A(new_n19596), .B(new_n19574), .Y(new_n19624));
  and_5  g17276(.A(new_n19624), .B(new_n9350), .Y(new_n19625));
  xnor_4 g17277(.A(new_n19624), .B(new_n9350), .Y(new_n19626));
  xor_4  g17278(.A(new_n19594), .B(new_n19576), .Y(new_n19627));
  and_5  g17279(.A(new_n19627), .B(new_n9354), .Y(new_n19628));
  xnor_4 g17280(.A(new_n19627), .B(new_n9354), .Y(new_n19629));
  xor_4  g17281(.A(new_n19592), .B(new_n19578), .Y(new_n19630));
  and_5  g17282(.A(new_n19630), .B(new_n9359), .Y(new_n19631));
  xnor_4 g17283(.A(new_n19630), .B(new_n9359), .Y(new_n19632));
  xor_4  g17284(.A(new_n19590), .B(new_n19580), .Y(new_n19633));
  and_5  g17285(.A(new_n19633), .B(new_n9364_1), .Y(new_n19634));
  xnor_4 g17286(.A(new_n19633), .B(new_n9364_1), .Y(new_n19635));
  xor_4  g17287(.A(new_n19588), .B(new_n19587), .Y(new_n19636));
  nor_5  g17288(.A(new_n19636), .B(new_n9370), .Y(new_n19637));
  xnor_4 g17289(.A(new_n19636), .B(new_n9370), .Y(new_n19638));
  xnor_4 g17290(.A(new_n19585), .B(new_n13147), .Y(new_n19639));
  and_5  g17291(.A(new_n19639), .B(new_n9373), .Y(new_n19640));
  xnor_4 g17292(.A(new_n10607), .B(new_n6596_1), .Y(new_n19641_1));
  nor_5  g17293(.A(new_n19641_1), .B(new_n9377), .Y(new_n19642));
  xnor_4 g17294(.A(new_n19639), .B(new_n9373), .Y(new_n19643));
  nor_5  g17295(.A(new_n19643), .B(new_n19642), .Y(new_n19644));
  nor_5  g17296(.A(new_n19644), .B(new_n19640), .Y(new_n19645));
  nor_5  g17297(.A(new_n19645), .B(new_n19638), .Y(new_n19646));
  nor_5  g17298(.A(new_n19646), .B(new_n19637), .Y(new_n19647));
  nor_5  g17299(.A(new_n19647), .B(new_n19635), .Y(new_n19648_1));
  nor_5  g17300(.A(new_n19648_1), .B(new_n19634), .Y(new_n19649));
  nor_5  g17301(.A(new_n19649), .B(new_n19632), .Y(new_n19650));
  nor_5  g17302(.A(new_n19650), .B(new_n19631), .Y(new_n19651));
  nor_5  g17303(.A(new_n19651), .B(new_n19629), .Y(new_n19652_1));
  nor_5  g17304(.A(new_n19652_1), .B(new_n19628), .Y(new_n19653));
  nor_5  g17305(.A(new_n19653), .B(new_n19626), .Y(new_n19654));
  nor_5  g17306(.A(new_n19654), .B(new_n19625), .Y(new_n19655));
  nor_5  g17307(.A(new_n19655), .B(new_n19623_1), .Y(new_n19656));
  nor_5  g17308(.A(new_n19656), .B(new_n19622), .Y(new_n19657));
  nor_5  g17309(.A(new_n19657), .B(new_n19620), .Y(new_n19658));
  nor_5  g17310(.A(new_n19658), .B(new_n19619), .Y(new_n19659));
  nor_5  g17311(.A(new_n19659), .B(new_n19617_1), .Y(new_n19660));
  nor_5  g17312(.A(new_n19660), .B(new_n19616), .Y(new_n19661));
  nor_5  g17313(.A(new_n19661), .B(new_n19614), .Y(new_n19662));
  or_5   g17314(.A(new_n19662), .B(new_n19613), .Y(new_n19663));
  not_8  g17315(.A(new_n19663), .Y(new_n19664_1));
  xnor_4 g17316(.A(new_n19664_1), .B(new_n18895), .Y(new_n19665));
  xnor_4 g17317(.A(new_n19665), .B(new_n19610), .Y(n6628));
  xnor_4 g17318(.A(new_n2835), .B(new_n2815), .Y(n6630));
  not_8  g17319(.A(n17911), .Y(new_n19668));
  xnor_4 g17320(.A(n25331), .B(new_n19668), .Y(new_n19669));
  nor_5  g17321(.A(n21997), .B(n18483), .Y(new_n19670));
  and_5  g17322(.A(new_n18983), .B(new_n18976), .Y(new_n19671));
  or_5   g17323(.A(new_n19671), .B(new_n19670), .Y(new_n19672));
  xor_4  g17324(.A(new_n19672), .B(new_n19669), .Y(new_n19673));
  xnor_4 g17325(.A(new_n19673), .B(new_n7487), .Y(new_n19674));
  nor_5  g17326(.A(new_n18984), .B(new_n7479), .Y(new_n19675));
  and_5  g17327(.A(new_n18994), .B(new_n18985), .Y(new_n19676));
  or_5   g17328(.A(new_n19676), .B(new_n19675), .Y(new_n19677));
  xor_4  g17329(.A(new_n19677), .B(new_n19674), .Y(new_n19678));
  xnor_4 g17330(.A(n14130), .B(n468), .Y(new_n19679));
  nor_5  g17331(.A(n16482), .B(new_n8280), .Y(new_n19680_1));
  xnor_4 g17332(.A(n16482), .B(n5400), .Y(new_n19681));
  nor_5  g17333(.A(new_n8284), .B(n9942), .Y(new_n19682));
  nor_5  g17334(.A(n25643), .B(new_n8353), .Y(new_n19683));
  xnor_4 g17335(.A(n25643), .B(n329), .Y(new_n19684));
  nor_5  g17336(.A(new_n13046), .B(n9557), .Y(new_n19685));
  xnor_4 g17337(.A(n24170), .B(n9557), .Y(new_n19686));
  nor_5  g17338(.A(new_n5106), .B(n2409), .Y(new_n19687));
  xnor_4 g17339(.A(n3136), .B(n2409), .Y(new_n19688));
  nor_5  g17340(.A(n8869), .B(new_n2359), .Y(new_n19689));
  and_5  g17341(.A(new_n18608), .B(new_n18605), .Y(new_n19690));
  or_5   g17342(.A(new_n19690), .B(new_n19689), .Y(new_n19691));
  and_5  g17343(.A(new_n19691), .B(new_n19688), .Y(new_n19692));
  nor_5  g17344(.A(new_n19692), .B(new_n19687), .Y(new_n19693));
  and_5  g17345(.A(new_n19693), .B(new_n19686), .Y(new_n19694));
  or_5   g17346(.A(new_n19694), .B(new_n19685), .Y(new_n19695));
  and_5  g17347(.A(new_n19695), .B(new_n19684), .Y(new_n19696));
  or_5   g17348(.A(new_n19696), .B(new_n19683), .Y(new_n19697));
  xnor_4 g17349(.A(n23923), .B(n9942), .Y(new_n19698));
  and_5  g17350(.A(new_n19698), .B(new_n19697), .Y(new_n19699));
  or_5   g17351(.A(new_n19699), .B(new_n19682), .Y(new_n19700));
  and_5  g17352(.A(new_n19700), .B(new_n19681), .Y(new_n19701_1));
  or_5   g17353(.A(new_n19701_1), .B(new_n19680_1), .Y(new_n19702));
  xor_4  g17354(.A(new_n19702), .B(new_n19679), .Y(new_n19703));
  xor_4  g17355(.A(new_n19703), .B(new_n19678), .Y(new_n19704));
  xor_4  g17356(.A(new_n19700), .B(new_n19681), .Y(new_n19705));
  nor_5  g17357(.A(new_n19705), .B(new_n18995), .Y(new_n19706));
  xnor_4 g17358(.A(new_n19705), .B(new_n18995), .Y(new_n19707));
  not_8  g17359(.A(new_n19707), .Y(new_n19708));
  xor_4  g17360(.A(new_n19698), .B(new_n19697), .Y(new_n19709));
  and_5  g17361(.A(new_n19709), .B(new_n18999_1), .Y(new_n19710));
  xor_4  g17362(.A(new_n19695), .B(new_n19684), .Y(new_n19711));
  nor_5  g17363(.A(new_n19711), .B(new_n18645), .Y(new_n19712));
  xnor_4 g17364(.A(new_n19711), .B(new_n18645), .Y(new_n19713));
  xnor_4 g17365(.A(new_n19693), .B(new_n19686), .Y(new_n19714));
  and_5  g17366(.A(new_n19714), .B(new_n18670), .Y(new_n19715));
  xnor_4 g17367(.A(new_n19714), .B(new_n18670), .Y(new_n19716));
  xor_4  g17368(.A(new_n19691), .B(new_n19688), .Y(new_n19717));
  and_5  g17369(.A(new_n19717), .B(new_n18672), .Y(new_n19718));
  xnor_4 g17370(.A(new_n19717), .B(new_n18672), .Y(new_n19719));
  and_5  g17371(.A(new_n18609), .B(new_n18676), .Y(new_n19720));
  and_5  g17372(.A(new_n18613), .B(new_n18610_1), .Y(new_n19721));
  nor_5  g17373(.A(new_n19721), .B(new_n19720), .Y(new_n19722));
  nor_5  g17374(.A(new_n19722), .B(new_n19719), .Y(new_n19723));
  nor_5  g17375(.A(new_n19723), .B(new_n19718), .Y(new_n19724));
  nor_5  g17376(.A(new_n19724), .B(new_n19716), .Y(new_n19725));
  nor_5  g17377(.A(new_n19725), .B(new_n19715), .Y(new_n19726));
  nor_5  g17378(.A(new_n19726), .B(new_n19713), .Y(new_n19727));
  nor_5  g17379(.A(new_n19727), .B(new_n19712), .Y(new_n19728));
  xnor_4 g17380(.A(new_n19709), .B(new_n19004), .Y(new_n19729));
  and_5  g17381(.A(new_n19729), .B(new_n19728), .Y(new_n19730));
  nor_5  g17382(.A(new_n19730), .B(new_n19710), .Y(new_n19731));
  and_5  g17383(.A(new_n19731), .B(new_n19708), .Y(new_n19732));
  nor_5  g17384(.A(new_n19732), .B(new_n19706), .Y(new_n19733));
  xor_4  g17385(.A(new_n19733), .B(new_n19704), .Y(n6634));
  xnor_4 g17386(.A(new_n6577), .B(new_n6563), .Y(n6652));
  xnor_4 g17387(.A(new_n12344), .B(new_n12331), .Y(n6655));
  xnor_4 g17388(.A(new_n11892), .B(new_n11874), .Y(n6669));
  xnor_4 g17389(.A(new_n9385), .B(new_n9367), .Y(n6671));
  xnor_4 g17390(.A(new_n13296), .B(new_n13279), .Y(n6673));
  and_5  g17391(.A(new_n19466), .B(new_n19460), .Y(new_n19740));
  or_5   g17392(.A(new_n11336), .B(new_n11793), .Y(new_n19741));
  nor_5  g17393(.A(new_n19464), .B(new_n19741), .Y(new_n19742));
  or_5   g17394(.A(new_n19742), .B(new_n19740), .Y(n6674));
  xnor_4 g17395(.A(new_n16215_1), .B(new_n16206_1), .Y(n6684));
  xor_4  g17396(.A(new_n12106), .B(new_n12061), .Y(n6706));
  xnor_4 g17397(.A(n12702), .B(n8614), .Y(new_n19746));
  nor_5  g17398(.A(n26797), .B(n15182), .Y(new_n19747));
  xnor_4 g17399(.A(n26797), .B(n15182), .Y(new_n19748));
  nor_5  g17400(.A(n27037), .B(n23913), .Y(new_n19749_1));
  xnor_4 g17401(.A(n27037), .B(n23913), .Y(new_n19750));
  nor_5  g17402(.A(n22554), .B(n8964), .Y(new_n19751));
  xnor_4 g17403(.A(n22554), .B(n8964), .Y(new_n19752));
  nor_5  g17404(.A(n20429), .B(n20151), .Y(new_n19753));
  xnor_4 g17405(.A(n20429), .B(n20151), .Y(new_n19754));
  nor_5  g17406(.A(n7693), .B(n3909), .Y(new_n19755));
  xnor_4 g17407(.A(n7693), .B(n3909), .Y(new_n19756_1));
  nor_5  g17408(.A(n23974), .B(n10405), .Y(new_n19757));
  xnor_4 g17409(.A(n23974), .B(new_n4021), .Y(new_n19758));
  nor_5  g17410(.A(new_n4106), .B(new_n8050), .Y(new_n19759));
  or_5   g17411(.A(n11302), .B(n2146), .Y(new_n19760));
  nor_5  g17412(.A(n22173), .B(n17090), .Y(new_n19761));
  nor_5  g17413(.A(new_n15353_1), .B(new_n15352), .Y(new_n19762));
  nor_5  g17414(.A(new_n19762), .B(new_n19761), .Y(new_n19763));
  and_5  g17415(.A(new_n19763), .B(new_n19760), .Y(new_n19764));
  nor_5  g17416(.A(new_n19764), .B(new_n19759), .Y(new_n19765));
  and_5  g17417(.A(new_n19765), .B(new_n19758), .Y(new_n19766));
  nor_5  g17418(.A(new_n19766), .B(new_n19757), .Y(new_n19767_1));
  nor_5  g17419(.A(new_n19767_1), .B(new_n19756_1), .Y(new_n19768));
  nor_5  g17420(.A(new_n19768), .B(new_n19755), .Y(new_n19769));
  nor_5  g17421(.A(new_n19769), .B(new_n19754), .Y(new_n19770_1));
  nor_5  g17422(.A(new_n19770_1), .B(new_n19753), .Y(new_n19771));
  nor_5  g17423(.A(new_n19771), .B(new_n19752), .Y(new_n19772));
  nor_5  g17424(.A(new_n19772), .B(new_n19751), .Y(new_n19773));
  nor_5  g17425(.A(new_n19773), .B(new_n19750), .Y(new_n19774));
  nor_5  g17426(.A(new_n19774), .B(new_n19749_1), .Y(new_n19775));
  nor_5  g17427(.A(new_n19775), .B(new_n19748), .Y(new_n19776));
  nor_5  g17428(.A(new_n19776), .B(new_n19747), .Y(new_n19777));
  xnor_4 g17429(.A(new_n19777), .B(new_n19746), .Y(new_n19778));
  nor_5  g17430(.A(new_n19778), .B(new_n6152), .Y(new_n19779));
  xnor_4 g17431(.A(new_n19778), .B(new_n6152), .Y(new_n19780_1));
  xnor_4 g17432(.A(new_n19775), .B(new_n19748), .Y(new_n19781));
  nor_5  g17433(.A(new_n19781), .B(new_n13645), .Y(new_n19782));
  xnor_4 g17434(.A(new_n19781), .B(new_n13645), .Y(new_n19783));
  xnor_4 g17435(.A(new_n19773), .B(new_n19750), .Y(new_n19784));
  nor_5  g17436(.A(new_n19784), .B(new_n13648), .Y(new_n19785));
  xnor_4 g17437(.A(new_n19784), .B(new_n13648), .Y(new_n19786));
  xnor_4 g17438(.A(new_n19771), .B(new_n19752), .Y(new_n19787));
  nor_5  g17439(.A(new_n19787), .B(new_n13651), .Y(new_n19788));
  xnor_4 g17440(.A(new_n19787), .B(new_n13651), .Y(new_n19789_1));
  xnor_4 g17441(.A(new_n19769), .B(new_n19754), .Y(new_n19790));
  nor_5  g17442(.A(new_n19790), .B(new_n6164), .Y(new_n19791));
  xnor_4 g17443(.A(new_n19790), .B(new_n6164), .Y(new_n19792_1));
  xnor_4 g17444(.A(new_n19767_1), .B(new_n19756_1), .Y(new_n19793));
  nor_5  g17445(.A(new_n19793), .B(new_n6167), .Y(new_n19794));
  xnor_4 g17446(.A(new_n19793), .B(new_n6167), .Y(new_n19795));
  xnor_4 g17447(.A(new_n19765), .B(new_n19758), .Y(new_n19796));
  not_8  g17448(.A(new_n19796), .Y(new_n19797));
  and_5  g17449(.A(new_n19797), .B(n20169), .Y(new_n19798_1));
  xnor_4 g17450(.A(new_n19797), .B(n20169), .Y(new_n19799));
  xnor_4 g17451(.A(n11302), .B(n2146), .Y(new_n19800));
  xnor_4 g17452(.A(new_n19800), .B(new_n19763), .Y(new_n19801));
  nor_5  g17453(.A(new_n19801), .B(new_n6173), .Y(new_n19802));
  xnor_4 g17454(.A(new_n19801), .B(n8285), .Y(new_n19803_1));
  and_5  g17455(.A(new_n15354), .B(new_n15351), .Y(new_n19804));
  or_5   g17456(.A(new_n19804), .B(new_n15350), .Y(new_n19805));
  and_5  g17457(.A(new_n19805), .B(new_n19803_1), .Y(new_n19806));
  nor_5  g17458(.A(new_n19806), .B(new_n19802), .Y(new_n19807));
  nor_5  g17459(.A(new_n19807), .B(new_n19799), .Y(new_n19808));
  nor_5  g17460(.A(new_n19808), .B(new_n19798_1), .Y(new_n19809));
  nor_5  g17461(.A(new_n19809), .B(new_n19795), .Y(new_n19810));
  nor_5  g17462(.A(new_n19810), .B(new_n19794), .Y(new_n19811));
  nor_5  g17463(.A(new_n19811), .B(new_n19792_1), .Y(new_n19812));
  nor_5  g17464(.A(new_n19812), .B(new_n19791), .Y(new_n19813));
  nor_5  g17465(.A(new_n19813), .B(new_n19789_1), .Y(new_n19814));
  nor_5  g17466(.A(new_n19814), .B(new_n19788), .Y(new_n19815));
  nor_5  g17467(.A(new_n19815), .B(new_n19786), .Y(new_n19816));
  nor_5  g17468(.A(new_n19816), .B(new_n19785), .Y(new_n19817));
  nor_5  g17469(.A(new_n19817), .B(new_n19783), .Y(new_n19818));
  nor_5  g17470(.A(new_n19818), .B(new_n19782), .Y(new_n19819));
  nor_5  g17471(.A(new_n19819), .B(new_n19780_1), .Y(new_n19820));
  nor_5  g17472(.A(new_n19820), .B(new_n19779), .Y(new_n19821));
  nor_5  g17473(.A(n12702), .B(n8614), .Y(new_n19822));
  nor_5  g17474(.A(new_n19777), .B(new_n19746), .Y(new_n19823));
  nor_5  g17475(.A(new_n19823), .B(new_n19822), .Y(new_n19824));
  xnor_4 g17476(.A(new_n19824), .B(new_n19821), .Y(new_n19825));
  and_5  g17477(.A(new_n19502), .B(new_n4477), .Y(new_n19826));
  and_5  g17478(.A(new_n19521), .B(new_n19503), .Y(new_n19827));
  nor_5  g17479(.A(new_n19827), .B(new_n19826), .Y(new_n19828));
  not_8  g17480(.A(new_n19828), .Y(new_n19829));
  not_8  g17481(.A(new_n19501), .Y(new_n19830));
  nor_5  g17482(.A(new_n19830), .B(n1536), .Y(new_n19831));
  xnor_4 g17483(.A(new_n19831), .B(new_n4538), .Y(new_n19832));
  xnor_4 g17484(.A(new_n19832), .B(new_n19829), .Y(new_n19833));
  xnor_4 g17485(.A(new_n19833), .B(new_n19825), .Y(new_n19834));
  xnor_4 g17486(.A(new_n19819), .B(new_n19780_1), .Y(new_n19835));
  nor_5  g17487(.A(new_n19835), .B(new_n19523_1), .Y(new_n19836));
  xnor_4 g17488(.A(new_n19835), .B(new_n19523_1), .Y(new_n19837));
  xnor_4 g17489(.A(new_n19817), .B(new_n19783), .Y(new_n19838));
  not_8  g17490(.A(new_n19838), .Y(new_n19839));
  and_5  g17491(.A(new_n19839), .B(new_n19542), .Y(new_n19840));
  xnor_4 g17492(.A(new_n19839), .B(new_n19542), .Y(new_n19841));
  xnor_4 g17493(.A(new_n19815), .B(new_n19786), .Y(new_n19842));
  not_8  g17494(.A(new_n19842), .Y(new_n19843));
  and_5  g17495(.A(new_n19843), .B(new_n19546), .Y(new_n19844));
  xnor_4 g17496(.A(new_n19843), .B(new_n19546), .Y(new_n19845));
  xnor_4 g17497(.A(new_n19813), .B(new_n19789_1), .Y(new_n19846));
  nor_5  g17498(.A(new_n19846), .B(new_n19550), .Y(new_n19847));
  xnor_4 g17499(.A(new_n19846), .B(new_n19550), .Y(new_n19848));
  xnor_4 g17500(.A(new_n19811), .B(new_n19792_1), .Y(new_n19849));
  nor_5  g17501(.A(new_n19849), .B(new_n13432), .Y(new_n19850));
  xnor_4 g17502(.A(new_n19849), .B(new_n13432), .Y(new_n19851));
  xnor_4 g17503(.A(new_n19809), .B(new_n19795), .Y(new_n19852));
  nor_5  g17504(.A(new_n19852), .B(new_n13454), .Y(new_n19853));
  xnor_4 g17505(.A(new_n19852), .B(new_n13454), .Y(new_n19854));
  xnor_4 g17506(.A(new_n19807), .B(new_n19799), .Y(new_n19855));
  nor_5  g17507(.A(new_n19855), .B(new_n13458), .Y(new_n19856));
  xor_4  g17508(.A(new_n19855), .B(new_n13458), .Y(new_n19857));
  xor_4  g17509(.A(new_n19805), .B(new_n19803_1), .Y(new_n19858));
  nor_5  g17510(.A(new_n19858), .B(new_n13462), .Y(new_n19859));
  and_5  g17511(.A(new_n15356), .B(new_n13466), .Y(new_n19860));
  nor_5  g17512(.A(new_n15357), .B(new_n15346), .Y(new_n19861));
  nor_5  g17513(.A(new_n19861), .B(new_n19860), .Y(new_n19862));
  xor_4  g17514(.A(new_n19858), .B(new_n13462), .Y(new_n19863));
  and_5  g17515(.A(new_n19863), .B(new_n19862), .Y(new_n19864));
  nor_5  g17516(.A(new_n19864), .B(new_n19859), .Y(new_n19865));
  and_5  g17517(.A(new_n19865), .B(new_n19857), .Y(new_n19866));
  nor_5  g17518(.A(new_n19866), .B(new_n19856), .Y(new_n19867));
  nor_5  g17519(.A(new_n19867), .B(new_n19854), .Y(new_n19868));
  nor_5  g17520(.A(new_n19868), .B(new_n19853), .Y(new_n19869));
  nor_5  g17521(.A(new_n19869), .B(new_n19851), .Y(new_n19870));
  nor_5  g17522(.A(new_n19870), .B(new_n19850), .Y(new_n19871));
  nor_5  g17523(.A(new_n19871), .B(new_n19848), .Y(new_n19872));
  nor_5  g17524(.A(new_n19872), .B(new_n19847), .Y(new_n19873_1));
  nor_5  g17525(.A(new_n19873_1), .B(new_n19845), .Y(new_n19874));
  nor_5  g17526(.A(new_n19874), .B(new_n19844), .Y(new_n19875));
  nor_5  g17527(.A(new_n19875), .B(new_n19841), .Y(new_n19876));
  nor_5  g17528(.A(new_n19876), .B(new_n19840), .Y(new_n19877));
  nor_5  g17529(.A(new_n19877), .B(new_n19837), .Y(new_n19878));
  nor_5  g17530(.A(new_n19878), .B(new_n19836), .Y(new_n19879));
  xnor_4 g17531(.A(new_n19879), .B(new_n19834), .Y(n6707));
  xnor_4 g17532(.A(new_n12872), .B(new_n12645), .Y(n6736));
  xnor_4 g17533(.A(n23895), .B(n5101), .Y(new_n19882));
  and_5  g17534(.A(new_n5456), .B(n16507), .Y(new_n19883));
  xnor_4 g17535(.A(n17351), .B(n16507), .Y(new_n19884));
  and_5  g17536(.A(n22470), .B(new_n5459), .Y(new_n19885));
  xnor_4 g17537(.A(n22470), .B(n11736), .Y(new_n19886));
  and_5  g17538(.A(new_n5462), .B(n19116), .Y(new_n19887));
  and_5  g17539(.A(new_n5465), .B(n6861), .Y(new_n19888));
  and_5  g17540(.A(new_n17531), .B(new_n17514), .Y(new_n19889));
  or_5   g17541(.A(new_n19889), .B(new_n19888), .Y(new_n19890));
  xnor_4 g17542(.A(n23200), .B(n19116), .Y(new_n19891));
  and_5  g17543(.A(new_n19891), .B(new_n19890), .Y(new_n19892));
  or_5   g17544(.A(new_n19892), .B(new_n19887), .Y(new_n19893));
  and_5  g17545(.A(new_n19893), .B(new_n19886), .Y(new_n19894));
  or_5   g17546(.A(new_n19894), .B(new_n19885), .Y(new_n19895));
  and_5  g17547(.A(new_n19895), .B(new_n19884), .Y(new_n19896));
  or_5   g17548(.A(new_n19896), .B(new_n19883), .Y(new_n19897));
  xor_4  g17549(.A(new_n19897), .B(new_n19882), .Y(new_n19898));
  not_8  g17550(.A(new_n17539), .Y(new_n19899));
  nor_5  g17551(.A(new_n19899), .B(n22660), .Y(new_n19900));
  not_8  g17552(.A(new_n19900), .Y(new_n19901));
  nor_5  g17553(.A(new_n19901), .B(n13490), .Y(new_n19902));
  not_8  g17554(.A(new_n19902), .Y(new_n19903));
  nor_5  g17555(.A(new_n19903), .B(n9655), .Y(new_n19904));
  not_8  g17556(.A(new_n19904), .Y(new_n19905_1));
  nor_5  g17557(.A(new_n19905_1), .B(n25345), .Y(new_n19906));
  xnor_4 g17558(.A(new_n19906), .B(n13494), .Y(new_n19907));
  xnor_4 g17559(.A(new_n19907), .B(n12650), .Y(new_n19908));
  xnor_4 g17560(.A(new_n19904), .B(n25345), .Y(new_n19909_1));
  nor_5  g17561(.A(new_n19909_1), .B(new_n5560), .Y(new_n19910));
  xnor_4 g17562(.A(new_n19909_1), .B(n10201), .Y(new_n19911_1));
  xnor_4 g17563(.A(new_n19902), .B(n9655), .Y(new_n19912));
  nor_5  g17564(.A(new_n19912), .B(new_n5564_1), .Y(new_n19913));
  xnor_4 g17565(.A(new_n19912), .B(new_n5564_1), .Y(new_n19914));
  xnor_4 g17566(.A(new_n19900), .B(n13490), .Y(new_n19915));
  nor_5  g17567(.A(new_n19915), .B(new_n5568), .Y(new_n19916_1));
  xnor_4 g17568(.A(new_n19915), .B(n18290), .Y(new_n19917));
  nor_5  g17569(.A(new_n17540), .B(new_n5572), .Y(new_n19918));
  and_5  g17570(.A(new_n17562), .B(new_n17541), .Y(new_n19919));
  or_5   g17571(.A(new_n19919), .B(new_n19918), .Y(new_n19920));
  and_5  g17572(.A(new_n19920), .B(new_n19917), .Y(new_n19921));
  nor_5  g17573(.A(new_n19921), .B(new_n19916_1), .Y(new_n19922_1));
  nor_5  g17574(.A(new_n19922_1), .B(new_n19914), .Y(new_n19923_1));
  or_5   g17575(.A(new_n19923_1), .B(new_n19913), .Y(new_n19924));
  and_5  g17576(.A(new_n19924), .B(new_n19911_1), .Y(new_n19925));
  or_5   g17577(.A(new_n19925), .B(new_n19910), .Y(new_n19926));
  xor_4  g17578(.A(new_n19926), .B(new_n19908), .Y(new_n19927));
  xnor_4 g17579(.A(new_n19927), .B(new_n15563), .Y(new_n19928));
  xor_4  g17580(.A(new_n19924), .B(new_n19911_1), .Y(new_n19929));
  nor_5  g17581(.A(new_n19929), .B(new_n15567), .Y(new_n19930_1));
  xnor_4 g17582(.A(new_n19922_1), .B(new_n19914), .Y(new_n19931));
  nor_5  g17583(.A(new_n19931), .B(new_n15574), .Y(new_n19932));
  xnor_4 g17584(.A(new_n19931), .B(new_n15572), .Y(new_n19933));
  xor_4  g17585(.A(new_n19920), .B(new_n19917), .Y(new_n19934));
  nor_5  g17586(.A(new_n19934), .B(new_n15577), .Y(new_n19935));
  xnor_4 g17587(.A(new_n19934), .B(new_n15577), .Y(new_n19936));
  nor_5  g17588(.A(new_n17563), .B(new_n15581), .Y(new_n19937));
  nor_5  g17589(.A(new_n17587), .B(new_n17564), .Y(new_n19938));
  nor_5  g17590(.A(new_n19938), .B(new_n19937), .Y(new_n19939));
  nor_5  g17591(.A(new_n19939), .B(new_n19936), .Y(new_n19940));
  nor_5  g17592(.A(new_n19940), .B(new_n19935), .Y(new_n19941_1));
  and_5  g17593(.A(new_n19941_1), .B(new_n19933), .Y(new_n19942));
  nor_5  g17594(.A(new_n19942), .B(new_n19932), .Y(new_n19943));
  xnor_4 g17595(.A(new_n19929), .B(new_n15569), .Y(new_n19944));
  and_5  g17596(.A(new_n19944), .B(new_n19943), .Y(new_n19945));
  nor_5  g17597(.A(new_n19945), .B(new_n19930_1), .Y(new_n19946));
  xnor_4 g17598(.A(new_n19946), .B(new_n19928), .Y(new_n19947));
  xnor_4 g17599(.A(new_n19947), .B(new_n19898), .Y(new_n19948));
  xor_4  g17600(.A(new_n19895), .B(new_n19884), .Y(new_n19949));
  xor_4  g17601(.A(new_n19944), .B(new_n19943), .Y(new_n19950));
  nor_5  g17602(.A(new_n19950), .B(new_n19949), .Y(new_n19951));
  xnor_4 g17603(.A(new_n19950), .B(new_n19949), .Y(new_n19952));
  xor_4  g17604(.A(new_n19893), .B(new_n19886), .Y(new_n19953));
  xnor_4 g17605(.A(new_n19941_1), .B(new_n19933), .Y(new_n19954));
  nor_5  g17606(.A(new_n19954), .B(new_n19953), .Y(new_n19955));
  not_8  g17607(.A(new_n19954), .Y(new_n19956));
  xnor_4 g17608(.A(new_n19956), .B(new_n19953), .Y(new_n19957));
  xor_4  g17609(.A(new_n19891), .B(new_n19890), .Y(new_n19958));
  xnor_4 g17610(.A(new_n19939), .B(new_n19936), .Y(new_n19959));
  not_8  g17611(.A(new_n19959), .Y(new_n19960));
  and_5  g17612(.A(new_n19960), .B(new_n19958), .Y(new_n19961));
  xnor_4 g17613(.A(new_n19959), .B(new_n19958), .Y(new_n19962));
  not_8  g17614(.A(new_n17588), .Y(new_n19963));
  and_5  g17615(.A(new_n19963), .B(new_n17532), .Y(new_n19964));
  and_5  g17616(.A(new_n17621), .B(new_n17589), .Y(new_n19965));
  or_5   g17617(.A(new_n19965), .B(new_n19964), .Y(new_n19966));
  and_5  g17618(.A(new_n19966), .B(new_n19962), .Y(new_n19967));
  nor_5  g17619(.A(new_n19967), .B(new_n19961), .Y(new_n19968_1));
  and_5  g17620(.A(new_n19968_1), .B(new_n19957), .Y(new_n19969));
  nor_5  g17621(.A(new_n19969), .B(new_n19955), .Y(new_n19970));
  nor_5  g17622(.A(new_n19970), .B(new_n19952), .Y(new_n19971));
  nor_5  g17623(.A(new_n19971), .B(new_n19951), .Y(new_n19972));
  xor_4  g17624(.A(new_n19972), .B(new_n19948), .Y(n6791));
  xnor_4 g17625(.A(new_n3709), .B(new_n3700), .Y(n6802));
  xnor_4 g17626(.A(new_n15917_1), .B(new_n15894), .Y(n6826));
  xnor_4 g17627(.A(new_n9972), .B(new_n9945), .Y(n6835));
  nor_5  g17628(.A(new_n17829), .B(new_n10030), .Y(new_n19977));
  xnor_4 g17629(.A(new_n17831), .B(new_n10030), .Y(new_n19978));
  nor_5  g17630(.A(new_n2925), .B(new_n17810), .Y(new_n19979));
  xnor_4 g17631(.A(new_n2925), .B(n22379), .Y(new_n19980));
  nor_5  g17632(.A(new_n2972), .B(new_n2850), .Y(new_n19981));
  xnor_4 g17633(.A(new_n2976), .B(new_n2850), .Y(new_n19982));
  nor_5  g17634(.A(new_n2979_1), .B(new_n2853_1), .Y(new_n19983));
  xnor_4 g17635(.A(new_n2980), .B(new_n2853_1), .Y(new_n19984));
  nor_5  g17636(.A(new_n2985_1), .B(new_n2856), .Y(new_n19985));
  nor_5  g17637(.A(new_n2990), .B(n5213), .Y(new_n19986));
  xnor_4 g17638(.A(new_n2990), .B(new_n2859), .Y(new_n19987));
  nor_5  g17639(.A(new_n2996), .B(n4665), .Y(new_n19988_1));
  xnor_4 g17640(.A(new_n2996), .B(new_n2862), .Y(new_n19989));
  nor_5  g17641(.A(new_n3002), .B(new_n2866), .Y(new_n19990));
  xnor_4 g17642(.A(new_n3002), .B(n19005), .Y(new_n19991));
  nor_5  g17643(.A(new_n3063), .B(new_n5287), .Y(new_n19992));
  nor_5  g17644(.A(new_n19992), .B(n4326), .Y(new_n19993));
  xnor_4 g17645(.A(new_n19992), .B(new_n2869), .Y(new_n19994));
  and_5  g17646(.A(new_n19994), .B(new_n3008), .Y(new_n19995));
  nor_5  g17647(.A(new_n19995), .B(new_n19993), .Y(new_n19996));
  and_5  g17648(.A(new_n19996), .B(new_n19991), .Y(new_n19997));
  nor_5  g17649(.A(new_n19997), .B(new_n19990), .Y(new_n19998));
  and_5  g17650(.A(new_n19998), .B(new_n19989), .Y(new_n19999));
  or_5   g17651(.A(new_n19999), .B(new_n19988_1), .Y(new_n20000));
  and_5  g17652(.A(new_n20000), .B(new_n19987), .Y(new_n20001));
  nor_5  g17653(.A(new_n20001), .B(new_n19986), .Y(new_n20002));
  xnor_4 g17654(.A(new_n2986), .B(new_n2856), .Y(new_n20003));
  and_5  g17655(.A(new_n20003), .B(new_n20002), .Y(new_n20004_1));
  or_5   g17656(.A(new_n20004_1), .B(new_n19985), .Y(new_n20005));
  and_5  g17657(.A(new_n20005), .B(new_n19984), .Y(new_n20006));
  or_5   g17658(.A(new_n20006), .B(new_n19983), .Y(new_n20007));
  and_5  g17659(.A(new_n20007), .B(new_n19982), .Y(new_n20008));
  or_5   g17660(.A(new_n20008), .B(new_n19981), .Y(new_n20009));
  and_5  g17661(.A(new_n20009), .B(new_n19980), .Y(new_n20010));
  or_5   g17662(.A(new_n20010), .B(new_n19979), .Y(new_n20011));
  and_5  g17663(.A(new_n20011), .B(new_n19978), .Y(new_n20012));
  nor_5  g17664(.A(new_n20012), .B(new_n19977), .Y(new_n20013_1));
  nor_5  g17665(.A(new_n20013_1), .B(new_n17823), .Y(new_n20014));
  xnor_4 g17666(.A(new_n20014), .B(new_n17498), .Y(new_n20015));
  xnor_4 g17667(.A(new_n20013_1), .B(new_n17823), .Y(new_n20016));
  and_5  g17668(.A(new_n20016), .B(new_n17500_1), .Y(new_n20017_1));
  xnor_4 g17669(.A(new_n20016), .B(new_n17500_1), .Y(new_n20018));
  xor_4  g17670(.A(new_n20011), .B(new_n19978), .Y(new_n20019));
  nor_5  g17671(.A(new_n20019), .B(new_n12670_1), .Y(new_n20020));
  xnor_4 g17672(.A(new_n20019), .B(new_n12670_1), .Y(new_n20021));
  xor_4  g17673(.A(new_n20009), .B(new_n19980), .Y(new_n20022));
  nor_5  g17674(.A(new_n20022), .B(new_n12698), .Y(new_n20023));
  xnor_4 g17675(.A(new_n20022), .B(new_n12698), .Y(new_n20024));
  not_8  g17676(.A(new_n6097), .Y(new_n20025));
  xor_4  g17677(.A(new_n20007), .B(new_n19982), .Y(new_n20026));
  nor_5  g17678(.A(new_n20026), .B(new_n20025), .Y(new_n20027));
  xnor_4 g17679(.A(new_n20026), .B(new_n20025), .Y(new_n20028));
  xor_4  g17680(.A(new_n20005), .B(new_n19984), .Y(new_n20029));
  nor_5  g17681(.A(new_n20029), .B(new_n12704), .Y(new_n20030));
  xnor_4 g17682(.A(new_n20029), .B(new_n12704), .Y(new_n20031));
  not_8  g17683(.A(new_n6107), .Y(new_n20032));
  xor_4  g17684(.A(new_n20003), .B(new_n20002), .Y(new_n20033_1));
  nor_5  g17685(.A(new_n20033_1), .B(new_n20032), .Y(new_n20034));
  xnor_4 g17686(.A(new_n20033_1), .B(new_n20032), .Y(new_n20035));
  xor_4  g17687(.A(new_n20000), .B(new_n19987), .Y(new_n20036_1));
  and_5  g17688(.A(new_n20036_1), .B(new_n6112), .Y(new_n20037));
  xnor_4 g17689(.A(new_n20036_1), .B(new_n6112), .Y(new_n20038));
  xnor_4 g17690(.A(new_n19998), .B(new_n19989), .Y(new_n20039));
  not_8  g17691(.A(new_n20039), .Y(new_n20040_1));
  and_5  g17692(.A(new_n20040_1), .B(new_n6116), .Y(new_n20041));
  xnor_4 g17693(.A(new_n20040_1), .B(new_n6116), .Y(new_n20042));
  xor_4  g17694(.A(new_n19996), .B(new_n19991), .Y(new_n20043));
  nor_5  g17695(.A(new_n20043), .B(new_n6121), .Y(new_n20044));
  xnor_4 g17696(.A(new_n20043), .B(new_n6121), .Y(new_n20045));
  xnor_4 g17697(.A(new_n19994), .B(new_n3009), .Y(new_n20046));
  and_5  g17698(.A(new_n20046), .B(new_n6132), .Y(new_n20047));
  nor_5  g17699(.A(new_n5795), .B(new_n5794), .Y(new_n20048));
  xnor_4 g17700(.A(new_n20046), .B(new_n6126), .Y(new_n20049));
  and_5  g17701(.A(new_n20049), .B(new_n20048), .Y(new_n20050));
  nor_5  g17702(.A(new_n20050), .B(new_n20047), .Y(new_n20051));
  nor_5  g17703(.A(new_n20051), .B(new_n20045), .Y(new_n20052));
  nor_5  g17704(.A(new_n20052), .B(new_n20044), .Y(new_n20053));
  nor_5  g17705(.A(new_n20053), .B(new_n20042), .Y(new_n20054));
  nor_5  g17706(.A(new_n20054), .B(new_n20041), .Y(new_n20055));
  nor_5  g17707(.A(new_n20055), .B(new_n20038), .Y(new_n20056));
  nor_5  g17708(.A(new_n20056), .B(new_n20037), .Y(new_n20057));
  nor_5  g17709(.A(new_n20057), .B(new_n20035), .Y(new_n20058));
  nor_5  g17710(.A(new_n20058), .B(new_n20034), .Y(new_n20059));
  nor_5  g17711(.A(new_n20059), .B(new_n20031), .Y(new_n20060));
  nor_5  g17712(.A(new_n20060), .B(new_n20030), .Y(new_n20061_1));
  nor_5  g17713(.A(new_n20061_1), .B(new_n20028), .Y(new_n20062));
  nor_5  g17714(.A(new_n20062), .B(new_n20027), .Y(new_n20063));
  nor_5  g17715(.A(new_n20063), .B(new_n20024), .Y(new_n20064));
  nor_5  g17716(.A(new_n20064), .B(new_n20023), .Y(new_n20065));
  nor_5  g17717(.A(new_n20065), .B(new_n20021), .Y(new_n20066));
  nor_5  g17718(.A(new_n20066), .B(new_n20020), .Y(new_n20067));
  nor_5  g17719(.A(new_n20067), .B(new_n20018), .Y(new_n20068));
  nor_5  g17720(.A(new_n20068), .B(new_n20017_1), .Y(new_n20069_1));
  xnor_4 g17721(.A(new_n20069_1), .B(new_n20015), .Y(n6853));
  xnor_4 g17722(.A(new_n14607), .B(new_n11042), .Y(new_n20071));
  nor_5  g17723(.A(new_n14612), .B(new_n11048), .Y(new_n20072));
  xnor_4 g17724(.A(new_n14610), .B(new_n11048), .Y(new_n20073));
  nor_5  g17725(.A(new_n11050), .B(new_n4194), .Y(new_n20074));
  nor_5  g17726(.A(new_n12750), .B(new_n12737), .Y(new_n20075));
  nor_5  g17727(.A(new_n20075), .B(new_n20074), .Y(new_n20076));
  and_5  g17728(.A(new_n20076), .B(new_n20073), .Y(new_n20077_1));
  or_5   g17729(.A(new_n20077_1), .B(new_n20072), .Y(new_n20078));
  xor_4  g17730(.A(new_n20078), .B(new_n20071), .Y(n6862));
  and_5  g17731(.A(n22253), .B(new_n7110), .Y(new_n20080));
  and_5  g17732(.A(new_n15520), .B(new_n15505), .Y(new_n20081));
  nor_5  g17733(.A(new_n20081), .B(new_n20080), .Y(new_n20082));
  not_8  g17734(.A(n25296), .Y(new_n20083));
  nor_5  g17735(.A(new_n20083), .B(n23717), .Y(new_n20084));
  and_5  g17736(.A(new_n11202), .B(new_n11187), .Y(new_n20085));
  nor_5  g17737(.A(new_n20085), .B(new_n20084), .Y(new_n20086_1));
  nor_5  g17738(.A(new_n20086_1), .B(new_n17984), .Y(new_n20087));
  and_5  g17739(.A(new_n11203), .B(new_n11186), .Y(new_n20088));
  nor_5  g17740(.A(new_n11225), .B(new_n11204), .Y(new_n20089));
  nor_5  g17741(.A(new_n20089), .B(new_n20088), .Y(new_n20090));
  xnor_4 g17742(.A(new_n20086_1), .B(new_n17984), .Y(new_n20091));
  nor_5  g17743(.A(new_n20091), .B(new_n20090), .Y(new_n20092));
  nor_5  g17744(.A(new_n20092), .B(new_n20087), .Y(new_n20093));
  and_5  g17745(.A(new_n20093), .B(new_n20082), .Y(new_n20094));
  not_8  g17746(.A(new_n11226), .Y(new_n20095));
  and_5  g17747(.A(new_n15521), .B(new_n20095), .Y(new_n20096_1));
  and_5  g17748(.A(new_n15541), .B(new_n15522), .Y(new_n20097));
  nor_5  g17749(.A(new_n20097), .B(new_n20096_1), .Y(new_n20098));
  nor_5  g17750(.A(new_n20098), .B(new_n20093), .Y(new_n20099));
  nor_5  g17751(.A(new_n20099), .B(new_n20094), .Y(new_n20100));
  xnor_4 g17752(.A(new_n20091), .B(new_n20090), .Y(new_n20101));
  not_8  g17753(.A(new_n20101), .Y(new_n20102));
  nor_5  g17754(.A(new_n20102), .B(new_n20082), .Y(new_n20103_1));
  not_8  g17755(.A(new_n20098), .Y(new_n20104));
  nor_5  g17756(.A(new_n20101), .B(new_n20104), .Y(new_n20105));
  nor_5  g17757(.A(new_n20105), .B(new_n20103_1), .Y(new_n20106));
  and_5  g17758(.A(new_n20106), .B(new_n20100), .Y(n6863));
  xnor_4 g17759(.A(new_n6147), .B(new_n6094), .Y(n6867));
  xnor_4 g17760(.A(new_n17448), .B(new_n17440_1), .Y(n6965));
  xnor_4 g17761(.A(new_n7419), .B(new_n7379), .Y(n6967));
  xor_4  g17762(.A(new_n14160), .B(new_n14113), .Y(n6975));
  xor_4  g17763(.A(new_n19440), .B(new_n19439), .Y(n6983));
  xnor_4 g17764(.A(new_n14586), .B(new_n11028), .Y(new_n20113));
  nor_5  g17765(.A(new_n14592), .B(new_n11030), .Y(new_n20114));
  xnor_4 g17766(.A(new_n14591), .B(new_n11033), .Y(new_n20115));
  nor_5  g17767(.A(new_n14596), .B(new_n11035), .Y(new_n20116));
  xnor_4 g17768(.A(new_n14596), .B(new_n11037), .Y(new_n20117));
  not_8  g17769(.A(new_n11039), .Y(new_n20118));
  nor_5  g17770(.A(new_n14603_1), .B(new_n20118), .Y(new_n20119));
  nor_5  g17771(.A(new_n14607), .B(new_n11044_1), .Y(new_n20120));
  and_5  g17772(.A(new_n20078), .B(new_n20071), .Y(new_n20121));
  or_5   g17773(.A(new_n20121), .B(new_n20120), .Y(new_n20122));
  xnor_4 g17774(.A(new_n14600), .B(new_n20118), .Y(new_n20123));
  and_5  g17775(.A(new_n20123), .B(new_n20122), .Y(new_n20124));
  nor_5  g17776(.A(new_n20124), .B(new_n20119), .Y(new_n20125));
  and_5  g17777(.A(new_n20125), .B(new_n20117), .Y(new_n20126_1));
  nor_5  g17778(.A(new_n20126_1), .B(new_n20116), .Y(new_n20127));
  nor_5  g17779(.A(new_n20127), .B(new_n20115), .Y(new_n20128));
  nor_5  g17780(.A(new_n20128), .B(new_n20114), .Y(new_n20129));
  xnor_4 g17781(.A(new_n20129), .B(new_n20113), .Y(n6985));
  xnor_4 g17782(.A(new_n14407), .B(new_n14369), .Y(n6998));
  not_8  g17783(.A(new_n8886), .Y(new_n20132));
  xnor_4 g17784(.A(new_n10992), .B(new_n20132), .Y(n7032));
  xnor_4 g17785(.A(new_n19299), .B(new_n19267), .Y(n7038));
  xnor_4 g17786(.A(new_n17277), .B(new_n17276), .Y(n7079));
  xnor_4 g17787(.A(new_n7408_1), .B(new_n7407), .Y(n7190));
  xnor_4 g17788(.A(new_n15476), .B(new_n15473), .Y(n7229));
  xnor_4 g17789(.A(new_n8562), .B(new_n8550_1), .Y(n7230));
  xnor_4 g17790(.A(new_n18582_1), .B(new_n18581), .Y(n7233));
  xnor_4 g17791(.A(new_n12979), .B(new_n12971), .Y(n7236));
  xnor_4 g17792(.A(new_n15806), .B(new_n6946), .Y(n7253));
  and_5  g17793(.A(new_n18929), .B(new_n10870), .Y(new_n20142));
  nor_5  g17794(.A(new_n18930), .B(n12507), .Y(new_n20143));
  and_5  g17795(.A(new_n18930), .B(n12507), .Y(new_n20144));
  nor_5  g17796(.A(new_n18934), .B(new_n20144), .Y(new_n20145));
  nor_5  g17797(.A(new_n20145), .B(new_n20143), .Y(new_n20146));
  nor_5  g17798(.A(new_n20146), .B(new_n20142), .Y(new_n20147));
  not_8  g17799(.A(new_n19375), .Y(new_n20148));
  nor_5  g17800(.A(new_n20148), .B(new_n13859), .Y(new_n20149_1));
  xnor_4 g17801(.A(new_n20149_1), .B(new_n13823), .Y(new_n20150));
  nor_5  g17802(.A(new_n20150), .B(new_n10095), .Y(new_n20151_1));
  xnor_4 g17803(.A(new_n20150), .B(new_n10054), .Y(new_n20152));
  nor_5  g17804(.A(new_n19376), .B(new_n10058), .Y(new_n20153));
  and_5  g17805(.A(new_n19415), .B(new_n19377), .Y(new_n20154));
  or_5   g17806(.A(new_n20154), .B(new_n20153), .Y(new_n20155));
  and_5  g17807(.A(new_n20155), .B(new_n20152), .Y(new_n20156));
  nor_5  g17808(.A(new_n20156), .B(new_n20151_1), .Y(new_n20157));
  xor_4  g17809(.A(new_n13822), .B(new_n13810), .Y(new_n20158));
  and_5  g17810(.A(new_n20149_1), .B(new_n20158), .Y(new_n20159));
  nor_5  g17811(.A(new_n20159), .B(new_n13869), .Y(new_n20160));
  and_5  g17812(.A(new_n20159), .B(new_n13866), .Y(new_n20161));
  nor_5  g17813(.A(new_n20161), .B(new_n20160), .Y(new_n20162));
  xnor_4 g17814(.A(new_n20162), .B(new_n10044), .Y(new_n20163));
  xnor_4 g17815(.A(new_n20163), .B(new_n20157), .Y(new_n20164));
  nor_5  g17816(.A(new_n20164), .B(new_n20147), .Y(new_n20165));
  not_8  g17817(.A(new_n20147), .Y(new_n20166));
  xnor_4 g17818(.A(new_n20164), .B(new_n20166), .Y(new_n20167));
  xor_4  g17819(.A(new_n20155), .B(new_n20152), .Y(new_n20168));
  nor_5  g17820(.A(new_n20168), .B(new_n18935), .Y(new_n20169_1));
  nor_5  g17821(.A(new_n19416), .B(new_n16280), .Y(new_n20170));
  and_5  g17822(.A(new_n19455), .B(new_n19417), .Y(new_n20171));
  nor_5  g17823(.A(new_n20171), .B(new_n20170), .Y(new_n20172));
  xnor_4 g17824(.A(new_n20168), .B(new_n18935), .Y(new_n20173));
  nor_5  g17825(.A(new_n20173), .B(new_n20172), .Y(new_n20174));
  nor_5  g17826(.A(new_n20174), .B(new_n20169_1), .Y(new_n20175));
  and_5  g17827(.A(new_n20175), .B(new_n20167), .Y(new_n20176));
  nor_5  g17828(.A(new_n20176), .B(new_n20165), .Y(new_n20177));
  not_8  g17829(.A(new_n20177), .Y(new_n20178));
  and_5  g17830(.A(new_n20162), .B(new_n10044), .Y(new_n20179_1));
  or_5   g17831(.A(new_n20162), .B(new_n10044), .Y(new_n20180));
  and_5  g17832(.A(new_n20180), .B(new_n20157), .Y(new_n20181));
  or_5   g17833(.A(new_n20181), .B(new_n20161), .Y(new_n20182));
  nor_5  g17834(.A(new_n20182), .B(new_n20179_1), .Y(new_n20183));
  xnor_4 g17835(.A(new_n20183), .B(new_n20178), .Y(n7256));
  not_8  g17836(.A(new_n15180_1), .Y(new_n20185));
  nor_5  g17837(.A(new_n12048), .B(n2416), .Y(new_n20186));
  xnor_4 g17838(.A(n22764), .B(n2416), .Y(new_n20187_1));
  not_8  g17839(.A(n26264), .Y(new_n20188));
  nor_5  g17840(.A(new_n20188), .B(n21905), .Y(new_n20189));
  and_5  g17841(.A(new_n19029), .B(new_n19015), .Y(new_n20190));
  or_5   g17842(.A(new_n20190), .B(new_n20189), .Y(new_n20191));
  and_5  g17843(.A(new_n20191), .B(new_n20187_1), .Y(new_n20192));
  nor_5  g17844(.A(new_n20192), .B(new_n20186), .Y(new_n20193));
  xor_4  g17845(.A(new_n20191), .B(new_n20187_1), .Y(new_n20194));
  and_5  g17846(.A(new_n20194), .B(new_n15184), .Y(new_n20195));
  xnor_4 g17847(.A(new_n20194), .B(new_n15182_1), .Y(new_n20196));
  and_5  g17848(.A(new_n19030), .B(new_n15189), .Y(new_n20197));
  and_5  g17849(.A(new_n19044_1), .B(new_n19031), .Y(new_n20198));
  or_5   g17850(.A(new_n20198), .B(new_n20197), .Y(new_n20199));
  and_5  g17851(.A(new_n20199), .B(new_n20196), .Y(new_n20200));
  nor_5  g17852(.A(new_n20200), .B(new_n20195), .Y(new_n20201));
  xnor_4 g17853(.A(new_n20201), .B(new_n20193), .Y(new_n20202));
  xnor_4 g17854(.A(new_n20202), .B(new_n20185), .Y(new_n20203));
  xnor_4 g17855(.A(new_n20203), .B(new_n19127), .Y(new_n20204));
  xor_4  g17856(.A(new_n20199), .B(new_n20196), .Y(new_n20205));
  nor_5  g17857(.A(new_n20205), .B(new_n19139), .Y(new_n20206));
  xnor_4 g17858(.A(new_n20205), .B(new_n19139), .Y(new_n20207));
  nor_5  g17859(.A(new_n19045), .B(new_n19014), .Y(new_n20208));
  nor_5  g17860(.A(new_n19059), .B(new_n19046), .Y(new_n20209));
  nor_5  g17861(.A(new_n20209), .B(new_n20208), .Y(new_n20210));
  nor_5  g17862(.A(new_n20210), .B(new_n20207), .Y(new_n20211));
  nor_5  g17863(.A(new_n20211), .B(new_n20206), .Y(new_n20212));
  xnor_4 g17864(.A(new_n20212), .B(new_n20204), .Y(n7268));
  not_8  g17865(.A(new_n10789), .Y(new_n20214));
  nor_5  g17866(.A(new_n20214), .B(n752), .Y(new_n20215));
  not_8  g17867(.A(new_n20215), .Y(new_n20216));
  nor_5  g17868(.A(new_n20216), .B(n2175), .Y(new_n20217));
  not_8  g17869(.A(new_n20217), .Y(new_n20218));
  nor_5  g17870(.A(new_n20218), .B(n13026), .Y(new_n20219));
  not_8  g17871(.A(new_n20219), .Y(new_n20220));
  nor_5  g17872(.A(new_n20220), .B(n23912), .Y(new_n20221));
  not_8  g17873(.A(n10514), .Y(new_n20222));
  xnor_4 g17874(.A(new_n20219), .B(n23912), .Y(new_n20223));
  nor_5  g17875(.A(new_n20223), .B(new_n20222), .Y(new_n20224));
  not_8  g17876(.A(new_n20223), .Y(new_n20225));
  xnor_4 g17877(.A(new_n20225), .B(new_n20222), .Y(new_n20226));
  xnor_4 g17878(.A(new_n20217), .B(n13026), .Y(new_n20227));
  nor_5  g17879(.A(new_n20227), .B(new_n11276), .Y(new_n20228));
  not_8  g17880(.A(new_n20227), .Y(new_n20229));
  xnor_4 g17881(.A(new_n20229), .B(new_n11276), .Y(new_n20230));
  xnor_4 g17882(.A(new_n20215), .B(n2175), .Y(new_n20231));
  nor_5  g17883(.A(new_n20231), .B(new_n11389), .Y(new_n20232));
  not_8  g17884(.A(new_n20231), .Y(new_n20233));
  xnor_4 g17885(.A(new_n20233), .B(new_n11389), .Y(new_n20234));
  nor_5  g17886(.A(new_n10790), .B(new_n10824), .Y(new_n20235_1));
  xnor_4 g17887(.A(new_n10790), .B(n20470), .Y(new_n20236));
  nor_5  g17888(.A(new_n10792_1), .B(new_n10837), .Y(new_n20237));
  xnor_4 g17889(.A(new_n10792_1), .B(n21222), .Y(new_n20238));
  not_8  g17890(.A(n9832), .Y(new_n20239));
  nor_5  g17891(.A(new_n10795), .B(new_n20239), .Y(new_n20240));
  xnor_4 g17892(.A(new_n10795), .B(n9832), .Y(new_n20241));
  nor_5  g17893(.A(new_n10798), .B(new_n9479), .Y(new_n20242));
  xnor_4 g17894(.A(new_n10798), .B(n1558), .Y(new_n20243));
  xnor_4 g17895(.A(new_n10782), .B(n5131), .Y(new_n20244));
  and_5  g17896(.A(new_n20244), .B(n21749), .Y(new_n20245));
  xnor_4 g17897(.A(new_n10800), .B(n21749), .Y(new_n20246));
  nor_5  g17898(.A(new_n10806), .B(new_n9487), .Y(new_n20247));
  nor_5  g17899(.A(new_n9485), .B(n15506), .Y(new_n20248));
  xnor_4 g17900(.A(new_n10805), .B(new_n9487), .Y(new_n20249));
  and_5  g17901(.A(new_n20249), .B(new_n20248), .Y(new_n20250_1));
  or_5   g17902(.A(new_n20250_1), .B(new_n20247), .Y(new_n20251));
  and_5  g17903(.A(new_n20251), .B(new_n20246), .Y(new_n20252));
  or_5   g17904(.A(new_n20252), .B(new_n20245), .Y(new_n20253));
  and_5  g17905(.A(new_n20253), .B(new_n20243), .Y(new_n20254));
  or_5   g17906(.A(new_n20254), .B(new_n20242), .Y(new_n20255));
  and_5  g17907(.A(new_n20255), .B(new_n20241), .Y(new_n20256));
  or_5   g17908(.A(new_n20256), .B(new_n20240), .Y(new_n20257));
  and_5  g17909(.A(new_n20257), .B(new_n20238), .Y(new_n20258));
  or_5   g17910(.A(new_n20258), .B(new_n20237), .Y(new_n20259_1));
  and_5  g17911(.A(new_n20259_1), .B(new_n20236), .Y(new_n20260));
  or_5   g17912(.A(new_n20260), .B(new_n20235_1), .Y(new_n20261));
  and_5  g17913(.A(new_n20261), .B(new_n20234), .Y(new_n20262));
  or_5   g17914(.A(new_n20262), .B(new_n20232), .Y(new_n20263));
  and_5  g17915(.A(new_n20263), .B(new_n20230), .Y(new_n20264));
  or_5   g17916(.A(new_n20264), .B(new_n20228), .Y(new_n20265));
  and_5  g17917(.A(new_n20265), .B(new_n20226), .Y(new_n20266));
  nor_5  g17918(.A(new_n20266), .B(new_n20224), .Y(new_n20267));
  and_5  g17919(.A(new_n20267), .B(new_n20221), .Y(new_n20268));
  xor_4  g17920(.A(new_n20265), .B(new_n20226), .Y(new_n20269));
  nor_5  g17921(.A(new_n20269), .B(n9872), .Y(new_n20270));
  not_8  g17922(.A(n9872), .Y(new_n20271));
  xnor_4 g17923(.A(new_n20269), .B(new_n20271), .Y(new_n20272));
  xor_4  g17924(.A(new_n20263), .B(new_n20230), .Y(new_n20273));
  nor_5  g17925(.A(new_n20273), .B(n5842), .Y(new_n20274));
  not_8  g17926(.A(n5842), .Y(new_n20275));
  xnor_4 g17927(.A(new_n20273), .B(new_n20275), .Y(new_n20276));
  xor_4  g17928(.A(new_n20261), .B(new_n20234), .Y(new_n20277));
  nor_5  g17929(.A(new_n20277), .B(n6379), .Y(new_n20278));
  not_8  g17930(.A(n6379), .Y(new_n20279_1));
  xnor_4 g17931(.A(new_n20277), .B(new_n20279_1), .Y(new_n20280));
  xor_4  g17932(.A(new_n20259_1), .B(new_n20236), .Y(new_n20281));
  nor_5  g17933(.A(new_n20281), .B(n2102), .Y(new_n20282));
  not_8  g17934(.A(n2102), .Y(new_n20283));
  xnor_4 g17935(.A(new_n20281), .B(new_n20283), .Y(new_n20284));
  xor_4  g17936(.A(new_n20257), .B(new_n20238), .Y(new_n20285));
  nor_5  g17937(.A(new_n20285), .B(n17954), .Y(new_n20286));
  xor_4  g17938(.A(new_n20255), .B(new_n20241), .Y(new_n20287_1));
  nor_5  g17939(.A(new_n20287_1), .B(n8256), .Y(new_n20288));
  not_8  g17940(.A(n8256), .Y(new_n20289));
  xnor_4 g17941(.A(new_n20287_1), .B(new_n20289), .Y(new_n20290));
  xor_4  g17942(.A(new_n20253), .B(new_n20243), .Y(new_n20291));
  nor_5  g17943(.A(new_n20291), .B(n24150), .Y(new_n20292));
  not_8  g17944(.A(n24150), .Y(new_n20293));
  xnor_4 g17945(.A(new_n20291), .B(new_n20293), .Y(new_n20294));
  xor_4  g17946(.A(new_n20251), .B(new_n20246), .Y(new_n20295));
  nor_5  g17947(.A(new_n20295), .B(n19584), .Y(new_n20296));
  not_8  g17948(.A(n19584), .Y(new_n20297));
  xnor_4 g17949(.A(new_n20295), .B(new_n20297), .Y(new_n20298));
  not_8  g17950(.A(n5060), .Y(new_n20299));
  xnor_4 g17951(.A(new_n20249), .B(new_n20248), .Y(new_n20300));
  nor_5  g17952(.A(new_n20300), .B(new_n20299), .Y(new_n20301_1));
  not_8  g17953(.A(new_n20300), .Y(new_n20302));
  or_5   g17954(.A(new_n20302), .B(n5060), .Y(new_n20303));
  xnor_4 g17955(.A(n21138), .B(n15506), .Y(new_n20304));
  and_5  g17956(.A(new_n20304), .B(n15332), .Y(new_n20305));
  and_5  g17957(.A(new_n20305), .B(new_n20303), .Y(new_n20306));
  nor_5  g17958(.A(new_n20306), .B(new_n20301_1), .Y(new_n20307));
  and_5  g17959(.A(new_n20307), .B(new_n20298), .Y(new_n20308));
  or_5   g17960(.A(new_n20308), .B(new_n20296), .Y(new_n20309));
  and_5  g17961(.A(new_n20309), .B(new_n20294), .Y(new_n20310));
  or_5   g17962(.A(new_n20310), .B(new_n20292), .Y(new_n20311));
  and_5  g17963(.A(new_n20311), .B(new_n20290), .Y(new_n20312));
  or_5   g17964(.A(new_n20312), .B(new_n20288), .Y(new_n20313));
  not_8  g17965(.A(n17954), .Y(new_n20314));
  xnor_4 g17966(.A(new_n20285), .B(new_n20314), .Y(new_n20315));
  and_5  g17967(.A(new_n20315), .B(new_n20313), .Y(new_n20316));
  or_5   g17968(.A(new_n20316), .B(new_n20286), .Y(new_n20317));
  and_5  g17969(.A(new_n20317), .B(new_n20284), .Y(new_n20318));
  or_5   g17970(.A(new_n20318), .B(new_n20282), .Y(new_n20319));
  and_5  g17971(.A(new_n20319), .B(new_n20280), .Y(new_n20320));
  or_5   g17972(.A(new_n20320), .B(new_n20278), .Y(new_n20321));
  and_5  g17973(.A(new_n20321), .B(new_n20276), .Y(new_n20322));
  or_5   g17974(.A(new_n20322), .B(new_n20274), .Y(new_n20323));
  and_5  g17975(.A(new_n20323), .B(new_n20272), .Y(new_n20324));
  nor_5  g17976(.A(new_n20324), .B(new_n20270), .Y(new_n20325));
  not_8  g17977(.A(new_n20325), .Y(new_n20326));
  and_5  g17978(.A(new_n20326), .B(new_n20268), .Y(new_n20327));
  or_5   g17979(.A(new_n20267), .B(new_n20221), .Y(new_n20328));
  nor_5  g17980(.A(new_n20328), .B(new_n20326), .Y(new_n20329));
  nor_5  g17981(.A(new_n20329), .B(new_n20327), .Y(new_n20330_1));
  xnor_4 g17982(.A(new_n20330_1), .B(new_n14356), .Y(new_n20331));
  not_8  g17983(.A(new_n20221), .Y(new_n20332));
  xnor_4 g17984(.A(new_n20267), .B(new_n20332), .Y(new_n20333_1));
  xnor_4 g17985(.A(new_n20333_1), .B(new_n20326), .Y(new_n20334));
  nor_5  g17986(.A(new_n20334), .B(new_n14361), .Y(new_n20335));
  xnor_4 g17987(.A(new_n20334), .B(new_n14361), .Y(new_n20336));
  xor_4  g17988(.A(new_n20323), .B(new_n20272), .Y(new_n20337));
  nor_5  g17989(.A(new_n20337), .B(new_n2655), .Y(new_n20338));
  xnor_4 g17990(.A(new_n20337), .B(new_n2655), .Y(new_n20339));
  xor_4  g17991(.A(new_n20321), .B(new_n20276), .Y(new_n20340));
  nor_5  g17992(.A(new_n20340), .B(new_n2786), .Y(new_n20341));
  xor_4  g17993(.A(new_n20319), .B(new_n20280), .Y(new_n20342));
  nor_5  g17994(.A(new_n20342), .B(new_n2792), .Y(new_n20343));
  xnor_4 g17995(.A(new_n20342), .B(new_n2792), .Y(new_n20344));
  xor_4  g17996(.A(new_n20317), .B(new_n20284), .Y(new_n20345));
  nor_5  g17997(.A(new_n20345), .B(new_n2797), .Y(new_n20346));
  xnor_4 g17998(.A(new_n20345), .B(new_n2797), .Y(new_n20347));
  xor_4  g17999(.A(new_n20315), .B(new_n20313), .Y(new_n20348));
  nor_5  g18000(.A(new_n20348), .B(new_n2801), .Y(new_n20349_1));
  xnor_4 g18001(.A(new_n20348), .B(new_n2801), .Y(new_n20350));
  not_8  g18002(.A(new_n2806), .Y(new_n20351));
  xor_4  g18003(.A(new_n20311), .B(new_n20290), .Y(new_n20352));
  nor_5  g18004(.A(new_n20352), .B(new_n20351), .Y(new_n20353));
  xnor_4 g18005(.A(new_n20352), .B(new_n20351), .Y(new_n20354));
  xor_4  g18006(.A(new_n20309), .B(new_n20294), .Y(new_n20355_1));
  nor_5  g18007(.A(new_n20355_1), .B(new_n2812), .Y(new_n20356));
  xnor_4 g18008(.A(new_n20355_1), .B(new_n2812), .Y(new_n20357));
  xor_4  g18009(.A(new_n20307), .B(new_n20298), .Y(new_n20358));
  nor_5  g18010(.A(new_n20358), .B(new_n2818), .Y(new_n20359_1));
  xnor_4 g18011(.A(new_n20358), .B(new_n2818), .Y(new_n20360));
  xnor_4 g18012(.A(new_n20302), .B(new_n20299), .Y(new_n20361));
  xnor_4 g18013(.A(new_n20361), .B(new_n20305), .Y(new_n20362));
  nor_5  g18014(.A(new_n20362), .B(new_n2824), .Y(new_n20363));
  xnor_4 g18015(.A(new_n20304), .B(new_n16103), .Y(new_n20364));
  nor_5  g18016(.A(new_n20364), .B(new_n2827), .Y(new_n20365));
  xnor_4 g18017(.A(new_n20362), .B(new_n2824), .Y(new_n20366_1));
  nor_5  g18018(.A(new_n20366_1), .B(new_n20365), .Y(new_n20367));
  nor_5  g18019(.A(new_n20367), .B(new_n20363), .Y(new_n20368));
  nor_5  g18020(.A(new_n20368), .B(new_n20360), .Y(new_n20369));
  nor_5  g18021(.A(new_n20369), .B(new_n20359_1), .Y(new_n20370));
  nor_5  g18022(.A(new_n20370), .B(new_n20357), .Y(new_n20371));
  nor_5  g18023(.A(new_n20371), .B(new_n20356), .Y(new_n20372));
  nor_5  g18024(.A(new_n20372), .B(new_n20354), .Y(new_n20373));
  nor_5  g18025(.A(new_n20373), .B(new_n20353), .Y(new_n20374));
  nor_5  g18026(.A(new_n20374), .B(new_n20350), .Y(new_n20375));
  nor_5  g18027(.A(new_n20375), .B(new_n20349_1), .Y(new_n20376));
  nor_5  g18028(.A(new_n20376), .B(new_n20347), .Y(new_n20377));
  nor_5  g18029(.A(new_n20377), .B(new_n20346), .Y(new_n20378));
  nor_5  g18030(.A(new_n20378), .B(new_n20344), .Y(new_n20379));
  nor_5  g18031(.A(new_n20379), .B(new_n20343), .Y(new_n20380));
  xnor_4 g18032(.A(new_n20340), .B(new_n2786), .Y(new_n20381));
  nor_5  g18033(.A(new_n20381), .B(new_n20380), .Y(new_n20382));
  nor_5  g18034(.A(new_n20382), .B(new_n20341), .Y(new_n20383));
  nor_5  g18035(.A(new_n20383), .B(new_n20339), .Y(new_n20384));
  nor_5  g18036(.A(new_n20384), .B(new_n20338), .Y(new_n20385_1));
  nor_5  g18037(.A(new_n20385_1), .B(new_n20336), .Y(new_n20386));
  nor_5  g18038(.A(new_n20386), .B(new_n20335), .Y(new_n20387));
  xnor_4 g18039(.A(new_n20387), .B(new_n20331), .Y(n7277));
  xor_4  g18040(.A(new_n13133), .B(new_n13126), .Y(n7280));
  xnor_4 g18041(.A(new_n5753), .B(new_n5728), .Y(n7298));
  xnor_4 g18042(.A(new_n18919_1), .B(new_n18910), .Y(n7308));
  xnor_4 g18043(.A(new_n19135), .B(new_n7242), .Y(new_n20392));
  nor_5  g18044(.A(new_n19141_1), .B(new_n7266), .Y(new_n20393));
  xnor_4 g18045(.A(new_n19138), .B(new_n7266), .Y(new_n20394));
  nor_5  g18046(.A(new_n14653), .B(new_n14628), .Y(new_n20395));
  nor_5  g18047(.A(new_n14680_1), .B(new_n14654), .Y(new_n20396));
  or_5   g18048(.A(new_n20396), .B(new_n20395), .Y(new_n20397));
  and_5  g18049(.A(new_n20397), .B(new_n20394), .Y(new_n20398));
  nor_5  g18050(.A(new_n20398), .B(new_n20393), .Y(new_n20399));
  xnor_4 g18051(.A(new_n20399), .B(new_n20392), .Y(new_n20400));
  not_8  g18052(.A(new_n20400), .Y(new_n20401));
  xnor_4 g18053(.A(new_n20401), .B(new_n19163_1), .Y(new_n20402_1));
  xor_4  g18054(.A(new_n20397), .B(new_n20394), .Y(new_n20403_1));
  nor_5  g18055(.A(new_n20403_1), .B(new_n19169), .Y(new_n20404));
  and_5  g18056(.A(new_n18560), .B(new_n14682), .Y(new_n20405));
  and_5  g18057(.A(new_n18590), .B(new_n18561), .Y(new_n20406));
  nor_5  g18058(.A(new_n20406), .B(new_n20405), .Y(new_n20407));
  xnor_4 g18059(.A(new_n20403_1), .B(new_n19169), .Y(new_n20408));
  not_8  g18060(.A(new_n20408), .Y(new_n20409_1));
  and_5  g18061(.A(new_n20409_1), .B(new_n20407), .Y(new_n20410));
  nor_5  g18062(.A(new_n20410), .B(new_n20404), .Y(new_n20411_1));
  xnor_4 g18063(.A(new_n20411_1), .B(new_n20402_1), .Y(n7313));
  xnor_4 g18064(.A(new_n3713), .B(new_n3689), .Y(n7346));
  xnor_4 g18065(.A(new_n20086_1), .B(new_n13735), .Y(new_n20414));
  nor_5  g18066(.A(new_n20086_1), .B(new_n13739), .Y(new_n20415));
  xnor_4 g18067(.A(new_n20086_1), .B(new_n13739), .Y(new_n20416));
  nor_5  g18068(.A(new_n13743), .B(new_n11203), .Y(new_n20417));
  xnor_4 g18069(.A(new_n13743), .B(new_n11203), .Y(new_n20418));
  nor_5  g18070(.A(new_n13747), .B(new_n11206), .Y(new_n20419));
  xnor_4 g18071(.A(new_n13747), .B(new_n11206), .Y(new_n20420));
  nor_5  g18072(.A(new_n13752), .B(new_n11210), .Y(new_n20421));
  nor_5  g18073(.A(new_n6551), .B(new_n6431_1), .Y(new_n20422));
  and_5  g18074(.A(new_n6583), .B(new_n6553), .Y(new_n20423));
  nor_5  g18075(.A(new_n20423), .B(new_n20422), .Y(new_n20424_1));
  xnor_4 g18076(.A(new_n13751), .B(new_n11210), .Y(new_n20425));
  and_5  g18077(.A(new_n20425), .B(new_n20424_1), .Y(new_n20426));
  nor_5  g18078(.A(new_n20426), .B(new_n20421), .Y(new_n20427));
  nor_5  g18079(.A(new_n20427), .B(new_n20420), .Y(new_n20428));
  nor_5  g18080(.A(new_n20428), .B(new_n20419), .Y(new_n20429_1));
  nor_5  g18081(.A(new_n20429_1), .B(new_n20418), .Y(new_n20430));
  nor_5  g18082(.A(new_n20430), .B(new_n20417), .Y(new_n20431));
  nor_5  g18083(.A(new_n20431), .B(new_n20416), .Y(new_n20432));
  nor_5  g18084(.A(new_n20432), .B(new_n20415), .Y(new_n20433));
  xor_4  g18085(.A(new_n20433), .B(new_n20414), .Y(n7349));
  xnor_4 g18086(.A(new_n20383), .B(new_n20339), .Y(n7363));
  nor_5  g18087(.A(n21839), .B(new_n8954), .Y(new_n20436_1));
  and_5  g18088(.A(new_n19113), .B(new_n19110), .Y(new_n20437));
  nor_5  g18089(.A(new_n20437), .B(new_n20436_1), .Y(new_n20438));
  xnor_4 g18090(.A(new_n20438), .B(new_n10099), .Y(new_n20439));
  nor_5  g18091(.A(new_n19114), .B(new_n10102), .Y(new_n20440));
  nor_5  g18092(.A(new_n19118), .B(new_n19115), .Y(new_n20441_1));
  nor_5  g18093(.A(new_n20441_1), .B(new_n20440), .Y(new_n20442));
  xnor_4 g18094(.A(new_n20442), .B(new_n20439), .Y(n7390));
  xnor_4 g18095(.A(new_n9045), .B(new_n9044), .Y(n7403));
  xnor_4 g18096(.A(new_n9219), .B(new_n9182_1), .Y(n7408));
  xnor_4 g18097(.A(new_n19449), .B(new_n19426), .Y(n7432));
  nor_5  g18098(.A(new_n17497), .B(new_n15098), .Y(new_n20447));
  nor_5  g18099(.A(new_n17507), .B(new_n17499), .Y(new_n20448));
  or_5   g18100(.A(new_n20448), .B(new_n20447), .Y(n7475));
  xnor_4 g18101(.A(new_n5209), .B(new_n5208), .Y(n7477));
  xnor_4 g18102(.A(new_n8899), .B(new_n8874), .Y(n7507));
  nor_5  g18103(.A(new_n11803), .B(new_n5453), .Y(new_n20452));
  xnor_4 g18104(.A(new_n11802), .B(new_n5453), .Y(new_n20453));
  nor_5  g18105(.A(new_n6863_1), .B(new_n5456), .Y(new_n20454));
  and_5  g18106(.A(new_n6908), .B(new_n6865), .Y(new_n20455_1));
  or_5   g18107(.A(new_n20455_1), .B(new_n20454), .Y(new_n20456));
  and_5  g18108(.A(new_n20456), .B(new_n20453), .Y(new_n20457));
  nor_5  g18109(.A(new_n20457), .B(new_n20452), .Y(new_n20458));
  xnor_4 g18110(.A(new_n20458), .B(new_n11851), .Y(new_n20459));
  xnor_4 g18111(.A(new_n20459), .B(new_n16853), .Y(new_n20460));
  xor_4  g18112(.A(new_n20456), .B(new_n20453), .Y(new_n20461));
  nor_5  g18113(.A(new_n20461), .B(new_n16857), .Y(new_n20462));
  xnor_4 g18114(.A(new_n20461), .B(new_n16857), .Y(new_n20463));
  nor_5  g18115(.A(new_n6909), .B(new_n6833), .Y(new_n20464));
  nor_5  g18116(.A(new_n6964), .B(new_n6910), .Y(new_n20465));
  nor_5  g18117(.A(new_n20465), .B(new_n20464), .Y(new_n20466));
  nor_5  g18118(.A(new_n20466), .B(new_n20463), .Y(new_n20467));
  nor_5  g18119(.A(new_n20467), .B(new_n20462), .Y(new_n20468));
  xnor_4 g18120(.A(new_n20468), .B(new_n20460), .Y(n7514));
  xnor_4 g18121(.A(new_n10767), .B(new_n10744), .Y(n7558));
  xnor_4 g18122(.A(new_n11886), .B(new_n11885), .Y(n7572));
  xnor_4 g18123(.A(new_n6274), .B(new_n4015), .Y(new_n20472));
  nor_5  g18124(.A(new_n6276_1), .B(new_n4021), .Y(new_n20473));
  and_5  g18125(.A(new_n19479), .B(new_n19470), .Y(new_n20474));
  or_5   g18126(.A(new_n20474), .B(new_n20473), .Y(new_n20475));
  xor_4  g18127(.A(new_n20475), .B(new_n20472), .Y(new_n20476));
  xnor_4 g18128(.A(new_n20476), .B(new_n9668), .Y(new_n20477));
  nor_5  g18129(.A(new_n19480), .B(new_n9673), .Y(new_n20478_1));
  nor_5  g18130(.A(new_n19492), .B(new_n19481), .Y(new_n20479));
  nor_5  g18131(.A(new_n20479), .B(new_n20478_1), .Y(new_n20480));
  xnor_4 g18132(.A(new_n20480), .B(new_n20477), .Y(n7575));
  xnor_4 g18133(.A(new_n20229), .B(new_n9600), .Y(new_n20482));
  nor_5  g18134(.A(new_n20233), .B(new_n9652), .Y(new_n20483));
  xnor_4 g18135(.A(new_n20233), .B(new_n9652), .Y(new_n20484));
  and_5  g18136(.A(new_n10790), .B(new_n9657), .Y(new_n20485));
  and_5  g18137(.A(new_n10822), .B(new_n10791), .Y(new_n20486));
  nor_5  g18138(.A(new_n20486), .B(new_n20485), .Y(new_n20487));
  nor_5  g18139(.A(new_n20487), .B(new_n20484), .Y(new_n20488));
  nor_5  g18140(.A(new_n20488), .B(new_n20483), .Y(new_n20489_1));
  xnor_4 g18141(.A(new_n20489_1), .B(new_n20482), .Y(new_n20490_1));
  xnor_4 g18142(.A(new_n20490_1), .B(new_n11384), .Y(new_n20491));
  xnor_4 g18143(.A(new_n20487), .B(new_n20484), .Y(new_n20492));
  nor_5  g18144(.A(new_n20492), .B(new_n11392), .Y(new_n20493));
  xnor_4 g18145(.A(new_n20492), .B(new_n11392), .Y(new_n20494));
  nor_5  g18146(.A(new_n10834_1), .B(new_n10823), .Y(new_n20495_1));
  nor_5  g18147(.A(new_n10868), .B(new_n10835), .Y(new_n20496));
  or_5   g18148(.A(new_n20496), .B(new_n20495_1), .Y(new_n20497));
  nor_5  g18149(.A(new_n20497), .B(new_n20494), .Y(new_n20498));
  nor_5  g18150(.A(new_n20498), .B(new_n20493), .Y(new_n20499));
  xor_4  g18151(.A(new_n20499), .B(new_n20491), .Y(n7585));
  not_8  g18152(.A(new_n19947), .Y(new_n20501));
  xnor_4 g18153(.A(new_n20501), .B(new_n7698_1), .Y(new_n20502));
  nor_5  g18154(.A(new_n19950), .B(new_n7705), .Y(new_n20503));
  xnor_4 g18155(.A(new_n19950), .B(new_n7705), .Y(new_n20504));
  nor_5  g18156(.A(new_n19954), .B(new_n7710), .Y(new_n20505));
  xnor_4 g18157(.A(new_n19956), .B(new_n7714), .Y(new_n20506));
  nor_5  g18158(.A(new_n19960), .B(new_n7717), .Y(new_n20507));
  xnor_4 g18159(.A(new_n19960), .B(new_n7717), .Y(new_n20508));
  nor_5  g18160(.A(new_n19963), .B(new_n7721_1), .Y(new_n20509));
  xnor_4 g18161(.A(new_n19963), .B(new_n7721_1), .Y(new_n20510));
  nor_5  g18162(.A(new_n17591), .B(new_n7725), .Y(new_n20511));
  xnor_4 g18163(.A(new_n17591), .B(new_n7725), .Y(new_n20512));
  nor_5  g18164(.A(new_n17594), .B(new_n7730), .Y(new_n20513));
  xnor_4 g18165(.A(new_n17595), .B(new_n7729), .Y(new_n20514));
  not_8  g18166(.A(new_n17599), .Y(new_n20515_1));
  nor_5  g18167(.A(new_n20515_1), .B(new_n7739), .Y(new_n20516));
  xnor_4 g18168(.A(new_n20515_1), .B(new_n7739), .Y(new_n20517));
  nor_5  g18169(.A(new_n17605), .B(new_n7748), .Y(new_n20518));
  nor_5  g18170(.A(new_n20518), .B(new_n7743), .Y(new_n20519));
  xnor_4 g18171(.A(new_n20518), .B(new_n7742), .Y(new_n20520));
  and_5  g18172(.A(new_n20520), .B(new_n17611), .Y(new_n20521));
  nor_5  g18173(.A(new_n20521), .B(new_n20519), .Y(new_n20522));
  nor_5  g18174(.A(new_n20522), .B(new_n20517), .Y(new_n20523));
  nor_5  g18175(.A(new_n20523), .B(new_n20516), .Y(new_n20524));
  nor_5  g18176(.A(new_n20524), .B(new_n20514), .Y(new_n20525));
  nor_5  g18177(.A(new_n20525), .B(new_n20513), .Y(new_n20526));
  nor_5  g18178(.A(new_n20526), .B(new_n20512), .Y(new_n20527));
  nor_5  g18179(.A(new_n20527), .B(new_n20511), .Y(new_n20528));
  nor_5  g18180(.A(new_n20528), .B(new_n20510), .Y(new_n20529));
  nor_5  g18181(.A(new_n20529), .B(new_n20509), .Y(new_n20530));
  nor_5  g18182(.A(new_n20530), .B(new_n20508), .Y(new_n20531));
  nor_5  g18183(.A(new_n20531), .B(new_n20507), .Y(new_n20532));
  nor_5  g18184(.A(new_n20532), .B(new_n20506), .Y(new_n20533_1));
  nor_5  g18185(.A(new_n20533_1), .B(new_n20505), .Y(new_n20534));
  nor_5  g18186(.A(new_n20534), .B(new_n20504), .Y(new_n20535));
  nor_5  g18187(.A(new_n20535), .B(new_n20503), .Y(new_n20536));
  xnor_4 g18188(.A(new_n20536), .B(new_n20502), .Y(n7588));
  not_8  g18189(.A(new_n6679), .Y(new_n20538));
  nor_5  g18190(.A(new_n20538), .B(n21832), .Y(new_n20539));
  not_8  g18191(.A(new_n20539), .Y(new_n20540));
  nor_5  g18192(.A(new_n20540), .B(n21753), .Y(new_n20541));
  not_8  g18193(.A(new_n20541), .Y(new_n20542));
  nor_5  g18194(.A(new_n20542), .B(n10739), .Y(new_n20543));
  not_8  g18195(.A(new_n20543), .Y(new_n20544));
  nor_5  g18196(.A(new_n20544), .B(n13074), .Y(new_n20545));
  xnor_4 g18197(.A(new_n20545), .B(n23463), .Y(new_n20546));
  not_8  g18198(.A(new_n20546), .Y(new_n20547));
  xnor_4 g18199(.A(new_n20547), .B(n23250), .Y(new_n20548));
  xnor_4 g18200(.A(new_n20543), .B(n13074), .Y(new_n20549));
  nor_5  g18201(.A(new_n20549), .B(n11455), .Y(new_n20550));
  not_8  g18202(.A(new_n20549), .Y(new_n20551));
  xnor_4 g18203(.A(new_n20551), .B(n11455), .Y(new_n20552));
  xnor_4 g18204(.A(new_n20541), .B(n10739), .Y(new_n20553));
  nor_5  g18205(.A(new_n20553), .B(n3945), .Y(new_n20554));
  xnor_4 g18206(.A(new_n20553), .B(new_n15602_1), .Y(new_n20555));
  xnor_4 g18207(.A(new_n20539), .B(n21753), .Y(new_n20556));
  nor_5  g18208(.A(new_n20556), .B(n5255), .Y(new_n20557));
  not_8  g18209(.A(new_n20556), .Y(new_n20558));
  xnor_4 g18210(.A(new_n20558), .B(n5255), .Y(new_n20559));
  nor_5  g18211(.A(new_n6680), .B(n21649), .Y(new_n20560));
  xnor_4 g18212(.A(new_n6680), .B(new_n5163), .Y(new_n20561));
  nor_5  g18213(.A(new_n6698), .B(n18274), .Y(new_n20562));
  nor_5  g18214(.A(new_n6711), .B(n3828), .Y(new_n20563));
  xnor_4 g18215(.A(new_n6712), .B(n3828), .Y(new_n20564));
  nor_5  g18216(.A(new_n6706_1), .B(n23842), .Y(new_n20565));
  or_5   g18217(.A(new_n15011_1), .B(new_n3116), .Y(new_n20566));
  xnor_4 g18218(.A(new_n6706_1), .B(new_n5172), .Y(new_n20567));
  and_5  g18219(.A(new_n20567), .B(new_n20566), .Y(new_n20568));
  or_5   g18220(.A(new_n20568), .B(new_n20565), .Y(new_n20569));
  and_5  g18221(.A(new_n20569), .B(new_n20564), .Y(new_n20570));
  or_5   g18222(.A(new_n20570), .B(new_n20563), .Y(new_n20571));
  xnor_4 g18223(.A(new_n6698), .B(new_n5166), .Y(new_n20572));
  and_5  g18224(.A(new_n20572), .B(new_n20571), .Y(new_n20573));
  or_5   g18225(.A(new_n20573), .B(new_n20562), .Y(new_n20574));
  and_5  g18226(.A(new_n20574), .B(new_n20561), .Y(new_n20575));
  or_5   g18227(.A(new_n20575), .B(new_n20560), .Y(new_n20576));
  and_5  g18228(.A(new_n20576), .B(new_n20559), .Y(new_n20577));
  or_5   g18229(.A(new_n20577), .B(new_n20557), .Y(new_n20578));
  and_5  g18230(.A(new_n20578), .B(new_n20555), .Y(new_n20579));
  or_5   g18231(.A(new_n20579), .B(new_n20554), .Y(new_n20580));
  and_5  g18232(.A(new_n20580), .B(new_n20552), .Y(new_n20581));
  or_5   g18233(.A(new_n20581), .B(new_n20550), .Y(new_n20582_1));
  xor_4  g18234(.A(new_n20582_1), .B(new_n20548), .Y(new_n20583));
  xnor_4 g18235(.A(new_n20583), .B(new_n14074), .Y(new_n20584));
  xor_4  g18236(.A(new_n20580), .B(new_n20552), .Y(new_n20585));
  and_5  g18237(.A(new_n20585), .B(new_n14108), .Y(new_n20586));
  xnor_4 g18238(.A(new_n20585), .B(new_n14112), .Y(new_n20587));
  xor_4  g18239(.A(new_n20578), .B(new_n20555), .Y(new_n20588));
  nor_5  g18240(.A(new_n20588), .B(new_n14116), .Y(new_n20589));
  xnor_4 g18241(.A(new_n20588), .B(new_n14115), .Y(new_n20590_1));
  xor_4  g18242(.A(new_n20576), .B(new_n20559), .Y(new_n20591));
  nor_5  g18243(.A(new_n20591), .B(new_n14122), .Y(new_n20592));
  xor_4  g18244(.A(new_n20574), .B(new_n20561), .Y(new_n20593));
  nor_5  g18245(.A(new_n20593), .B(new_n14125), .Y(new_n20594));
  xor_4  g18246(.A(new_n20572), .B(new_n20571), .Y(new_n20595));
  nor_5  g18247(.A(new_n20595), .B(new_n14130_1), .Y(new_n20596));
  xnor_4 g18248(.A(new_n20595), .B(new_n14129), .Y(new_n20597));
  xor_4  g18249(.A(new_n20569), .B(new_n20564), .Y(new_n20598));
  nor_5  g18250(.A(new_n20598), .B(new_n14136_1), .Y(new_n20599));
  xnor_4 g18251(.A(new_n20598), .B(new_n14135), .Y(new_n20600));
  nor_5  g18252(.A(new_n20567), .B(new_n14140), .Y(new_n20601));
  xor_4  g18253(.A(new_n20567), .B(new_n20566), .Y(new_n20602_1));
  nor_5  g18254(.A(new_n20602_1), .B(new_n14139), .Y(new_n20603));
  xnor_4 g18255(.A(n21654), .B(n2387), .Y(new_n20604_1));
  nor_5  g18256(.A(new_n20604_1), .B(new_n14146), .Y(new_n20605));
  nor_5  g18257(.A(new_n20605), .B(new_n20603), .Y(new_n20606));
  nor_5  g18258(.A(new_n20606), .B(new_n20601), .Y(new_n20607));
  and_5  g18259(.A(new_n20607), .B(new_n20600), .Y(new_n20608));
  or_5   g18260(.A(new_n20608), .B(new_n20599), .Y(new_n20609_1));
  and_5  g18261(.A(new_n20609_1), .B(new_n20597), .Y(new_n20610));
  nor_5  g18262(.A(new_n20610), .B(new_n20596), .Y(new_n20611));
  xnor_4 g18263(.A(new_n20593), .B(new_n14125), .Y(new_n20612));
  nor_5  g18264(.A(new_n20612), .B(new_n20611), .Y(new_n20613));
  or_5   g18265(.A(new_n20613), .B(new_n20594), .Y(new_n20614));
  xnor_4 g18266(.A(new_n20591), .B(new_n14120), .Y(new_n20615));
  and_5  g18267(.A(new_n20615), .B(new_n20614), .Y(new_n20616));
  or_5   g18268(.A(new_n20616), .B(new_n20592), .Y(new_n20617));
  and_5  g18269(.A(new_n20617), .B(new_n20590_1), .Y(new_n20618));
  nor_5  g18270(.A(new_n20618), .B(new_n20589), .Y(new_n20619));
  and_5  g18271(.A(new_n20619), .B(new_n20587), .Y(new_n20620));
  nor_5  g18272(.A(new_n20620), .B(new_n20586), .Y(new_n20621));
  xor_4  g18273(.A(new_n20621), .B(new_n20584), .Y(n7598));
  xnor_4 g18274(.A(new_n17505), .B(new_n17502), .Y(n7607));
  xnor_4 g18275(.A(new_n5016), .B(new_n4991), .Y(n7610));
  xnor_4 g18276(.A(new_n3377), .B(new_n3366_1), .Y(n7616));
  xnor_4 g18277(.A(n10514), .B(n6105), .Y(new_n20626));
  nor_5  g18278(.A(n18649), .B(n3795), .Y(new_n20627));
  xnor_4 g18279(.A(n18649), .B(n3795), .Y(new_n20628));
  nor_5  g18280(.A(n25464), .B(n6218), .Y(new_n20629_1));
  xnor_4 g18281(.A(n25464), .B(n6218), .Y(new_n20630));
  nor_5  g18282(.A(n20470), .B(n4590), .Y(new_n20631));
  xnor_4 g18283(.A(n20470), .B(n4590), .Y(new_n20632));
  nor_5  g18284(.A(n26752), .B(n21222), .Y(new_n20633));
  xnor_4 g18285(.A(n26752), .B(n21222), .Y(new_n20634));
  nor_5  g18286(.A(n9832), .B(n6513), .Y(new_n20635));
  xnor_4 g18287(.A(n9832), .B(new_n6334), .Y(new_n20636));
  nor_5  g18288(.A(new_n6336), .B(new_n9479), .Y(new_n20637));
  or_5   g18289(.A(n3918), .B(n1558), .Y(new_n20638));
  nor_5  g18290(.A(n21749), .B(n919), .Y(new_n20639));
  nor_5  g18291(.A(new_n16100), .B(new_n16095), .Y(new_n20640));
  nor_5  g18292(.A(new_n20640), .B(new_n20639), .Y(new_n20641));
  and_5  g18293(.A(new_n20641), .B(new_n20638), .Y(new_n20642));
  nor_5  g18294(.A(new_n20642), .B(new_n20637), .Y(new_n20643));
  and_5  g18295(.A(new_n20643), .B(new_n20636), .Y(new_n20644));
  nor_5  g18296(.A(new_n20644), .B(new_n20635), .Y(new_n20645));
  nor_5  g18297(.A(new_n20645), .B(new_n20634), .Y(new_n20646));
  nor_5  g18298(.A(new_n20646), .B(new_n20633), .Y(new_n20647));
  nor_5  g18299(.A(new_n20647), .B(new_n20632), .Y(new_n20648));
  nor_5  g18300(.A(new_n20648), .B(new_n20631), .Y(new_n20649));
  nor_5  g18301(.A(new_n20649), .B(new_n20630), .Y(new_n20650));
  nor_5  g18302(.A(new_n20650), .B(new_n20629_1), .Y(new_n20651));
  nor_5  g18303(.A(new_n20651), .B(new_n20628), .Y(new_n20652));
  nor_5  g18304(.A(new_n20652), .B(new_n20627), .Y(new_n20653));
  xnor_4 g18305(.A(new_n20653), .B(new_n20626), .Y(new_n20654));
  nor_5  g18306(.A(new_n20654), .B(new_n20271), .Y(new_n20655));
  xnor_4 g18307(.A(new_n20654), .B(new_n20271), .Y(new_n20656));
  xnor_4 g18308(.A(new_n20651), .B(new_n20628), .Y(new_n20657));
  nor_5  g18309(.A(new_n20657), .B(new_n20275), .Y(new_n20658_1));
  xnor_4 g18310(.A(new_n20657), .B(new_n20275), .Y(new_n20659));
  xnor_4 g18311(.A(new_n20649), .B(new_n20630), .Y(new_n20660));
  nor_5  g18312(.A(new_n20660), .B(new_n20279_1), .Y(new_n20661_1));
  xnor_4 g18313(.A(new_n20660), .B(new_n20279_1), .Y(new_n20662));
  xnor_4 g18314(.A(new_n20647), .B(new_n20632), .Y(new_n20663));
  nor_5  g18315(.A(new_n20663), .B(new_n20283), .Y(new_n20664));
  xnor_4 g18316(.A(new_n20663), .B(new_n20283), .Y(new_n20665));
  xnor_4 g18317(.A(new_n20645), .B(new_n20634), .Y(new_n20666));
  nor_5  g18318(.A(new_n20666), .B(new_n20314), .Y(new_n20667));
  xnor_4 g18319(.A(new_n20666), .B(new_n20314), .Y(new_n20668));
  xnor_4 g18320(.A(new_n20643), .B(new_n20636), .Y(new_n20669));
  nor_5  g18321(.A(new_n20669), .B(new_n20289), .Y(new_n20670));
  xnor_4 g18322(.A(new_n20669), .B(new_n20289), .Y(new_n20671));
  xnor_4 g18323(.A(n3918), .B(n1558), .Y(new_n20672));
  xnor_4 g18324(.A(new_n20672), .B(new_n20641), .Y(new_n20673_1));
  nor_5  g18325(.A(new_n20673_1), .B(new_n20293), .Y(new_n20674));
  xnor_4 g18326(.A(new_n20673_1), .B(n24150), .Y(new_n20675));
  nor_5  g18327(.A(new_n16101), .B(new_n20297), .Y(new_n20676));
  and_5  g18328(.A(new_n16110_1), .B(new_n16102), .Y(new_n20677));
  or_5   g18329(.A(new_n20677), .B(new_n20676), .Y(new_n20678_1));
  and_5  g18330(.A(new_n20678_1), .B(new_n20675), .Y(new_n20679));
  nor_5  g18331(.A(new_n20679), .B(new_n20674), .Y(new_n20680_1));
  nor_5  g18332(.A(new_n20680_1), .B(new_n20671), .Y(new_n20681));
  nor_5  g18333(.A(new_n20681), .B(new_n20670), .Y(new_n20682));
  nor_5  g18334(.A(new_n20682), .B(new_n20668), .Y(new_n20683));
  nor_5  g18335(.A(new_n20683), .B(new_n20667), .Y(new_n20684));
  nor_5  g18336(.A(new_n20684), .B(new_n20665), .Y(new_n20685_1));
  nor_5  g18337(.A(new_n20685_1), .B(new_n20664), .Y(new_n20686));
  nor_5  g18338(.A(new_n20686), .B(new_n20662), .Y(new_n20687));
  nor_5  g18339(.A(new_n20687), .B(new_n20661_1), .Y(new_n20688));
  nor_5  g18340(.A(new_n20688), .B(new_n20659), .Y(new_n20689));
  nor_5  g18341(.A(new_n20689), .B(new_n20658_1), .Y(new_n20690));
  nor_5  g18342(.A(new_n20690), .B(new_n20656), .Y(new_n20691_1));
  nor_5  g18343(.A(new_n20691_1), .B(new_n20655), .Y(new_n20692));
  nor_5  g18344(.A(n10514), .B(n6105), .Y(new_n20693));
  nor_5  g18345(.A(new_n20653), .B(new_n20626), .Y(new_n20694));
  nor_5  g18346(.A(new_n20694), .B(new_n20693), .Y(new_n20695));
  nor_5  g18347(.A(new_n20695), .B(new_n20692), .Y(new_n20696_1));
  xnor_4 g18348(.A(new_n20696_1), .B(new_n15335), .Y(new_n20697));
  xnor_4 g18349(.A(new_n20695), .B(new_n20692), .Y(new_n20698));
  nor_5  g18350(.A(new_n20698), .B(new_n15227), .Y(new_n20699));
  xnor_4 g18351(.A(new_n20698), .B(new_n15227), .Y(new_n20700_1));
  xnor_4 g18352(.A(new_n20690), .B(new_n20656), .Y(new_n20701));
  nor_5  g18353(.A(new_n20701), .B(new_n15270), .Y(new_n20702));
  xnor_4 g18354(.A(new_n20701), .B(new_n15270), .Y(new_n20703));
  xnor_4 g18355(.A(new_n20688), .B(new_n20659), .Y(new_n20704_1));
  nor_5  g18356(.A(new_n20704_1), .B(new_n15274), .Y(new_n20705_1));
  xnor_4 g18357(.A(new_n20704_1), .B(new_n15274), .Y(new_n20706));
  xnor_4 g18358(.A(new_n20686), .B(new_n20662), .Y(new_n20707));
  nor_5  g18359(.A(new_n20707), .B(new_n15278), .Y(new_n20708));
  xnor_4 g18360(.A(new_n20707), .B(new_n15278), .Y(new_n20709_1));
  xnor_4 g18361(.A(new_n20684), .B(new_n20665), .Y(new_n20710));
  nor_5  g18362(.A(new_n20710), .B(new_n15282), .Y(new_n20711));
  xnor_4 g18363(.A(new_n20710), .B(new_n15282), .Y(new_n20712));
  xnor_4 g18364(.A(new_n20682), .B(new_n20668), .Y(new_n20713_1));
  nor_5  g18365(.A(new_n20713_1), .B(new_n15286), .Y(new_n20714));
  xnor_4 g18366(.A(new_n20713_1), .B(new_n15286), .Y(new_n20715));
  xnor_4 g18367(.A(new_n20680_1), .B(new_n20671), .Y(new_n20716));
  nor_5  g18368(.A(new_n20716), .B(new_n15291), .Y(new_n20717));
  xnor_4 g18369(.A(new_n20716), .B(new_n15291), .Y(new_n20718));
  xor_4  g18370(.A(new_n20678_1), .B(new_n20675), .Y(new_n20719));
  and_5  g18371(.A(new_n20719), .B(new_n15296), .Y(new_n20720));
  xnor_4 g18372(.A(new_n20719), .B(new_n15296), .Y(new_n20721));
  nor_5  g18373(.A(new_n16111), .B(new_n15301), .Y(new_n20722_1));
  nor_5  g18374(.A(new_n16119), .B(new_n16112), .Y(new_n20723_1));
  nor_5  g18375(.A(new_n20723_1), .B(new_n20722_1), .Y(new_n20724));
  nor_5  g18376(.A(new_n20724), .B(new_n20721), .Y(new_n20725));
  nor_5  g18377(.A(new_n20725), .B(new_n20720), .Y(new_n20726));
  nor_5  g18378(.A(new_n20726), .B(new_n20718), .Y(new_n20727));
  nor_5  g18379(.A(new_n20727), .B(new_n20717), .Y(new_n20728));
  nor_5  g18380(.A(new_n20728), .B(new_n20715), .Y(new_n20729));
  nor_5  g18381(.A(new_n20729), .B(new_n20714), .Y(new_n20730));
  nor_5  g18382(.A(new_n20730), .B(new_n20712), .Y(new_n20731));
  nor_5  g18383(.A(new_n20731), .B(new_n20711), .Y(new_n20732));
  nor_5  g18384(.A(new_n20732), .B(new_n20709_1), .Y(new_n20733));
  nor_5  g18385(.A(new_n20733), .B(new_n20708), .Y(new_n20734));
  nor_5  g18386(.A(new_n20734), .B(new_n20706), .Y(new_n20735));
  nor_5  g18387(.A(new_n20735), .B(new_n20705_1), .Y(new_n20736));
  nor_5  g18388(.A(new_n20736), .B(new_n20703), .Y(new_n20737));
  nor_5  g18389(.A(new_n20737), .B(new_n20702), .Y(new_n20738));
  nor_5  g18390(.A(new_n20738), .B(new_n20700_1), .Y(new_n20739));
  nor_5  g18391(.A(new_n20739), .B(new_n20699), .Y(new_n20740));
  xnor_4 g18392(.A(new_n20740), .B(new_n20697), .Y(n7630));
  nor_5  g18393(.A(new_n18324), .B(new_n18300), .Y(new_n20742));
  nor_5  g18394(.A(new_n18333), .B(new_n18325), .Y(new_n20743));
  nor_5  g18395(.A(new_n20743), .B(new_n20742), .Y(n7643));
  xnor_4 g18396(.A(new_n12010), .B(new_n11987), .Y(n7647));
  xnor_4 g18397(.A(new_n9974), .B(new_n9941), .Y(n7679));
  xnor_4 g18398(.A(new_n19651), .B(new_n19629), .Y(n7686));
  xnor_4 g18399(.A(new_n17857), .B(new_n17816), .Y(new_n20748_1));
  xnor_4 g18400(.A(new_n20748_1), .B(new_n17855_1), .Y(n7698));
  xnor_4 g18401(.A(new_n18921), .B(new_n18906), .Y(n7708));
  not_8  g18402(.A(n3324), .Y(new_n20751));
  xnor_4 g18403(.A(new_n17831), .B(new_n20751), .Y(new_n20752));
  nor_5  g18404(.A(new_n2925), .B(new_n19668), .Y(new_n20753));
  xnor_4 g18405(.A(new_n2925), .B(n17911), .Y(new_n20754));
  nor_5  g18406(.A(new_n2976), .B(n21997), .Y(new_n20755));
  xnor_4 g18407(.A(new_n2976), .B(new_n18472), .Y(new_n20756));
  nor_5  g18408(.A(new_n2980), .B(n25119), .Y(new_n20757));
  and_5  g18409(.A(new_n8526_1), .B(new_n8502), .Y(new_n20758));
  or_5   g18410(.A(new_n20758), .B(new_n20757), .Y(new_n20759));
  and_5  g18411(.A(new_n20759), .B(new_n20756), .Y(new_n20760));
  nor_5  g18412(.A(new_n20760), .B(new_n20755), .Y(new_n20761_1));
  and_5  g18413(.A(new_n20761_1), .B(new_n20754), .Y(new_n20762));
  nor_5  g18414(.A(new_n20762), .B(new_n20753), .Y(new_n20763));
  xnor_4 g18415(.A(new_n20763), .B(new_n20752), .Y(new_n20764));
  xnor_4 g18416(.A(new_n6023), .B(new_n4907), .Y(new_n20765));
  nor_5  g18417(.A(new_n6029), .B(n2858), .Y(new_n20766));
  and_5  g18418(.A(new_n15882), .B(new_n15874), .Y(new_n20767));
  nor_5  g18419(.A(new_n20767), .B(new_n20766), .Y(new_n20768));
  xnor_4 g18420(.A(new_n20768), .B(new_n20765), .Y(new_n20769));
  xnor_4 g18421(.A(new_n20769), .B(new_n20764), .Y(new_n20770));
  not_8  g18422(.A(new_n15883), .Y(new_n20771));
  xor_4  g18423(.A(new_n20761_1), .B(new_n20754), .Y(new_n20772));
  nor_5  g18424(.A(new_n20772), .B(new_n20771), .Y(new_n20773));
  xnor_4 g18425(.A(new_n20772), .B(new_n20771), .Y(new_n20774_1));
  xor_4  g18426(.A(new_n20759), .B(new_n20756), .Y(new_n20775));
  and_5  g18427(.A(new_n20775), .B(new_n15885_1), .Y(new_n20776));
  xnor_4 g18428(.A(new_n20775), .B(new_n15885_1), .Y(new_n20777));
  nor_5  g18429(.A(new_n8527), .B(new_n8500), .Y(new_n20778));
  nor_5  g18430(.A(new_n8570), .B(new_n8528), .Y(new_n20779));
  nor_5  g18431(.A(new_n20779), .B(new_n20778), .Y(new_n20780));
  nor_5  g18432(.A(new_n20780), .B(new_n20777), .Y(new_n20781));
  nor_5  g18433(.A(new_n20781), .B(new_n20776), .Y(new_n20782));
  nor_5  g18434(.A(new_n20782), .B(new_n20774_1), .Y(new_n20783));
  nor_5  g18435(.A(new_n20783), .B(new_n20773), .Y(new_n20784));
  xnor_4 g18436(.A(new_n20784), .B(new_n20770), .Y(n7780));
  nor_5  g18437(.A(new_n2603), .B(new_n4471), .Y(new_n20786));
  xnor_4 g18438(.A(new_n2603), .B(new_n4471), .Y(new_n20787));
  nor_5  g18439(.A(new_n2607), .B(new_n4431), .Y(new_n20788_1));
  nor_5  g18440(.A(new_n9598_1), .B(new_n9569), .Y(new_n20789));
  nor_5  g18441(.A(new_n20789), .B(new_n20788_1), .Y(new_n20790));
  nor_5  g18442(.A(new_n20790), .B(new_n20787), .Y(new_n20791));
  nor_5  g18443(.A(new_n20791), .B(new_n20786), .Y(new_n20792));
  xnor_4 g18444(.A(new_n20792), .B(new_n14355), .Y(new_n20793));
  not_8  g18445(.A(new_n20793), .Y(new_n20794_1));
  nor_5  g18446(.A(new_n16940), .B(new_n10052), .Y(new_n20795_1));
  xnor_4 g18447(.A(new_n16939), .B(new_n10052), .Y(new_n20796));
  and_5  g18448(.A(new_n9611), .B(new_n2723), .Y(new_n20797));
  and_5  g18449(.A(new_n9648_1), .B(new_n9612), .Y(new_n20798));
  or_5   g18450(.A(new_n20798), .B(new_n20797), .Y(new_n20799));
  and_5  g18451(.A(new_n20799), .B(new_n20796), .Y(new_n20800));
  nor_5  g18452(.A(new_n20800), .B(new_n20795_1), .Y(new_n20801));
  not_8  g18453(.A(new_n20801), .Y(new_n20802));
  and_5  g18454(.A(new_n16938), .B(new_n4312), .Y(new_n20803_1));
  xnor_4 g18455(.A(new_n20803_1), .B(new_n10049), .Y(new_n20804));
  xnor_4 g18456(.A(new_n20804), .B(new_n20802), .Y(new_n20805));
  xnor_4 g18457(.A(new_n20805), .B(new_n20794_1), .Y(new_n20806));
  xor_4  g18458(.A(new_n20790), .B(new_n20787), .Y(new_n20807));
  xor_4  g18459(.A(new_n20799), .B(new_n20796), .Y(new_n20808));
  nor_5  g18460(.A(new_n20808), .B(new_n20807), .Y(new_n20809));
  xnor_4 g18461(.A(new_n20808), .B(new_n20807), .Y(new_n20810));
  nor_5  g18462(.A(new_n9649), .B(new_n9599), .Y(new_n20811));
  and_5  g18463(.A(new_n9703), .B(new_n9650), .Y(new_n20812));
  nor_5  g18464(.A(new_n20812), .B(new_n20811), .Y(new_n20813));
  nor_5  g18465(.A(new_n20813), .B(new_n20810), .Y(new_n20814));
  nor_5  g18466(.A(new_n20814), .B(new_n20809), .Y(new_n20815));
  xnor_4 g18467(.A(new_n20815), .B(new_n20806), .Y(n7794));
  xnor_4 g18468(.A(new_n17118), .B(new_n17113), .Y(n7811));
  xor_4  g18469(.A(new_n17066), .B(new_n17061), .Y(n7830));
  xnor_4 g18470(.A(new_n20532), .B(new_n20506), .Y(n7834));
  xnor_4 g18471(.A(new_n10862), .B(new_n10850), .Y(n7884));
  xnor_4 g18472(.A(new_n3070), .B(new_n3069), .Y(n7937));
  xnor_4 g18473(.A(new_n3082), .B(new_n3037), .Y(n7943));
  xor_4  g18474(.A(new_n9697), .B(new_n9666), .Y(n7950));
  xnor_4 g18475(.A(new_n19167), .B(new_n15180_1), .Y(new_n20824));
  nor_5  g18476(.A(new_n19170), .B(new_n15184), .Y(new_n20825));
  nor_5  g18477(.A(new_n19173), .B(new_n15189), .Y(new_n20826_1));
  xnor_4 g18478(.A(new_n19173), .B(new_n15189), .Y(new_n20827));
  nor_5  g18479(.A(new_n15192), .B(new_n14886), .Y(new_n20828));
  nor_5  g18480(.A(new_n14979), .B(new_n14933), .Y(new_n20829));
  nor_5  g18481(.A(new_n20829), .B(new_n20828), .Y(new_n20830));
  nor_5  g18482(.A(new_n20830), .B(new_n20827), .Y(new_n20831));
  nor_5  g18483(.A(new_n20831), .B(new_n20826_1), .Y(new_n20832));
  xnor_4 g18484(.A(new_n19181), .B(new_n15182_1), .Y(new_n20833));
  nor_5  g18485(.A(new_n20833), .B(new_n20832), .Y(new_n20834));
  nor_5  g18486(.A(new_n20834), .B(new_n20825), .Y(new_n20835));
  xor_4  g18487(.A(new_n20835), .B(new_n20824), .Y(n7959));
  xnor_4 g18488(.A(new_n17122), .B(new_n17109), .Y(n7968));
  xnor_4 g18489(.A(new_n18071_1), .B(new_n18070), .Y(n7992));
  xnor_4 g18490(.A(new_n12681), .B(n9554), .Y(new_n20839));
  nor_5  g18491(.A(new_n12685), .B(new_n7773_1), .Y(new_n20840));
  xnor_4 g18492(.A(new_n12687), .B(new_n7773_1), .Y(new_n20841));
  nor_5  g18493(.A(new_n10450), .B(n18227), .Y(new_n20842));
  and_5  g18494(.A(new_n17094), .B(new_n17082), .Y(new_n20843));
  nor_5  g18495(.A(new_n20843), .B(new_n20842), .Y(new_n20844));
  and_5  g18496(.A(new_n20844), .B(new_n20841), .Y(new_n20845));
  nor_5  g18497(.A(new_n20845), .B(new_n20840), .Y(new_n20846));
  xnor_4 g18498(.A(new_n20846), .B(new_n20839), .Y(new_n20847));
  xnor_4 g18499(.A(new_n20847), .B(new_n18231), .Y(new_n20848));
  xnor_4 g18500(.A(new_n20844), .B(new_n20841), .Y(new_n20849));
  nor_5  g18501(.A(new_n20849), .B(new_n18235), .Y(new_n20850));
  not_8  g18502(.A(new_n20849), .Y(new_n20851));
  xnor_4 g18503(.A(new_n20851), .B(new_n18236), .Y(new_n20852));
  nor_5  g18504(.A(new_n18240), .B(new_n17096), .Y(new_n20853));
  xnor_4 g18505(.A(new_n18241_1), .B(new_n17095_1), .Y(new_n20854));
  nor_5  g18506(.A(new_n18245), .B(new_n17100), .Y(new_n20855));
  xnor_4 g18507(.A(new_n18246), .B(new_n17099), .Y(new_n20856));
  and_5  g18508(.A(new_n18251), .B(new_n17104_1), .Y(new_n20857));
  xnor_4 g18509(.A(new_n18251), .B(new_n17104_1), .Y(new_n20858));
  nor_5  g18510(.A(new_n12769), .B(new_n17107), .Y(new_n20859));
  nor_5  g18511(.A(new_n12774), .B(new_n12771), .Y(new_n20860));
  nor_5  g18512(.A(new_n20860), .B(new_n20859), .Y(new_n20861));
  nor_5  g18513(.A(new_n20861), .B(new_n20858), .Y(new_n20862));
  nor_5  g18514(.A(new_n20862), .B(new_n20857), .Y(new_n20863));
  nor_5  g18515(.A(new_n20863), .B(new_n20856), .Y(new_n20864));
  nor_5  g18516(.A(new_n20864), .B(new_n20855), .Y(new_n20865));
  nor_5  g18517(.A(new_n20865), .B(new_n20854), .Y(new_n20866));
  nor_5  g18518(.A(new_n20866), .B(new_n20853), .Y(new_n20867));
  nor_5  g18519(.A(new_n20867), .B(new_n20852), .Y(new_n20868));
  nor_5  g18520(.A(new_n20868), .B(new_n20850), .Y(new_n20869_1));
  xnor_4 g18521(.A(new_n20869_1), .B(new_n20848), .Y(n7999));
  xnor_4 g18522(.A(new_n17725), .B(new_n17712), .Y(n8027));
  nor_5  g18523(.A(new_n20792), .B(new_n14355), .Y(new_n20872));
  not_8  g18524(.A(new_n20872), .Y(new_n20873));
  nor_5  g18525(.A(new_n6244), .B(new_n6198), .Y(new_n20874));
  xnor_4 g18526(.A(new_n6244), .B(n8614), .Y(new_n20875));
  nor_5  g18527(.A(new_n6250), .B(new_n6215), .Y(new_n20876));
  nor_5  g18528(.A(new_n6257), .B(n27037), .Y(new_n20877));
  xnor_4 g18529(.A(new_n6256_1), .B(n27037), .Y(new_n20878));
  nor_5  g18530(.A(new_n6304), .B(n8964), .Y(new_n20879_1));
  xnor_4 g18531(.A(new_n6304), .B(new_n6222), .Y(new_n20880));
  nor_5  g18532(.A(new_n6268), .B(new_n6227), .Y(new_n20881));
  nor_5  g18533(.A(new_n6273), .B(new_n4015), .Y(new_n20882));
  and_5  g18534(.A(new_n20475), .B(new_n20472), .Y(new_n20883));
  or_5   g18535(.A(new_n20883), .B(new_n20882), .Y(new_n20884));
  xnor_4 g18536(.A(new_n6269), .B(new_n6227), .Y(new_n20885));
  and_5  g18537(.A(new_n20885), .B(new_n20884), .Y(new_n20886));
  nor_5  g18538(.A(new_n20886), .B(new_n20881), .Y(new_n20887));
  and_5  g18539(.A(new_n20887), .B(new_n20880), .Y(new_n20888));
  or_5   g18540(.A(new_n20888), .B(new_n20879_1), .Y(new_n20889));
  and_5  g18541(.A(new_n20889), .B(new_n20878), .Y(new_n20890));
  nor_5  g18542(.A(new_n20890), .B(new_n20877), .Y(new_n20891));
  xnor_4 g18543(.A(new_n6251), .B(new_n6215), .Y(new_n20892));
  and_5  g18544(.A(new_n20892), .B(new_n20891), .Y(new_n20893));
  or_5   g18545(.A(new_n20893), .B(new_n20876), .Y(new_n20894));
  and_5  g18546(.A(new_n20894), .B(new_n20875), .Y(new_n20895));
  nor_5  g18547(.A(new_n20895), .B(new_n20874), .Y(new_n20896));
  nor_5  g18548(.A(new_n20896), .B(new_n6242), .Y(new_n20897));
  nor_5  g18549(.A(new_n20897), .B(new_n20873), .Y(new_n20898));
  and_5  g18550(.A(new_n20897), .B(new_n20873), .Y(new_n20899));
  xnor_4 g18551(.A(new_n20896), .B(new_n6197), .Y(new_n20900));
  nor_5  g18552(.A(new_n20900), .B(new_n20793), .Y(new_n20901));
  xnor_4 g18553(.A(new_n20900), .B(new_n20793), .Y(new_n20902));
  not_8  g18554(.A(new_n20807), .Y(new_n20903));
  xor_4  g18555(.A(new_n20894), .B(new_n20875), .Y(new_n20904));
  nor_5  g18556(.A(new_n20904), .B(new_n20903), .Y(new_n20905));
  xnor_4 g18557(.A(new_n20904), .B(new_n20903), .Y(new_n20906));
  xor_4  g18558(.A(new_n20892), .B(new_n20891), .Y(new_n20907));
  nor_5  g18559(.A(new_n20907), .B(new_n9600), .Y(new_n20908));
  xnor_4 g18560(.A(new_n20907), .B(new_n9600), .Y(new_n20909));
  xor_4  g18561(.A(new_n20889), .B(new_n20878), .Y(new_n20910));
  and_5  g18562(.A(new_n20910), .B(new_n9651), .Y(new_n20911));
  xnor_4 g18563(.A(new_n20910), .B(new_n9651), .Y(new_n20912));
  xnor_4 g18564(.A(new_n20887), .B(new_n20880), .Y(new_n20913));
  nor_5  g18565(.A(new_n20913), .B(new_n9660), .Y(new_n20914));
  xnor_4 g18566(.A(new_n20913), .B(new_n9660), .Y(new_n20915_1));
  xor_4  g18567(.A(new_n20885), .B(new_n20884), .Y(new_n20916));
  nor_5  g18568(.A(new_n20916), .B(new_n9663), .Y(new_n20917));
  xnor_4 g18569(.A(new_n20916), .B(new_n9663), .Y(new_n20918));
  nor_5  g18570(.A(new_n20476), .B(new_n9668), .Y(new_n20919));
  nor_5  g18571(.A(new_n20480), .B(new_n20477), .Y(new_n20920));
  nor_5  g18572(.A(new_n20920), .B(new_n20919), .Y(new_n20921));
  nor_5  g18573(.A(new_n20921), .B(new_n20918), .Y(new_n20922));
  nor_5  g18574(.A(new_n20922), .B(new_n20917), .Y(new_n20923_1));
  nor_5  g18575(.A(new_n20923_1), .B(new_n20915_1), .Y(new_n20924));
  nor_5  g18576(.A(new_n20924), .B(new_n20914), .Y(new_n20925));
  nor_5  g18577(.A(new_n20925), .B(new_n20912), .Y(new_n20926));
  nor_5  g18578(.A(new_n20926), .B(new_n20911), .Y(new_n20927));
  nor_5  g18579(.A(new_n20927), .B(new_n20909), .Y(new_n20928));
  nor_5  g18580(.A(new_n20928), .B(new_n20908), .Y(new_n20929_1));
  nor_5  g18581(.A(new_n20929_1), .B(new_n20906), .Y(new_n20930));
  nor_5  g18582(.A(new_n20930), .B(new_n20905), .Y(new_n20931));
  nor_5  g18583(.A(new_n20931), .B(new_n20902), .Y(new_n20932));
  nor_5  g18584(.A(new_n20932), .B(new_n20901), .Y(new_n20933));
  nor_5  g18585(.A(new_n20933), .B(new_n20899), .Y(new_n20934));
  or_5   g18586(.A(new_n20934), .B(new_n20898), .Y(n8031));
  and_5  g18587(.A(new_n16939), .B(n22626), .Y(new_n20936_1));
  nor_5  g18588(.A(new_n16939), .B(n22626), .Y(new_n20937));
  nor_5  g18589(.A(new_n16949), .B(new_n20937), .Y(new_n20938));
  or_5   g18590(.A(new_n20938), .B(new_n20803_1), .Y(new_n20939));
  nor_5  g18591(.A(new_n20939), .B(new_n20936_1), .Y(new_n20940));
  not_8  g18592(.A(new_n20940), .Y(new_n20941));
  nor_5  g18593(.A(new_n20941), .B(new_n19325), .Y(new_n20942));
  xnor_4 g18594(.A(new_n20941), .B(new_n19325), .Y(new_n20943));
  nor_5  g18595(.A(new_n16950), .B(new_n16936), .Y(new_n20944));
  not_8  g18596(.A(new_n16977), .Y(new_n20945));
  nor_5  g18597(.A(new_n20945), .B(new_n16951_1), .Y(new_n20946_1));
  nor_5  g18598(.A(new_n20946_1), .B(new_n20944), .Y(new_n20947));
  nor_5  g18599(.A(new_n20947), .B(new_n20943), .Y(new_n20948));
  nor_5  g18600(.A(new_n20948), .B(new_n20942), .Y(new_n20949));
  not_8  g18601(.A(new_n20949), .Y(new_n20950));
  or_5   g18602(.A(new_n16992), .B(n9554), .Y(new_n20951));
  and_5  g18603(.A(new_n17022), .B(new_n20951), .Y(new_n20952));
  and_5  g18604(.A(new_n16992), .B(n9554), .Y(new_n20953));
  or_5   g18605(.A(new_n20953), .B(new_n19605), .Y(new_n20954));
  nor_5  g18606(.A(new_n20954), .B(new_n20952), .Y(new_n20955));
  nor_5  g18607(.A(new_n20955), .B(new_n20950), .Y(new_n20956));
  not_8  g18608(.A(new_n20955), .Y(new_n20957));
  xnor_4 g18609(.A(new_n20957), .B(new_n20950), .Y(new_n20958));
  xnor_4 g18610(.A(new_n20947), .B(new_n20943), .Y(new_n20959));
  not_8  g18611(.A(new_n20959), .Y(new_n20960));
  nor_5  g18612(.A(new_n20960), .B(new_n20957), .Y(new_n20961));
  xnor_4 g18613(.A(new_n20960), .B(new_n20957), .Y(new_n20962));
  nor_5  g18614(.A(new_n17023), .B(new_n16978), .Y(new_n20963));
  nor_5  g18615(.A(new_n17080), .B(new_n17025), .Y(new_n20964));
  nor_5  g18616(.A(new_n20964), .B(new_n20963), .Y(new_n20965));
  nor_5  g18617(.A(new_n20965), .B(new_n20962), .Y(new_n20966));
  or_5   g18618(.A(new_n20966), .B(new_n20961), .Y(new_n20967));
  and_5  g18619(.A(new_n20967), .B(new_n20958), .Y(new_n20968));
  nor_5  g18620(.A(new_n20968), .B(new_n20956), .Y(n8042));
  nor_5  g18621(.A(new_n9910), .B(new_n9817), .Y(new_n20970));
  nor_5  g18622(.A(new_n9986), .B(new_n9911), .Y(new_n20971));
  or_5   g18623(.A(new_n20971), .B(new_n20970), .Y(n8095));
  nor_5  g18624(.A(new_n17625), .B(n4306), .Y(new_n20973));
  xnor_4 g18625(.A(n23166), .B(n4306), .Y(new_n20974));
  nor_5  g18626(.A(new_n9079), .B(n3279), .Y(new_n20975));
  xnor_4 g18627(.A(n10577), .B(n3279), .Y(new_n20976));
  nor_5  g18628(.A(n13914), .B(new_n9082), .Y(new_n20977));
  xnor_4 g18629(.A(n13914), .B(n6381), .Y(new_n20978));
  nor_5  g18630(.A(n14702), .B(new_n9085), .Y(new_n20979));
  and_5  g18631(.A(new_n19072), .B(new_n19061), .Y(new_n20980));
  or_5   g18632(.A(new_n20980), .B(new_n20979), .Y(new_n20981));
  and_5  g18633(.A(new_n20981), .B(new_n20978), .Y(new_n20982));
  or_5   g18634(.A(new_n20982), .B(new_n20977), .Y(new_n20983));
  and_5  g18635(.A(new_n20983), .B(new_n20976), .Y(new_n20984));
  or_5   g18636(.A(new_n20984), .B(new_n20975), .Y(new_n20985));
  and_5  g18637(.A(new_n20985), .B(new_n20974), .Y(new_n20986_1));
  nor_5  g18638(.A(new_n20986_1), .B(new_n20973), .Y(new_n20987));
  xnor_4 g18639(.A(new_n20987), .B(new_n8953), .Y(new_n20988));
  xor_4  g18640(.A(new_n20985), .B(new_n20974), .Y(new_n20989));
  nor_5  g18641(.A(new_n20989), .B(new_n8999), .Y(new_n20990));
  xnor_4 g18642(.A(new_n20989), .B(new_n8999), .Y(new_n20991));
  xor_4  g18643(.A(new_n20983), .B(new_n20976), .Y(new_n20992));
  nor_5  g18644(.A(new_n20992), .B(new_n9003_1), .Y(new_n20993));
  xnor_4 g18645(.A(new_n20992), .B(new_n9003_1), .Y(new_n20994));
  xor_4  g18646(.A(new_n20981), .B(new_n20978), .Y(new_n20995));
  nor_5  g18647(.A(new_n20995), .B(new_n9007), .Y(new_n20996));
  xnor_4 g18648(.A(new_n20995), .B(new_n9007), .Y(new_n20997));
  not_8  g18649(.A(new_n20997), .Y(new_n20998));
  and_5  g18650(.A(new_n19073), .B(new_n9011), .Y(new_n20999));
  and_5  g18651(.A(new_n19088), .B(new_n19074), .Y(new_n21000));
  nor_5  g18652(.A(new_n21000), .B(new_n20999), .Y(new_n21001));
  and_5  g18653(.A(new_n21001), .B(new_n20998), .Y(new_n21002));
  nor_5  g18654(.A(new_n21002), .B(new_n20996), .Y(new_n21003));
  nor_5  g18655(.A(new_n21003), .B(new_n20994), .Y(new_n21004));
  nor_5  g18656(.A(new_n21004), .B(new_n20993), .Y(new_n21005));
  nor_5  g18657(.A(new_n21005), .B(new_n20991), .Y(new_n21006));
  nor_5  g18658(.A(new_n21006), .B(new_n20990), .Y(new_n21007));
  xnor_4 g18659(.A(new_n21007), .B(new_n20988), .Y(n8103));
  xnor_4 g18660(.A(new_n18467_1), .B(new_n18456), .Y(n8109));
  nor_5  g18661(.A(new_n18896), .B(new_n18878), .Y(new_n21010));
  nor_5  g18662(.A(new_n18925), .B(new_n18897), .Y(new_n21011));
  or_5   g18663(.A(new_n21011), .B(new_n21010), .Y(n8127));
  xnor_4 g18664(.A(new_n16483), .B(new_n16480), .Y(n8130));
  nor_5  g18665(.A(n8856), .B(new_n3087), .Y(new_n21014));
  xnor_4 g18666(.A(n8856), .B(n4319), .Y(new_n21015));
  nor_5  g18667(.A(new_n11610), .B(n14130), .Y(new_n21016));
  xnor_4 g18668(.A(n23463), .B(n14130), .Y(new_n21017_1));
  nor_5  g18669(.A(n16482), .B(new_n3095), .Y(new_n21018));
  xnor_4 g18670(.A(n16482), .B(n13074), .Y(new_n21019));
  nor_5  g18671(.A(new_n3099), .B(n9942), .Y(new_n21020));
  and_5  g18672(.A(new_n2379), .B(new_n2349), .Y(new_n21021));
  or_5   g18673(.A(new_n21021), .B(new_n21020), .Y(new_n21022));
  and_5  g18674(.A(new_n21022), .B(new_n21019), .Y(new_n21023));
  or_5   g18675(.A(new_n21023), .B(new_n21018), .Y(new_n21024));
  and_5  g18676(.A(new_n21024), .B(new_n21017_1), .Y(new_n21025));
  or_5   g18677(.A(new_n21025), .B(new_n21016), .Y(new_n21026));
  and_5  g18678(.A(new_n21026), .B(new_n21015), .Y(new_n21027));
  nor_5  g18679(.A(new_n21027), .B(new_n21014), .Y(new_n21028));
  xnor_4 g18680(.A(new_n21028), .B(new_n7547), .Y(new_n21029));
  nor_5  g18681(.A(new_n21028), .B(new_n7550), .Y(new_n21030));
  xnor_4 g18682(.A(new_n21028), .B(new_n7550), .Y(new_n21031));
  xor_4  g18683(.A(new_n21026), .B(new_n21015), .Y(new_n21032));
  nor_5  g18684(.A(new_n21032), .B(new_n7554), .Y(new_n21033));
  xnor_4 g18685(.A(new_n21032), .B(new_n7554), .Y(new_n21034_1));
  xor_4  g18686(.A(new_n21024), .B(new_n21017_1), .Y(new_n21035));
  nor_5  g18687(.A(new_n21035), .B(new_n7558_1), .Y(new_n21036));
  xnor_4 g18688(.A(new_n21035), .B(new_n7558_1), .Y(new_n21037));
  not_8  g18689(.A(new_n21037), .Y(new_n21038));
  xor_4  g18690(.A(new_n21022), .B(new_n21019), .Y(new_n21039));
  and_5  g18691(.A(new_n21039), .B(new_n7562), .Y(new_n21040));
  xnor_4 g18692(.A(new_n21039), .B(new_n7562), .Y(new_n21041));
  and_5  g18693(.A(new_n2501), .B(new_n2380), .Y(new_n21042));
  and_5  g18694(.A(new_n2540), .B(new_n2502), .Y(new_n21043));
  nor_5  g18695(.A(new_n21043), .B(new_n21042), .Y(new_n21044));
  nor_5  g18696(.A(new_n21044), .B(new_n21041), .Y(new_n21045));
  nor_5  g18697(.A(new_n21045), .B(new_n21040), .Y(new_n21046_1));
  and_5  g18698(.A(new_n21046_1), .B(new_n21038), .Y(new_n21047));
  nor_5  g18699(.A(new_n21047), .B(new_n21036), .Y(new_n21048));
  nor_5  g18700(.A(new_n21048), .B(new_n21034_1), .Y(new_n21049));
  nor_5  g18701(.A(new_n21049), .B(new_n21033), .Y(new_n21050));
  nor_5  g18702(.A(new_n21050), .B(new_n21031), .Y(new_n21051));
  nor_5  g18703(.A(new_n21051), .B(new_n21030), .Y(new_n21052));
  xnor_4 g18704(.A(new_n21052), .B(new_n21029), .Y(n8135));
  xnor_4 g18705(.A(new_n7586), .B(new_n2529), .Y(n8139));
  not_8  g18706(.A(new_n17865), .Y(new_n21055));
  nor_5  g18707(.A(new_n21055), .B(n3018), .Y(new_n21056));
  not_8  g18708(.A(new_n21056), .Y(new_n21057));
  nor_5  g18709(.A(new_n21057), .B(n26660), .Y(new_n21058));
  xnor_4 g18710(.A(new_n21058), .B(n13783), .Y(new_n21059));
  xnor_4 g18711(.A(new_n21059), .B(new_n2981), .Y(new_n21060));
  xnor_4 g18712(.A(new_n21056), .B(n26660), .Y(new_n21061));
  and_5  g18713(.A(new_n21061), .B(new_n2987), .Y(new_n21062_1));
  xnor_4 g18714(.A(new_n21061), .B(new_n2987), .Y(new_n21063));
  and_5  g18715(.A(new_n17866), .B(new_n2992), .Y(new_n21064));
  and_5  g18716(.A(new_n17884), .B(new_n17867), .Y(new_n21065));
  nor_5  g18717(.A(new_n21065), .B(new_n21064), .Y(new_n21066));
  nor_5  g18718(.A(new_n21066), .B(new_n21063), .Y(new_n21067));
  nor_5  g18719(.A(new_n21067), .B(new_n21062_1), .Y(new_n21068));
  xor_4  g18720(.A(new_n21068), .B(new_n21060), .Y(new_n21069));
  xnor_4 g18721(.A(new_n21069), .B(new_n6918), .Y(new_n21070));
  xor_4  g18722(.A(new_n21066), .B(new_n21063), .Y(new_n21071));
  nor_5  g18723(.A(new_n21071), .B(new_n6923), .Y(new_n21072));
  xnor_4 g18724(.A(new_n21071), .B(new_n6923), .Y(new_n21073));
  nor_5  g18725(.A(new_n17885), .B(new_n6926), .Y(new_n21074));
  nor_5  g18726(.A(new_n17903), .B(new_n17886), .Y(new_n21075));
  nor_5  g18727(.A(new_n21075), .B(new_n21074), .Y(new_n21076));
  nor_5  g18728(.A(new_n21076), .B(new_n21073), .Y(new_n21077));
  nor_5  g18729(.A(new_n21077), .B(new_n21072), .Y(new_n21078_1));
  xnor_4 g18730(.A(new_n21078_1), .B(new_n21070), .Y(n8148));
  xor_4  g18731(.A(new_n17284), .B(new_n17283), .Y(n8149));
  xnor_4 g18732(.A(new_n3920), .B(new_n3903), .Y(n8159));
  xnor_4 g18733(.A(new_n11560), .B(new_n2552), .Y(n8179));
  xnor_4 g18734(.A(new_n14616), .B(new_n14613), .Y(n8215));
  xnor_4 g18735(.A(new_n18465), .B(new_n18458), .Y(n8267));
  xnor_4 g18736(.A(new_n19488), .B(new_n19487), .Y(n8276));
  not_8  g18737(.A(new_n21058), .Y(new_n21086));
  nor_5  g18738(.A(new_n21086), .B(n13783), .Y(new_n21087));
  not_8  g18739(.A(new_n21087), .Y(new_n21088));
  nor_5  g18740(.A(new_n21088), .B(n1654), .Y(new_n21089));
  not_8  g18741(.A(new_n21089), .Y(new_n21090));
  nor_5  g18742(.A(new_n21090), .B(n14440), .Y(new_n21091));
  xnor_4 g18743(.A(new_n21091), .B(n22626), .Y(new_n21092));
  nor_5  g18744(.A(new_n21092), .B(new_n14785), .Y(new_n21093_1));
  xnor_4 g18745(.A(new_n21092), .B(new_n14785), .Y(new_n21094_1));
  xnor_4 g18746(.A(new_n21089), .B(n14440), .Y(new_n21095_1));
  nor_5  g18747(.A(new_n21095_1), .B(new_n2969), .Y(new_n21096));
  xnor_4 g18748(.A(new_n21095_1), .B(new_n2969), .Y(new_n21097));
  xnor_4 g18749(.A(new_n21087), .B(n1654), .Y(new_n21098));
  and_5  g18750(.A(new_n21098), .B(new_n2973), .Y(new_n21099));
  and_5  g18751(.A(new_n21059), .B(new_n2981), .Y(new_n21100));
  nor_5  g18752(.A(new_n21068), .B(new_n21060), .Y(new_n21101));
  nor_5  g18753(.A(new_n21101), .B(new_n21100), .Y(new_n21102));
  xnor_4 g18754(.A(new_n21098), .B(new_n2973), .Y(new_n21103));
  nor_5  g18755(.A(new_n21103), .B(new_n21102), .Y(new_n21104));
  or_5   g18756(.A(new_n21104), .B(new_n21099), .Y(new_n21105));
  nor_5  g18757(.A(new_n21105), .B(new_n21097), .Y(new_n21106));
  nor_5  g18758(.A(new_n21106), .B(new_n21096), .Y(new_n21107));
  nor_5  g18759(.A(new_n21107), .B(new_n21094_1), .Y(new_n21108));
  nor_5  g18760(.A(new_n21108), .B(new_n21093_1), .Y(new_n21109));
  not_8  g18761(.A(new_n21091), .Y(new_n21110));
  nor_5  g18762(.A(new_n21110), .B(n22626), .Y(new_n21111));
  xnor_4 g18763(.A(new_n21111), .B(new_n14810), .Y(new_n21112));
  xnor_4 g18764(.A(new_n21112), .B(new_n21109), .Y(new_n21113));
  nor_5  g18765(.A(new_n21113), .B(new_n16852), .Y(new_n21114));
  xnor_4 g18766(.A(new_n21113), .B(new_n16852), .Y(new_n21115));
  xor_4  g18767(.A(new_n21107), .B(new_n21094_1), .Y(new_n21116));
  and_5  g18768(.A(new_n21116), .B(new_n16857), .Y(new_n21117));
  xnor_4 g18769(.A(new_n21116), .B(new_n16857), .Y(new_n21118));
  xor_4  g18770(.A(new_n21105), .B(new_n21097), .Y(new_n21119));
  and_5  g18771(.A(new_n21119), .B(new_n6833), .Y(new_n21120));
  xor_4  g18772(.A(new_n21103), .B(new_n21102), .Y(new_n21121));
  nor_5  g18773(.A(new_n21121), .B(new_n6913), .Y(new_n21122));
  xnor_4 g18774(.A(new_n21121), .B(new_n6913), .Y(new_n21123_1));
  nor_5  g18775(.A(new_n21069), .B(new_n6918), .Y(new_n21124));
  nor_5  g18776(.A(new_n21078_1), .B(new_n21070), .Y(new_n21125));
  nor_5  g18777(.A(new_n21125), .B(new_n21124), .Y(new_n21126));
  nor_5  g18778(.A(new_n21126), .B(new_n21123_1), .Y(new_n21127));
  nor_5  g18779(.A(new_n21127), .B(new_n21122), .Y(new_n21128));
  xnor_4 g18780(.A(new_n21119), .B(new_n6833), .Y(new_n21129));
  nor_5  g18781(.A(new_n21129), .B(new_n21128), .Y(new_n21130));
  nor_5  g18782(.A(new_n21130), .B(new_n21120), .Y(new_n21131));
  nor_5  g18783(.A(new_n21131), .B(new_n21118), .Y(new_n21132));
  nor_5  g18784(.A(new_n21132), .B(new_n21117), .Y(new_n21133));
  nor_5  g18785(.A(new_n21133), .B(new_n21115), .Y(new_n21134_1));
  nor_5  g18786(.A(new_n21134_1), .B(new_n21114), .Y(new_n21135));
  and_5  g18787(.A(new_n21135), .B(new_n16797), .Y(new_n21136));
  or_5   g18788(.A(new_n21111), .B(new_n14811), .Y(new_n21137));
  nor_5  g18789(.A(new_n21137), .B(new_n21109), .Y(new_n21138_1));
  or_5   g18790(.A(new_n21135), .B(new_n16797), .Y(new_n21139));
  and_5  g18791(.A(new_n21111), .B(new_n14811), .Y(new_n21140));
  and_5  g18792(.A(new_n21140), .B(new_n21109), .Y(new_n21141));
  nor_5  g18793(.A(new_n21141), .B(new_n21139), .Y(new_n21142));
  nor_5  g18794(.A(new_n21142), .B(new_n21138_1), .Y(new_n21143));
  nor_5  g18795(.A(new_n21143), .B(new_n21136), .Y(n8288));
  xnor_4 g18796(.A(new_n11147), .B(new_n7400), .Y(n8306));
  xor_4  g18797(.A(new_n7910), .B(new_n7857), .Y(n8320));
  xnor_4 g18798(.A(new_n12298), .B(new_n12279), .Y(n8321));
  xnor_4 g18799(.A(new_n16066), .B(new_n16053), .Y(n8339));
  xnor_4 g18800(.A(new_n9053), .B(new_n9009), .Y(n8376));
  not_8  g18801(.A(new_n10134), .Y(new_n21150));
  xnor_4 g18802(.A(new_n18769), .B(new_n21150), .Y(n8408));
  xnor_4 g18803(.A(new_n14145), .B(new_n14144), .Y(n8417));
  xnor_4 g18804(.A(new_n12722), .B(new_n12709), .Y(n8432));
  nor_5  g18805(.A(new_n10049), .B(new_n10045), .Y(new_n21154_1));
  and_5  g18806(.A(new_n10098), .B(new_n10051), .Y(new_n21155));
  nor_5  g18807(.A(new_n21155), .B(new_n21154_1), .Y(new_n21156));
  not_8  g18808(.A(new_n21156), .Y(new_n21157_1));
  and_5  g18809(.A(new_n21157_1), .B(new_n10028), .Y(new_n21158));
  nor_5  g18810(.A(new_n10099), .B(new_n10028), .Y(new_n21159));
  nor_5  g18811(.A(new_n10163), .B(new_n10100), .Y(new_n21160));
  nor_5  g18812(.A(new_n21160), .B(new_n21159), .Y(new_n21161));
  nor_5  g18813(.A(new_n21161), .B(new_n21158), .Y(new_n21162));
  nor_5  g18814(.A(new_n21157_1), .B(new_n10028), .Y(new_n21163));
  nor_5  g18815(.A(new_n21163), .B(new_n21160), .Y(new_n21164));
  nor_5  g18816(.A(new_n21164), .B(new_n21162), .Y(n8453));
  xnor_4 g18817(.A(new_n15345_1), .B(new_n13470), .Y(n8480));
  xnor_4 g18818(.A(new_n16219_1), .B(new_n16200), .Y(n8489));
  xnor_4 g18819(.A(new_n21048), .B(new_n21034_1), .Y(n8505));
  xnor_4 g18820(.A(new_n19184), .B(new_n19168), .Y(n8510));
  xnor_4 g18821(.A(new_n12002), .B(new_n8631), .Y(n8519));
  xnor_4 g18822(.A(new_n9689_1), .B(new_n9688), .Y(n8535));
  xnor_4 g18823(.A(new_n18917), .B(new_n18914), .Y(n8550));
  xnor_4 g18824(.A(new_n20051), .B(new_n20045), .Y(n8563));
  xnor_4 g18825(.A(new_n13131), .B(new_n13130), .Y(n8594));
  xnor_4 g18826(.A(new_n6954), .B(new_n6934), .Y(n8608));
  xnor_4 g18827(.A(new_n4585), .B(new_n4584), .Y(n8620));
  xnor_4 g18828(.A(new_n7423), .B(new_n7371), .Y(n8637));
  xnor_4 g18829(.A(new_n16870), .B(new_n16869), .Y(n8662));
  xnor_4 g18830(.A(new_n18512), .B(new_n18503), .Y(n8716));
  xnor_4 g18831(.A(new_n7861), .B(new_n7858), .Y(new_n21180));
  xnor_4 g18832(.A(new_n21180), .B(new_n7908), .Y(n8744));
  nor_5  g18833(.A(new_n12681), .B(new_n7772), .Y(new_n21182_1));
  or_5   g18834(.A(new_n20845), .B(new_n20840), .Y(new_n21183));
  and_5  g18835(.A(new_n21183), .B(new_n20839), .Y(new_n21184));
  nor_5  g18836(.A(new_n21184), .B(new_n21182_1), .Y(new_n21185));
  xnor_4 g18837(.A(new_n21185), .B(new_n15096), .Y(new_n21186));
  nor_5  g18838(.A(new_n6022_1), .B(new_n4907), .Y(new_n21187));
  and_5  g18839(.A(new_n20768), .B(new_n20765), .Y(new_n21188));
  nor_5  g18840(.A(new_n21188), .B(new_n21187), .Y(new_n21189));
  xnor_4 g18841(.A(new_n21189), .B(new_n17495), .Y(new_n21190));
  xnor_4 g18842(.A(new_n21190), .B(new_n21186), .Y(new_n21191));
  not_8  g18843(.A(new_n20769), .Y(new_n21192));
  not_8  g18844(.A(new_n20847), .Y(new_n21193_1));
  nor_5  g18845(.A(new_n21193_1), .B(new_n21192), .Y(new_n21194));
  xnor_4 g18846(.A(new_n20847), .B(new_n21192), .Y(new_n21195));
  nor_5  g18847(.A(new_n20851), .B(new_n20771), .Y(new_n21196));
  xnor_4 g18848(.A(new_n20851), .B(new_n15883), .Y(new_n21197));
  nor_5  g18849(.A(new_n17096), .B(new_n15885_1), .Y(new_n21198));
  nor_5  g18850(.A(new_n17128), .B(new_n17097), .Y(new_n21199));
  nor_5  g18851(.A(new_n21199), .B(new_n21198), .Y(new_n21200));
  and_5  g18852(.A(new_n21200), .B(new_n21197), .Y(new_n21201));
  nor_5  g18853(.A(new_n21201), .B(new_n21196), .Y(new_n21202));
  and_5  g18854(.A(new_n21202), .B(new_n21195), .Y(new_n21203_1));
  nor_5  g18855(.A(new_n21203_1), .B(new_n21194), .Y(new_n21204));
  xnor_4 g18856(.A(new_n21204), .B(new_n21191), .Y(n8803));
  and_5  g18857(.A(new_n19906), .B(new_n5500), .Y(new_n21206));
  nor_5  g18858(.A(new_n19907), .B(new_n5610), .Y(new_n21207));
  and_5  g18859(.A(new_n19926), .B(new_n19908), .Y(new_n21208));
  nor_5  g18860(.A(new_n21208), .B(new_n21207), .Y(new_n21209));
  xnor_4 g18861(.A(new_n21209), .B(new_n21206), .Y(new_n21210));
  nor_5  g18862(.A(n16544), .B(n4319), .Y(new_n21211));
  or_5   g18863(.A(new_n15561), .B(new_n15544), .Y(new_n21212));
  and_5  g18864(.A(new_n21212), .B(new_n15543), .Y(new_n21213));
  nor_5  g18865(.A(new_n21213), .B(new_n21211), .Y(new_n21214));
  xnor_4 g18866(.A(new_n21214), .B(new_n21210), .Y(new_n21215));
  nor_5  g18867(.A(new_n19927), .B(new_n15563), .Y(new_n21216));
  nor_5  g18868(.A(new_n19946), .B(new_n19928), .Y(new_n21217));
  nor_5  g18869(.A(new_n21217), .B(new_n21216), .Y(new_n21218));
  xnor_4 g18870(.A(new_n21218), .B(new_n21215), .Y(new_n21219));
  not_8  g18871(.A(new_n21219), .Y(new_n21220));
  xnor_4 g18872(.A(new_n21220), .B(new_n7695), .Y(new_n21221));
  nor_5  g18873(.A(new_n20501), .B(new_n7698_1), .Y(new_n21222_1));
  nor_5  g18874(.A(new_n20536), .B(new_n20502), .Y(new_n21223));
  nor_5  g18875(.A(new_n21223), .B(new_n21222_1), .Y(new_n21224));
  xnor_4 g18876(.A(new_n21224), .B(new_n21221), .Y(n8809));
  nor_5  g18877(.A(new_n21189), .B(new_n17496), .Y(new_n21226_1));
  not_8  g18878(.A(new_n21226_1), .Y(new_n21227));
  nor_5  g18879(.A(new_n17831), .B(n3324), .Y(new_n21228));
  and_5  g18880(.A(new_n20763), .B(new_n20752), .Y(new_n21229));
  nor_5  g18881(.A(new_n21229), .B(new_n21228), .Y(new_n21230));
  and_5  g18882(.A(new_n21230), .B(new_n17825), .Y(new_n21231));
  xnor_4 g18883(.A(new_n21231), .B(new_n21227), .Y(new_n21232));
  not_8  g18884(.A(new_n21190), .Y(new_n21233));
  xnor_4 g18885(.A(new_n21230), .B(new_n17823), .Y(new_n21234));
  nor_5  g18886(.A(new_n21234), .B(new_n21233), .Y(new_n21235));
  xnor_4 g18887(.A(new_n21234), .B(new_n21233), .Y(new_n21236));
  nor_5  g18888(.A(new_n20769), .B(new_n20764), .Y(new_n21237));
  nor_5  g18889(.A(new_n20784), .B(new_n20770), .Y(new_n21238_1));
  nor_5  g18890(.A(new_n21238_1), .B(new_n21237), .Y(new_n21239));
  nor_5  g18891(.A(new_n21239), .B(new_n21236), .Y(new_n21240));
  nor_5  g18892(.A(new_n21240), .B(new_n21235), .Y(new_n21241));
  xnor_4 g18893(.A(new_n21241), .B(new_n21232), .Y(n8821));
  xnor_4 g18894(.A(new_n15315), .B(new_n15314), .Y(n8824));
  xor_4  g18895(.A(new_n17446), .B(new_n17445), .Y(n8849));
  xnor_4 g18896(.A(new_n13582), .B(new_n13574), .Y(n8861));
  xnor_4 g18897(.A(n22442), .B(n8856), .Y(new_n21246));
  nor_5  g18898(.A(n14130), .B(new_n8273), .Y(new_n21247));
  and_5  g18899(.A(new_n19702), .B(new_n19679), .Y(new_n21248));
  or_5   g18900(.A(new_n21248), .B(new_n21247), .Y(new_n21249));
  xor_4  g18901(.A(new_n21249), .B(new_n21246), .Y(new_n21250));
  xnor_4 g18902(.A(n3324), .B(new_n7179), .Y(new_n21251));
  nor_5  g18903(.A(n25331), .B(n17911), .Y(new_n21252));
  and_5  g18904(.A(new_n19672), .B(new_n19669), .Y(new_n21253));
  or_5   g18905(.A(new_n21253), .B(new_n21252), .Y(new_n21254_1));
  xor_4  g18906(.A(new_n21254_1), .B(new_n21251), .Y(new_n21255));
  xnor_4 g18907(.A(new_n21255), .B(new_n7522), .Y(new_n21256));
  nor_5  g18908(.A(new_n19673), .B(new_n7488), .Y(new_n21257));
  and_5  g18909(.A(new_n19677), .B(new_n19674), .Y(new_n21258));
  nor_5  g18910(.A(new_n21258), .B(new_n21257), .Y(new_n21259));
  xnor_4 g18911(.A(new_n21259), .B(new_n21256), .Y(new_n21260));
  xnor_4 g18912(.A(new_n21260), .B(new_n21250), .Y(new_n21261));
  and_5  g18913(.A(new_n19703), .B(new_n19678), .Y(new_n21262));
  and_5  g18914(.A(new_n19733), .B(new_n19704), .Y(new_n21263));
  or_5   g18915(.A(new_n21263), .B(new_n21262), .Y(new_n21264));
  xor_4  g18916(.A(new_n21264), .B(new_n21261), .Y(n8862));
  xor_4  g18917(.A(new_n13476), .B(new_n13475), .Y(n8884));
  not_8  g18918(.A(new_n17910), .Y(new_n21267));
  xnor_4 g18919(.A(new_n18681), .B(new_n21267), .Y(n8909));
  xnor_4 g18920(.A(new_n11578), .B(new_n11537), .Y(n8911));
  xnor_4 g18921(.A(new_n11088), .B(new_n11087), .Y(n8971));
  xnor_4 g18922(.A(new_n20929_1), .B(new_n20906), .Y(n8982));
  xnor_4 g18923(.A(new_n5441), .B(new_n5425), .Y(n8993));
  xor_4  g18924(.A(new_n14154), .B(new_n14153), .Y(n9012));
  nor_5  g18925(.A(new_n19824), .B(new_n19821), .Y(new_n21274));
  or_5   g18926(.A(new_n19831), .B(new_n4453), .Y(new_n21275));
  nor_5  g18927(.A(new_n21275), .B(new_n19829), .Y(new_n21276_1));
  xnor_4 g18928(.A(new_n21276_1), .B(new_n21274), .Y(new_n21277));
  nor_5  g18929(.A(new_n19833), .B(new_n19825), .Y(new_n21278));
  nor_5  g18930(.A(new_n19879), .B(new_n19834), .Y(new_n21279));
  nor_5  g18931(.A(new_n21279), .B(new_n21278), .Y(new_n21280));
  xnor_4 g18932(.A(new_n21280), .B(new_n21277), .Y(n9032));
  xor_4  g18933(.A(new_n15808), .B(new_n15807), .Y(n9042));
  xnor_4 g18934(.A(new_n17074), .B(new_n17043), .Y(n9046));
  xnor_4 g18935(.A(new_n8200), .B(new_n8142), .Y(n9047));
  xnor_4 g18936(.A(new_n15035), .B(new_n15034), .Y(n9104));
  nor_5  g18937(.A(new_n20201), .B(new_n20193), .Y(new_n21286));
  nor_5  g18938(.A(new_n21286), .B(new_n20185), .Y(new_n21287_1));
  and_5  g18939(.A(new_n20201), .B(new_n20193), .Y(new_n21288));
  nor_5  g18940(.A(new_n21288), .B(new_n15180_1), .Y(new_n21289));
  nor_5  g18941(.A(new_n21289), .B(new_n21287_1), .Y(new_n21290));
  not_8  g18942(.A(new_n21290), .Y(new_n21291));
  xnor_4 g18943(.A(new_n21291), .B(new_n19127), .Y(new_n21292));
  nor_5  g18944(.A(new_n20203), .B(new_n19127), .Y(new_n21293));
  nor_5  g18945(.A(new_n20212), .B(new_n20204), .Y(new_n21294));
  nor_5  g18946(.A(new_n21294), .B(new_n21293), .Y(new_n21295));
  xor_4  g18947(.A(new_n21295), .B(new_n21292), .Y(n9129));
  xnor_4 g18948(.A(new_n18858_1), .B(new_n18827), .Y(n9146));
  xnor_4 g18949(.A(new_n8631), .B(new_n6702), .Y(n9164));
  xor_4  g18950(.A(new_n12647), .B(new_n12646), .Y(n9166));
  xnor_4 g18951(.A(new_n17842), .B(new_n17815), .Y(new_n21300));
  xnor_4 g18952(.A(new_n21300), .B(new_n17853), .Y(n9182));
  xnor_4 g18953(.A(new_n7168), .B(new_n7136), .Y(n9191));
  xnor_4 g18954(.A(new_n11583), .B(new_n11528), .Y(n9217));
  xor_4  g18955(.A(new_n15969), .B(new_n15968), .Y(n9220));
  xnor_4 g18956(.A(new_n18848), .B(new_n18842), .Y(n9261));
  xnor_4 g18957(.A(n22626), .B(n3324), .Y(new_n21306));
  nor_5  g18958(.A(new_n19668), .B(n14440), .Y(new_n21307));
  and_5  g18959(.A(new_n18491), .B(new_n18471), .Y(new_n21308));
  or_5   g18960(.A(new_n21308), .B(new_n21307), .Y(new_n21309));
  xor_4  g18961(.A(new_n21309), .B(new_n21306), .Y(new_n21310));
  and_5  g18962(.A(new_n21310), .B(new_n17846), .Y(new_n21311));
  xnor_4 g18963(.A(new_n21310), .B(new_n17846), .Y(new_n21312));
  and_5  g18964(.A(new_n18492), .B(new_n3032), .Y(new_n21313));
  and_5  g18965(.A(new_n18518), .B(new_n18493), .Y(new_n21314));
  nor_5  g18966(.A(new_n21314), .B(new_n21313), .Y(new_n21315));
  nor_5  g18967(.A(new_n21315), .B(new_n21312), .Y(new_n21316));
  nor_5  g18968(.A(new_n21316), .B(new_n21311), .Y(new_n21317_1));
  not_8  g18969(.A(new_n21317_1), .Y(new_n21318));
  nor_5  g18970(.A(n22626), .B(new_n20751), .Y(new_n21319));
  and_5  g18971(.A(new_n21309), .B(new_n21306), .Y(new_n21320));
  nor_5  g18972(.A(new_n21320), .B(new_n21319), .Y(new_n21321));
  xnor_4 g18973(.A(new_n21321), .B(new_n17842), .Y(new_n21322));
  xnor_4 g18974(.A(new_n21322), .B(new_n21318), .Y(n9287));
  xor_4  g18975(.A(new_n13974), .B(new_n13965), .Y(n9308));
  xnor_4 g18976(.A(new_n5020_1), .B(new_n4983), .Y(n9344));
  xnor_4 g18977(.A(new_n3711), .B(new_n3694), .Y(n9364));
  or_5   g18978(.A(new_n21321), .B(new_n17841), .Y(new_n21327));
  nor_5  g18979(.A(new_n21327), .B(new_n21317_1), .Y(new_n21328));
  and_5  g18980(.A(new_n21328), .B(new_n17839), .Y(new_n21329));
  and_5  g18981(.A(new_n21321), .B(new_n17841), .Y(new_n21330));
  and_5  g18982(.A(new_n21330), .B(new_n21317_1), .Y(new_n21331));
  and_5  g18983(.A(new_n21331), .B(new_n17857), .Y(new_n21332));
  or_5   g18984(.A(new_n21332), .B(new_n21329), .Y(n9371));
  xnor_4 g18985(.A(new_n10135), .B(new_n21150), .Y(n9382));
  xor_4  g18986(.A(new_n20967), .B(new_n20958), .Y(n9403));
  xnor_4 g18987(.A(new_n12653), .B(new_n12628), .Y(n9419));
  xnor_4 g18988(.A(new_n20732), .B(new_n20709_1), .Y(n9423));
  xnor_4 g18989(.A(new_n18514), .B(new_n18499), .Y(n9430));
  xnor_4 g18990(.A(n25120), .B(n23272), .Y(new_n21339));
  and_5  g18991(.A(new_n4361), .B(n8363), .Y(new_n21340));
  xnor_4 g18992(.A(n11481), .B(n8363), .Y(new_n21341));
  and_5  g18993(.A(new_n4365), .B(n14680), .Y(new_n21342));
  and_5  g18994(.A(new_n15485), .B(new_n15482), .Y(new_n21343));
  or_5   g18995(.A(new_n21343), .B(new_n21342), .Y(new_n21344));
  and_5  g18996(.A(new_n21344), .B(new_n21341), .Y(new_n21345));
  or_5   g18997(.A(new_n21345), .B(new_n21340), .Y(new_n21346));
  xor_4  g18998(.A(new_n21346), .B(new_n21339), .Y(new_n21347));
  xnor_4 g18999(.A(new_n21347), .B(new_n16950), .Y(new_n21348));
  xor_4  g19000(.A(new_n21344), .B(new_n21341), .Y(new_n21349_1));
  and_5  g19001(.A(new_n21349_1), .B(new_n16974), .Y(new_n21350));
  xnor_4 g19002(.A(new_n21349_1), .B(new_n16974), .Y(new_n21351));
  and_5  g19003(.A(new_n15492), .B(new_n15486), .Y(new_n21352));
  nor_5  g19004(.A(new_n15496_1), .B(new_n15493), .Y(new_n21353));
  nor_5  g19005(.A(new_n21353), .B(new_n21352), .Y(new_n21354));
  nor_5  g19006(.A(new_n21354), .B(new_n21351), .Y(new_n21355));
  nor_5  g19007(.A(new_n21355), .B(new_n21350), .Y(new_n21356));
  xor_4  g19008(.A(new_n21356), .B(new_n21348), .Y(new_n21357));
  xnor_4 g19009(.A(new_n21357), .B(new_n17024), .Y(new_n21358));
  xor_4  g19010(.A(new_n21354), .B(new_n21351), .Y(new_n21359));
  nor_5  g19011(.A(new_n21359), .B(new_n17026), .Y(new_n21360));
  xnor_4 g19012(.A(new_n21359), .B(new_n17026), .Y(new_n21361));
  nor_5  g19013(.A(new_n17032), .B(new_n15498), .Y(new_n21362));
  xnor_4 g19014(.A(new_n17032), .B(new_n15498), .Y(new_n21363));
  nor_5  g19015(.A(new_n17039), .B(new_n10576), .Y(new_n21364));
  xnor_4 g19016(.A(new_n17039), .B(new_n10576), .Y(new_n21365_1));
  nor_5  g19017(.A(new_n17048), .B(new_n10578), .Y(new_n21366));
  xnor_4 g19018(.A(new_n17048), .B(new_n10578), .Y(new_n21367_1));
  nor_5  g19019(.A(new_n17054), .B(new_n10582), .Y(new_n21368));
  and_5  g19020(.A(new_n14764), .B(new_n10584), .Y(new_n21369));
  nor_5  g19021(.A(new_n14777), .B(new_n14765), .Y(new_n21370));
  nor_5  g19022(.A(new_n21370), .B(new_n21369), .Y(new_n21371));
  xnor_4 g19023(.A(new_n17051), .B(new_n10600), .Y(new_n21372));
  nor_5  g19024(.A(new_n21372), .B(new_n21371), .Y(new_n21373));
  or_5   g19025(.A(new_n21373), .B(new_n21368), .Y(new_n21374));
  nor_5  g19026(.A(new_n21374), .B(new_n21367_1), .Y(new_n21375));
  nor_5  g19027(.A(new_n21375), .B(new_n21366), .Y(new_n21376));
  nor_5  g19028(.A(new_n21376), .B(new_n21365_1), .Y(new_n21377));
  nor_5  g19029(.A(new_n21377), .B(new_n21364), .Y(new_n21378));
  nor_5  g19030(.A(new_n21378), .B(new_n21363), .Y(new_n21379));
  nor_5  g19031(.A(new_n21379), .B(new_n21362), .Y(new_n21380));
  nor_5  g19032(.A(new_n21380), .B(new_n21361), .Y(new_n21381));
  or_5   g19033(.A(new_n21381), .B(new_n21360), .Y(new_n21382));
  xor_4  g19034(.A(new_n21382), .B(new_n21358), .Y(n9435));
  xnor_4 g19035(.A(new_n15919), .B(new_n15891), .Y(n9451));
  xnor_4 g19036(.A(n12657), .B(n10763), .Y(new_n21385));
  nor_5  g19037(.A(n17077), .B(new_n2890), .Y(new_n21386));
  and_5  g19038(.A(new_n18974), .B(new_n18967), .Y(new_n21387));
  or_5   g19039(.A(new_n21387), .B(new_n21386), .Y(new_n21388));
  xor_4  g19040(.A(new_n21388), .B(new_n21385), .Y(new_n21389));
  xnor_4 g19041(.A(new_n21389), .B(new_n19678), .Y(new_n21390));
  nor_5  g19042(.A(new_n18995), .B(new_n18975), .Y(new_n21391));
  and_5  g19043(.A(new_n19007), .B(new_n18997), .Y(new_n21392));
  nor_5  g19044(.A(new_n21392), .B(new_n21391), .Y(new_n21393));
  xnor_4 g19045(.A(new_n21393), .B(new_n21390), .Y(n9458));
  nor_5  g19046(.A(n12507), .B(new_n10030), .Y(new_n21395));
  xnor_4 g19047(.A(n12507), .B(n11220), .Y(new_n21396_1));
  nor_5  g19048(.A(new_n17810), .B(n15077), .Y(new_n21397));
  and_5  g19049(.A(new_n14702_1), .B(new_n14683), .Y(new_n21398_1));
  or_5   g19050(.A(new_n21398_1), .B(new_n21397), .Y(new_n21399_1));
  and_5  g19051(.A(new_n21399_1), .B(new_n21396_1), .Y(new_n21400));
  nor_5  g19052(.A(new_n21400), .B(new_n21395), .Y(new_n21401));
  not_8  g19053(.A(new_n21401), .Y(new_n21402));
  xnor_4 g19054(.A(new_n21402), .B(new_n20401), .Y(new_n21403));
  xor_4  g19055(.A(new_n21399_1), .B(new_n21396_1), .Y(new_n21404_1));
  nor_5  g19056(.A(new_n21404_1), .B(new_n20403_1), .Y(new_n21405));
  xnor_4 g19057(.A(new_n21404_1), .B(new_n20403_1), .Y(new_n21406));
  nor_5  g19058(.A(new_n14703), .B(new_n14682), .Y(new_n21407));
  nor_5  g19059(.A(new_n14734_1), .B(new_n14704_1), .Y(new_n21408));
  nor_5  g19060(.A(new_n21408), .B(new_n21407), .Y(new_n21409));
  nor_5  g19061(.A(new_n21409), .B(new_n21406), .Y(new_n21410));
  nor_5  g19062(.A(new_n21410), .B(new_n21405), .Y(new_n21411));
  xnor_4 g19063(.A(new_n21411), .B(new_n21403), .Y(n9459));
  xnor_4 g19064(.A(new_n14977_1), .B(new_n14976), .Y(n9508));
  xnor_4 g19065(.A(new_n12657_1), .B(new_n12619), .Y(n9552));
  xnor_4 g19066(.A(new_n4588_1), .B(new_n4587), .Y(n9556));
  xnor_4 g19067(.A(new_n11060), .B(new_n8832), .Y(n9558));
  xnor_4 g19068(.A(new_n20604_1), .B(new_n14145), .Y(n9616));
  xnor_4 g19069(.A(new_n8566), .B(new_n8539), .Y(n9622));
  xnor_4 g19070(.A(new_n16412), .B(new_n16397), .Y(n9626));
  xnor_4 g19071(.A(new_n4594), .B(new_n4576), .Y(n9633));
  not_8  g19072(.A(n23272), .Y(new_n21421));
  and_5  g19073(.A(n25120), .B(new_n21421), .Y(new_n21422));
  and_5  g19074(.A(new_n21346), .B(new_n21339), .Y(new_n21423));
  nor_5  g19075(.A(new_n21423), .B(new_n21422), .Y(new_n21424));
  not_8  g19076(.A(new_n21424), .Y(new_n21425));
  nor_5  g19077(.A(new_n21425), .B(new_n20941), .Y(new_n21426));
  xnor_4 g19078(.A(new_n21424), .B(new_n20941), .Y(new_n21427));
  and_5  g19079(.A(new_n21347), .B(new_n16950), .Y(new_n21428));
  nor_5  g19080(.A(new_n21356), .B(new_n21348), .Y(new_n21429));
  nor_5  g19081(.A(new_n21429), .B(new_n21428), .Y(new_n21430));
  and_5  g19082(.A(new_n21430), .B(new_n21427), .Y(new_n21431));
  nor_5  g19083(.A(new_n21431), .B(new_n21426), .Y(new_n21432));
  not_8  g19084(.A(new_n21432), .Y(new_n21433));
  nor_5  g19085(.A(new_n21433), .B(new_n5542), .Y(new_n21434));
  xnor_4 g19086(.A(new_n21433), .B(new_n10165_1), .Y(new_n21435));
  xnor_4 g19087(.A(new_n21430), .B(new_n21427), .Y(new_n21436));
  not_8  g19088(.A(new_n21436), .Y(new_n21437));
  nor_5  g19089(.A(new_n21437), .B(new_n10165_1), .Y(new_n21438));
  xnor_4 g19090(.A(new_n21437), .B(new_n10165_1), .Y(new_n21439));
  nor_5  g19091(.A(new_n21357), .B(new_n5544), .Y(new_n21440));
  and_5  g19092(.A(new_n21359), .B(new_n5619), .Y(new_n21441));
  xnor_4 g19093(.A(new_n21359), .B(new_n5619), .Y(new_n21442));
  nor_5  g19094(.A(new_n15497), .B(new_n5626), .Y(new_n21443));
  nor_5  g19095(.A(new_n15502), .B(new_n15499), .Y(new_n21444));
  nor_5  g19096(.A(new_n21444), .B(new_n21443), .Y(new_n21445));
  nor_5  g19097(.A(new_n21445), .B(new_n21442), .Y(new_n21446_1));
  or_5   g19098(.A(new_n21446_1), .B(new_n21441), .Y(new_n21447));
  xnor_4 g19099(.A(new_n21357), .B(new_n5544), .Y(new_n21448));
  nor_5  g19100(.A(new_n21448), .B(new_n21447), .Y(new_n21449));
  or_5   g19101(.A(new_n21449), .B(new_n21440), .Y(new_n21450));
  nor_5  g19102(.A(new_n21450), .B(new_n21439), .Y(new_n21451));
  or_5   g19103(.A(new_n21451), .B(new_n21438), .Y(new_n21452));
  and_5  g19104(.A(new_n21452), .B(new_n21435), .Y(new_n21453));
  nor_5  g19105(.A(new_n21453), .B(new_n21434), .Y(n9635));
  xnor_4 g19106(.A(new_n19208), .B(new_n19205), .Y(n9648));
  xnor_4 g19107(.A(new_n16081), .B(new_n5003), .Y(n9689));
  xnor_4 g19108(.A(new_n10765), .B(new_n10747), .Y(n9695));
  xnor_4 g19109(.A(new_n7600), .B(new_n7560), .Y(n9699));
  xnor_4 g19110(.A(new_n16500), .B(new_n14513), .Y(new_n21459));
  nor_5  g19111(.A(new_n16503), .B(new_n14513), .Y(new_n21460));
  nor_5  g19112(.A(new_n15975), .B(new_n15937), .Y(new_n21461));
  nor_5  g19113(.A(new_n21461), .B(new_n21460), .Y(new_n21462));
  xor_4  g19114(.A(new_n21462), .B(new_n21459), .Y(n9726));
  xnor_4 g19115(.A(new_n13142), .B(new_n9963), .Y(n9753));
  xnor_4 g19116(.A(new_n3379), .B(new_n3360), .Y(n9761));
  xnor_4 g19117(.A(new_n9978), .B(new_n9931), .Y(n9763));
  xnor_4 g19118(.A(new_n13473), .B(new_n13472), .Y(n9767));
  xnor_4 g19119(.A(new_n13628), .B(new_n13376), .Y(n9771));
  xor_4  g19120(.A(new_n21044), .B(new_n21041), .Y(n9778));
  xnor_4 g19121(.A(new_n15705), .B(new_n15696), .Y(n9783));
  xnor_4 g19122(.A(new_n6735), .B(new_n6733), .Y(n9803));
  and_5  g19123(.A(new_n20545), .B(new_n11610), .Y(new_n21472_1));
  and_5  g19124(.A(new_n21472_1), .B(new_n3087), .Y(new_n21473));
  xnor_4 g19125(.A(new_n21472_1), .B(n4319), .Y(new_n21474));
  not_8  g19126(.A(new_n21474), .Y(new_n21475));
  nor_5  g19127(.A(new_n21475), .B(new_n17789), .Y(new_n21476));
  nor_5  g19128(.A(new_n21474), .B(new_n17788), .Y(new_n21477));
  nor_5  g19129(.A(new_n20547), .B(new_n17793), .Y(new_n21478));
  and_5  g19130(.A(new_n20547), .B(new_n17793), .Y(new_n21479));
  and_5  g19131(.A(new_n20549), .B(new_n16564), .Y(new_n21480));
  or_5   g19132(.A(new_n20549), .B(new_n16564), .Y(new_n21481));
  nor_5  g19133(.A(new_n20553), .B(new_n16567), .Y(new_n21482));
  nor_5  g19134(.A(new_n20558), .B(new_n16570), .Y(new_n21483));
  xnor_4 g19135(.A(new_n20556), .B(new_n16571), .Y(new_n21484));
  and_5  g19136(.A(new_n6696), .B(new_n6680), .Y(new_n21485));
  nor_5  g19137(.A(new_n6720), .B(new_n6697), .Y(new_n21486));
  nor_5  g19138(.A(new_n21486), .B(new_n21485), .Y(new_n21487));
  nor_5  g19139(.A(new_n21487), .B(new_n21484), .Y(new_n21488));
  nor_5  g19140(.A(new_n21488), .B(new_n21483), .Y(new_n21489_1));
  xor_4  g19141(.A(new_n20553), .B(new_n16567), .Y(new_n21490));
  and_5  g19142(.A(new_n21490), .B(new_n21489_1), .Y(new_n21491));
  nor_5  g19143(.A(new_n21491), .B(new_n21482), .Y(new_n21492));
  and_5  g19144(.A(new_n21492), .B(new_n21481), .Y(new_n21493));
  nor_5  g19145(.A(new_n21493), .B(new_n21480), .Y(new_n21494));
  nor_5  g19146(.A(new_n21494), .B(new_n21479), .Y(new_n21495));
  nor_5  g19147(.A(new_n21495), .B(new_n21478), .Y(new_n21496));
  nor_5  g19148(.A(new_n21496), .B(new_n21477), .Y(new_n21497));
  nor_5  g19149(.A(new_n21497), .B(new_n21476), .Y(new_n21498));
  xnor_4 g19150(.A(new_n21498), .B(new_n17784_1), .Y(new_n21499));
  xnor_4 g19151(.A(new_n21499), .B(new_n21473), .Y(new_n21500));
  nor_5  g19152(.A(new_n21500), .B(new_n3327), .Y(new_n21501));
  xnor_4 g19153(.A(new_n21500), .B(new_n3327), .Y(new_n21502));
  xnor_4 g19154(.A(new_n21474), .B(new_n17789), .Y(new_n21503));
  xnor_4 g19155(.A(new_n21503), .B(new_n21496), .Y(new_n21504));
  nor_5  g19156(.A(new_n21504), .B(new_n3334), .Y(new_n21505));
  xnor_4 g19157(.A(new_n21504), .B(new_n3334), .Y(new_n21506));
  xnor_4 g19158(.A(new_n20546), .B(new_n17793), .Y(new_n21507));
  xnor_4 g19159(.A(new_n21507), .B(new_n21494), .Y(new_n21508));
  nor_5  g19160(.A(new_n21508), .B(new_n3338), .Y(new_n21509));
  xnor_4 g19161(.A(new_n21508), .B(new_n3338), .Y(new_n21510));
  xnor_4 g19162(.A(new_n20549), .B(new_n16564), .Y(new_n21511));
  xnor_4 g19163(.A(new_n21511), .B(new_n21492), .Y(new_n21512));
  nor_5  g19164(.A(new_n21512), .B(new_n3342), .Y(new_n21513));
  xnor_4 g19165(.A(new_n21512), .B(new_n3342), .Y(new_n21514));
  xnor_4 g19166(.A(new_n21490), .B(new_n21489_1), .Y(new_n21515));
  nor_5  g19167(.A(new_n21515), .B(new_n3346), .Y(new_n21516));
  xnor_4 g19168(.A(new_n21515), .B(new_n3346), .Y(new_n21517));
  xor_4  g19169(.A(new_n21487), .B(new_n21484), .Y(new_n21518));
  nor_5  g19170(.A(new_n21518), .B(new_n3350), .Y(new_n21519));
  xnor_4 g19171(.A(new_n21518), .B(new_n3350), .Y(new_n21520));
  nor_5  g19172(.A(new_n6721), .B(new_n3354), .Y(new_n21521));
  nor_5  g19173(.A(new_n6742), .B(new_n6722), .Y(new_n21522));
  nor_5  g19174(.A(new_n21522), .B(new_n21521), .Y(new_n21523));
  nor_5  g19175(.A(new_n21523), .B(new_n21520), .Y(new_n21524));
  nor_5  g19176(.A(new_n21524), .B(new_n21519), .Y(new_n21525_1));
  nor_5  g19177(.A(new_n21525_1), .B(new_n21517), .Y(new_n21526));
  nor_5  g19178(.A(new_n21526), .B(new_n21516), .Y(new_n21527));
  nor_5  g19179(.A(new_n21527), .B(new_n21514), .Y(new_n21528));
  nor_5  g19180(.A(new_n21528), .B(new_n21513), .Y(new_n21529));
  nor_5  g19181(.A(new_n21529), .B(new_n21510), .Y(new_n21530));
  nor_5  g19182(.A(new_n21530), .B(new_n21509), .Y(new_n21531));
  nor_5  g19183(.A(new_n21531), .B(new_n21506), .Y(new_n21532));
  nor_5  g19184(.A(new_n21532), .B(new_n21505), .Y(new_n21533));
  nor_5  g19185(.A(new_n21533), .B(new_n21502), .Y(new_n21534));
  nor_5  g19186(.A(new_n21534), .B(new_n21501), .Y(new_n21535));
  not_8  g19187(.A(new_n21498), .Y(new_n21536));
  nor_5  g19188(.A(new_n21536), .B(new_n17784_1), .Y(new_n21537));
  xnor_4 g19189(.A(new_n21473), .B(new_n17744), .Y(new_n21538_1));
  and_5  g19190(.A(new_n21538_1), .B(new_n21537), .Y(new_n21539));
  nor_5  g19191(.A(new_n21538_1), .B(new_n21498), .Y(new_n21540));
  nor_5  g19192(.A(new_n21540), .B(new_n21539), .Y(new_n21541));
  and_5  g19193(.A(new_n21541), .B(new_n21535), .Y(new_n21542));
  or_5   g19194(.A(new_n21473), .B(new_n17745), .Y(new_n21543));
  nor_5  g19195(.A(new_n21543), .B(new_n21536), .Y(new_n21544));
  xor_4  g19196(.A(new_n21544), .B(new_n21542), .Y(n9833));
  not_8  g19197(.A(new_n17217), .Y(new_n21546));
  nor_5  g19198(.A(new_n21546), .B(n13775), .Y(new_n21547));
  and_5  g19199(.A(new_n21547), .B(new_n8646), .Y(new_n21548));
  and_5  g19200(.A(new_n21548), .B(new_n11842_1), .Y(new_n21549_1));
  or_5   g19201(.A(new_n21549_1), .B(new_n17781), .Y(new_n21550));
  xnor_4 g19202(.A(new_n21548), .B(n25972), .Y(new_n21551));
  and_5  g19203(.A(new_n21551), .B(new_n17760), .Y(new_n21552));
  xnor_4 g19204(.A(new_n21551), .B(new_n17760), .Y(new_n21553));
  xnor_4 g19205(.A(new_n21547), .B(n21915), .Y(new_n21554));
  and_5  g19206(.A(new_n21554), .B(new_n17765), .Y(new_n21555));
  xnor_4 g19207(.A(new_n21554), .B(new_n17764), .Y(new_n21556));
  and_5  g19208(.A(new_n17218), .B(new_n16534), .Y(new_n21557));
  and_5  g19209(.A(new_n17248), .B(new_n17219_1), .Y(new_n21558));
  or_5   g19210(.A(new_n21558), .B(new_n21557), .Y(new_n21559));
  and_5  g19211(.A(new_n21559), .B(new_n21556), .Y(new_n21560));
  nor_5  g19212(.A(new_n21560), .B(new_n21555), .Y(new_n21561));
  nor_5  g19213(.A(new_n21561), .B(new_n21553), .Y(new_n21562));
  nor_5  g19214(.A(new_n21562), .B(new_n21552), .Y(new_n21563));
  not_8  g19215(.A(new_n21563), .Y(new_n21564));
  nor_5  g19216(.A(new_n21564), .B(new_n21550), .Y(new_n21565));
  not_8  g19217(.A(new_n17251_1), .Y(new_n21566));
  nor_5  g19218(.A(new_n21566), .B(n3710), .Y(new_n21567));
  and_5  g19219(.A(new_n21567), .B(new_n8789), .Y(new_n21568));
  and_5  g19220(.A(new_n21568), .B(new_n8719), .Y(new_n21569));
  xnor_4 g19221(.A(new_n21569), .B(new_n16496), .Y(new_n21570));
  xnor_4 g19222(.A(new_n21568), .B(n12507), .Y(new_n21571));
  nor_5  g19223(.A(new_n21571), .B(new_n12818), .Y(new_n21572));
  xnor_4 g19224(.A(new_n21567), .B(n15077), .Y(new_n21573));
  nor_5  g19225(.A(new_n21573), .B(new_n5304), .Y(new_n21574));
  xnor_4 g19226(.A(new_n21573), .B(new_n5304), .Y(new_n21575));
  and_5  g19227(.A(new_n17252), .B(new_n5341), .Y(new_n21576));
  and_5  g19228(.A(new_n17256), .B(new_n17253), .Y(new_n21577));
  nor_5  g19229(.A(new_n21577), .B(new_n21576), .Y(new_n21578));
  not_8  g19230(.A(new_n21578), .Y(new_n21579));
  nor_5  g19231(.A(new_n21579), .B(new_n21575), .Y(new_n21580));
  nor_5  g19232(.A(new_n21580), .B(new_n21574), .Y(new_n21581));
  xnor_4 g19233(.A(new_n21571), .B(new_n12818), .Y(new_n21582));
  nor_5  g19234(.A(new_n21582), .B(new_n21581), .Y(new_n21583));
  nor_5  g19235(.A(new_n21583), .B(new_n21572), .Y(new_n21584));
  xnor_4 g19236(.A(new_n21584), .B(new_n21570), .Y(new_n21585));
  xnor_4 g19237(.A(new_n21549_1), .B(new_n17782), .Y(new_n21586));
  xnor_4 g19238(.A(new_n21586), .B(new_n21564), .Y(new_n21587));
  nor_5  g19239(.A(new_n21587), .B(new_n21585), .Y(new_n21588));
  xnor_4 g19240(.A(new_n21587), .B(new_n21585), .Y(new_n21589));
  xnor_4 g19241(.A(new_n21561), .B(new_n21553), .Y(new_n21590));
  xnor_4 g19242(.A(new_n21582), .B(new_n21581), .Y(new_n21591));
  not_8  g19243(.A(new_n21591), .Y(new_n21592));
  and_5  g19244(.A(new_n21592), .B(new_n21590), .Y(new_n21593));
  xnor_4 g19245(.A(new_n21592), .B(new_n21590), .Y(new_n21594));
  xnor_4 g19246(.A(new_n21578), .B(new_n21575), .Y(new_n21595));
  not_8  g19247(.A(new_n21595), .Y(new_n21596));
  xor_4  g19248(.A(new_n21559), .B(new_n21556), .Y(new_n21597));
  nor_5  g19249(.A(new_n21597), .B(new_n21596), .Y(new_n21598));
  xnor_4 g19250(.A(new_n21597), .B(new_n21596), .Y(new_n21599_1));
  nor_5  g19251(.A(new_n17257), .B(new_n17249), .Y(new_n21600));
  nor_5  g19252(.A(new_n17291), .B(new_n17258), .Y(new_n21601));
  nor_5  g19253(.A(new_n21601), .B(new_n21600), .Y(new_n21602));
  nor_5  g19254(.A(new_n21602), .B(new_n21599_1), .Y(new_n21603));
  nor_5  g19255(.A(new_n21603), .B(new_n21598), .Y(new_n21604));
  nor_5  g19256(.A(new_n21604), .B(new_n21594), .Y(new_n21605));
  nor_5  g19257(.A(new_n21605), .B(new_n21593), .Y(new_n21606));
  nor_5  g19258(.A(new_n21606), .B(new_n21589), .Y(new_n21607));
  or_5   g19259(.A(new_n21607), .B(new_n21588), .Y(new_n21608));
  and_5  g19260(.A(new_n21608), .B(new_n21565), .Y(new_n21609));
  xor_4  g19261(.A(new_n21608), .B(new_n21565), .Y(new_n21610));
  or_5   g19262(.A(new_n21569), .B(new_n15927), .Y(new_n21611));
  nor_5  g19263(.A(new_n21584), .B(new_n21611), .Y(new_n21612));
  not_8  g19264(.A(new_n21612), .Y(new_n21613));
  nor_5  g19265(.A(new_n21613), .B(new_n21610), .Y(new_n21614));
  or_5   g19266(.A(new_n21614), .B(new_n21609), .Y(n9838));
  xnor_4 g19267(.A(new_n19357_1), .B(new_n19354_1), .Y(n9867));
  nor_5  g19268(.A(new_n18935), .B(new_n5686), .Y(new_n21617));
  and_5  g19269(.A(new_n18939), .B(new_n18936), .Y(new_n21618));
  nor_5  g19270(.A(new_n21618), .B(new_n21617), .Y(new_n21619));
  nor_5  g19271(.A(new_n21619), .B(new_n20166), .Y(new_n21620));
  xnor_4 g19272(.A(new_n21619), .B(new_n20147), .Y(new_n21621));
  nor_5  g19273(.A(new_n21621), .B(new_n8134), .Y(new_n21622));
  nor_5  g19274(.A(new_n18940_1), .B(new_n18928), .Y(new_n21623));
  nor_5  g19275(.A(new_n18944), .B(new_n18941), .Y(new_n21624));
  nor_5  g19276(.A(new_n21624), .B(new_n21623), .Y(new_n21625));
  xnor_4 g19277(.A(new_n21621), .B(new_n8134), .Y(new_n21626));
  nor_5  g19278(.A(new_n21626), .B(new_n21625), .Y(new_n21627));
  nor_5  g19279(.A(new_n21627), .B(new_n21622), .Y(new_n21628_1));
  nor_5  g19280(.A(new_n21628_1), .B(new_n21620), .Y(new_n21629));
  nor_5  g19281(.A(new_n21629), .B(new_n8028), .Y(n9890));
  xor_4  g19282(.A(new_n17801), .B(new_n17792), .Y(n9917));
  xnor_4 g19283(.A(new_n20427), .B(new_n20420), .Y(n9919));
  xnor_4 g19284(.A(new_n17970), .B(new_n17957), .Y(n9938));
  xnor_4 g19285(.A(new_n17613), .B(new_n17612), .Y(n9946));
  xnor_4 g19286(.A(n21784), .B(new_n4907), .Y(new_n21635));
  nor_5  g19287(.A(n5521), .B(n2858), .Y(new_n21636));
  xnor_4 g19288(.A(n5521), .B(n2858), .Y(new_n21637_1));
  nor_5  g19289(.A(n11926), .B(n2659), .Y(new_n21638));
  xnor_4 g19290(.A(n11926), .B(n2659), .Y(new_n21639));
  nor_5  g19291(.A(n24327), .B(n4325), .Y(new_n21640));
  xnor_4 g19292(.A(n24327), .B(new_n5991), .Y(new_n21641));
  nor_5  g19293(.A(new_n4922), .B(new_n14435), .Y(new_n21642));
  or_5   g19294(.A(n22198), .B(n5337), .Y(new_n21643));
  nor_5  g19295(.A(n20826), .B(n626), .Y(new_n21644));
  and_5  g19296(.A(new_n12793), .B(new_n12790), .Y(new_n21645_1));
  nor_5  g19297(.A(new_n21645_1), .B(new_n21644), .Y(new_n21646));
  and_5  g19298(.A(new_n21646), .B(new_n21643), .Y(new_n21647));
  nor_5  g19299(.A(new_n21647), .B(new_n21642), .Y(new_n21648));
  and_5  g19300(.A(new_n21648), .B(new_n21641), .Y(new_n21649_1));
  nor_5  g19301(.A(new_n21649_1), .B(new_n21640), .Y(new_n21650));
  nor_5  g19302(.A(new_n21650), .B(new_n21639), .Y(new_n21651));
  nor_5  g19303(.A(new_n21651), .B(new_n21638), .Y(new_n21652));
  nor_5  g19304(.A(new_n21652), .B(new_n21637_1), .Y(new_n21653));
  or_5   g19305(.A(new_n21653), .B(new_n21636), .Y(new_n21654_1));
  xor_4  g19306(.A(new_n21654_1), .B(new_n21635), .Y(new_n21655));
  xnor_4 g19307(.A(new_n21655), .B(new_n4837), .Y(new_n21656));
  xnor_4 g19308(.A(new_n21652), .B(new_n21637_1), .Y(new_n21657));
  nor_5  g19309(.A(new_n21657), .B(new_n4841), .Y(new_n21658));
  xnor_4 g19310(.A(new_n21657), .B(new_n4841), .Y(new_n21659));
  xnor_4 g19311(.A(new_n21650), .B(new_n21639), .Y(new_n21660));
  nor_5  g19312(.A(new_n21660), .B(new_n4845), .Y(new_n21661));
  xnor_4 g19313(.A(new_n21648), .B(new_n21641), .Y(new_n21662));
  nor_5  g19314(.A(new_n21662), .B(new_n4850_1), .Y(new_n21663));
  not_8  g19315(.A(new_n21662), .Y(new_n21664));
  xnor_4 g19316(.A(new_n21664), .B(new_n4850_1), .Y(new_n21665_1));
  xnor_4 g19317(.A(n22198), .B(n5337), .Y(new_n21666));
  xnor_4 g19318(.A(new_n21666), .B(new_n21646), .Y(new_n21667));
  nor_5  g19319(.A(new_n21667), .B(new_n4854), .Y(new_n21668));
  and_5  g19320(.A(new_n12795), .B(new_n12789), .Y(new_n21669));
  nor_5  g19321(.A(new_n12796), .B(new_n4861), .Y(new_n21670));
  nor_5  g19322(.A(new_n21670), .B(new_n21669), .Y(new_n21671));
  xor_4  g19323(.A(new_n21667), .B(new_n4854), .Y(new_n21672));
  and_5  g19324(.A(new_n21672), .B(new_n21671), .Y(new_n21673));
  or_5   g19325(.A(new_n21673), .B(new_n21668), .Y(new_n21674_1));
  and_5  g19326(.A(new_n21674_1), .B(new_n21665_1), .Y(new_n21675));
  nor_5  g19327(.A(new_n21675), .B(new_n21663), .Y(new_n21676));
  xnor_4 g19328(.A(new_n21660), .B(new_n4845), .Y(new_n21677));
  nor_5  g19329(.A(new_n21677), .B(new_n21676), .Y(new_n21678));
  nor_5  g19330(.A(new_n21678), .B(new_n21661), .Y(new_n21679));
  nor_5  g19331(.A(new_n21679), .B(new_n21659), .Y(new_n21680_1));
  nor_5  g19332(.A(new_n21680_1), .B(new_n21658), .Y(new_n21681));
  xnor_4 g19333(.A(new_n21681), .B(new_n21656), .Y(new_n21682));
  xnor_4 g19334(.A(new_n21682), .B(new_n17137), .Y(new_n21683));
  xnor_4 g19335(.A(new_n21679), .B(new_n21659), .Y(new_n21684));
  nor_5  g19336(.A(new_n21684), .B(new_n16464), .Y(new_n21685_1));
  xnor_4 g19337(.A(new_n21684), .B(new_n16464), .Y(new_n21686));
  xnor_4 g19338(.A(new_n21677), .B(new_n21676), .Y(new_n21687_1));
  nor_5  g19339(.A(new_n21687_1), .B(new_n16469), .Y(new_n21688));
  xnor_4 g19340(.A(new_n21687_1), .B(new_n16469), .Y(new_n21689));
  xor_4  g19341(.A(new_n21674_1), .B(new_n21665_1), .Y(new_n21690));
  and_5  g19342(.A(new_n21690), .B(new_n3771), .Y(new_n21691));
  xnor_4 g19343(.A(new_n21690), .B(new_n3772), .Y(new_n21692));
  xor_4  g19344(.A(new_n21672), .B(new_n21671), .Y(new_n21693));
  nor_5  g19345(.A(new_n21693), .B(new_n3775), .Y(new_n21694));
  and_5  g19346(.A(new_n12797), .B(new_n3782), .Y(new_n21695));
  and_5  g19347(.A(new_n12806), .B(new_n12798), .Y(new_n21696));
  nor_5  g19348(.A(new_n21696), .B(new_n21695), .Y(new_n21697));
  xnor_4 g19349(.A(new_n21693), .B(new_n3775), .Y(new_n21698));
  nor_5  g19350(.A(new_n21698), .B(new_n21697), .Y(new_n21699));
  nor_5  g19351(.A(new_n21699), .B(new_n21694), .Y(new_n21700));
  and_5  g19352(.A(new_n21700), .B(new_n21692), .Y(new_n21701));
  nor_5  g19353(.A(new_n21701), .B(new_n21691), .Y(new_n21702));
  nor_5  g19354(.A(new_n21702), .B(new_n21689), .Y(new_n21703));
  nor_5  g19355(.A(new_n21703), .B(new_n21688), .Y(new_n21704));
  nor_5  g19356(.A(new_n21704), .B(new_n21686), .Y(new_n21705));
  nor_5  g19357(.A(new_n21705), .B(new_n21685_1), .Y(new_n21706));
  xor_4  g19358(.A(new_n21706), .B(new_n21683), .Y(n9968));
  nor_5  g19359(.A(new_n20093), .B(new_n13678), .Y(new_n21708));
  xor_4  g19360(.A(new_n20093), .B(new_n13678), .Y(new_n21709));
  nor_5  g19361(.A(new_n20102), .B(new_n13678), .Y(new_n21710));
  xnor_4 g19362(.A(new_n20101), .B(new_n13678), .Y(new_n21711));
  and_5  g19363(.A(new_n20095), .B(new_n11169), .Y(new_n21712));
  and_5  g19364(.A(new_n11267), .B(new_n11227), .Y(new_n21713));
  nor_5  g19365(.A(new_n21713), .B(new_n21712), .Y(new_n21714));
  and_5  g19366(.A(new_n21714), .B(new_n21711), .Y(new_n21715));
  nor_5  g19367(.A(new_n21715), .B(new_n21710), .Y(new_n21716));
  and_5  g19368(.A(new_n21716), .B(new_n21709), .Y(new_n21717_1));
  nor_5  g19369(.A(new_n21717_1), .B(new_n21708), .Y(n10009));
  xnor_4 g19370(.A(new_n20813), .B(new_n20810), .Y(n10010));
  and_5  g19371(.A(new_n14513), .B(new_n10955), .Y(new_n21720));
  and_5  g19372(.A(new_n14544), .B(new_n14515), .Y(new_n21721));
  nor_5  g19373(.A(new_n21721), .B(new_n21720), .Y(new_n21722));
  not_8  g19374(.A(new_n21722), .Y(new_n21723));
  nor_5  g19375(.A(new_n21723), .B(new_n14586), .Y(new_n21724));
  xnor_4 g19376(.A(new_n21722), .B(new_n14586), .Y(new_n21725));
  and_5  g19377(.A(new_n14586), .B(new_n14545), .Y(new_n21726));
  and_5  g19378(.A(new_n14626), .B(new_n14587), .Y(new_n21727));
  or_5   g19379(.A(new_n21727), .B(new_n21726), .Y(new_n21728));
  and_5  g19380(.A(new_n21728), .B(new_n21725), .Y(new_n21729));
  nor_5  g19381(.A(new_n21729), .B(new_n21724), .Y(n10019));
  xnor_4 g19382(.A(new_n14411), .B(new_n14363), .Y(n10021));
  xor_4  g19383(.A(new_n9563), .B(new_n9553), .Y(n10055));
  xnor_4 g19384(.A(new_n10603), .B(new_n10581), .Y(n10101));
  xnor_4 g19385(.A(new_n4602), .B(new_n4556), .Y(n10111));
  nor_5  g19386(.A(n16544), .B(new_n20751), .Y(new_n21735_1));
  xnor_4 g19387(.A(n16544), .B(n3324), .Y(new_n21736));
  nor_5  g19388(.A(new_n19668), .B(n6814), .Y(new_n21737));
  xnor_4 g19389(.A(n17911), .B(n6814), .Y(new_n21738));
  nor_5  g19390(.A(new_n18472), .B(n19701), .Y(new_n21739));
  xnor_4 g19391(.A(n21997), .B(n19701), .Y(new_n21740));
  nor_5  g19392(.A(new_n8501), .B(n23529), .Y(new_n21741));
  xnor_4 g19393(.A(n25119), .B(n23529), .Y(new_n21742));
  nor_5  g19394(.A(n24620), .B(new_n8503), .Y(new_n21743));
  xnor_4 g19395(.A(n24620), .B(n1163), .Y(new_n21744));
  nor_5  g19396(.A(new_n8506), .B(n5211), .Y(new_n21745));
  or_5   g19397(.A(n18537), .B(new_n8968), .Y(new_n21746));
  nor_5  g19398(.A(new_n8971_1), .B(n7057), .Y(new_n21747));
  and_5  g19399(.A(new_n9451_1), .B(new_n9442), .Y(new_n21748));
  nor_5  g19400(.A(new_n21748), .B(new_n21747), .Y(new_n21749_1));
  and_5  g19401(.A(new_n21749_1), .B(new_n21746), .Y(new_n21750_1));
  or_5   g19402(.A(new_n21750_1), .B(new_n21745), .Y(new_n21751));
  and_5  g19403(.A(new_n21751), .B(new_n21744), .Y(new_n21752));
  or_5   g19404(.A(new_n21752), .B(new_n21743), .Y(new_n21753_1));
  and_5  g19405(.A(new_n21753_1), .B(new_n21742), .Y(new_n21754));
  or_5   g19406(.A(new_n21754), .B(new_n21741), .Y(new_n21755));
  and_5  g19407(.A(new_n21755), .B(new_n21740), .Y(new_n21756));
  or_5   g19408(.A(new_n21756), .B(new_n21739), .Y(new_n21757));
  and_5  g19409(.A(new_n21757), .B(new_n21738), .Y(new_n21758));
  or_5   g19410(.A(new_n21758), .B(new_n21737), .Y(new_n21759));
  and_5  g19411(.A(new_n21759), .B(new_n21736), .Y(new_n21760));
  nor_5  g19412(.A(new_n21760), .B(new_n21735_1), .Y(new_n21761));
  not_8  g19413(.A(new_n21761), .Y(new_n21762));
  xnor_4 g19414(.A(new_n21762), .B(new_n20950), .Y(new_n21763));
  nor_5  g19415(.A(new_n21762), .B(new_n20960), .Y(new_n21764));
  nor_5  g19416(.A(new_n21761), .B(new_n20959), .Y(new_n21765_1));
  xor_4  g19417(.A(new_n21759), .B(new_n21736), .Y(new_n21766));
  nor_5  g19418(.A(new_n21766), .B(new_n16979), .Y(new_n21767));
  xnor_4 g19419(.A(new_n21766), .B(new_n16979), .Y(new_n21768));
  xor_4  g19420(.A(new_n21757), .B(new_n21738), .Y(new_n21769));
  nor_5  g19421(.A(new_n21769), .B(new_n17027), .Y(new_n21770));
  xnor_4 g19422(.A(new_n21769), .B(new_n17027), .Y(new_n21771));
  xor_4  g19423(.A(new_n21755), .B(new_n21740), .Y(new_n21772));
  nor_5  g19424(.A(new_n21772), .B(new_n17034), .Y(new_n21773));
  xnor_4 g19425(.A(new_n21772), .B(new_n17034), .Y(new_n21774));
  xor_4  g19426(.A(new_n21753_1), .B(new_n21742), .Y(new_n21775));
  nor_5  g19427(.A(new_n21775), .B(new_n17041), .Y(new_n21776));
  xnor_4 g19428(.A(new_n21775), .B(new_n17041), .Y(new_n21777));
  xor_4  g19429(.A(new_n21751), .B(new_n21744), .Y(new_n21778));
  nor_5  g19430(.A(new_n21778), .B(new_n17046), .Y(new_n21779_1));
  xnor_4 g19431(.A(n18537), .B(n5211), .Y(new_n21780));
  xnor_4 g19432(.A(new_n21780), .B(new_n21749_1), .Y(new_n21781));
  nor_5  g19433(.A(new_n21781), .B(new_n17055), .Y(new_n21782));
  xnor_4 g19434(.A(new_n21781), .B(new_n17052), .Y(new_n21783));
  and_5  g19435(.A(new_n9452), .B(new_n9441), .Y(new_n21784_1));
  and_5  g19436(.A(new_n9473), .B(new_n9453), .Y(new_n21785));
  or_5   g19437(.A(new_n21785), .B(new_n21784_1), .Y(new_n21786));
  and_5  g19438(.A(new_n21786), .B(new_n21783), .Y(new_n21787));
  nor_5  g19439(.A(new_n21787), .B(new_n21782), .Y(new_n21788));
  xnor_4 g19440(.A(new_n21778), .B(new_n17045), .Y(new_n21789));
  and_5  g19441(.A(new_n21789), .B(new_n21788), .Y(new_n21790));
  nor_5  g19442(.A(new_n21790), .B(new_n21779_1), .Y(new_n21791));
  nor_5  g19443(.A(new_n21791), .B(new_n21777), .Y(new_n21792));
  nor_5  g19444(.A(new_n21792), .B(new_n21776), .Y(new_n21793));
  nor_5  g19445(.A(new_n21793), .B(new_n21774), .Y(new_n21794));
  nor_5  g19446(.A(new_n21794), .B(new_n21773), .Y(new_n21795));
  nor_5  g19447(.A(new_n21795), .B(new_n21771), .Y(new_n21796));
  nor_5  g19448(.A(new_n21796), .B(new_n21770), .Y(new_n21797));
  nor_5  g19449(.A(new_n21797), .B(new_n21768), .Y(new_n21798));
  nor_5  g19450(.A(new_n21798), .B(new_n21767), .Y(new_n21799));
  not_8  g19451(.A(new_n21799), .Y(new_n21800_1));
  nor_5  g19452(.A(new_n21800_1), .B(new_n21765_1), .Y(new_n21801));
  nor_5  g19453(.A(new_n21801), .B(new_n21764), .Y(new_n21802));
  xnor_4 g19454(.A(new_n21802), .B(new_n21763), .Y(n10165));
  xnor_4 g19455(.A(new_n12874), .B(new_n12873_1), .Y(n10236));
  xnor_4 g19456(.A(new_n14285), .B(new_n14263), .Y(n10239));
  xnor_4 g19457(.A(new_n6415), .B(new_n6375_1), .Y(n10244));
  xnor_4 g19458(.A(new_n17901), .B(new_n17889_1), .Y(n10261));
  xnor_4 g19459(.A(new_n15539_1), .B(new_n15525), .Y(n10262));
  xnor_4 g19460(.A(new_n16714), .B(new_n16713), .Y(n10287));
  nor_5  g19461(.A(new_n21185), .B(new_n15096), .Y(new_n21810));
  xnor_4 g19462(.A(new_n21227), .B(new_n21810), .Y(new_n21811));
  nor_5  g19463(.A(new_n21190), .B(new_n21186), .Y(new_n21812));
  nor_5  g19464(.A(new_n21204), .B(new_n21191), .Y(new_n21813));
  nor_5  g19465(.A(new_n21813), .B(new_n21812), .Y(new_n21814));
  xnor_4 g19466(.A(new_n21814), .B(new_n21811), .Y(n10295));
  xnor_4 g19467(.A(new_n14725), .B(new_n14722), .Y(n10321));
  xnor_4 g19468(.A(new_n14287), .B(new_n14260), .Y(n10326));
  xor_4  g19469(.A(new_n2833), .B(new_n2820), .Y(n10327));
  xnor_4 g19470(.A(new_n20102), .B(new_n20082), .Y(new_n21819));
  xnor_4 g19471(.A(new_n21819), .B(new_n20104), .Y(n10330));
  xnor_4 g19472(.A(new_n20736), .B(new_n20703), .Y(n10340));
  xnor_4 g19473(.A(new_n16711), .B(new_n16708), .Y(new_n21822));
  xnor_4 g19474(.A(new_n21822), .B(new_n16716), .Y(n10345));
  nor_5  g19475(.A(new_n13919), .B(new_n4897), .Y(new_n21824));
  nor_5  g19476(.A(new_n18896), .B(new_n21824), .Y(new_n21825));
  not_8  g19477(.A(new_n4902), .Y(new_n21826));
  nor_5  g19478(.A(new_n18899), .B(new_n21826), .Y(new_n21827));
  xnor_4 g19479(.A(new_n18899), .B(new_n21826), .Y(new_n21828));
  and_5  g19480(.A(new_n18904), .B(new_n4904), .Y(new_n21829));
  xnor_4 g19481(.A(new_n18904), .B(new_n4904), .Y(new_n21830));
  and_5  g19482(.A(new_n18908), .B(new_n4910), .Y(new_n21831));
  xnor_4 g19483(.A(new_n18908), .B(new_n4910), .Y(new_n21832_1));
  and_5  g19484(.A(new_n18912), .B(new_n4914), .Y(new_n21833));
  xnor_4 g19485(.A(new_n18912), .B(new_n4914), .Y(new_n21834));
  nor_5  g19486(.A(new_n9351), .B(new_n4920), .Y(new_n21835));
  xnor_4 g19487(.A(new_n9351), .B(new_n4920), .Y(new_n21836));
  nor_5  g19488(.A(new_n9355), .B(new_n4925_1), .Y(new_n21837));
  xnor_4 g19489(.A(new_n9355), .B(new_n4925_1), .Y(new_n21838));
  nor_5  g19490(.A(new_n9360), .B(new_n4930), .Y(new_n21839_1));
  xnor_4 g19491(.A(new_n9360), .B(new_n4930), .Y(new_n21840));
  nor_5  g19492(.A(new_n9365), .B(new_n4950), .Y(new_n21841));
  xnor_4 g19493(.A(new_n9365), .B(new_n4950), .Y(new_n21842));
  nor_5  g19494(.A(new_n9370), .B(new_n4936), .Y(new_n21843));
  xnor_4 g19495(.A(new_n9370), .B(new_n4936), .Y(new_n21844));
  nor_5  g19496(.A(new_n9376), .B(new_n4943), .Y(new_n21845));
  and_5  g19497(.A(new_n21845), .B(new_n9373), .Y(new_n21846));
  xnor_4 g19498(.A(new_n21845), .B(new_n9380_1), .Y(new_n21847));
  and_5  g19499(.A(new_n21847), .B(new_n4940), .Y(new_n21848));
  nor_5  g19500(.A(new_n21848), .B(new_n21846), .Y(new_n21849));
  nor_5  g19501(.A(new_n21849), .B(new_n21844), .Y(new_n21850));
  nor_5  g19502(.A(new_n21850), .B(new_n21843), .Y(new_n21851));
  nor_5  g19503(.A(new_n21851), .B(new_n21842), .Y(new_n21852));
  nor_5  g19504(.A(new_n21852), .B(new_n21841), .Y(new_n21853));
  nor_5  g19505(.A(new_n21853), .B(new_n21840), .Y(new_n21854));
  nor_5  g19506(.A(new_n21854), .B(new_n21839_1), .Y(new_n21855));
  nor_5  g19507(.A(new_n21855), .B(new_n21838), .Y(new_n21856));
  nor_5  g19508(.A(new_n21856), .B(new_n21837), .Y(new_n21857));
  nor_5  g19509(.A(new_n21857), .B(new_n21836), .Y(new_n21858));
  nor_5  g19510(.A(new_n21858), .B(new_n21835), .Y(new_n21859));
  nor_5  g19511(.A(new_n21859), .B(new_n21834), .Y(new_n21860));
  nor_5  g19512(.A(new_n21860), .B(new_n21833), .Y(new_n21861));
  nor_5  g19513(.A(new_n21861), .B(new_n21832_1), .Y(new_n21862));
  nor_5  g19514(.A(new_n21862), .B(new_n21831), .Y(new_n21863));
  nor_5  g19515(.A(new_n21863), .B(new_n21830), .Y(new_n21864));
  nor_5  g19516(.A(new_n21864), .B(new_n21829), .Y(new_n21865));
  nor_5  g19517(.A(new_n21865), .B(new_n21828), .Y(new_n21866));
  nor_5  g19518(.A(new_n21866), .B(new_n21827), .Y(new_n21867));
  xnor_4 g19519(.A(new_n18895), .B(new_n21824), .Y(new_n21868));
  and_5  g19520(.A(new_n21868), .B(new_n21867), .Y(new_n21869));
  nor_5  g19521(.A(new_n21869), .B(new_n21825), .Y(n10356));
  xor_4  g19522(.A(new_n19447), .B(new_n19446), .Y(n10385));
  nor_5  g19523(.A(new_n19664_1), .B(new_n18895), .Y(new_n21872));
  or_5   g19524(.A(new_n19663), .B(new_n18896), .Y(new_n21873));
  and_5  g19525(.A(new_n21873), .B(new_n19609), .Y(new_n21874_1));
  nor_5  g19526(.A(new_n21874_1), .B(new_n21872), .Y(new_n21875));
  nor_5  g19527(.A(new_n21875), .B(new_n19607), .Y(n10387));
  xnor_4 g19528(.A(new_n19867), .B(new_n19854), .Y(n10388));
  xnor_4 g19529(.A(new_n15325), .B(new_n15280), .Y(n10390));
  xnor_4 g19530(.A(new_n9461), .B(new_n9460_1), .Y(n10404));
  xnor_4 g19531(.A(new_n15703), .B(new_n15700), .Y(n10409));
  xnor_4 g19532(.A(new_n15907), .B(new_n8557), .Y(n10420));
  xnor_4 g19533(.A(new_n17894), .B(new_n6946), .Y(n10432));
  xnor_4 g19534(.A(new_n20903), .B(new_n20225), .Y(new_n21883));
  nor_5  g19535(.A(new_n20229), .B(new_n9600), .Y(new_n21884));
  nor_5  g19536(.A(new_n20489_1), .B(new_n20482), .Y(new_n21885));
  nor_5  g19537(.A(new_n21885), .B(new_n21884), .Y(new_n21886));
  xnor_4 g19538(.A(new_n21886), .B(new_n21883), .Y(new_n21887));
  xnor_4 g19539(.A(new_n21887), .B(new_n11380), .Y(new_n21888));
  nor_5  g19540(.A(new_n20490_1), .B(new_n11384), .Y(new_n21889));
  nor_5  g19541(.A(new_n20499), .B(new_n20491), .Y(new_n21890));
  nor_5  g19542(.A(new_n21890), .B(new_n21889), .Y(new_n21891));
  xor_4  g19543(.A(new_n21891), .B(new_n21888), .Y(n10484));
  xnor_4 g19544(.A(new_n11256), .B(new_n11243), .Y(n10489));
  xnor_4 g19545(.A(new_n13288), .B(new_n3641), .Y(n10525));
  xor_4  g19546(.A(new_n17271), .B(new_n11992), .Y(new_n21895));
  xnor_4 g19547(.A(new_n21895), .B(new_n17279), .Y(n10540));
  xnor_4 g19548(.A(new_n15816_1), .B(new_n15792), .Y(n10561));
  xnor_4 g19549(.A(new_n15329), .B(new_n15272), .Y(n10564));
  xnor_4 g19550(.A(new_n9963), .B(new_n9961), .Y(n10588));
  xnor_4 g19551(.A(new_n9966), .B(new_n9964), .Y(n10595));
  xor_4  g19552(.A(new_n20609_1), .B(new_n20597), .Y(n10617));
  xnor_4 g19553(.A(new_n12310), .B(new_n12254), .Y(n10628));
  xnor_4 g19554(.A(new_n10549), .B(new_n5726), .Y(new_n21903));
  nor_5  g19555(.A(new_n10558), .B(new_n5729), .Y(new_n21904));
  xnor_4 g19556(.A(new_n10557), .B(new_n5730), .Y(new_n21905_1));
  and_5  g19557(.A(new_n10561_1), .B(new_n5734), .Y(new_n21906));
  xnor_4 g19558(.A(new_n10561_1), .B(new_n5734), .Y(new_n21907));
  nor_5  g19559(.A(new_n5769), .B(new_n5739), .Y(new_n21908));
  nor_5  g19560(.A(new_n21908), .B(new_n5779), .Y(new_n21909));
  xnor_4 g19561(.A(new_n21908), .B(new_n5779), .Y(new_n21910));
  nor_5  g19562(.A(new_n21910), .B(new_n5746), .Y(new_n21911));
  nor_5  g19563(.A(new_n21911), .B(new_n21909), .Y(new_n21912));
  nor_5  g19564(.A(new_n21912), .B(new_n21907), .Y(new_n21913));
  nor_5  g19565(.A(new_n21913), .B(new_n21906), .Y(new_n21914));
  nor_5  g19566(.A(new_n21914), .B(new_n21905_1), .Y(new_n21915_1));
  nor_5  g19567(.A(new_n21915_1), .B(new_n21904), .Y(new_n21916));
  xnor_4 g19568(.A(new_n21916), .B(new_n21903), .Y(n10647));
  nor_5  g19569(.A(new_n19318), .B(new_n8333), .Y(new_n21918));
  not_8  g19570(.A(new_n21918), .Y(new_n21919));
  nor_5  g19571(.A(new_n19344), .B(new_n3582_1), .Y(new_n21920));
  and_5  g19572(.A(new_n3661), .B(new_n3599), .Y(new_n21921));
  or_5   g19573(.A(new_n21921), .B(new_n19343), .Y(new_n21922));
  or_5   g19574(.A(new_n21922), .B(new_n21920), .Y(new_n21923));
  nor_5  g19575(.A(new_n21923), .B(new_n13257), .Y(new_n21924));
  xnor_4 g19576(.A(new_n21924), .B(new_n21919), .Y(new_n21925));
  not_8  g19577(.A(new_n8340), .Y(new_n21926));
  xor_4  g19578(.A(new_n21923), .B(new_n13257), .Y(new_n21927));
  nor_5  g19579(.A(new_n21927), .B(new_n21926), .Y(new_n21928));
  nor_5  g19580(.A(new_n3662), .B(new_n3535), .Y(new_n21929));
  nor_5  g19581(.A(new_n3723), .B(new_n3663), .Y(new_n21930));
  nor_5  g19582(.A(new_n21930), .B(new_n21929), .Y(new_n21931));
  xnor_4 g19583(.A(new_n21927), .B(new_n8340), .Y(new_n21932));
  and_5  g19584(.A(new_n21932), .B(new_n21931), .Y(new_n21933));
  nor_5  g19585(.A(new_n21933), .B(new_n21928), .Y(new_n21934_1));
  xnor_4 g19586(.A(new_n21934_1), .B(new_n21925), .Y(n10653));
  xnor_4 g19587(.A(new_n9033), .B(new_n9032_1), .Y(n10692));
  xnor_4 g19588(.A(new_n14463), .B(new_n4302), .Y(n10694));
  xnor_4 g19589(.A(new_n19731), .B(new_n19708), .Y(n10701));
  xnor_4 g19590(.A(new_n6137), .B(new_n6118), .Y(n10756));
  not_8  g19591(.A(n6659), .Y(new_n21940));
  nor_5  g19592(.A(new_n21940), .B(n5101), .Y(new_n21941));
  and_5  g19593(.A(new_n15670), .B(new_n15666), .Y(new_n21942));
  nor_5  g19594(.A(new_n21942), .B(new_n21941), .Y(new_n21943_1));
  not_8  g19595(.A(new_n21943_1), .Y(new_n21944));
  not_8  g19596(.A(n13419), .Y(new_n21945));
  and_5  g19597(.A(new_n15671), .B(new_n21945), .Y(new_n21946));
  nor_5  g19598(.A(new_n15671), .B(new_n21945), .Y(new_n21947));
  not_8  g19599(.A(n4967), .Y(new_n21948));
  and_5  g19600(.A(new_n15626), .B(new_n21948), .Y(new_n21949));
  nor_5  g19601(.A(new_n15626), .B(new_n21948), .Y(new_n21950));
  nor_5  g19602(.A(new_n18822), .B(new_n21950), .Y(new_n21951));
  nor_5  g19603(.A(new_n21951), .B(new_n21949), .Y(new_n21952));
  nor_5  g19604(.A(new_n21952), .B(new_n21947), .Y(new_n21953));
  nor_5  g19605(.A(new_n21953), .B(new_n21946), .Y(new_n21954));
  and_5  g19606(.A(new_n21954), .B(new_n21944), .Y(new_n21955));
  xnor_4 g19607(.A(new_n21955), .B(new_n3197), .Y(new_n21956));
  xnor_4 g19608(.A(new_n21954), .B(new_n21943_1), .Y(new_n21957_1));
  and_5  g19609(.A(new_n21957_1), .B(new_n3329), .Y(new_n21958));
  xnor_4 g19610(.A(new_n21957_1), .B(new_n3329), .Y(new_n21959));
  xnor_4 g19611(.A(new_n21952), .B(new_n15672), .Y(new_n21960_1));
  nor_5  g19612(.A(new_n21960_1), .B(new_n3215), .Y(new_n21961));
  xnor_4 g19613(.A(new_n21960_1), .B(new_n3215), .Y(new_n21962));
  nor_5  g19614(.A(new_n18823), .B(new_n3224), .Y(new_n21963));
  nor_5  g19615(.A(new_n18860), .B(new_n18824), .Y(new_n21964));
  or_5   g19616(.A(new_n21964), .B(new_n21963), .Y(new_n21965));
  nor_5  g19617(.A(new_n21965), .B(new_n21962), .Y(new_n21966));
  nor_5  g19618(.A(new_n21966), .B(new_n21961), .Y(new_n21967));
  nor_5  g19619(.A(new_n21967), .B(new_n21959), .Y(new_n21968));
  nor_5  g19620(.A(new_n21968), .B(new_n21958), .Y(new_n21969));
  xnor_4 g19621(.A(new_n21969), .B(new_n21956), .Y(n10775));
  xnor_4 g19622(.A(new_n20522), .B(new_n20517), .Y(n10780));
  xnor_4 g19623(.A(n17095), .B(new_n16134), .Y(new_n21972));
  nor_5  g19624(.A(n22591), .B(n22274), .Y(new_n21973));
  or_5   g19625(.A(new_n9532), .B(new_n4122), .Y(new_n21974));
  xnor_4 g19626(.A(n22591), .B(new_n4118), .Y(new_n21975));
  and_5  g19627(.A(new_n21975), .B(new_n21974), .Y(new_n21976_1));
  or_5   g19628(.A(new_n21976_1), .B(new_n21973), .Y(new_n21977));
  xor_4  g19629(.A(new_n21977), .B(new_n21972), .Y(new_n21978));
  xnor_4 g19630(.A(new_n21978), .B(n21749), .Y(new_n21979));
  nor_5  g19631(.A(new_n8912), .B(new_n9485), .Y(new_n21980));
  nor_5  g19632(.A(new_n21980), .B(n7769), .Y(new_n21981_1));
  xor_4  g19633(.A(new_n21975), .B(new_n21974), .Y(new_n21982));
  xnor_4 g19634(.A(new_n21980), .B(new_n9487), .Y(new_n21983));
  not_8  g19635(.A(new_n21983), .Y(new_n21984));
  nor_5  g19636(.A(new_n21984), .B(new_n21982), .Y(new_n21985));
  nor_5  g19637(.A(new_n21985), .B(new_n21981_1), .Y(new_n21986_1));
  xnor_4 g19638(.A(new_n21986_1), .B(new_n21979), .Y(new_n21987));
  xnor_4 g19639(.A(new_n21987), .B(new_n18061_1), .Y(new_n21988));
  xnor_4 g19640(.A(new_n21983), .B(new_n21982), .Y(new_n21989));
  and_5  g19641(.A(new_n21989), .B(new_n18065), .Y(new_n21990));
  nor_5  g19642(.A(new_n8913), .B(new_n18068), .Y(new_n21991));
  xnor_4 g19643(.A(new_n21989), .B(new_n18064), .Y(new_n21992));
  and_5  g19644(.A(new_n21992), .B(new_n21991), .Y(new_n21993_1));
  or_5   g19645(.A(new_n21993_1), .B(new_n21990), .Y(new_n21994));
  xor_4  g19646(.A(new_n21994), .B(new_n21988), .Y(n10817));
  not_8  g19647(.A(new_n21210), .Y(new_n21996));
  and_5  g19648(.A(new_n21214), .B(new_n21996), .Y(new_n21997_1));
  and_5  g19649(.A(new_n21209), .B(new_n21206), .Y(new_n21998));
  nor_5  g19650(.A(new_n21214), .B(new_n21996), .Y(new_n21999));
  nor_5  g19651(.A(new_n21218), .B(new_n21999), .Y(new_n22000));
  or_5   g19652(.A(new_n22000), .B(new_n21998), .Y(new_n22001));
  nor_5  g19653(.A(new_n22001), .B(new_n21997_1), .Y(new_n22002));
  nor_5  g19654(.A(new_n22002), .B(new_n7694), .Y(new_n22003));
  nor_5  g19655(.A(new_n21219), .B(new_n7694), .Y(new_n22004));
  nor_5  g19656(.A(new_n21224), .B(new_n21221), .Y(new_n22005));
  nor_5  g19657(.A(new_n22005), .B(new_n22004), .Y(new_n22006));
  not_8  g19658(.A(new_n22002), .Y(new_n22007));
  xnor_4 g19659(.A(new_n22007), .B(new_n7694), .Y(new_n22008));
  and_5  g19660(.A(new_n22008), .B(new_n22006), .Y(new_n22009));
  nor_5  g19661(.A(new_n22009), .B(new_n22003), .Y(n10834));
  xor_4  g19662(.A(new_n21452), .B(new_n21435), .Y(n10851));
  xnor_4 g19663(.A(new_n21003), .B(new_n20994), .Y(n10874));
  xor_4  g19664(.A(new_n21628_1), .B(new_n21620), .Y(new_n22013));
  xnor_4 g19665(.A(new_n22013), .B(new_n8028), .Y(n10924));
  nor_5  g19666(.A(new_n11025_1), .B(new_n11021), .Y(new_n22015));
  and_5  g19667(.A(new_n11090), .B(new_n11027), .Y(new_n22016_1));
  nor_5  g19668(.A(new_n22016_1), .B(new_n22015), .Y(n10943));
  xnor_4 g19669(.A(new_n11785), .B(new_n11752), .Y(n10961));
  xnor_4 g19670(.A(new_n10499), .B(new_n10487), .Y(n11005));
  xnor_4 g19671(.A(new_n20782), .B(new_n20774_1), .Y(n11023));
  nor_5  g19672(.A(new_n17749_1), .B(new_n7263), .Y(new_n22021));
  xnor_4 g19673(.A(new_n17749_1), .B(new_n7263), .Y(new_n22022));
  nor_5  g19674(.A(new_n17751), .B(new_n7269), .Y(new_n22023));
  xnor_4 g19675(.A(new_n17751), .B(new_n7269), .Y(new_n22024));
  nor_5  g19676(.A(new_n16518), .B(new_n14657), .Y(new_n22025));
  xnor_4 g19677(.A(new_n16518), .B(new_n14657), .Y(new_n22026));
  and_5  g19678(.A(new_n11951), .B(new_n7278), .Y(new_n22027_1));
  nor_5  g19679(.A(new_n11976), .B(new_n11952), .Y(new_n22028));
  nor_5  g19680(.A(new_n22028), .B(new_n22027_1), .Y(new_n22029));
  nor_5  g19681(.A(new_n22029), .B(new_n22026), .Y(new_n22030));
  or_5   g19682(.A(new_n22030), .B(new_n22025), .Y(new_n22031));
  nor_5  g19683(.A(new_n22031), .B(new_n22024), .Y(new_n22032));
  nor_5  g19684(.A(new_n22032), .B(new_n22023), .Y(new_n22033));
  nor_5  g19685(.A(new_n22033), .B(new_n22022), .Y(new_n22034));
  nor_5  g19686(.A(new_n22034), .B(new_n22021), .Y(new_n22035));
  or_5   g19687(.A(new_n22035), .B(new_n7241), .Y(new_n22036));
  nor_5  g19688(.A(new_n22036), .B(new_n17776), .Y(new_n22037));
  not_8  g19689(.A(new_n21585), .Y(new_n22038));
  xnor_4 g19690(.A(new_n22035), .B(new_n7241), .Y(new_n22039));
  xnor_4 g19691(.A(new_n22039), .B(new_n17776), .Y(new_n22040));
  and_5  g19692(.A(new_n22040), .B(new_n22038), .Y(new_n22041));
  xnor_4 g19693(.A(new_n22040), .B(new_n22038), .Y(new_n22042));
  xnor_4 g19694(.A(new_n22033), .B(new_n22022), .Y(new_n22043_1));
  nor_5  g19695(.A(new_n22043_1), .B(new_n21591), .Y(new_n22044));
  xnor_4 g19696(.A(new_n22043_1), .B(new_n21591), .Y(new_n22045));
  xnor_4 g19697(.A(new_n22031), .B(new_n22024), .Y(new_n22046));
  nor_5  g19698(.A(new_n22046), .B(new_n21596), .Y(new_n22047));
  xnor_4 g19699(.A(new_n22046), .B(new_n21596), .Y(new_n22048));
  xor_4  g19700(.A(new_n22029), .B(new_n22026), .Y(new_n22049));
  nor_5  g19701(.A(new_n22049), .B(new_n17257), .Y(new_n22050_1));
  xnor_4 g19702(.A(new_n22049), .B(new_n17257), .Y(new_n22051));
  nor_5  g19703(.A(new_n11977), .B(new_n11946), .Y(new_n22052));
  nor_5  g19704(.A(new_n12014), .B(new_n11978), .Y(new_n22053));
  nor_5  g19705(.A(new_n22053), .B(new_n22052), .Y(new_n22054));
  nor_5  g19706(.A(new_n22054), .B(new_n22051), .Y(new_n22055));
  nor_5  g19707(.A(new_n22055), .B(new_n22050_1), .Y(new_n22056));
  nor_5  g19708(.A(new_n22056), .B(new_n22048), .Y(new_n22057));
  nor_5  g19709(.A(new_n22057), .B(new_n22047), .Y(new_n22058));
  nor_5  g19710(.A(new_n22058), .B(new_n22045), .Y(new_n22059));
  nor_5  g19711(.A(new_n22059), .B(new_n22044), .Y(new_n22060));
  nor_5  g19712(.A(new_n22060), .B(new_n22042), .Y(new_n22061));
  or_5   g19713(.A(new_n22061), .B(new_n22041), .Y(new_n22062));
  and_5  g19714(.A(new_n22062), .B(new_n22037), .Y(new_n22063_1));
  xor_4  g19715(.A(new_n22062), .B(new_n22037), .Y(new_n22064));
  nor_5  g19716(.A(new_n22064), .B(new_n21613), .Y(new_n22065));
  or_5   g19717(.A(new_n22065), .B(new_n22063_1), .Y(n11025));
  xnor_4 g19718(.A(new_n16154), .B(n21915), .Y(new_n22067));
  nor_5  g19719(.A(new_n16157), .B(new_n6836), .Y(new_n22068_1));
  xnor_4 g19720(.A(new_n16157), .B(n13775), .Y(new_n22069));
  nor_5  g19721(.A(new_n16160), .B(new_n6839), .Y(new_n22070));
  xnor_4 g19722(.A(new_n16160), .B(n1293), .Y(new_n22071));
  nor_5  g19723(.A(new_n16163), .B(new_n6842), .Y(new_n22072_1));
  and_5  g19724(.A(new_n18704), .B(new_n18701), .Y(new_n22073));
  or_5   g19725(.A(new_n22073), .B(new_n22072_1), .Y(new_n22074));
  and_5  g19726(.A(new_n22074), .B(new_n22071), .Y(new_n22075));
  or_5   g19727(.A(new_n22075), .B(new_n22070), .Y(new_n22076_1));
  and_5  g19728(.A(new_n22076_1), .B(new_n22069), .Y(new_n22077));
  or_5   g19729(.A(new_n22077), .B(new_n22068_1), .Y(new_n22078));
  xor_4  g19730(.A(new_n22078), .B(new_n22067), .Y(new_n22079));
  not_8  g19731(.A(new_n18707), .Y(new_n22080));
  nor_5  g19732(.A(new_n22080), .B(n26752), .Y(new_n22081));
  not_8  g19733(.A(new_n22081), .Y(new_n22082));
  nor_5  g19734(.A(new_n22082), .B(n4590), .Y(new_n22083));
  not_8  g19735(.A(new_n22083), .Y(new_n22084));
  nor_5  g19736(.A(new_n22084), .B(n25464), .Y(new_n22085));
  xnor_4 g19737(.A(new_n22085), .B(n3795), .Y(new_n22086));
  xnor_4 g19738(.A(new_n22086), .B(new_n8788), .Y(new_n22087));
  xnor_4 g19739(.A(new_n22083), .B(n25464), .Y(new_n22088));
  nor_5  g19740(.A(new_n22088), .B(new_n8795), .Y(new_n22089));
  xnor_4 g19741(.A(new_n22088), .B(new_n8795), .Y(new_n22090_1));
  xnor_4 g19742(.A(new_n22081), .B(n4590), .Y(new_n22091));
  nor_5  g19743(.A(new_n22091), .B(new_n8801), .Y(new_n22092));
  xnor_4 g19744(.A(new_n22091), .B(new_n8801), .Y(new_n22093));
  nor_5  g19745(.A(new_n18708_1), .B(new_n8807), .Y(new_n22094));
  nor_5  g19746(.A(new_n18712), .B(new_n18709), .Y(new_n22095));
  nor_5  g19747(.A(new_n22095), .B(new_n22094), .Y(new_n22096));
  nor_5  g19748(.A(new_n22096), .B(new_n22093), .Y(new_n22097));
  nor_5  g19749(.A(new_n22097), .B(new_n22092), .Y(new_n22098));
  nor_5  g19750(.A(new_n22098), .B(new_n22090_1), .Y(new_n22099));
  nor_5  g19751(.A(new_n22099), .B(new_n22089), .Y(new_n22100));
  xnor_4 g19752(.A(new_n22100), .B(new_n22087), .Y(new_n22101));
  xnor_4 g19753(.A(new_n22101), .B(new_n22079), .Y(new_n22102));
  xor_4  g19754(.A(new_n22076_1), .B(new_n22069), .Y(new_n22103));
  xnor_4 g19755(.A(new_n22098), .B(new_n22090_1), .Y(new_n22104));
  nor_5  g19756(.A(new_n22104), .B(new_n22103), .Y(new_n22105));
  xnor_4 g19757(.A(new_n22104), .B(new_n22103), .Y(new_n22106));
  xor_4  g19758(.A(new_n22074), .B(new_n22071), .Y(new_n22107_1));
  xnor_4 g19759(.A(new_n22096), .B(new_n22093), .Y(new_n22108));
  nor_5  g19760(.A(new_n22108), .B(new_n22107_1), .Y(new_n22109));
  xnor_4 g19761(.A(new_n22108), .B(new_n22107_1), .Y(new_n22110));
  nor_5  g19762(.A(new_n18713), .B(new_n18705), .Y(new_n22111));
  nor_5  g19763(.A(new_n18717), .B(new_n18714), .Y(new_n22112));
  nor_5  g19764(.A(new_n22112), .B(new_n22111), .Y(new_n22113_1));
  nor_5  g19765(.A(new_n22113_1), .B(new_n22110), .Y(new_n22114));
  nor_5  g19766(.A(new_n22114), .B(new_n22109), .Y(new_n22115));
  nor_5  g19767(.A(new_n22115), .B(new_n22106), .Y(new_n22116));
  nor_5  g19768(.A(new_n22116), .B(new_n22105), .Y(new_n22117));
  xnor_4 g19769(.A(new_n22117), .B(new_n22102), .Y(n11063));
  xnor_4 g19770(.A(new_n19865), .B(new_n19857), .Y(n11078));
  xnor_4 g19771(.A(new_n20524), .B(new_n20514), .Y(n11080));
  xnor_4 g19772(.A(new_n13584), .B(new_n13571), .Y(n11094));
  xnor_4 g19773(.A(new_n21789), .B(new_n21788), .Y(n11101));
  xnor_4 g19774(.A(new_n20602_1), .B(new_n14139), .Y(new_n22123));
  xnor_4 g19775(.A(new_n22123), .B(new_n20605), .Y(n11103));
  xnor_4 g19776(.A(new_n6581), .B(new_n6556_1), .Y(n11120));
  xor_4  g19777(.A(new_n5010), .B(new_n5007), .Y(n11127));
  xnor_4 g19778(.A(new_n14728), .B(new_n14727), .Y(n11132));
  xnor_4 g19779(.A(new_n11083), .B(new_n11038), .Y(n11134));
  xnor_4 g19780(.A(new_n3707), .B(new_n3706), .Y(n11138));
  xnor_4 g19781(.A(new_n10391), .B(new_n10381), .Y(n11182));
  xnor_4 g19782(.A(new_n13594), .B(new_n13556), .Y(n11234));
  xnor_4 g19783(.A(new_n21186), .B(new_n18226), .Y(new_n22132));
  nor_5  g19784(.A(new_n21193_1), .B(new_n18230), .Y(new_n22133));
  nor_5  g19785(.A(new_n20869_1), .B(new_n20848), .Y(new_n22134));
  nor_5  g19786(.A(new_n22134), .B(new_n22133), .Y(new_n22135));
  xnor_4 g19787(.A(new_n22135), .B(new_n22132), .Y(n11245));
  xnor_4 g19788(.A(new_n8641), .B(new_n8627), .Y(n11261));
  xnor_4 g19789(.A(new_n22115), .B(new_n22106), .Y(n11275));
  nand_5 g19790(.A(new_n13310), .B(new_n13251), .Y(n11290));
  xnor_4 g19791(.A(new_n9381), .B(new_n9379), .Y(n11313));
  xnor_4 g19792(.A(new_n16494), .B(new_n15936_1), .Y(new_n22141));
  xnor_4 g19793(.A(new_n22141), .B(new_n16508), .Y(n11325));
  xnor_4 g19794(.A(new_n13636), .B(new_n13635), .Y(n11326));
  xnor_4 g19795(.A(new_n16724), .B(new_n16692), .Y(n11330));
  xnor_4 g19796(.A(new_n11077), .B(new_n11049), .Y(n11347));
  xnor_4 g19797(.A(new_n21849), .B(new_n21844), .Y(n11348));
  xnor_4 g19798(.A(new_n14838), .B(new_n14830), .Y(n11352));
  nor_5  g19799(.A(new_n8271), .B(n3324), .Y(new_n22148));
  xnor_4 g19800(.A(n22442), .B(n3324), .Y(new_n22149));
  nor_5  g19801(.A(n17911), .B(new_n8273), .Y(new_n22150_1));
  nor_5  g19802(.A(n21997), .B(new_n8280), .Y(new_n22151));
  and_5  g19803(.A(new_n16915), .B(new_n16908), .Y(new_n22152));
  or_5   g19804(.A(new_n22152), .B(new_n22151), .Y(new_n22153));
  xnor_4 g19805(.A(n17911), .B(n468), .Y(new_n22154));
  and_5  g19806(.A(new_n22154), .B(new_n22153), .Y(new_n22155));
  or_5   g19807(.A(new_n22155), .B(new_n22150_1), .Y(new_n22156));
  and_5  g19808(.A(new_n22156), .B(new_n22149), .Y(new_n22157_1));
  nor_5  g19809(.A(new_n22157_1), .B(new_n22148), .Y(new_n22158));
  not_8  g19810(.A(new_n22158), .Y(new_n22159));
  and_5  g19811(.A(new_n17425), .B(new_n17419), .Y(new_n22160));
  nor_5  g19812(.A(new_n22160), .B(new_n7649), .Y(new_n22161));
  nor_5  g19813(.A(new_n17425), .B(new_n17419), .Y(new_n22162));
  nor_5  g19814(.A(new_n22162), .B(new_n7650), .Y(new_n22163));
  nor_5  g19815(.A(new_n22163), .B(new_n22161), .Y(new_n22164));
  xnor_4 g19816(.A(new_n22164), .B(new_n22159), .Y(new_n22165));
  nor_5  g19817(.A(new_n22159), .B(new_n17427), .Y(new_n22166));
  nor_5  g19818(.A(new_n22158), .B(new_n17428), .Y(new_n22167));
  xor_4  g19819(.A(new_n22156), .B(new_n22149), .Y(new_n22168));
  nor_5  g19820(.A(new_n22168), .B(new_n17430), .Y(new_n22169));
  xnor_4 g19821(.A(new_n22168), .B(new_n17430), .Y(new_n22170));
  not_8  g19822(.A(new_n22170), .Y(new_n22171));
  xor_4  g19823(.A(new_n22154), .B(new_n22153), .Y(new_n22172));
  and_5  g19824(.A(new_n22172), .B(new_n17433), .Y(new_n22173_1));
  xnor_4 g19825(.A(new_n22172), .B(new_n17432_1), .Y(new_n22174));
  and_5  g19826(.A(new_n16916), .B(new_n17436_1), .Y(new_n22175));
  and_5  g19827(.A(new_n16927), .B(new_n16917), .Y(new_n22176));
  or_5   g19828(.A(new_n22176), .B(new_n22175), .Y(new_n22177));
  and_5  g19829(.A(new_n22177), .B(new_n22174), .Y(new_n22178));
  nor_5  g19830(.A(new_n22178), .B(new_n22173_1), .Y(new_n22179));
  and_5  g19831(.A(new_n22179), .B(new_n22171), .Y(new_n22180));
  nor_5  g19832(.A(new_n22180), .B(new_n22169), .Y(new_n22181));
  not_8  g19833(.A(new_n22181), .Y(new_n22182));
  nor_5  g19834(.A(new_n22182), .B(new_n22167), .Y(new_n22183));
  nor_5  g19835(.A(new_n22183), .B(new_n22166), .Y(new_n22184));
  xnor_4 g19836(.A(new_n22184), .B(new_n22165), .Y(n11375));
  xnor_4 g19837(.A(new_n12337), .B(new_n7158), .Y(n11379));
  nor_5  g19838(.A(new_n11795), .B(n2570), .Y(new_n22187));
  and_5  g19839(.A(new_n16151), .B(new_n16122), .Y(new_n22188));
  nor_5  g19840(.A(new_n22188), .B(new_n22187), .Y(new_n22189));
  xnor_4 g19841(.A(new_n22189), .B(new_n11846), .Y(new_n22190));
  nor_5  g19842(.A(new_n16152), .B(new_n11802), .Y(new_n22191));
  nor_5  g19843(.A(new_n16188), .B(new_n16153), .Y(new_n22192));
  or_5   g19844(.A(new_n22192), .B(new_n22191), .Y(new_n22193));
  xor_4  g19845(.A(new_n22193), .B(new_n22190), .Y(new_n22194));
  xnor_4 g19846(.A(new_n22194), .B(new_n6356_1), .Y(new_n22195));
  nor_5  g19847(.A(new_n16189), .B(new_n6361), .Y(new_n22196));
  nor_5  g19848(.A(new_n16225), .B(new_n16190), .Y(new_n22197));
  nor_5  g19849(.A(new_n22197), .B(new_n22196), .Y(new_n22198_1));
  xnor_4 g19850(.A(new_n22198_1), .B(new_n22195), .Y(n11386));
  xnor_4 g19851(.A(new_n18850), .B(new_n18839), .Y(n11391));
  xnor_4 g19852(.A(new_n20833), .B(new_n20832), .Y(n11398));
  xnor_4 g19853(.A(new_n12644), .B(new_n12643), .Y(n11403));
  xnor_4 g19854(.A(new_n12087), .B(new_n12082), .Y(n11419));
  xnor_4 g19855(.A(new_n18690_1), .B(new_n18675), .Y(n11439));
  xnor_4 g19856(.A(new_n11325_1), .B(n2570), .Y(new_n22205));
  nor_5  g19857(.A(n19033), .B(n17037), .Y(new_n22206));
  xnor_4 g19858(.A(n19033), .B(n17037), .Y(new_n22207));
  nor_5  g19859(.A(n5386), .B(n655), .Y(new_n22208));
  xnor_4 g19860(.A(n5386), .B(n655), .Y(new_n22209));
  nor_5  g19861(.A(n26191), .B(n18145), .Y(new_n22210));
  xnor_4 g19862(.A(n26191), .B(n18145), .Y(new_n22211));
  nor_5  g19863(.A(n26512), .B(n10712), .Y(new_n22212));
  xnor_4 g19864(.A(n26512), .B(n10712), .Y(new_n22213_1));
  nor_5  g19865(.A(n25126), .B(n19575), .Y(new_n22214));
  xnor_4 g19866(.A(n25126), .B(new_n15732), .Y(new_n22215));
  and_5  g19867(.A(n19608), .B(n15378), .Y(new_n22216));
  or_5   g19868(.A(n19608), .B(n15378), .Y(new_n22217));
  nor_5  g19869(.A(n17095), .B(n1689), .Y(new_n22218));
  and_5  g19870(.A(new_n21977), .B(new_n21972), .Y(new_n22219));
  nor_5  g19871(.A(new_n22219), .B(new_n22218), .Y(new_n22220));
  and_5  g19872(.A(new_n22220), .B(new_n22217), .Y(new_n22221));
  nor_5  g19873(.A(new_n22221), .B(new_n22216), .Y(new_n22222));
  and_5  g19874(.A(new_n22222), .B(new_n22215), .Y(new_n22223));
  nor_5  g19875(.A(new_n22223), .B(new_n22214), .Y(new_n22224));
  nor_5  g19876(.A(new_n22224), .B(new_n22213_1), .Y(new_n22225));
  nor_5  g19877(.A(new_n22225), .B(new_n22212), .Y(new_n22226));
  nor_5  g19878(.A(new_n22226), .B(new_n22211), .Y(new_n22227));
  nor_5  g19879(.A(new_n22227), .B(new_n22210), .Y(new_n22228));
  nor_5  g19880(.A(new_n22228), .B(new_n22209), .Y(new_n22229));
  nor_5  g19881(.A(new_n22229), .B(new_n22208), .Y(new_n22230));
  nor_5  g19882(.A(new_n22230), .B(new_n22207), .Y(new_n22231));
  or_5   g19883(.A(new_n22231), .B(new_n22206), .Y(new_n22232));
  xor_4  g19884(.A(new_n22232), .B(new_n22205), .Y(new_n22233));
  nor_5  g19885(.A(new_n22233), .B(n10514), .Y(new_n22234));
  xnor_4 g19886(.A(new_n22233), .B(new_n20222), .Y(new_n22235));
  xnor_4 g19887(.A(new_n22230), .B(new_n22207), .Y(new_n22236));
  nor_5  g19888(.A(new_n22236), .B(new_n11276), .Y(new_n22237));
  xnor_4 g19889(.A(new_n22236), .B(new_n11276), .Y(new_n22238));
  xnor_4 g19890(.A(new_n22228), .B(new_n22209), .Y(new_n22239));
  nor_5  g19891(.A(new_n22239), .B(new_n11389), .Y(new_n22240));
  xnor_4 g19892(.A(new_n22239), .B(new_n11389), .Y(new_n22241));
  xnor_4 g19893(.A(new_n22226), .B(new_n22211), .Y(new_n22242));
  nor_5  g19894(.A(new_n22242), .B(new_n10824), .Y(new_n22243));
  xnor_4 g19895(.A(new_n22242), .B(new_n10824), .Y(new_n22244));
  xnor_4 g19896(.A(new_n22224), .B(new_n22213_1), .Y(new_n22245));
  nor_5  g19897(.A(new_n22245), .B(new_n10837), .Y(new_n22246));
  xnor_4 g19898(.A(new_n22245), .B(new_n10837), .Y(new_n22247));
  xnor_4 g19899(.A(new_n22222), .B(new_n22215), .Y(new_n22248));
  nor_5  g19900(.A(new_n22248), .B(new_n20239), .Y(new_n22249));
  xnor_4 g19901(.A(new_n22248), .B(n9832), .Y(new_n22250));
  xnor_4 g19902(.A(n19608), .B(new_n15736), .Y(new_n22251));
  xnor_4 g19903(.A(new_n22251), .B(new_n22220), .Y(new_n22252));
  nor_5  g19904(.A(new_n22252), .B(n1558), .Y(new_n22253_1));
  xnor_4 g19905(.A(new_n22252), .B(new_n9479), .Y(new_n22254));
  nor_5  g19906(.A(new_n21978), .B(n21749), .Y(new_n22255));
  nor_5  g19907(.A(new_n21986_1), .B(new_n21979), .Y(new_n22256));
  or_5   g19908(.A(new_n22256), .B(new_n22255), .Y(new_n22257));
  and_5  g19909(.A(new_n22257), .B(new_n22254), .Y(new_n22258));
  nor_5  g19910(.A(new_n22258), .B(new_n22253_1), .Y(new_n22259));
  and_5  g19911(.A(new_n22259), .B(new_n22250), .Y(new_n22260));
  nor_5  g19912(.A(new_n22260), .B(new_n22249), .Y(new_n22261));
  nor_5  g19913(.A(new_n22261), .B(new_n22247), .Y(new_n22262));
  nor_5  g19914(.A(new_n22262), .B(new_n22246), .Y(new_n22263));
  nor_5  g19915(.A(new_n22263), .B(new_n22244), .Y(new_n22264));
  nor_5  g19916(.A(new_n22264), .B(new_n22243), .Y(new_n22265));
  nor_5  g19917(.A(new_n22265), .B(new_n22241), .Y(new_n22266));
  nor_5  g19918(.A(new_n22266), .B(new_n22240), .Y(new_n22267));
  nor_5  g19919(.A(new_n22267), .B(new_n22238), .Y(new_n22268));
  nor_5  g19920(.A(new_n22268), .B(new_n22237), .Y(new_n22269));
  and_5  g19921(.A(new_n22269), .B(new_n22235), .Y(new_n22270_1));
  nor_5  g19922(.A(new_n22270_1), .B(new_n22234), .Y(new_n22271));
  nor_5  g19923(.A(n7569), .B(n2570), .Y(new_n22272));
  and_5  g19924(.A(new_n22232), .B(new_n22205), .Y(new_n22273));
  or_5   g19925(.A(new_n22273), .B(new_n22272), .Y(new_n22274_1));
  xor_4  g19926(.A(new_n22274_1), .B(new_n22271), .Y(new_n22275));
  not_8  g19927(.A(new_n22085), .Y(new_n22276));
  nor_5  g19928(.A(new_n22276), .B(n3795), .Y(new_n22277));
  not_8  g19929(.A(new_n22277), .Y(new_n22278));
  nor_5  g19930(.A(new_n22278), .B(n6105), .Y(new_n22279));
  xnor_4 g19931(.A(new_n22279), .B(new_n11026), .Y(new_n22280));
  xnor_4 g19932(.A(new_n22277), .B(n6105), .Y(new_n22281));
  nor_5  g19933(.A(new_n22281), .B(new_n8718), .Y(new_n22282));
  xnor_4 g19934(.A(new_n22281), .B(new_n11032), .Y(new_n22283_1));
  nor_5  g19935(.A(new_n22086), .B(new_n8788), .Y(new_n22284));
  nor_5  g19936(.A(new_n22100), .B(new_n22087), .Y(new_n22285));
  or_5   g19937(.A(new_n22285), .B(new_n22284), .Y(new_n22286));
  and_5  g19938(.A(new_n22286), .B(new_n22283_1), .Y(new_n22287));
  nor_5  g19939(.A(new_n22287), .B(new_n22282), .Y(new_n22288));
  xnor_4 g19940(.A(new_n22288), .B(new_n22280), .Y(new_n22289));
  not_8  g19941(.A(new_n22289), .Y(new_n22290_1));
  xnor_4 g19942(.A(new_n22290_1), .B(new_n22275), .Y(new_n22291));
  xnor_4 g19943(.A(new_n22269), .B(new_n22235), .Y(new_n22292));
  nor_5  g19944(.A(new_n22285), .B(new_n22284), .Y(new_n22293));
  xnor_4 g19945(.A(new_n22293), .B(new_n22283_1), .Y(new_n22294));
  and_5  g19946(.A(new_n22294), .B(new_n22292), .Y(new_n22295));
  xnor_4 g19947(.A(new_n22294), .B(new_n22292), .Y(new_n22296));
  xnor_4 g19948(.A(new_n22267), .B(new_n22238), .Y(new_n22297));
  nor_5  g19949(.A(new_n22297), .B(new_n22101), .Y(new_n22298));
  xnor_4 g19950(.A(new_n22297), .B(new_n22101), .Y(new_n22299));
  xnor_4 g19951(.A(new_n22265), .B(new_n22241), .Y(new_n22300));
  nor_5  g19952(.A(new_n22300), .B(new_n22104), .Y(new_n22301));
  xnor_4 g19953(.A(new_n22300), .B(new_n22104), .Y(new_n22302));
  xnor_4 g19954(.A(new_n22263), .B(new_n22244), .Y(new_n22303));
  nor_5  g19955(.A(new_n22303), .B(new_n22108), .Y(new_n22304));
  xnor_4 g19956(.A(new_n22303), .B(new_n22108), .Y(new_n22305));
  xnor_4 g19957(.A(new_n22261), .B(new_n22247), .Y(new_n22306));
  nor_5  g19958(.A(new_n22306), .B(new_n18713), .Y(new_n22307));
  xnor_4 g19959(.A(new_n22306), .B(new_n18713), .Y(new_n22308));
  xnor_4 g19960(.A(new_n22259), .B(new_n22250), .Y(new_n22309_1));
  nor_5  g19961(.A(new_n22309_1), .B(new_n18039), .Y(new_n22310));
  xnor_4 g19962(.A(new_n22309_1), .B(new_n18039), .Y(new_n22311_1));
  xor_4  g19963(.A(new_n22257), .B(new_n22254), .Y(new_n22312));
  nor_5  g19964(.A(new_n22312), .B(new_n18057), .Y(new_n22313));
  not_8  g19965(.A(new_n18061_1), .Y(new_n22314));
  nor_5  g19966(.A(new_n21987), .B(new_n22314), .Y(new_n22315));
  and_5  g19967(.A(new_n21994), .B(new_n21988), .Y(new_n22316));
  nor_5  g19968(.A(new_n22316), .B(new_n22315), .Y(new_n22317_1));
  xnor_4 g19969(.A(new_n22312), .B(new_n18057), .Y(new_n22318));
  not_8  g19970(.A(new_n22318), .Y(new_n22319));
  and_5  g19971(.A(new_n22319), .B(new_n22317_1), .Y(new_n22320));
  nor_5  g19972(.A(new_n22320), .B(new_n22313), .Y(new_n22321));
  nor_5  g19973(.A(new_n22321), .B(new_n22311_1), .Y(new_n22322));
  nor_5  g19974(.A(new_n22322), .B(new_n22310), .Y(new_n22323));
  nor_5  g19975(.A(new_n22323), .B(new_n22308), .Y(new_n22324));
  nor_5  g19976(.A(new_n22324), .B(new_n22307), .Y(new_n22325));
  nor_5  g19977(.A(new_n22325), .B(new_n22305), .Y(new_n22326));
  nor_5  g19978(.A(new_n22326), .B(new_n22304), .Y(new_n22327));
  nor_5  g19979(.A(new_n22327), .B(new_n22302), .Y(new_n22328));
  nor_5  g19980(.A(new_n22328), .B(new_n22301), .Y(new_n22329));
  nor_5  g19981(.A(new_n22329), .B(new_n22299), .Y(new_n22330));
  nor_5  g19982(.A(new_n22330), .B(new_n22298), .Y(new_n22331));
  nor_5  g19983(.A(new_n22331), .B(new_n22296), .Y(new_n22332_1));
  nor_5  g19984(.A(new_n22332_1), .B(new_n22295), .Y(new_n22333));
  xnor_4 g19985(.A(new_n22333), .B(new_n22291), .Y(n11462));
  xnor_4 g19986(.A(new_n19871), .B(new_n19848), .Y(n11470));
  xnor_4 g19987(.A(new_n15157), .B(new_n15143), .Y(n11472));
  xnor_4 g19988(.A(new_n18533), .B(new_n7323), .Y(new_n22337));
  xnor_4 g19989(.A(new_n22337), .B(new_n18547), .Y(n11496));
  xnor_4 g19990(.A(new_n19655), .B(new_n19623_1), .Y(n11506));
  xnor_4 g19991(.A(new_n21349_1), .B(new_n5710), .Y(new_n22340));
  nor_5  g19992(.A(new_n15486), .B(new_n5714), .Y(new_n22341_1));
  xnor_4 g19993(.A(new_n15486), .B(new_n5714), .Y(new_n22342));
  nor_5  g19994(.A(new_n10526), .B(new_n5718), .Y(new_n22343));
  xnor_4 g19995(.A(new_n10526), .B(new_n5718), .Y(new_n22344));
  nor_5  g19996(.A(new_n10544), .B(new_n5722), .Y(new_n22345));
  xnor_4 g19997(.A(new_n10544), .B(new_n5722), .Y(new_n22346));
  nor_5  g19998(.A(new_n10549), .B(new_n5726), .Y(new_n22347));
  nor_5  g19999(.A(new_n21916), .B(new_n21903), .Y(new_n22348));
  nor_5  g20000(.A(new_n22348), .B(new_n22347), .Y(new_n22349));
  nor_5  g20001(.A(new_n22349), .B(new_n22346), .Y(new_n22350));
  nor_5  g20002(.A(new_n22350), .B(new_n22345), .Y(new_n22351));
  nor_5  g20003(.A(new_n22351), .B(new_n22344), .Y(new_n22352));
  nor_5  g20004(.A(new_n22352), .B(new_n22343), .Y(new_n22353_1));
  nor_5  g20005(.A(new_n22353_1), .B(new_n22342), .Y(new_n22354));
  nor_5  g20006(.A(new_n22354), .B(new_n22341_1), .Y(new_n22355));
  xnor_4 g20007(.A(new_n22355), .B(new_n22340), .Y(n11515));
  xnor_4 g20008(.A(new_n20534), .B(new_n20504), .Y(n11538));
  xnor_4 g20009(.A(new_n18331), .B(new_n18330), .Y(n11548));
  xnor_4 g20010(.A(new_n18577), .B(new_n18572_1), .Y(n11564));
  nor_5  g20011(.A(new_n8271), .B(n8856), .Y(new_n22360));
  and_5  g20012(.A(new_n21249), .B(new_n21246), .Y(new_n22361));
  nor_5  g20013(.A(new_n22361), .B(new_n22360), .Y(new_n22362));
  nor_5  g20014(.A(n3324), .B(n2272), .Y(new_n22363));
  and_5  g20015(.A(new_n21254_1), .B(new_n21251), .Y(new_n22364));
  nor_5  g20016(.A(new_n22364), .B(new_n22363), .Y(new_n22365));
  nor_5  g20017(.A(new_n22365), .B(new_n7500), .Y(new_n22366));
  nor_5  g20018(.A(new_n21255), .B(new_n7522), .Y(new_n22367));
  nor_5  g20019(.A(new_n21259), .B(new_n21256), .Y(new_n22368));
  nor_5  g20020(.A(new_n22368), .B(new_n22367), .Y(new_n22369));
  xnor_4 g20021(.A(new_n22365), .B(new_n7499), .Y(new_n22370));
  and_5  g20022(.A(new_n22370), .B(new_n22369), .Y(new_n22371));
  nor_5  g20023(.A(new_n22371), .B(new_n22366), .Y(new_n22372));
  not_8  g20024(.A(new_n22372), .Y(new_n22373));
  xnor_4 g20025(.A(new_n22373), .B(new_n22362), .Y(new_n22374));
  xnor_4 g20026(.A(new_n22370), .B(new_n22369), .Y(new_n22375));
  nor_5  g20027(.A(new_n22375), .B(new_n22362), .Y(new_n22376));
  not_8  g20028(.A(new_n22375), .Y(new_n22377));
  xnor_4 g20029(.A(new_n22377), .B(new_n22362), .Y(new_n22378));
  not_8  g20030(.A(new_n21260), .Y(new_n22379_1));
  and_5  g20031(.A(new_n22379_1), .B(new_n21250), .Y(new_n22380));
  and_5  g20032(.A(new_n21264), .B(new_n21261), .Y(new_n22381));
  nor_5  g20033(.A(new_n22381), .B(new_n22380), .Y(new_n22382));
  and_5  g20034(.A(new_n22382), .B(new_n22378), .Y(new_n22383));
  nor_5  g20035(.A(new_n22383), .B(new_n22376), .Y(new_n22384));
  xnor_4 g20036(.A(new_n22384), .B(new_n22374), .Y(n11591));
  or_5   g20037(.A(new_n8327), .B(new_n8320_1), .Y(new_n22386));
  nor_5  g20038(.A(new_n21926), .B(new_n8329), .Y(new_n22387));
  nor_5  g20039(.A(new_n8340), .B(new_n8328), .Y(new_n22388));
  nor_5  g20040(.A(new_n8391), .B(new_n22388), .Y(new_n22389));
  or_5   g20041(.A(new_n22389), .B(new_n21918), .Y(new_n22390));
  nor_5  g20042(.A(new_n22390), .B(new_n22387), .Y(new_n22391));
  and_5  g20043(.A(new_n22391), .B(new_n22386), .Y(n11607));
  xnor_4 g20044(.A(new_n18274_1), .B(new_n18249), .Y(n11647));
  xor_4  g20045(.A(new_n22177), .B(new_n22174), .Y(n11674));
  xnor_4 g20046(.A(new_n19155), .B(new_n20185), .Y(new_n22395));
  nor_5  g20047(.A(new_n19167), .B(new_n20185), .Y(new_n22396));
  and_5  g20048(.A(new_n20835), .B(new_n20824), .Y(new_n22397));
  or_5   g20049(.A(new_n22397), .B(new_n22396), .Y(new_n22398));
  xor_4  g20050(.A(new_n22398), .B(new_n22395), .Y(n11682));
  xor_4  g20051(.A(new_n21450), .B(new_n21439), .Y(n11710));
  xnor_4 g20052(.A(new_n13588), .B(new_n13565), .Y(n11712));
  xnor_4 g20053(.A(new_n21131), .B(new_n21118), .Y(n11724));
  xnor_4 g20054(.A(new_n17721_1), .B(new_n17720), .Y(n11741));
  not_8  g20055(.A(new_n3064), .Y(new_n22404));
  xnor_4 g20056(.A(new_n17476), .B(new_n22404), .Y(n11770));
  xnor_4 g20057(.A(new_n8378), .B(new_n8377), .Y(n11771));
  xnor_4 g20058(.A(new_n18440), .B(new_n18411), .Y(n11818));
  xnor_4 g20059(.A(new_n21912), .B(new_n21907), .Y(n11837));
  not_8  g20060(.A(new_n15833), .Y(new_n22409));
  nor_5  g20061(.A(new_n22409), .B(n7026), .Y(new_n22410));
  xnor_4 g20062(.A(new_n22410), .B(n2743), .Y(new_n22411));
  and_5  g20063(.A(new_n22411), .B(new_n5914), .Y(new_n22412));
  xnor_4 g20064(.A(new_n22411), .B(new_n5915), .Y(new_n22413));
  and_5  g20065(.A(new_n15834), .B(new_n5919), .Y(new_n22414));
  and_5  g20066(.A(new_n15872), .B(new_n15835), .Y(new_n22415));
  or_5   g20067(.A(new_n22415), .B(new_n22414), .Y(new_n22416));
  and_5  g20068(.A(new_n22416), .B(new_n22413), .Y(new_n22417));
  nor_5  g20069(.A(new_n22417), .B(new_n22412), .Y(new_n22418));
  not_8  g20070(.A(new_n22418), .Y(new_n22419));
  and_5  g20071(.A(new_n22410), .B(new_n13254), .Y(new_n22420));
  xnor_4 g20072(.A(new_n22420), .B(new_n13193), .Y(new_n22421));
  xnor_4 g20073(.A(new_n22421), .B(new_n22419), .Y(new_n22422));
  xnor_4 g20074(.A(new_n22422), .B(new_n21190), .Y(new_n22423));
  xor_4  g20075(.A(new_n22416), .B(new_n22413), .Y(new_n22424));
  nor_5  g20076(.A(new_n22424), .B(new_n21192), .Y(new_n22425));
  xnor_4 g20077(.A(new_n22424), .B(new_n21192), .Y(new_n22426));
  nor_5  g20078(.A(new_n15883), .B(new_n15873), .Y(new_n22427));
  nor_5  g20079(.A(new_n15923), .B(new_n15884_1), .Y(new_n22428));
  nor_5  g20080(.A(new_n22428), .B(new_n22427), .Y(new_n22429));
  nor_5  g20081(.A(new_n22429), .B(new_n22426), .Y(new_n22430));
  nor_5  g20082(.A(new_n22430), .B(new_n22425), .Y(new_n22431));
  xnor_4 g20083(.A(new_n22431), .B(new_n22423), .Y(n11842));
  xnor_4 g20084(.A(new_n15451), .B(new_n15434), .Y(n11843));
  xnor_4 g20085(.A(new_n18075), .B(new_n18059_1), .Y(n11905));
  xnor_4 g20086(.A(new_n11251), .B(new_n11246), .Y(n11965));
  xnor_4 g20087(.A(new_n17966), .B(new_n17963_1), .Y(n12000));
  xor_4  g20088(.A(new_n15996), .B(new_n15993), .Y(n12003));
  xnor_4 g20089(.A(new_n16577), .B(new_n16576), .Y(n12011));
  xnor_4 g20090(.A(new_n17070_1), .B(new_n17056), .Y(n12072));
  xor_4  g20091(.A(new_n10601), .B(new_n10599), .Y(n12131));
  xor_4  g20092(.A(new_n15971), .B(new_n15941), .Y(n12146));
  xnor_4 g20093(.A(new_n16213), .B(new_n16210), .Y(n12157));
  xnor_4 g20094(.A(new_n10159), .B(new_n10108), .Y(n12158));
  xnor_4 g20095(.A(new_n21529), .B(new_n21510), .Y(n12179));
  xnor_4 g20096(.A(new_n6417), .B(new_n6370), .Y(n12192));
  xnor_4 g20097(.A(new_n21851), .B(new_n21842), .Y(n12223));
  xnor_4 g20098(.A(new_n10157), .B(new_n10112), .Y(n12225));
  xnor_4 g20099(.A(new_n21914), .B(new_n21905_1), .Y(n12228));
  xnor_4 g20100(.A(new_n13129), .B(new_n7199), .Y(n12235));
  xnor_4 g20101(.A(new_n9047_1), .B(new_n9021), .Y(n12302));
  xnor_4 g20102(.A(new_n16359), .B(new_n16331), .Y(n12304));
  xnor_4 g20103(.A(n19196), .B(n1742), .Y(new_n22452));
  nor_5  g20104(.A(new_n11812), .B(n4858), .Y(new_n22453));
  xnor_4 g20105(.A(n23586), .B(n4858), .Y(new_n22454));
  nor_5  g20106(.A(new_n15238), .B(n8244), .Y(new_n22455));
  xnor_4 g20107(.A(n21226), .B(n8244), .Y(new_n22456));
  nor_5  g20108(.A(n9493), .B(new_n6170), .Y(new_n22457));
  nor_5  g20109(.A(n20036), .B(new_n12132), .Y(new_n22458));
  and_5  g20110(.A(new_n19095), .B(new_n19090), .Y(new_n22459));
  nor_5  g20111(.A(new_n22459), .B(new_n22458), .Y(new_n22460));
  xnor_4 g20112(.A(n9493), .B(n4426), .Y(new_n22461));
  and_5  g20113(.A(new_n22461), .B(new_n22460), .Y(new_n22462));
  or_5   g20114(.A(new_n22462), .B(new_n22457), .Y(new_n22463));
  and_5  g20115(.A(new_n22463), .B(new_n22456), .Y(new_n22464));
  or_5   g20116(.A(new_n22464), .B(new_n22455), .Y(new_n22465));
  and_5  g20117(.A(new_n22465), .B(new_n22454), .Y(new_n22466));
  or_5   g20118(.A(new_n22466), .B(new_n22453), .Y(new_n22467_1));
  xor_4  g20119(.A(new_n22467_1), .B(new_n22452), .Y(new_n22468));
  xnor_4 g20120(.A(new_n22468), .B(new_n19050), .Y(new_n22469));
  xor_4  g20121(.A(new_n22465), .B(new_n22454), .Y(new_n22470_1));
  nor_5  g20122(.A(new_n22470_1), .B(new_n17704), .Y(new_n22471));
  xnor_4 g20123(.A(new_n22470_1), .B(new_n17704), .Y(new_n22472));
  xor_4  g20124(.A(new_n22463), .B(new_n22456), .Y(new_n22473));
  nor_5  g20125(.A(new_n22473), .B(new_n17706), .Y(new_n22474));
  xnor_4 g20126(.A(new_n22473), .B(new_n17706), .Y(new_n22475));
  xnor_4 g20127(.A(new_n22461), .B(new_n22460), .Y(new_n22476));
  and_5  g20128(.A(new_n22476), .B(new_n17711), .Y(new_n22477));
  xnor_4 g20129(.A(new_n22476), .B(new_n17711), .Y(new_n22478));
  and_5  g20130(.A(new_n19096), .B(new_n17713), .Y(new_n22479));
  nor_5  g20131(.A(new_n19105), .B(new_n19097), .Y(new_n22480));
  nor_5  g20132(.A(new_n22480), .B(new_n22479), .Y(new_n22481));
  nor_5  g20133(.A(new_n22481), .B(new_n22478), .Y(new_n22482));
  nor_5  g20134(.A(new_n22482), .B(new_n22477), .Y(new_n22483));
  nor_5  g20135(.A(new_n22483), .B(new_n22475), .Y(new_n22484_1));
  nor_5  g20136(.A(new_n22484_1), .B(new_n22474), .Y(new_n22485));
  nor_5  g20137(.A(new_n22485), .B(new_n22472), .Y(new_n22486));
  nor_5  g20138(.A(new_n22486), .B(new_n22471), .Y(new_n22487));
  xnor_4 g20139(.A(new_n22487), .B(new_n22469), .Y(n12324));
  xnor_4 g20140(.A(new_n20830), .B(new_n20827), .Y(n12325));
  xor_4  g20141(.A(new_n10393), .B(new_n10377), .Y(n12329));
  xnor_4 g20142(.A(new_n8639), .B(new_n8638_1), .Y(n12330));
  xnor_4 g20143(.A(new_n5759), .B(new_n5716), .Y(n12346));
  xnor_4 g20144(.A(new_n7592), .B(new_n7573), .Y(n12349));
  xnor_4 g20145(.A(new_n18846), .B(new_n18845), .Y(n12364));
  nor_5  g20146(.A(new_n21424), .B(new_n5699), .Y(new_n22495));
  xnor_4 g20147(.A(new_n21425), .B(new_n5699), .Y(new_n22496));
  nor_5  g20148(.A(new_n21424), .B(new_n5702), .Y(new_n22497));
  xnor_4 g20149(.A(new_n21424), .B(new_n5702), .Y(new_n22498));
  nor_5  g20150(.A(new_n21347), .B(new_n5706), .Y(new_n22499));
  xnor_4 g20151(.A(new_n21347), .B(new_n5706), .Y(new_n22500));
  nor_5  g20152(.A(new_n21349_1), .B(new_n5710), .Y(new_n22501));
  nor_5  g20153(.A(new_n22355), .B(new_n22340), .Y(new_n22502));
  nor_5  g20154(.A(new_n22502), .B(new_n22501), .Y(new_n22503));
  nor_5  g20155(.A(new_n22503), .B(new_n22500), .Y(new_n22504));
  nor_5  g20156(.A(new_n22504), .B(new_n22499), .Y(new_n22505));
  nor_5  g20157(.A(new_n22505), .B(new_n22498), .Y(new_n22506));
  nor_5  g20158(.A(new_n22506), .B(new_n22497), .Y(new_n22507));
  and_5  g20159(.A(new_n22507), .B(new_n22496), .Y(new_n22508));
  nor_5  g20160(.A(new_n22508), .B(new_n22495), .Y(n12383));
  xnor_4 g20161(.A(new_n8558), .B(new_n8557), .Y(n12397));
  xor_4  g20162(.A(new_n16718), .B(new_n16706), .Y(n12408));
  nor_5  g20163(.A(new_n19155), .B(new_n15180_1), .Y(new_n22512));
  and_5  g20164(.A(new_n22398), .B(new_n22395), .Y(new_n22513));
  nor_5  g20165(.A(new_n22513), .B(new_n22512), .Y(n12449));
  xnor_4 g20166(.A(new_n20619), .B(new_n20587), .Y(n12461));
  not_8  g20167(.A(new_n16797), .Y(new_n22516));
  nor_5  g20168(.A(new_n20458), .B(new_n11846), .Y(new_n22517));
  nor_5  g20169(.A(new_n22517), .B(new_n22516), .Y(new_n22518));
  and_5  g20170(.A(new_n22517), .B(new_n22516), .Y(new_n22519));
  nor_5  g20171(.A(new_n20459), .B(new_n16853), .Y(new_n22520));
  nor_5  g20172(.A(new_n20468), .B(new_n20460), .Y(new_n22521));
  nor_5  g20173(.A(new_n22521), .B(new_n22520), .Y(new_n22522));
  nor_5  g20174(.A(new_n22522), .B(new_n22519), .Y(new_n22523));
  or_5   g20175(.A(new_n22523), .B(new_n22518), .Y(n12462));
  xor_4  g20176(.A(new_n21541), .B(new_n21535), .Y(n12467));
  nor_5  g20177(.A(new_n15563), .B(n3324), .Y(new_n22526));
  or_5   g20178(.A(new_n15595), .B(new_n15568), .Y(new_n22527));
  and_5  g20179(.A(new_n22527), .B(new_n15565), .Y(new_n22528));
  nor_5  g20180(.A(new_n22528), .B(new_n22526), .Y(new_n22529));
  not_8  g20181(.A(new_n22529), .Y(new_n22530));
  nor_5  g20182(.A(new_n22530), .B(new_n21214), .Y(new_n22531));
  nor_5  g20183(.A(new_n15672), .B(new_n15665), .Y(new_n22532));
  nor_5  g20184(.A(new_n15671), .B(n13419), .Y(new_n22533_1));
  nor_5  g20185(.A(new_n22533_1), .B(new_n22532), .Y(new_n22534));
  not_8  g20186(.A(new_n22534), .Y(new_n22535));
  nor_5  g20187(.A(new_n22535), .B(new_n21944), .Y(new_n22536));
  xnor_4 g20188(.A(new_n22529), .B(new_n21214), .Y(new_n22537));
  xnor_4 g20189(.A(new_n22535), .B(new_n21943_1), .Y(new_n22538));
  nor_5  g20190(.A(new_n22538), .B(new_n22537), .Y(new_n22539));
  xnor_4 g20191(.A(new_n22538), .B(new_n22537), .Y(new_n22540));
  not_8  g20192(.A(new_n22540), .Y(new_n22541));
  nor_5  g20193(.A(new_n15673), .B(new_n15597), .Y(new_n22542));
  and_5  g20194(.A(new_n15715), .B(new_n15674), .Y(new_n22543));
  nor_5  g20195(.A(new_n22543), .B(new_n22542), .Y(new_n22544));
  and_5  g20196(.A(new_n22544), .B(new_n22541), .Y(new_n22545));
  nor_5  g20197(.A(new_n22545), .B(new_n22539), .Y(new_n22546));
  xor_4  g20198(.A(new_n22546), .B(new_n22536), .Y(new_n22547));
  xnor_4 g20199(.A(new_n22547), .B(new_n22531), .Y(n12469));
  xnor_4 g20200(.A(new_n10866), .B(new_n10842), .Y(n12515));
  nor_5  g20201(.A(new_n11795), .B(n5140), .Y(new_n22550));
  xnor_4 g20202(.A(n10250), .B(n5140), .Y(new_n22551));
  nor_5  g20203(.A(new_n6155), .B(n6204), .Y(new_n22552));
  xnor_4 g20204(.A(n7674), .B(n6204), .Y(new_n22553));
  nor_5  g20205(.A(new_n6158), .B(n3349), .Y(new_n22554_1));
  xnor_4 g20206(.A(n6397), .B(n3349), .Y(new_n22555));
  nor_5  g20207(.A(new_n6161), .B(n1742), .Y(new_n22556));
  and_5  g20208(.A(new_n22467_1), .B(new_n22452), .Y(new_n22557));
  or_5   g20209(.A(new_n22557), .B(new_n22556), .Y(new_n22558));
  and_5  g20210(.A(new_n22558), .B(new_n22555), .Y(new_n22559));
  or_5   g20211(.A(new_n22559), .B(new_n22554_1), .Y(new_n22560));
  and_5  g20212(.A(new_n22560), .B(new_n22553), .Y(new_n22561));
  or_5   g20213(.A(new_n22561), .B(new_n22552), .Y(new_n22562));
  and_5  g20214(.A(new_n22562), .B(new_n22551), .Y(new_n22563));
  nor_5  g20215(.A(new_n22563), .B(new_n22550), .Y(new_n22564));
  xnor_4 g20216(.A(new_n22564), .B(new_n21291), .Y(new_n22565));
  and_5  g20217(.A(new_n22564), .B(new_n20203), .Y(new_n22566));
  or_5   g20218(.A(new_n22564), .B(new_n20203), .Y(new_n22567));
  xor_4  g20219(.A(new_n22562), .B(new_n22551), .Y(new_n22568));
  nor_5  g20220(.A(new_n22568), .B(new_n20205), .Y(new_n22569));
  xnor_4 g20221(.A(new_n22568), .B(new_n20205), .Y(new_n22570));
  xor_4  g20222(.A(new_n22560), .B(new_n22553), .Y(new_n22571));
  nor_5  g20223(.A(new_n22571), .B(new_n19045), .Y(new_n22572));
  xnor_4 g20224(.A(new_n22571), .B(new_n19045), .Y(new_n22573));
  xor_4  g20225(.A(new_n22558), .B(new_n22555), .Y(new_n22574));
  nor_5  g20226(.A(new_n22574), .B(new_n19047), .Y(new_n22575));
  xnor_4 g20227(.A(new_n22574), .B(new_n19047), .Y(new_n22576));
  nor_5  g20228(.A(new_n22468), .B(new_n19050), .Y(new_n22577));
  nor_5  g20229(.A(new_n22487), .B(new_n22469), .Y(new_n22578));
  nor_5  g20230(.A(new_n22578), .B(new_n22577), .Y(new_n22579));
  nor_5  g20231(.A(new_n22579), .B(new_n22576), .Y(new_n22580));
  nor_5  g20232(.A(new_n22580), .B(new_n22575), .Y(new_n22581));
  nor_5  g20233(.A(new_n22581), .B(new_n22573), .Y(new_n22582));
  nor_5  g20234(.A(new_n22582), .B(new_n22572), .Y(new_n22583));
  nor_5  g20235(.A(new_n22583), .B(new_n22570), .Y(new_n22584_1));
  nor_5  g20236(.A(new_n22584_1), .B(new_n22569), .Y(new_n22585));
  and_5  g20237(.A(new_n22585), .B(new_n22567), .Y(new_n22586));
  nor_5  g20238(.A(new_n22586), .B(new_n22566), .Y(new_n22587));
  xnor_4 g20239(.A(new_n22587), .B(new_n22565), .Y(n12516));
  xnor_4 g20240(.A(new_n7410), .B(new_n7397), .Y(n12540));
  xnor_4 g20241(.A(new_n11565), .B(new_n11564_1), .Y(n12545));
  xnor_4 g20242(.A(new_n19869), .B(new_n19851), .Y(n12552));
  xnor_4 g20243(.A(new_n8190), .B(new_n8167), .Y(n12566));
  xnor_4 g20244(.A(new_n13091), .B(new_n13075), .Y(n12569));
  xnor_4 g20245(.A(new_n6421), .B(new_n6359), .Y(n12607));
  xnor_4 g20246(.A(new_n9984), .B(new_n9916), .Y(n12620));
  xnor_4 g20247(.A(new_n3717), .B(new_n3679_1), .Y(n12621));
  xnor_4 g20248(.A(new_n17896), .B(new_n17895), .Y(n12654));
  xnor_4 g20249(.A(new_n19098), .B(new_n14745), .Y(n12665));
  xnor_4 g20250(.A(new_n16753), .B(new_n16743_1), .Y(n12670));
  xnor_4 g20251(.A(new_n7581), .B(new_n2522), .Y(n12707));
  xnor_4 g20252(.A(new_n7161), .B(new_n7149_1), .Y(n12725));
  xnor_4 g20253(.A(new_n15713), .B(new_n15680), .Y(n12727));
  xor_4  g20254(.A(new_n9695_1), .B(new_n9671), .Y(n12740));
  xor_4  g20255(.A(new_n20173), .B(new_n20172), .Y(n12742));
  xnor_4 g20256(.A(new_n20364), .B(new_n2826_1), .Y(n12746));
  xor_4  g20257(.A(new_n9205), .B(new_n9204), .Y(n12756));
  xnor_4 g20258(.A(new_n7174), .B(new_n7124), .Y(n12783));
  xnor_4 g20259(.A(new_n22564), .B(new_n20203), .Y(new_n22608));
  xnor_4 g20260(.A(new_n22608), .B(new_n22585), .Y(n12801));
  xnor_4 g20261(.A(new_n17380), .B(new_n17377), .Y(n12812));
  xnor_4 g20262(.A(new_n15921), .B(new_n15888), .Y(n12816));
  nor_5  g20263(.A(new_n16936), .B(n6659), .Y(new_n22612));
  and_5  g20264(.A(new_n17949), .B(new_n17929), .Y(new_n22613));
  nor_5  g20265(.A(new_n22613), .B(new_n22612), .Y(new_n22614));
  not_8  g20266(.A(new_n22614), .Y(new_n22615));
  nor_5  g20267(.A(new_n22615), .B(new_n19325), .Y(new_n22616));
  xnor_4 g20268(.A(new_n22615), .B(new_n19324), .Y(new_n22617));
  nor_5  g20269(.A(new_n22617), .B(new_n22537), .Y(new_n22618));
  xnor_4 g20270(.A(new_n22617), .B(new_n22537), .Y(new_n22619_1));
  and_5  g20271(.A(new_n17950), .B(new_n15597), .Y(new_n22620_1));
  nor_5  g20272(.A(new_n17974), .B(new_n17951), .Y(new_n22621));
  nor_5  g20273(.A(new_n22621), .B(new_n22620_1), .Y(new_n22622));
  nor_5  g20274(.A(new_n22622), .B(new_n22619_1), .Y(new_n22623_1));
  nor_5  g20275(.A(new_n22623_1), .B(new_n22618), .Y(new_n22624));
  nor_5  g20276(.A(new_n22624), .B(new_n22616), .Y(new_n22625));
  nor_5  g20277(.A(new_n22625), .B(new_n22531), .Y(n12843));
  xnor_4 g20278(.A(new_n20409_1), .B(new_n20407), .Y(n12864));
  nor_5  g20279(.A(new_n21655), .B(new_n4839), .Y(new_n22628));
  and_5  g20280(.A(new_n21681), .B(new_n21656), .Y(new_n22629));
  nor_5  g20281(.A(new_n22629), .B(new_n22628), .Y(new_n22630));
  nor_5  g20282(.A(n21784), .B(n3740), .Y(new_n22631_1));
  and_5  g20283(.A(new_n21654_1), .B(new_n21635), .Y(new_n22632));
  nor_5  g20284(.A(new_n22632), .B(new_n22631_1), .Y(new_n22633));
  xnor_4 g20285(.A(new_n22633), .B(new_n4901), .Y(new_n22634));
  xnor_4 g20286(.A(new_n22634), .B(new_n22630), .Y(new_n22635));
  not_8  g20287(.A(new_n22635), .Y(new_n22636));
  nor_5  g20288(.A(new_n22636), .B(new_n18323_1), .Y(new_n22637));
  nor_5  g20289(.A(new_n21682), .B(new_n17136), .Y(new_n22638));
  and_5  g20290(.A(new_n21706), .B(new_n21683), .Y(new_n22639));
  or_5   g20291(.A(new_n22639), .B(new_n22638), .Y(new_n22640));
  xnor_4 g20292(.A(new_n22636), .B(new_n18322), .Y(new_n22641));
  and_5  g20293(.A(new_n22641), .B(new_n22640), .Y(new_n22642));
  nor_5  g20294(.A(new_n22642), .B(new_n22637), .Y(new_n22643));
  and_5  g20295(.A(new_n22633), .B(new_n13919), .Y(new_n22644));
  nor_5  g20296(.A(new_n22633), .B(new_n13919), .Y(new_n22645));
  nor_5  g20297(.A(new_n22645), .B(new_n22630), .Y(new_n22646));
  nor_5  g20298(.A(new_n22646), .B(new_n22644), .Y(new_n22647));
  and_5  g20299(.A(new_n22647), .B(new_n22643), .Y(n12865));
  xnor_4 g20300(.A(new_n12724), .B(new_n12707_1), .Y(n12870));
  xnor_4 g20301(.A(new_n20372), .B(new_n20354), .Y(n12873));
  not_8  g20302(.A(new_n21810), .Y(new_n22651));
  nor_5  g20303(.A(new_n22651), .B(new_n18143_1), .Y(new_n22652));
  xnor_4 g20304(.A(new_n21810), .B(new_n18144), .Y(new_n22653));
  nor_5  g20305(.A(new_n21186), .B(new_n18226), .Y(new_n22654));
  nor_5  g20306(.A(new_n22135), .B(new_n22132), .Y(new_n22655));
  nor_5  g20307(.A(new_n22655), .B(new_n22654), .Y(new_n22656));
  nor_5  g20308(.A(new_n22656), .B(new_n22653), .Y(new_n22657));
  or_5   g20309(.A(new_n22657), .B(new_n22652), .Y(n12904));
  xor_4  g20310(.A(new_n10398), .B(new_n10397), .Y(n12941));
  xnor_4 g20311(.A(new_n11137), .B(new_n11129), .Y(n12942));
  xnor_4 g20312(.A(new_n5844), .B(new_n5846), .Y(new_n22661));
  xnor_4 g20313(.A(new_n22661), .B(new_n5849), .Y(n12978));
  xnor_4 g20314(.A(new_n9709), .B(new_n7887), .Y(n12980));
  not_8  g20315(.A(new_n6568), .Y(new_n22664));
  xnor_4 g20316(.A(new_n22664), .B(new_n4711), .Y(n12985));
  xnor_4 g20317(.A(new_n14289), .B(new_n14257), .Y(n12987));
  nor_5  g20318(.A(n11220), .B(new_n12808), .Y(new_n22667));
  and_5  g20319(.A(new_n16431), .B(new_n16416), .Y(new_n22668));
  nor_5  g20320(.A(new_n22668), .B(new_n22667), .Y(new_n22669));
  xnor_4 g20321(.A(new_n22669), .B(new_n14546_1), .Y(new_n22670));
  and_5  g20322(.A(new_n16432), .B(new_n14589), .Y(new_n22671));
  and_5  g20323(.A(new_n16452), .B(new_n16433_1), .Y(new_n22672));
  nor_5  g20324(.A(new_n22672), .B(new_n22671), .Y(new_n22673));
  xnor_4 g20325(.A(new_n22673), .B(new_n22670), .Y(n12992));
  nor_5  g20326(.A(new_n21474), .B(n6659), .Y(new_n22675));
  nor_5  g20327(.A(new_n20546), .B(n23250), .Y(new_n22676));
  and_5  g20328(.A(new_n20582_1), .B(new_n20548), .Y(new_n22677));
  nor_5  g20329(.A(new_n22677), .B(new_n22676), .Y(new_n22678));
  nor_5  g20330(.A(new_n21475), .B(new_n21940), .Y(new_n22679));
  nor_5  g20331(.A(new_n22679), .B(new_n22678), .Y(new_n22680));
  nor_5  g20332(.A(new_n22680), .B(new_n22675), .Y(new_n22681));
  nor_5  g20333(.A(new_n22681), .B(new_n21473), .Y(new_n22682));
  not_8  g20334(.A(new_n22682), .Y(new_n22683));
  xnor_4 g20335(.A(new_n22683), .B(new_n19336), .Y(new_n22684));
  xnor_4 g20336(.A(new_n21475), .B(n6659), .Y(new_n22685));
  xnor_4 g20337(.A(new_n22685), .B(new_n22678), .Y(new_n22686));
  nor_5  g20338(.A(new_n22686), .B(new_n19349), .Y(new_n22687));
  nor_5  g20339(.A(new_n20583), .B(new_n14075), .Y(new_n22688));
  and_5  g20340(.A(new_n20621), .B(new_n20584), .Y(new_n22689));
  or_5   g20341(.A(new_n22689), .B(new_n22688), .Y(new_n22690));
  xnor_4 g20342(.A(new_n22686), .B(new_n19350), .Y(new_n22691));
  and_5  g20343(.A(new_n22691), .B(new_n22690), .Y(new_n22692));
  nor_5  g20344(.A(new_n22692), .B(new_n22687), .Y(new_n22693));
  xnor_4 g20345(.A(new_n22693), .B(new_n22684), .Y(n13005));
  xnor_4 g20346(.A(new_n19438), .B(new_n16307), .Y(n13043));
  xnor_4 g20347(.A(new_n17455), .B(new_n17454), .Y(n13048));
  xnor_4 g20348(.A(new_n15113), .B(new_n15112), .Y(n13054));
  xnor_4 g20349(.A(new_n17615), .B(new_n17603), .Y(n13082));
  xnor_4 g20350(.A(new_n7166), .B(new_n7140), .Y(n13096));
  xnor_4 g20351(.A(new_n17617), .B(new_n17598), .Y(n13116));
  xnor_4 g20352(.A(new_n19453), .B(new_n19420), .Y(n13122));
  xnor_4 g20353(.A(new_n6403), .B(new_n6402), .Y(n13141));
  xor_4  g20354(.A(new_n19289), .B(new_n19282_1), .Y(n13144));
  xnor_4 g20355(.A(new_n19875), .B(new_n19841), .Y(n13168));
  xnor_4 g20356(.A(new_n20528), .B(new_n20510), .Y(n13198));
  xnor_4 g20357(.A(new_n14283), .B(new_n14266), .Y(n13199));
  xnor_4 g20358(.A(new_n14397), .B(new_n14385), .Y(n13204));
  xnor_4 g20359(.A(new_n10150), .B(new_n10123), .Y(n13209));
  xnor_4 g20360(.A(new_n19086), .B(new_n19077), .Y(n13270));
  xnor_4 g20361(.A(new_n12983), .B(new_n12962), .Y(n13273));
  xnor_4 g20362(.A(new_n21531), .B(new_n21506), .Y(n13285));
  xnor_4 g20363(.A(new_n20927), .B(new_n20909), .Y(n13338));
  xnor_4 g20364(.A(new_n7904), .B(new_n7873), .Y(n13407));
  xnor_4 g20365(.A(new_n5432), .B(new_n4264), .Y(new_n22714_1));
  xnor_4 g20366(.A(new_n22714_1), .B(new_n15955), .Y(n13409));
  xnor_4 g20367(.A(new_n5445), .B(new_n5416), .Y(n13456));
  nor_5  g20368(.A(new_n20872), .B(new_n20221), .Y(new_n22717));
  nor_5  g20369(.A(new_n20903), .B(new_n20225), .Y(new_n22718));
  nor_5  g20370(.A(new_n21886), .B(new_n21883), .Y(new_n22719));
  nor_5  g20371(.A(new_n22719), .B(new_n22718), .Y(new_n22720));
  or_5   g20372(.A(new_n20793), .B(new_n20221), .Y(new_n22721));
  and_5  g20373(.A(new_n22721), .B(new_n22720), .Y(new_n22722));
  and_5  g20374(.A(new_n22722), .B(new_n22717), .Y(new_n22723));
  xnor_4 g20375(.A(new_n20794_1), .B(new_n20332), .Y(new_n22724));
  xnor_4 g20376(.A(new_n22724), .B(new_n22720), .Y(new_n22725));
  and_5  g20377(.A(new_n22725), .B(new_n11288), .Y(new_n22726));
  xnor_4 g20378(.A(new_n22725), .B(new_n11288), .Y(new_n22727));
  nor_5  g20379(.A(new_n21887), .B(new_n11380), .Y(new_n22728));
  nor_5  g20380(.A(new_n21891), .B(new_n21888), .Y(new_n22729));
  or_5   g20381(.A(new_n22729), .B(new_n22728), .Y(new_n22730));
  nor_5  g20382(.A(new_n22730), .B(new_n22727), .Y(new_n22731));
  nor_5  g20383(.A(new_n22731), .B(new_n22726), .Y(new_n22732));
  xnor_4 g20384(.A(new_n20873), .B(new_n20221), .Y(new_n22733));
  and_5  g20385(.A(new_n22733), .B(new_n22720), .Y(new_n22734));
  nor_5  g20386(.A(new_n22733), .B(new_n22722), .Y(new_n22735));
  nor_5  g20387(.A(new_n22735), .B(new_n22734), .Y(new_n22736));
  nor_5  g20388(.A(new_n22736), .B(new_n22732), .Y(new_n22737));
  or_5   g20389(.A(new_n22737), .B(new_n22723), .Y(n13457));
  xnor_4 g20390(.A(new_n12039), .B(new_n12031), .Y(n13477));
  xnor_4 g20391(.A(new_n12349_1), .B(new_n12348), .Y(n13484));
  xnor_4 g20392(.A(new_n20059), .B(new_n20031), .Y(n13486));
  xnor_4 g20393(.A(new_n21437), .B(new_n20957), .Y(new_n22742));
  and_5  g20394(.A(new_n21357), .B(new_n17024), .Y(new_n22743));
  nor_5  g20395(.A(new_n21382), .B(new_n21358), .Y(new_n22744));
  nor_5  g20396(.A(new_n22744), .B(new_n22743), .Y(new_n22745));
  xor_4  g20397(.A(new_n22745), .B(new_n22742), .Y(n13487));
  xnor_4 g20398(.A(new_n5213_1), .B(new_n5194), .Y(n13500));
  xor_4  g20399(.A(new_n4592), .B(new_n4590_1), .Y(n13501));
  xnor_4 g20400(.A(new_n6409), .B(new_n6388), .Y(n13506));
  xnor_4 g20401(.A(new_n6135), .B(new_n6124), .Y(n13548));
  xnor_4 g20402(.A(new_n22325), .B(new_n22305), .Y(n13551));
  xnor_4 g20403(.A(new_n5014), .B(new_n4995), .Y(n13602));
  xnor_4 g20404(.A(new_n17120), .B(new_n17111), .Y(n13626));
  xnor_4 g20405(.A(new_n8186), .B(new_n8177), .Y(n13683));
  xnor_4 g20406(.A(new_n19657), .B(new_n19620), .Y(n13710));
  xnor_4 g20407(.A(new_n19293), .B(new_n19276), .Y(n13722));
  xnor_4 g20408(.A(new_n13925), .B(new_n13870), .Y(new_n22757));
  xnor_4 g20409(.A(new_n22757), .B(new_n13992), .Y(n13754));
  xor_4  g20410(.A(new_n2839), .B(new_n2805), .Y(n13764));
  xnor_4 g20411(.A(new_n14142), .B(new_n14139), .Y(new_n22760));
  xnor_4 g20412(.A(new_n22760), .B(new_n14147_1), .Y(n13798));
  xnor_4 g20413(.A(new_n17124), .B(new_n17106_1), .Y(n13835));
  xnor_4 g20414(.A(new_n15537), .B(new_n15535), .Y(n13850));
  xnor_4 g20415(.A(new_n17605), .B(new_n7888), .Y(n13922));
  xnor_4 g20416(.A(new_n19057), .B(new_n19049), .Y(n13923));
  xnor_4 g20417(.A(new_n11570), .B(new_n11569), .Y(n14004));
  xnor_4 g20418(.A(new_n11787), .B(new_n11748), .Y(n14036));
  xnor_4 g20419(.A(new_n21005), .B(new_n20991), .Y(n14059));
  xor_4  g20420(.A(new_n16925), .B(new_n16922), .Y(n14081));
  xnor_4 g20421(.A(new_n18543), .B(new_n18540), .Y(n14095));
  xnor_4 g20422(.A(new_n6728), .B(new_n11603), .Y(n14107));
  xnor_4 g20423(.A(new_n8901), .B(new_n8870), .Y(n14121));
  xnor_4 g20424(.A(new_n12002), .B(new_n12000_1), .Y(n14126));
  xnor_4 g20425(.A(new_n19297), .B(new_n19270_1), .Y(n14136));
  not_8  g20426(.A(new_n22669), .Y(new_n22775));
  nor_5  g20427(.A(new_n22775), .B(new_n14546_1), .Y(new_n22776));
  nor_5  g20428(.A(new_n22669), .B(new_n14545), .Y(new_n22777));
  nor_5  g20429(.A(new_n22673), .B(new_n22777), .Y(new_n22778));
  nor_5  g20430(.A(new_n22778), .B(new_n22776), .Y(new_n22779_1));
  xnor_4 g20431(.A(new_n22775), .B(new_n21723), .Y(new_n22780));
  xnor_4 g20432(.A(new_n22780), .B(new_n22779_1), .Y(n14147));
  xnor_4 g20433(.A(new_n20738), .B(new_n20700_1), .Y(n14174));
  xnor_4 g20434(.A(new_n16221), .B(new_n16197), .Y(n14190));
  xnor_4 g20435(.A(new_n5443_1), .B(new_n5420), .Y(n14211));
  xnor_4 g20436(.A(new_n16407_1), .B(new_n16404), .Y(n14222));
  xnor_4 g20437(.A(new_n13306), .B(new_n13262), .Y(n14267));
  xnor_4 g20438(.A(new_n5749), .B(new_n5738), .Y(n14271));
  xnor_4 g20439(.A(new_n9383), .B(new_n9372_1), .Y(n14277));
  xnor_4 g20440(.A(new_n8373), .B(new_n8372), .Y(n14294));
  xnor_4 g20441(.A(new_n22331), .B(new_n22296), .Y(n14310));
  xnor_4 g20442(.A(new_n22349), .B(new_n22346), .Y(n14326));
  xnor_4 g20443(.A(new_n12306), .B(new_n12262), .Y(n14342));
  xnor_4 g20444(.A(new_n18073), .B(new_n18063), .Y(n14353));
  and_5  g20445(.A(new_n20987), .B(new_n11593), .Y(new_n22794));
  nor_5  g20446(.A(new_n20987), .B(new_n8953), .Y(new_n22795));
  nor_5  g20447(.A(new_n21007), .B(new_n20988), .Y(new_n22796));
  nor_5  g20448(.A(new_n22796), .B(new_n22795), .Y(new_n22797));
  nor_5  g20449(.A(new_n22797), .B(new_n22794), .Y(new_n22798));
  nor_5  g20450(.A(new_n20987), .B(new_n11593), .Y(new_n22799));
  nor_5  g20451(.A(new_n22799), .B(new_n22796), .Y(new_n22800));
  nor_5  g20452(.A(new_n22800), .B(new_n22798), .Y(n14364));
  xor_4  g20453(.A(new_n21445), .B(new_n21442), .Y(n14375));
  xnor_4 g20454(.A(new_n21859), .B(new_n21834), .Y(n14412));
  or_5   g20455(.A(new_n17339), .B(new_n6240), .Y(new_n22804));
  nor_5  g20456(.A(new_n17363), .B(new_n22804), .Y(new_n22805));
  xnor_4 g20457(.A(new_n22805), .B(new_n11524), .Y(new_n22806));
  and_5  g20458(.A(new_n17364), .B(new_n17331), .Y(new_n22807));
  nor_5  g20459(.A(new_n17388), .B(new_n17365), .Y(new_n22808));
  nor_5  g20460(.A(new_n22808), .B(new_n22807), .Y(new_n22809));
  not_8  g20461(.A(new_n22809), .Y(new_n22810));
  xnor_4 g20462(.A(new_n22810), .B(new_n22806), .Y(n14414));
  xnor_4 g20463(.A(new_n15310), .B(new_n15308), .Y(n14457));
  xnor_4 g20464(.A(new_n5018), .B(new_n4987), .Y(n14464));
  xnor_4 g20465(.A(new_n10864), .B(new_n10846), .Y(n14471));
  nor_5  g20466(.A(new_n19324), .B(new_n8339_1), .Y(new_n22815));
  nor_5  g20467(.A(new_n19334), .B(new_n19326), .Y(new_n22816));
  nor_5  g20468(.A(new_n22816), .B(new_n22815), .Y(new_n22817));
  not_8  g20469(.A(new_n22817), .Y(new_n22818));
  xnor_4 g20470(.A(new_n22818), .B(new_n22682), .Y(new_n22819_1));
  nor_5  g20471(.A(new_n22683), .B(new_n19335), .Y(new_n22820));
  nor_5  g20472(.A(new_n22682), .B(new_n19336), .Y(new_n22821));
  nor_5  g20473(.A(new_n22693), .B(new_n22821), .Y(new_n22822));
  nor_5  g20474(.A(new_n22822), .B(new_n22820), .Y(new_n22823));
  xnor_4 g20475(.A(new_n22823), .B(new_n22819_1), .Y(n14475));
  xnor_4 g20476(.A(new_n12294), .B(new_n12293), .Y(n14541));
  nor_5  g20477(.A(new_n21231), .B(new_n21227), .Y(new_n22826));
  nor_5  g20478(.A(new_n21241), .B(new_n21232), .Y(new_n22827));
  or_5   g20479(.A(new_n22827), .B(new_n22826), .Y(n14546));
  xnor_4 g20480(.A(new_n11065), .B(new_n11064), .Y(n14547));
  xnor_4 g20481(.A(new_n12651), .B(new_n12632), .Y(n14593));
  xnor_4 g20482(.A(new_n9387), .B(new_n9362), .Y(n14636));
  xnor_4 g20483(.A(new_n22485), .B(new_n22472), .Y(n14701));
  xnor_4 g20484(.A(new_n12089), .B(new_n12080), .Y(n14734));
  xnor_4 g20485(.A(new_n7172), .B(new_n7128), .Y(n14746));
  xnor_4 g20486(.A(new_n9687), .B(new_n9685), .Y(n14763));
  xnor_4 g20487(.A(new_n22056), .B(new_n22048), .Y(n14772));
  xnor_4 g20488(.A(new_n21448), .B(new_n21447), .Y(n14801));
  xnor_4 g20489(.A(new_n21050), .B(new_n21031), .Y(n14819));
  xnor_4 g20490(.A(new_n14405), .B(new_n14373), .Y(n14827));
  xnor_4 g20491(.A(new_n20466), .B(new_n20463), .Y(n14839));
  xnor_4 g20492(.A(new_n17116), .B(new_n17115), .Y(n14849));
  nor_5  g20493(.A(new_n20330_1), .B(new_n14356), .Y(new_n22842));
  nor_5  g20494(.A(new_n20387), .B(new_n20331), .Y(new_n22843_1));
  nor_5  g20495(.A(new_n22843_1), .B(new_n22842), .Y(new_n22844));
  nor_5  g20496(.A(new_n22844), .B(new_n20327), .Y(n14891));
  xnor_4 g20497(.A(new_n6532), .B(new_n15341), .Y(n14931));
  and_5  g20498(.A(new_n22805), .B(new_n11524), .Y(new_n22847));
  and_5  g20499(.A(new_n22810), .B(new_n22847), .Y(new_n22848));
  or_5   g20500(.A(new_n22805), .B(new_n11524), .Y(new_n22849));
  nor_5  g20501(.A(new_n22810), .B(new_n22849), .Y(new_n22850));
  or_5   g20502(.A(new_n22850), .B(new_n22848), .Y(n14944));
  xnor_4 g20503(.A(new_n18069), .B(new_n8911_1), .Y(n14977));
  xnor_4 g20504(.A(new_n12659), .B(new_n12614), .Y(n14989));
  xnor_4 g20505(.A(new_n10760), .B(new_n10752), .Y(n15002));
  xnor_4 g20506(.A(new_n21910), .B(new_n5746), .Y(n15004));
  xnor_4 g20507(.A(new_n9051), .B(new_n9013), .Y(n15011));
  xor_4  g20508(.A(new_n21965), .B(new_n21962), .Y(n15019));
  nor_5  g20509(.A(new_n15098), .B(new_n15090), .Y(new_n22858_1));
  nor_5  g20510(.A(new_n15119), .B(new_n15099), .Y(new_n22859));
  or_5   g20511(.A(new_n22859), .B(new_n22858_1), .Y(n15031));
  xnor_4 g20512(.A(new_n17606), .B(new_n17604), .Y(n15033));
  xnor_4 g20513(.A(new_n11884), .B(new_n7200), .Y(n15052));
  xnor_4 g20514(.A(new_n19210), .B(new_n19201), .Y(n15082));
  xnor_4 g20515(.A(new_n8188), .B(new_n8171), .Y(n15094));
  xor_4  g20516(.A(new_n11624), .B(new_n11621), .Y(n15118));
  xnor_4 g20517(.A(new_n22656), .B(new_n22653), .Y(n15128));
  xnor_4 g20518(.A(new_n18444_1), .B(new_n18405_1), .Y(n15139));
  xnor_4 g20519(.A(new_n16500), .B(new_n16495), .Y(new_n22868));
  xnor_4 g20520(.A(new_n22868), .B(new_n16510), .Y(n15145));
  xnor_4 g20521(.A(new_n14624), .B(new_n14594), .Y(n15165));
  xnor_4 g20522(.A(new_n15032), .B(new_n5081), .Y(n15176));
  xor_4  g20523(.A(new_n19863), .B(new_n19862), .Y(n15180));
  xnor_4 g20524(.A(new_n15973), .B(new_n15939), .Y(n15205));
  not_8  g20525(.A(new_n5436), .Y(new_n22874));
  xnor_4 g20526(.A(new_n22874), .B(new_n4266_1), .Y(n15230));
  xor_4  g20527(.A(new_n16749), .B(new_n16748), .Y(n15255));
  xnor_4 g20528(.A(new_n9699_1), .B(new_n9661), .Y(n15275));
  xnor_4 g20529(.A(new_n13766), .B(new_n13763), .Y(n15300));
  or_5   g20530(.A(new_n22420), .B(new_n13194), .Y(new_n22879_1));
  nor_5  g20531(.A(new_n22879_1), .B(new_n22419), .Y(new_n22880));
  and_5  g20532(.A(new_n22420), .B(new_n13194), .Y(new_n22881));
  and_5  g20533(.A(new_n22881), .B(new_n22419), .Y(new_n22882));
  nor_5  g20534(.A(new_n22882), .B(new_n22880), .Y(new_n22883));
  xnor_4 g20535(.A(new_n22883), .B(new_n21227), .Y(new_n22884));
  nor_5  g20536(.A(new_n22422), .B(new_n21190), .Y(new_n22885));
  nor_5  g20537(.A(new_n22431), .B(new_n22423), .Y(new_n22886));
  nor_5  g20538(.A(new_n22886), .B(new_n22885), .Y(new_n22887));
  not_8  g20539(.A(new_n22887), .Y(new_n22888));
  xnor_4 g20540(.A(new_n22888), .B(new_n22884), .Y(n15307));
  xnor_4 g20541(.A(new_n19659), .B(new_n19617_1), .Y(n15327));
  xnor_4 g20542(.A(new_n19645), .B(new_n19638), .Y(n15345));
  xnor_4 g20543(.A(new_n12649), .B(new_n12638), .Y(n15353));
  xor_4  g20544(.A(new_n22507), .B(new_n22496), .Y(n15366));
  xnor_4 g20545(.A(new_n22647), .B(new_n22643), .Y(n15382));
  xnor_4 g20546(.A(new_n9211), .B(new_n9194), .Y(n15407));
  not_8  g20547(.A(new_n13377), .Y(new_n22896));
  xnor_4 g20548(.A(new_n14962), .B(new_n22896), .Y(n15428));
  and_5  g20549(.A(new_n22274_1), .B(new_n22271), .Y(new_n22898));
  and_5  g20550(.A(new_n22290_1), .B(new_n22275), .Y(new_n22899));
  nor_5  g20551(.A(new_n22333), .B(new_n22291), .Y(new_n22900));
  nor_5  g20552(.A(new_n22900), .B(new_n22899), .Y(new_n22901));
  nor_5  g20553(.A(new_n22901), .B(new_n22898), .Y(new_n22902));
  or_5   g20554(.A(new_n22279), .B(new_n11025_1), .Y(new_n22903_1));
  nor_5  g20555(.A(new_n22288), .B(new_n22903_1), .Y(new_n22904));
  not_8  g20556(.A(new_n22904), .Y(new_n22905));
  nor_5  g20557(.A(new_n22905), .B(new_n22898), .Y(new_n22906));
  nor_5  g20558(.A(new_n22906), .B(new_n22900), .Y(new_n22907_1));
  nor_5  g20559(.A(new_n22907_1), .B(new_n22902), .Y(n15435));
  or_5   g20560(.A(new_n21924), .B(new_n21919), .Y(new_n22909));
  nor_5  g20561(.A(new_n21934_1), .B(new_n22909), .Y(new_n22910_1));
  and_5  g20562(.A(new_n21924), .B(new_n21919), .Y(new_n22911));
  and_5  g20563(.A(new_n21934_1), .B(new_n22911), .Y(new_n22912));
  or_5   g20564(.A(new_n22912), .B(new_n22910_1), .Y(n15438));
  xnor_4 g20565(.A(new_n22327), .B(new_n22302), .Y(n15465));
  xnor_4 g20566(.A(new_n8556), .B(new_n6665), .Y(n15467));
  xnor_4 g20567(.A(new_n7914), .B(new_n7843), .Y(n15470));
  xnor_4 g20568(.A(new_n14409), .B(new_n14366), .Y(n15477));
  xnor_4 g20569(.A(new_n22581), .B(new_n22573), .Y(n15481));
  xnor_4 g20570(.A(new_n14836), .B(new_n14833), .Y(n15496));
  xnor_4 g20571(.A(new_n12012), .B(new_n11983), .Y(n15501));
  xnor_4 g20572(.A(new_n18545), .B(new_n18537_1), .Y(n15555));
  xnor_4 g20573(.A(new_n20867), .B(new_n20852), .Y(n15558));
  nor_5  g20574(.A(new_n21226_1), .B(new_n22651), .Y(new_n22923));
  nor_5  g20575(.A(new_n21814), .B(new_n21811), .Y(new_n22924));
  or_5   g20576(.A(new_n22924), .B(new_n22923), .Y(n15559));
  and_5  g20577(.A(new_n5453), .B(n5101), .Y(new_n22926));
  and_5  g20578(.A(new_n19897), .B(new_n19882), .Y(new_n22927));
  nor_5  g20579(.A(new_n22927), .B(new_n22926), .Y(new_n22928));
  not_8  g20580(.A(new_n22928), .Y(new_n22929));
  nor_5  g20581(.A(new_n22929), .B(new_n22007), .Y(new_n22930));
  and_5  g20582(.A(new_n20501), .B(new_n19898), .Y(new_n22931));
  and_5  g20583(.A(new_n19972), .B(new_n19948), .Y(new_n22932));
  nor_5  g20584(.A(new_n22932), .B(new_n22931), .Y(new_n22933));
  nor_5  g20585(.A(new_n22928), .B(new_n21219), .Y(new_n22934));
  nor_5  g20586(.A(new_n22934), .B(new_n22933), .Y(new_n22935));
  and_5  g20587(.A(new_n22935), .B(new_n22007), .Y(new_n22936));
  nor_5  g20588(.A(new_n22929), .B(new_n21219), .Y(new_n22937));
  nor_5  g20589(.A(new_n22937), .B(new_n22935), .Y(new_n22938));
  or_5   g20590(.A(new_n22938), .B(new_n22936), .Y(new_n22939_1));
  nor_5  g20591(.A(new_n22939_1), .B(new_n22930), .Y(n15570));
  xnor_4 g20592(.A(new_n12312), .B(new_n12250), .Y(n15573));
  xnor_4 g20593(.A(new_n11581), .B(new_n11580_1), .Y(n15588));
  xnor_4 g20594(.A(new_n21046_1), .B(new_n21038), .Y(n15590));
  xnor_4 g20595(.A(new_n21604), .B(new_n21594), .Y(n15598));
  xnor_4 g20596(.A(new_n9389), .B(new_n9357), .Y(n15614));
  xnor_4 g20597(.A(new_n22060), .B(new_n22042), .Y(n15662));
  xnor_4 g20598(.A(new_n3383), .B(new_n3352), .Y(n15716));
  xnor_4 g20599(.A(new_n14291), .B(new_n14254), .Y(n15749));
  xnor_4 g20600(.A(new_n18463), .B(new_n18460), .Y(n15762));
  xnor_4 g20601(.A(new_n7889), .B(new_n7887), .Y(n15793));
  xnor_4 g20602(.A(new_n21853), .B(new_n21840), .Y(n15812));
  xnor_4 g20603(.A(new_n12308), .B(new_n12258), .Y(n15815));
  xnor_4 g20604(.A(new_n8370), .B(new_n8369), .Y(n15816));
  xnor_4 g20605(.A(new_n11890), .B(new_n11878), .Y(n15831));
  xnor_4 g20606(.A(new_n9561), .B(new_n9559), .Y(n15846));
  xnor_4 g20607(.A(new_n8428), .B(new_n8427), .Y(n15859));
  nor_5  g20608(.A(new_n8079), .B(new_n21421), .Y(new_n22957));
  and_5  g20609(.A(new_n19539_1), .B(new_n19524), .Y(new_n22958));
  nor_5  g20610(.A(new_n22958), .B(new_n22957), .Y(new_n22959));
  nor_5  g20611(.A(new_n22959), .B(new_n8075), .Y(new_n22960));
  xnor_4 g20612(.A(new_n22960), .B(new_n21276_1), .Y(new_n22961));
  xnor_4 g20613(.A(new_n22959), .B(new_n8074), .Y(new_n22962));
  nor_5  g20614(.A(new_n22962), .B(new_n19833), .Y(new_n22963));
  nor_5  g20615(.A(new_n19540), .B(new_n19523_1), .Y(new_n22964));
  nor_5  g20616(.A(new_n19562), .B(new_n19541), .Y(new_n22965));
  nor_5  g20617(.A(new_n22965), .B(new_n22964), .Y(new_n22966));
  xnor_4 g20618(.A(new_n22962), .B(new_n19833), .Y(new_n22967));
  nor_5  g20619(.A(new_n22967), .B(new_n22966), .Y(new_n22968));
  nor_5  g20620(.A(new_n22968), .B(new_n22963), .Y(new_n22969));
  xnor_4 g20621(.A(new_n22969), .B(new_n22961), .Y(n15869));
  xnor_4 g20622(.A(new_n18588), .B(new_n18563), .Y(n15885));
  not_8  g20623(.A(new_n20696_1), .Y(new_n22972));
  and_5  g20624(.A(new_n22972), .B(new_n15335), .Y(new_n22973));
  and_5  g20625(.A(new_n20740), .B(new_n22973), .Y(new_n22974));
  and_5  g20626(.A(new_n20739), .B(new_n20696_1), .Y(new_n22975));
  or_5   g20627(.A(new_n22975), .B(new_n22974), .Y(n15889));
  xnor_4 g20628(.A(new_n18575), .B(new_n13634), .Y(n15917));
  xnor_4 g20629(.A(new_n13628), .B(new_n13627), .Y(n15922));
  not_8  g20630(.A(new_n7150), .Y(new_n22979));
  xnor_4 g20631(.A(new_n7151), .B(new_n22979), .Y(n15947));
  and_5  g20632(.A(new_n19135), .B(new_n7241), .Y(new_n22981));
  and_5  g20633(.A(new_n20399), .B(new_n20392), .Y(new_n22982));
  nor_5  g20634(.A(new_n22982), .B(new_n22981), .Y(new_n22983));
  not_8  g20635(.A(new_n22983), .Y(new_n22984));
  xnor_4 g20636(.A(new_n22984), .B(new_n19163_1), .Y(new_n22985));
  nor_5  g20637(.A(new_n20400), .B(new_n19162), .Y(new_n22986));
  nor_5  g20638(.A(new_n20411_1), .B(new_n20402_1), .Y(new_n22987));
  nor_5  g20639(.A(new_n22987), .B(new_n22986), .Y(new_n22988));
  xor_4  g20640(.A(new_n22988), .B(new_n22985), .Y(n15956));
  xor_4  g20641(.A(new_n13398), .B(new_n13395), .Y(n15958));
  nor_5  g20642(.A(new_n16781), .B(new_n12059), .Y(new_n22991));
  and_5  g20643(.A(new_n16781), .B(new_n12063), .Y(new_n22992));
  nor_5  g20644(.A(new_n22992), .B(new_n22991), .Y(new_n22993));
  nor_5  g20645(.A(new_n16776), .B(new_n12059), .Y(new_n22994));
  or_5   g20646(.A(new_n16778), .B(new_n22994), .Y(new_n22995));
  nor_5  g20647(.A(new_n22995), .B(new_n22993), .Y(n15986));
  xnor_4 g20648(.A(new_n22429), .B(new_n22426), .Y(n16013));
  nor_5  g20649(.A(new_n21401), .B(new_n20400), .Y(new_n22998_1));
  nor_5  g20650(.A(new_n21402), .B(new_n20401), .Y(new_n22999));
  nor_5  g20651(.A(new_n21411), .B(new_n22999), .Y(new_n23000));
  nor_5  g20652(.A(new_n23000), .B(new_n22998_1), .Y(new_n23001));
  xnor_4 g20653(.A(new_n22984), .B(new_n21401), .Y(new_n23002));
  xnor_4 g20654(.A(new_n23002), .B(new_n23001), .Y(n16060));
  nor_5  g20655(.A(new_n16152), .B(new_n11842_1), .Y(new_n23004));
  xnor_4 g20656(.A(new_n16152), .B(n25972), .Y(new_n23005));
  nor_5  g20657(.A(new_n16154), .B(new_n8646), .Y(new_n23006_1));
  and_5  g20658(.A(new_n22078), .B(new_n22067), .Y(new_n23007_1));
  or_5   g20659(.A(new_n23007_1), .B(new_n23006_1), .Y(new_n23008));
  and_5  g20660(.A(new_n23008), .B(new_n23005), .Y(new_n23009_1));
  nor_5  g20661(.A(new_n23009_1), .B(new_n23004), .Y(new_n23010));
  nor_5  g20662(.A(new_n23010), .B(new_n22189), .Y(new_n23011));
  xnor_4 g20663(.A(new_n23010), .B(new_n22189), .Y(new_n23012));
  and_5  g20664(.A(new_n23012), .B(new_n22290_1), .Y(new_n23013));
  xnor_4 g20665(.A(new_n23012), .B(new_n22290_1), .Y(new_n23014_1));
  not_8  g20666(.A(new_n22294), .Y(new_n23015));
  xor_4  g20667(.A(new_n23008), .B(new_n23005), .Y(new_n23016));
  nor_5  g20668(.A(new_n23016), .B(new_n23015), .Y(new_n23017));
  xnor_4 g20669(.A(new_n23016), .B(new_n23015), .Y(new_n23018));
  nor_5  g20670(.A(new_n22101), .B(new_n22079), .Y(new_n23019));
  nor_5  g20671(.A(new_n22117), .B(new_n22102), .Y(new_n23020));
  nor_5  g20672(.A(new_n23020), .B(new_n23019), .Y(new_n23021));
  nor_5  g20673(.A(new_n23021), .B(new_n23018), .Y(new_n23022));
  nor_5  g20674(.A(new_n23022), .B(new_n23017), .Y(new_n23023));
  nor_5  g20675(.A(new_n23023), .B(new_n23014_1), .Y(new_n23024));
  nor_5  g20676(.A(new_n23024), .B(new_n23013), .Y(new_n23025));
  xnor_4 g20677(.A(new_n23025), .B(new_n23011), .Y(new_n23026));
  xnor_4 g20678(.A(new_n23026), .B(new_n22905), .Y(n16062));
  xnor_4 g20679(.A(new_n22505), .B(new_n22498), .Y(n16068));
  xnor_4 g20680(.A(new_n22730), .B(new_n22727), .Y(n16080));
  and_5  g20681(.A(new_n22194), .B(new_n6356_1), .Y(new_n23030));
  nor_5  g20682(.A(new_n22198_1), .B(new_n22195), .Y(new_n23031));
  nor_5  g20683(.A(new_n23031), .B(new_n23030), .Y(new_n23032));
  nor_5  g20684(.A(new_n22189), .B(new_n11851), .Y(new_n23033));
  and_5  g20685(.A(new_n22193), .B(new_n22190), .Y(new_n23034));
  nor_5  g20686(.A(new_n23034), .B(new_n23033), .Y(new_n23035_1));
  xnor_4 g20687(.A(new_n23035_1), .B(new_n23032), .Y(n16098));
  xnor_4 g20688(.A(new_n17325), .B(new_n17317), .Y(n16110));
  xnor_4 g20689(.A(new_n14974), .B(new_n14945), .Y(n16142));
  xnor_4 g20690(.A(new_n16353), .B(new_n16341), .Y(n16185));
  xnor_4 g20691(.A(new_n12346_1), .B(new_n12329_1), .Y(n16196));
  xnor_4 g20692(.A(new_n20425), .B(new_n20424_1), .Y(n16206));
  xor_4  g20693(.A(new_n20497), .B(new_n20494), .Y(n16215));
  xnor_4 g20694(.A(new_n18688), .B(new_n18680), .Y(n16218));
  xnor_4 g20695(.A(new_n3913), .B(new_n3912), .Y(n16219));
  xnor_4 g20696(.A(new_n6950), .B(new_n6949), .Y(n16230));
  xor_4  g20697(.A(new_n8425), .B(new_n8417_1), .Y(n16243));
  xnor_4 g20698(.A(new_n17068_1), .B(new_n17059), .Y(n16275));
  xnor_4 g20699(.A(new_n10153), .B(new_n10152), .Y(n16279));
  nor_5  g20700(.A(new_n20014), .B(new_n17498), .Y(new_n23049));
  nor_5  g20701(.A(new_n20069_1), .B(new_n20015), .Y(new_n23050));
  or_5   g20702(.A(new_n23050), .B(new_n23049), .Y(n16322));
  xnor_4 g20703(.A(new_n17076), .B(new_n17036), .Y(n16327));
  xnor_4 g20704(.A(new_n20863), .B(new_n20856), .Y(n16350));
  xnor_4 g20705(.A(new_n6666), .B(new_n6665), .Y(n16367));
  xnor_4 g20706(.A(new_n18785), .B(new_n18784), .Y(n16379));
  xnor_4 g20707(.A(new_n19649), .B(new_n19632), .Y(n16398));
  xnor_4 g20708(.A(new_n13385), .B(new_n13383), .Y(n16406));
  xnor_4 g20709(.A(new_n21606), .B(new_n21589), .Y(n16407));
  xnor_4 g20710(.A(new_n23023), .B(new_n23014_1), .Y(n16419));
  xnor_4 g20711(.A(new_n8387), .B(new_n8347), .Y(n16424));
  xnor_4 g20712(.A(new_n13739), .B(new_n13673), .Y(new_n23061));
  xnor_4 g20713(.A(new_n23061), .B(new_n13779), .Y(n16428));
  xnor_4 g20714(.A(new_n11906), .B(new_n11849), .Y(n16433));
  xnor_4 g20715(.A(new_n11902), .B(new_n11857), .Y(n16440));
  xnor_4 g20716(.A(new_n17327), .B(new_n17313), .Y(n16445));
  xnor_4 g20717(.A(new_n13988), .B(new_n13936), .Y(n16460));
  xnor_4 g20718(.A(new_n19558), .B(new_n19549), .Y(n16481));
  nor_5  g20719(.A(new_n14586), .B(new_n11021), .Y(new_n23068_1));
  nor_5  g20720(.A(new_n14586), .B(new_n11028), .Y(new_n23069));
  nor_5  g20721(.A(new_n20129), .B(new_n20113), .Y(new_n23070));
  nor_5  g20722(.A(new_n23070), .B(new_n23069), .Y(new_n23071));
  xor_4  g20723(.A(new_n14586), .B(new_n11021), .Y(new_n23072));
  and_5  g20724(.A(new_n23072), .B(new_n23071), .Y(new_n23073));
  nor_5  g20725(.A(new_n23073), .B(new_n23068_1), .Y(n16493));
  xnor_4 g20726(.A(new_n4754), .B(new_n4728), .Y(n16506));
  xnor_4 g20727(.A(new_n12716), .B(new_n12715), .Y(n16516));
  xor_4  g20728(.A(new_n21698), .B(new_n21697), .Y(n16517));
  xnor_4 g20729(.A(new_n15444), .B(new_n15443), .Y(n16527));
  xnor_4 g20730(.A(new_n10753), .B(new_n9156), .Y(n16554));
  xnor_4 g20731(.A(new_n6130), .B(new_n5793), .Y(n16583));
  xnor_4 g20732(.A(new_n21156), .B(new_n10028), .Y(new_n23081));
  xnor_4 g20733(.A(new_n23081), .B(new_n21161), .Y(n16584));
  xnor_4 g20734(.A(new_n18854), .B(new_n18833), .Y(n16589));
  xor_4  g20735(.A(new_n19182), .B(new_n19180), .Y(n16596));
  xnor_4 g20736(.A(new_n21865), .B(new_n21828), .Y(n16617));
  xnor_4 g20737(.A(new_n7596), .B(new_n7567), .Y(n16630));
  xnor_4 g20738(.A(new_n21847), .B(new_n4940), .Y(n16640));
  xnor_4 g20739(.A(new_n2522), .B(new_n2521), .Y(n16656));
  xnor_4 g20740(.A(new_n6962), .B(new_n6915), .Y(n16674));
  xnor_4 g20741(.A(new_n13986), .B(new_n13940), .Y(n16682));
  xnor_4 g20742(.A(new_n21793), .B(new_n21774), .Y(n16684));
  xnor_4 g20743(.A(new_n10497), .B(new_n10493), .Y(n16688));
  xnor_4 g20744(.A(new_n6405), .B(new_n6397_1), .Y(n16733));
  xnor_4 g20745(.A(new_n7900), .B(new_n7898), .Y(n16798));
  xnor_4 g20746(.A(new_n16448), .B(new_n16447), .Y(n16834));
  xnor_4 g20747(.A(new_n3080), .B(new_n3041), .Y(n16837));
  xnor_4 g20748(.A(new_n21409), .B(new_n21406), .Y(n16841));
  xnor_4 g20749(.A(new_n5086), .B(new_n5085), .Y(n16885));
  xnor_4 g20750(.A(new_n8202), .B(new_n8137), .Y(n16905));
  nor_5  g20751(.A(new_n21331), .B(new_n21328), .Y(new_n23100));
  xnor_4 g20752(.A(new_n23100), .B(new_n17839), .Y(n16951));
  xor_4  g20753(.A(new_n15959), .B(new_n15950), .Y(n16954));
  xnor_4 g20754(.A(new_n8368), .B(new_n3704), .Y(n16989));
  xnor_4 g20755(.A(new_n18787), .B(new_n18757), .Y(n17006));
  xnor_4 g20756(.A(new_n13290), .B(new_n13289), .Y(n17068));
  xnor_4 g20757(.A(new_n14964), .B(new_n14963), .Y(n17070));
  xnor_4 g20758(.A(new_n20065), .B(new_n20021), .Y(n17075));
  xnor_4 g20759(.A(new_n16720), .B(new_n16702), .Y(n17084));
  xnor_4 g20760(.A(new_n4747_1), .B(new_n4746), .Y(n17104));
  xnor_4 g20761(.A(new_n13093), .B(new_n13070), .Y(n17106));
  xor_4  g20762(.A(new_n9691), .B(new_n9681), .Y(n17119));
  xnor_4 g20763(.A(new_n12987_1), .B(new_n12954), .Y(n17130));
  xnor_4 g20764(.A(new_n22323), .B(new_n22308), .Y(n17138));
  xnor_4 g20765(.A(new_n21700), .B(new_n21692), .Y(n17163));
  xor_4  g20766(.A(new_n19729), .B(new_n19728), .Y(n17168));
  xnor_4 g20767(.A(new_n11405), .B(new_n11397), .Y(n17202));
  xor_4  g20768(.A(new_n19005_1), .B(new_n19003), .Y(n17219));
  xnor_4 g20769(.A(new_n18276), .B(new_n18244), .Y(n17232));
  xnor_4 g20770(.A(new_n15072), .B(new_n15069), .Y(n17236));
  xor_4  g20771(.A(new_n10403), .B(new_n10402), .Y(n17243));
  xnor_4 g20772(.A(new_n11072), .B(new_n11056_1), .Y(n17263));
  nor_5  g20773(.A(new_n19162), .B(new_n19155), .Y(new_n23122));
  and_5  g20774(.A(new_n19186), .B(new_n19164_1), .Y(new_n23123));
  nor_5  g20775(.A(new_n23123), .B(new_n23122), .Y(n17285));
  xnor_4 g20776(.A(new_n11574), .B(new_n11546), .Y(n17320));
  xnor_4 g20777(.A(new_n2843), .B(new_n2795), .Y(n17337));
  xnor_4 g20778(.A(new_n21525_1), .B(new_n21517), .Y(n17344));
  xnor_4 g20779(.A(new_n21533), .B(new_n21502), .Y(n17359));
  xnor_4 g20780(.A(new_n13969), .B(new_n13143), .Y(n17387));
  xnor_4 g20781(.A(new_n5083), .B(new_n5081), .Y(n17391));
  xnor_4 g20782(.A(new_n18782_1), .B(new_n18762), .Y(n17392));
  xnor_4 g20783(.A(new_n21795), .B(new_n21771), .Y(n17421));
  xnor_4 g20784(.A(new_n12037), .B(new_n6571), .Y(n17432));
  xnor_4 g20785(.A(new_n20730), .B(new_n20712), .Y(n17436));
  xnor_4 g20786(.A(new_n22979), .B(new_n4710), .Y(n17440));
  xnor_4 g20787(.A(new_n8458), .B(new_n5794), .Y(n17450));
  nor_5  g20788(.A(new_n18553), .B(new_n7362), .Y(new_n23137));
  nor_5  g20789(.A(new_n7361), .B(new_n7322), .Y(new_n23138));
  nor_5  g20790(.A(new_n7362), .B(new_n7323), .Y(new_n23139));
  nor_5  g20791(.A(new_n7427), .B(new_n23139), .Y(new_n23140));
  nor_5  g20792(.A(new_n23140), .B(new_n23138), .Y(new_n23141));
  nor_5  g20793(.A(new_n23141), .B(new_n23137), .Y(new_n23142));
  nor_5  g20794(.A(new_n18552), .B(new_n7361), .Y(new_n23143));
  nor_5  g20795(.A(new_n23143), .B(new_n23140), .Y(new_n23144));
  nor_5  g20796(.A(new_n23144), .B(new_n23142), .Y(n17461));
  xor_4  g20797(.A(new_n22691), .B(new_n22690), .Y(n17466));
  xnor_4 g20798(.A(new_n13304), .B(new_n13265), .Y(n17493));
  xor_4  g20799(.A(new_n21200), .B(new_n21197), .Y(n17500));
  xnor_4 g20800(.A(new_n22054), .B(new_n22051), .Y(n17524));
  xnor_4 g20801(.A(new_n5757), .B(new_n5720), .Y(n17529));
  xnor_4 g20802(.A(new_n14770), .B(new_n10592), .Y(new_n23151));
  xnor_4 g20803(.A(new_n23151), .B(new_n14773), .Y(n17557));
  xnor_4 g20804(.A(new_n16361), .B(new_n16328), .Y(n17583));
  xnor_4 g20805(.A(new_n13978), .B(new_n13956), .Y(n17592));
  xnor_4 g20806(.A(new_n8375), .B(new_n8362), .Y(n17638));
  xnor_4 g20807(.A(new_n19560), .B(new_n19545), .Y(n17687));
  xnor_4 g20808(.A(new_n13592), .B(new_n13559), .Y(n17721));
  xnor_4 g20809(.A(new_n21380), .B(new_n21361), .Y(n17735));
  and_5  g20810(.A(new_n20803_1), .B(new_n10050), .Y(new_n23159));
  and_5  g20811(.A(new_n23159), .B(new_n20802), .Y(new_n23160_1));
  or_5   g20812(.A(new_n20803_1), .B(new_n10050), .Y(new_n23161));
  nor_5  g20813(.A(new_n23161), .B(new_n20802), .Y(new_n23162));
  nor_5  g20814(.A(new_n23162), .B(new_n23160_1), .Y(new_n23163));
  and_5  g20815(.A(new_n23163), .B(new_n20872), .Y(new_n23164));
  or_5   g20816(.A(new_n23163), .B(new_n20872), .Y(new_n23165));
  nor_5  g20817(.A(new_n20805), .B(new_n20794_1), .Y(new_n23166_1));
  nor_5  g20818(.A(new_n20815), .B(new_n20806), .Y(new_n23167));
  nor_5  g20819(.A(new_n23167), .B(new_n23166_1), .Y(new_n23168));
  and_5  g20820(.A(new_n23168), .B(new_n23165), .Y(new_n23169));
  or_5   g20821(.A(new_n23169), .B(new_n23160_1), .Y(new_n23170));
  nor_5  g20822(.A(new_n23170), .B(new_n23164), .Y(n17738));
  xor_4  g20823(.A(new_n15153), .B(new_n15150), .Y(n17746));
  xnor_4 g20824(.A(new_n22481), .B(new_n22478), .Y(n17749));
  xnor_4 g20825(.A(new_n18436), .B(new_n18417), .Y(n17820));
  xnor_4 g20826(.A(new_n13976), .B(new_n13961), .Y(n17855));
  and_5  g20827(.A(new_n13919), .B(new_n4897), .Y(new_n23176));
  and_5  g20828(.A(new_n4965), .B(new_n23176), .Y(new_n23177));
  not_8  g20829(.A(new_n21824), .Y(new_n23178));
  nor_5  g20830(.A(new_n4965), .B(new_n23178), .Y(new_n23179));
  nor_5  g20831(.A(new_n23179), .B(new_n23177), .Y(new_n23180));
  and_5  g20832(.A(new_n4966_1), .B(new_n4796), .Y(new_n23181));
  and_5  g20833(.A(new_n5028), .B(new_n4967_1), .Y(new_n23182));
  or_5   g20834(.A(new_n23182), .B(new_n23181), .Y(new_n23183));
  and_5  g20835(.A(new_n23183), .B(new_n23180), .Y(new_n23184));
  nor_5  g20836(.A(new_n23184), .B(new_n23177), .Y(n17877));
  xnor_4 g20837(.A(new_n15332_1), .B(new_n15331), .Y(n17889));
  and_5  g20838(.A(new_n22372), .B(new_n22362), .Y(new_n23187));
  nor_5  g20839(.A(new_n22384), .B(new_n23187), .Y(new_n23188));
  nor_5  g20840(.A(new_n22372), .B(new_n22362), .Y(new_n23189));
  nor_5  g20841(.A(new_n22383), .B(new_n23189), .Y(new_n23190));
  nor_5  g20842(.A(new_n23190), .B(new_n23188), .Y(n17912));
  xor_4  g20843(.A(new_n21786), .B(new_n21783), .Y(n17927));
  xnor_4 g20844(.A(new_n21857), .B(new_n21836), .Y(n17931));
  xnor_4 g20845(.A(new_n7892), .B(new_n7891), .Y(n17948));
  xor_4  g20846(.A(new_n15533), .B(new_n15530), .Y(n17956));
  nor_5  g20847(.A(new_n12667), .B(new_n12442), .Y(new_n23196));
  not_8  g20848(.A(new_n12592), .Y(new_n23197));
  nor_5  g20849(.A(new_n23197), .B(new_n12442), .Y(new_n23198));
  nor_5  g20850(.A(new_n12666), .B(new_n23198), .Y(new_n23199));
  nor_5  g20851(.A(new_n23199), .B(new_n23196), .Y(n17963));
  not_8  g20852(.A(new_n12948), .Y(new_n23201));
  nor_5  g20853(.A(n25494), .B(new_n21940), .Y(new_n23202));
  and_5  g20854(.A(new_n17308), .B(new_n17293), .Y(new_n23203));
  nor_5  g20855(.A(new_n23203), .B(new_n23202), .Y(new_n23204));
  and_5  g20856(.A(new_n23204), .B(new_n23201), .Y(new_n23205));
  nor_5  g20857(.A(new_n23204), .B(new_n12952), .Y(new_n23206));
  xnor_4 g20858(.A(new_n23204), .B(new_n12951), .Y(new_n23207));
  and_5  g20859(.A(new_n17309), .B(new_n12956_1), .Y(new_n23208));
  and_5  g20860(.A(new_n17329), .B(new_n17310), .Y(new_n23209));
  nor_5  g20861(.A(new_n23209), .B(new_n23208), .Y(new_n23210));
  and_5  g20862(.A(new_n23210), .B(new_n23207), .Y(new_n23211));
  nor_5  g20863(.A(new_n23211), .B(new_n23206), .Y(new_n23212));
  nor_5  g20864(.A(new_n23212), .B(new_n23205), .Y(new_n23213));
  nor_5  g20865(.A(new_n23204), .B(new_n23201), .Y(new_n23214));
  nor_5  g20866(.A(new_n23214), .B(new_n23211), .Y(new_n23215));
  nor_5  g20867(.A(new_n23215), .B(new_n23213), .Y(n17976));
  xnor_4 g20868(.A(new_n7170), .B(new_n7132), .Y(n17998));
  xnor_4 g20869(.A(new_n14391), .B(new_n2827), .Y(n18025));
  xnor_4 g20870(.A(new_n20381), .B(new_n20380), .Y(n18043));
  xnor_4 g20871(.A(new_n21714), .B(new_n21711), .Y(n18045));
  xnor_4 g20872(.A(new_n3918_1), .B(new_n3907), .Y(n18059));
  xnor_4 g20873(.A(new_n20063), .B(new_n20024), .Y(n18061));
  xnor_4 g20874(.A(new_n3391), .B(new_n3336), .Y(n18071));
  xnor_4 g20875(.A(new_n9982), .B(new_n9921), .Y(n18143));
  xnor_4 g20876(.A(new_n21202), .B(new_n21195), .Y(n18152));
  xnor_4 g20877(.A(new_n7588_1), .B(new_n7580), .Y(n18193));
  xnor_4 g20878(.A(new_n11615_1), .B(new_n13392), .Y(new_n23227));
  xnor_4 g20879(.A(new_n23227), .B(new_n11628), .Y(n18232));
  xnor_4 g20880(.A(new_n16722_1), .B(new_n16697), .Y(n18238));
  xnor_4 g20881(.A(new_n18265), .B(new_n18262), .Y(n18241));
  xnor_4 g20882(.A(new_n20726), .B(new_n20718), .Y(n18254));
  xnor_4 g20883(.A(new_n21378), .B(new_n21363), .Y(n18288));
  xnor_4 g20884(.A(new_n12104), .B(new_n12066), .Y(n18301));
  xnor_4 g20885(.A(new_n21702), .B(new_n21689), .Y(n18304));
  xnor_4 g20886(.A(new_n13308), .B(new_n13259), .Y(n18310));
  xnor_4 g20887(.A(new_n6669_1), .B(new_n6667), .Y(n18311));
  xnor_4 g20888(.A(new_n17452), .B(new_n17435), .Y(n18323));
  xnor_4 g20889(.A(new_n5447), .B(new_n5411), .Y(n18332));
  xor_4  g20890(.A(new_n21868), .B(new_n21867), .Y(n18343));
  xnor_4 g20891(.A(new_n19084), .B(new_n19081_1), .Y(n18350));
  xnor_4 g20892(.A(new_n17899), .B(new_n17898), .Y(n18362));
  xnor_4 g20893(.A(new_n5024_1), .B(new_n4975), .Y(n18377));
  xnor_4 g20894(.A(new_n4102), .B(new_n4082), .Y(n18405));
  xnor_4 g20895(.A(new_n16579), .B(new_n16569), .Y(n18414));
  xnor_4 g20896(.A(new_n14471_1), .B(new_n14462), .Y(n18418));
  xnor_4 g20897(.A(new_n8196), .B(new_n8152), .Y(n18437));
  xnor_4 g20898(.A(new_n19877), .B(new_n19837), .Y(n18439));
  xnor_4 g20899(.A(new_n11135), .B(new_n11134_1), .Y(n18445));
  xnor_4 g20900(.A(new_n6960), .B(new_n6920), .Y(n18467));
  xnor_4 g20901(.A(new_n18282), .B(new_n18229), .Y(n18482));
  xnor_4 g20902(.A(new_n18586), .B(new_n18565), .Y(n18509));
  xnor_4 g20903(.A(new_n13804), .B(new_n9039), .Y(n18513));
  xnor_4 g20904(.A(new_n14972), .B(new_n14970), .Y(n18515));
  xnor_4 g20905(.A(new_n15814), .B(new_n15795), .Y(n18572));
  and_5  g20906(.A(new_n23025), .B(new_n23011), .Y(new_n23255));
  nor_5  g20907(.A(new_n23255), .B(new_n22905), .Y(new_n23256));
  nor_5  g20908(.A(new_n23025), .B(new_n23011), .Y(new_n23257));
  nor_5  g20909(.A(new_n23257), .B(new_n22904), .Y(new_n23258));
  nor_5  g20910(.A(new_n23258), .B(new_n23256), .Y(n18574));
  xnor_4 g20911(.A(new_n20861), .B(new_n20858), .Y(n18576));
  xnor_4 g20912(.A(new_n22179), .B(new_n22171), .Y(n18582));
  xnor_4 g20913(.A(new_n19647), .B(new_n19635), .Y(n18583));
  xnor_4 g20914(.A(new_n20049), .B(new_n20048), .Y(n18610));
  xor_4  g20915(.A(new_n21728), .B(new_n21725), .Y(n18635));
  xnor_4 g20916(.A(new_n6740), .B(new_n6739), .Y(n18653));
  xnor_4 g20917(.A(new_n3721), .B(new_n3669), .Y(n18679));
  xnor_4 g20918(.A(new_n20175), .B(new_n20167), .Y(n18693));
  xnor_4 g20919(.A(new_n3078), .B(new_n3045), .Y(n18708));
  xnor_4 g20920(.A(new_n22517), .B(new_n22516), .Y(new_n23269));
  xnor_4 g20921(.A(new_n23269), .B(new_n22522), .Y(n18721));
  xnor_4 g20922(.A(new_n18442), .B(new_n18408), .Y(n18725));
  xnor_4 g20923(.A(new_n20530), .B(new_n20508), .Y(n18751));
  xnor_4 g20924(.A(new_n16355), .B(new_n16338), .Y(n18780));
  xnor_4 g20925(.A(new_n19303), .B(new_n19260), .Y(n18782));
  not_8  g20926(.A(new_n7547), .Y(new_n23275));
  and_5  g20927(.A(new_n23275), .B(new_n7469), .Y(new_n23276));
  nor_5  g20928(.A(new_n7606), .B(new_n23276), .Y(new_n23277));
  nor_5  g20929(.A(new_n23275), .B(new_n7469), .Y(new_n23278));
  nor_5  g20930(.A(new_n7605), .B(new_n23278), .Y(new_n23279));
  nor_5  g20931(.A(new_n23279), .B(new_n23277), .Y(n18802));
  xor_4  g20932(.A(new_n10860), .B(new_n10859), .Y(n18830));
  xor_4  g20933(.A(new_n12746_1), .B(new_n12741), .Y(n18831));
  xnor_4 g20934(.A(new_n11888), .B(new_n11881), .Y(n18843));
  xnor_4 g20935(.A(new_n3074), .B(new_n3056), .Y(n18858));
  xnor_4 g20936(.A(new_n9970), .B(new_n9950), .Y(n18859));
  xnor_4 g20937(.A(new_n17078), .B(new_n17029), .Y(n18864));
  xnor_4 g20938(.A(new_n4608), .B(new_n4541), .Y(n18865));
  xnor_4 g20939(.A(new_n21129), .B(new_n21128), .Y(n18886));
  xnor_4 g20940(.A(new_n16351), .B(new_n16350_1), .Y(n18887));
  xnor_4 g20941(.A(new_n8903), .B(new_n8866), .Y(n18919));
  xnor_4 g20942(.A(new_n12296), .B(new_n12284), .Y(n18940));
  xor_4  g20943(.A(new_n22641), .B(new_n22640), .Y(n18945));
  xnor_4 g20944(.A(new_n22353_1), .B(new_n22342), .Y(n18970));
  xnor_4 g20945(.A(new_n16776), .B(new_n12064), .Y(new_n23294));
  xnor_4 g20946(.A(new_n23294), .B(new_n16781), .Y(n18977));
  xnor_4 g20947(.A(new_n15074), .B(new_n15065), .Y(n18982));
  xor_4  g20948(.A(new_n20615), .B(new_n20614), .Y(n18999));
  xnor_4 g20949(.A(new_n5763), .B(new_n5708), .Y(n19044));
  xor_4  g20950(.A(new_n14775), .B(new_n14768), .Y(n19125));
  xnor_4 g20951(.A(new_n5761), .B(new_n5712), .Y(n19141));
  xnor_4 g20952(.A(new_n17185), .B(new_n13933), .Y(new_n23301));
  nor_5  g20953(.A(new_n17188), .B(new_n13938), .Y(new_n23302));
  xnor_4 g20954(.A(new_n17188), .B(new_n13938), .Y(new_n23303));
  nor_5  g20955(.A(new_n17193), .B(new_n13941), .Y(new_n23304_1));
  nor_5  g20956(.A(new_n18469), .B(new_n18454), .Y(new_n23305_1));
  nor_5  g20957(.A(new_n23305_1), .B(new_n23304_1), .Y(new_n23306));
  nor_5  g20958(.A(new_n23306), .B(new_n23303), .Y(new_n23307));
  nor_5  g20959(.A(new_n23307), .B(new_n23302), .Y(new_n23308));
  xnor_4 g20960(.A(new_n23308), .B(new_n23301), .Y(n19164));
  xnor_4 g20961(.A(new_n8383), .B(new_n8382), .Y(n19174));
  xnor_4 g20962(.A(new_n20780), .B(new_n20777), .Y(n19176));
  xnor_4 g20963(.A(new_n21704), .B(new_n21686), .Y(n19202));
  xnor_4 g20964(.A(new_n19968_1), .B(new_n19957), .Y(n19220));
  xor_4  g20965(.A(new_n7912), .B(new_n7850), .Y(n19221));
  xnor_4 g20966(.A(new_n11254), .B(new_n11253), .Y(n19223));
  xor_4  g20967(.A(new_n17064), .B(new_n17063), .Y(n19224));
  xnor_4 g20968(.A(new_n15478), .B(new_n15469), .Y(n19233));
  xnor_4 g20969(.A(new_n12730), .B(new_n12700), .Y(n19244));
  xnor_4 g20970(.A(new_n8905), .B(new_n8862_1), .Y(n19314));
  xnor_4 g20971(.A(new_n10763_1), .B(new_n10762), .Y(n19315));
  xnor_4 g20972(.A(new_n13300), .B(new_n13272), .Y(n19323));
  xnor_4 g20973(.A(new_n21523), .B(new_n21520), .Y(n19333));
  nor_5  g20974(.A(new_n17634), .B(new_n17177), .Y(new_n23323));
  nor_5  g20975(.A(new_n23323), .B(new_n9910), .Y(new_n23324));
  nor_5  g20976(.A(new_n17183), .B(new_n9914), .Y(new_n23325));
  nor_5  g20977(.A(new_n17204), .B(new_n17184), .Y(new_n23326));
  nor_5  g20978(.A(new_n23326), .B(new_n23325), .Y(new_n23327));
  not_8  g20979(.A(new_n23323), .Y(new_n23328));
  xnor_4 g20980(.A(new_n23328), .B(new_n9910), .Y(new_n23329));
  and_5  g20981(.A(new_n23329), .B(new_n23327), .Y(new_n23330));
  nor_5  g20982(.A(new_n23330), .B(new_n23324), .Y(n19348));
  xnor_4 g20983(.A(new_n16734), .B(new_n16670), .Y(n19354));
  xnor_4 g20984(.A(new_n11079), .B(new_n11045), .Y(n19367));
  xnor_4 g20985(.A(new_n18923), .B(new_n18902), .Y(n19385));
  xnor_4 g20986(.A(new_n16849), .B(new_n16797), .Y(new_n23335));
  xnor_4 g20987(.A(new_n23335), .B(new_n16878), .Y(n19389));
  xnor_4 g20988(.A(new_n16223_1), .B(new_n16193), .Y(n19401));
  xor_4  g20989(.A(new_n21967), .B(new_n21959), .Y(n19414));
  xnor_4 g20990(.A(new_n19103), .B(new_n17721_1), .Y(n19424));
  xnor_4 g20991(.A(new_n21133), .B(new_n21115), .Y(n19450));
  nor_5  g20992(.A(new_n23328), .B(new_n13870), .Y(new_n23341_1));
  xnor_4 g20993(.A(new_n23328), .B(new_n13870), .Y(new_n23342_1));
  nor_5  g20994(.A(new_n17183), .B(new_n13928), .Y(new_n23343));
  xnor_4 g20995(.A(new_n17183), .B(new_n13928), .Y(new_n23344));
  nor_5  g20996(.A(new_n17185), .B(new_n13933), .Y(new_n23345));
  nor_5  g20997(.A(new_n23308), .B(new_n23301), .Y(new_n23346));
  nor_5  g20998(.A(new_n23346), .B(new_n23345), .Y(new_n23347));
  nor_5  g20999(.A(new_n23347), .B(new_n23344), .Y(new_n23348));
  nor_5  g21000(.A(new_n23348), .B(new_n23343), .Y(new_n23349));
  nor_5  g21001(.A(new_n23349), .B(new_n23342_1), .Y(new_n23350));
  or_5   g21002(.A(new_n23350), .B(new_n23341_1), .Y(n19458));
  xnor_4 g21003(.A(new_n15155), .B(new_n15146_1), .Y(n19467));
  xnor_4 g21004(.A(new_n8198), .B(new_n8147), .Y(n19496));
  xor_4  g21005(.A(new_n15115), .B(new_n15107), .Y(n19523));
  xnor_4 g21006(.A(new_n4600), .B(new_n4561), .Y(n19570));
  xnor_4 g21007(.A(new_n12006), .B(new_n11996), .Y(n19602));
  xnor_4 g21008(.A(new_n12339), .B(new_n12334), .Y(n19617));
  xnor_4 g21009(.A(new_n13590), .B(new_n13562), .Y(n19623));
  xor_4  g21010(.A(new_n22008), .B(new_n22006), .Y(n19641));
  xnor_4 g21011(.A(new_n21797), .B(new_n21768), .Y(n19648));
  xnor_4 g21012(.A(new_n15812_1), .B(new_n15799), .Y(n19664));
  xnor_4 g21013(.A(new_n19726), .B(new_n19713), .Y(n19736));
  nor_5  g21014(.A(new_n21969), .B(new_n21955), .Y(new_n23363));
  nor_5  g21015(.A(new_n21955), .B(new_n3197), .Y(new_n23364));
  nor_5  g21016(.A(new_n21968), .B(new_n23364), .Y(new_n23365));
  nor_5  g21017(.A(new_n23365), .B(new_n23363), .Y(n19749));
  xnor_4 g21018(.A(new_n14840), .B(new_n14827_1), .Y(n19756));
  xnor_4 g21019(.A(new_n12004), .B(new_n12003_1), .Y(n19767));
  xor_4  g21020(.A(new_n3330), .B(new_n3327), .Y(new_n23369_1));
  xnor_4 g21021(.A(new_n23369_1), .B(new_n3393), .Y(n19780));
  xnor_4 g21022(.A(new_n22544), .B(new_n22541), .Y(n19792));
  xnor_4 g21023(.A(new_n20370), .B(new_n20357), .Y(n19798));
  xor_4  g21024(.A(new_n16445_1), .B(new_n16442), .Y(n19873));
  nor_5  g21025(.A(new_n18313), .B(new_n18294), .Y(new_n23374));
  not_8  g21026(.A(new_n18300), .Y(new_n23375));
  nor_5  g21027(.A(new_n23375), .B(new_n18294), .Y(new_n23376));
  nor_5  g21028(.A(new_n18312), .B(new_n23376), .Y(new_n23377));
  nor_5  g21029(.A(new_n23377), .B(new_n23374), .Y(n19909));
  xnor_4 g21030(.A(new_n19724), .B(new_n19716), .Y(n19916));
  xnor_4 g21031(.A(new_n20374), .B(new_n20350), .Y(n19923));
  xnor_4 g21032(.A(new_n18789), .B(new_n18754), .Y(n19930));
  xnor_4 g21033(.A(new_n6423), .B(new_n6317), .Y(n19968));
  xnor_4 g21034(.A(new_n19291), .B(new_n19279), .Y(n19988));
  and_5  g21035(.A(new_n21157_1), .B(new_n20438), .Y(new_n23384));
  nor_5  g21036(.A(new_n20438), .B(new_n10099), .Y(new_n23385));
  nor_5  g21037(.A(new_n20442), .B(new_n20439), .Y(new_n23386));
  nor_5  g21038(.A(new_n23386), .B(new_n23385), .Y(new_n23387));
  nor_5  g21039(.A(new_n23387), .B(new_n23384), .Y(new_n23388));
  nor_5  g21040(.A(new_n21157_1), .B(new_n20438), .Y(new_n23389));
  nor_5  g21041(.A(new_n23389), .B(new_n23386), .Y(new_n23390));
  nor_5  g21042(.A(new_n23390), .B(new_n23388), .Y(n20004));
  xnor_4 g21043(.A(new_n20526), .B(new_n20512), .Y(n20017));
  xnor_4 g21044(.A(new_n18278), .B(new_n18239), .Y(n20033));
  xnor_4 g21045(.A(new_n13771), .B(new_n13770), .Y(n20061));
  xnor_4 g21046(.A(new_n17851), .B(new_n17848), .Y(n20069));
  nor_5  g21047(.A(new_n14357), .B(new_n14346), .Y(new_n23396));
  nor_5  g21048(.A(new_n14413), .B(new_n14358), .Y(new_n23397));
  or_5   g21049(.A(new_n23397), .B(new_n23396), .Y(n20086));
  xnor_4 g21050(.A(new_n19178), .B(new_n19175), .Y(n20096));
  xnor_4 g21051(.A(new_n13292), .B(new_n13285_1), .Y(n20103));
  xnor_4 g21052(.A(new_n11576), .B(new_n11542), .Y(n20126));
  xnor_4 g21053(.A(new_n20931), .B(new_n20902), .Y(n20149));
  xnor_4 g21054(.A(new_n11900), .B(new_n11861), .Y(n20187));
  xnor_4 g21055(.A(new_n17289), .B(new_n17261), .Y(n20279));
  and_5  g21056(.A(new_n22164), .B(new_n22158), .Y(new_n23405));
  nor_5  g21057(.A(new_n22167), .B(new_n23405), .Y(new_n23406));
  nor_5  g21058(.A(new_n22182), .B(new_n22164), .Y(new_n23407));
  nor_5  g21059(.A(new_n22181), .B(new_n17427), .Y(new_n23408));
  nor_5  g21060(.A(new_n23408), .B(new_n23407), .Y(new_n23409));
  and_5  g21061(.A(new_n23409), .B(new_n23406), .Y(n20287));
  xnor_4 g21062(.A(new_n20210), .B(new_n20207), .Y(n20301));
  nor_5  g21063(.A(new_n8204), .B(new_n8133), .Y(new_n23412));
  nor_5  g21064(.A(new_n23412), .B(new_n8028), .Y(n20330));
  xnor_4 g21065(.A(new_n11896), .B(new_n11868), .Y(n20333));
  and_5  g21066(.A(new_n10346), .B(new_n10210), .Y(new_n23415));
  and_5  g21067(.A(new_n10410), .B(new_n23415), .Y(new_n23416));
  or_5   g21068(.A(new_n10346), .B(new_n10210), .Y(new_n23417));
  nor_5  g21069(.A(new_n10410), .B(new_n23417), .Y(new_n23418));
  or_5   g21070(.A(new_n23418), .B(new_n23416), .Y(n20355));
  xnor_4 g21071(.A(new_n8418), .B(new_n5201), .Y(n20366));
  xnor_4 g21072(.A(new_n18956), .B(new_n18953), .Y(n20388));
  xnor_4 g21073(.A(new_n21855), .B(new_n21838), .Y(n20402));
  xnor_4 g21074(.A(new_n15319), .B(new_n15293), .Y(n20403));
  xnor_4 g21075(.A(new_n22404), .B(new_n3062), .Y(n20424));
  xnor_4 g21076(.A(new_n20053), .B(new_n20042), .Y(n20436));
  xor_4  g21077(.A(new_n8184), .B(new_n8182), .Y(n20441));
  xnor_4 g21078(.A(new_n7604), .B(new_n7552), .Y(n20445));
  xnor_4 g21079(.A(new_n5026_1), .B(new_n4971), .Y(n20450));
  xnor_4 g21080(.A(new_n16367_1), .B(new_n16365), .Y(n20490));
  xor_4  g21081(.A(new_n19966), .B(new_n19962), .Y(n20495));
  and_5  g21082(.A(new_n15337), .B(new_n15335), .Y(new_n23431));
  and_5  g21083(.A(new_n23431), .B(new_n15334), .Y(new_n23432));
  or_5   g21084(.A(new_n15337), .B(new_n15335), .Y(new_n23433_1));
  nor_5  g21085(.A(new_n23433_1), .B(new_n15334), .Y(new_n23434_1));
  or_5   g21086(.A(new_n23434_1), .B(new_n23432), .Y(n20515));
  nor_5  g21087(.A(new_n22546), .B(new_n22536), .Y(new_n23436));
  nor_5  g21088(.A(new_n23436), .B(new_n22531), .Y(n20533));
  xnor_4 g21089(.A(new_n17723), .B(new_n17716), .Y(n20582));
  xnor_4 g21090(.A(new_n19451), .B(new_n19423), .Y(n20590));
  xnor_4 g21091(.A(new_n3375), .B(new_n3373), .Y(n20602));
  xnor_4 g21092(.A(new_n16348), .B(new_n16347), .Y(n20609));
  xnor_4 g21093(.A(new_n6575), .B(new_n6567_1), .Y(n20623));
  xnor_4 g21094(.A(new_n20385_1), .B(new_n20336), .Y(n20629));
  xnor_4 g21095(.A(new_n13768), .B(new_n13759), .Y(n20661));
  xnor_4 g21096(.A(new_n8463), .B(new_n8461), .Y(n20673));
  xnor_4 g21097(.A(new_n20378), .B(new_n20344), .Y(n20678));
  nor_5  g21098(.A(new_n14816), .B(new_n11793), .Y(new_n23447));
  nor_5  g21099(.A(new_n14847), .B(new_n23447), .Y(new_n23448));
  and_5  g21100(.A(new_n14816), .B(new_n11793), .Y(new_n23449));
  or_5   g21101(.A(new_n23449), .B(new_n14813), .Y(new_n23450_1));
  nor_5  g21102(.A(new_n23450_1), .B(new_n23448), .Y(n20680));
  xnor_4 g21103(.A(new_n6401), .B(new_n4157), .Y(n20685));
  xnor_4 g21104(.A(new_n23204), .B(new_n12948), .Y(new_n23453));
  xnor_4 g21105(.A(new_n23453), .B(new_n23212), .Y(n20691));
  xnor_4 g21106(.A(new_n15810), .B(new_n15802), .Y(n20696));
  xnor_4 g21107(.A(new_n22321), .B(new_n22311_1), .Y(n20704));
  xor_4  g21108(.A(new_n21372), .B(new_n21371), .Y(n20705));
  xnor_4 g21109(.A(new_n9980), .B(new_n9926_1), .Y(n20709));
  xnor_4 g21110(.A(new_n14732), .B(new_n14708), .Y(n20713));
  xnor_4 g21111(.A(new_n8634), .B(new_n8633), .Y(n20722));
  not_8  g21112(.A(new_n19347), .Y(new_n23461));
  nor_5  g21113(.A(new_n22817), .B(new_n23461), .Y(new_n23462));
  nor_5  g21114(.A(new_n19347), .B(new_n19336), .Y(new_n23463_1));
  nor_5  g21115(.A(new_n23461), .B(new_n19335), .Y(new_n23464));
  nor_5  g21116(.A(new_n19359), .B(new_n23464), .Y(new_n23465));
  nor_5  g21117(.A(new_n23465), .B(new_n23463_1), .Y(new_n23466));
  nor_5  g21118(.A(new_n23466), .B(new_n23462), .Y(new_n23467));
  nor_5  g21119(.A(new_n22818), .B(new_n19347), .Y(new_n23468));
  nor_5  g21120(.A(new_n23468), .B(new_n23465), .Y(new_n23469));
  nor_5  g21121(.A(new_n23469), .B(new_n23467), .Y(n20723));
  xnor_4 g21122(.A(new_n22159), .B(new_n17428), .Y(new_n23471_1));
  xnor_4 g21123(.A(new_n23471_1), .B(new_n22182), .Y(n20748));
  xor_4  g21124(.A(new_n5439_1), .B(new_n5429), .Y(n20761));
  xnor_4 g21125(.A(new_n20061_1), .B(new_n20028), .Y(n20774));
  xnor_4 g21126(.A(new_n23349), .B(new_n23342_1), .Y(n20788));
  nor_5  g21127(.A(new_n22669), .B(new_n21722), .Y(new_n23476));
  nor_5  g21128(.A(new_n23476), .B(new_n22779_1), .Y(new_n23477));
  nor_5  g21129(.A(new_n22775), .B(new_n21723), .Y(new_n23478));
  nor_5  g21130(.A(new_n23478), .B(new_n22778), .Y(new_n23479));
  nor_5  g21131(.A(new_n23479), .B(new_n23477), .Y(n20795));
  xnor_4 g21132(.A(new_n20093), .B(new_n20082), .Y(new_n23481));
  and_5  g21133(.A(new_n20102), .B(new_n20082), .Y(new_n23482));
  nor_5  g21134(.A(new_n23482), .B(new_n20104), .Y(new_n23483));
  nor_5  g21135(.A(new_n23483), .B(new_n20103_1), .Y(new_n23484));
  xnor_4 g21136(.A(new_n23484), .B(new_n23481), .Y(n20803));
  xor_4  g21137(.A(new_n23183), .B(new_n23180), .Y(n20869));
  xnor_4 g21138(.A(new_n22483), .B(new_n22475), .Y(n20879));
  xnor_4 g21139(.A(new_n6411), .B(new_n6384), .Y(n20915));
  xnor_4 g21140(.A(n19282), .B(n2160), .Y(new_n23489));
  nor_5  g21141(.A(n12657), .B(new_n11674_1), .Y(new_n23490));
  and_5  g21142(.A(new_n21388), .B(new_n21385), .Y(new_n23491));
  or_5   g21143(.A(new_n23491), .B(new_n23490), .Y(new_n23492));
  xor_4  g21144(.A(new_n23492), .B(new_n23489), .Y(new_n23493_1));
  nor_5  g21145(.A(new_n23493_1), .B(new_n22379_1), .Y(new_n23494));
  nor_5  g21146(.A(new_n21389), .B(new_n19678), .Y(new_n23495));
  nor_5  g21147(.A(new_n21393), .B(new_n21390), .Y(new_n23496));
  nor_5  g21148(.A(new_n23496), .B(new_n23495), .Y(new_n23497));
  xnor_4 g21149(.A(new_n23493_1), .B(new_n22379_1), .Y(new_n23498));
  nor_5  g21150(.A(new_n23498), .B(new_n23497), .Y(new_n23499));
  nor_5  g21151(.A(new_n23499), .B(new_n23494), .Y(new_n23500));
  not_8  g21152(.A(new_n23500), .Y(new_n23501));
  nor_5  g21153(.A(n19282), .B(new_n12808), .Y(new_n23502));
  and_5  g21154(.A(new_n23492), .B(new_n23489), .Y(new_n23503));
  nor_5  g21155(.A(new_n23503), .B(new_n23502), .Y(new_n23504));
  and_5  g21156(.A(new_n23504), .B(new_n22377), .Y(new_n23505));
  and_5  g21157(.A(new_n23505), .B(new_n23501), .Y(new_n23506));
  and_5  g21158(.A(new_n23506), .B(new_n22372), .Y(new_n23507));
  or_5   g21159(.A(new_n23504), .B(new_n22377), .Y(new_n23508));
  nor_5  g21160(.A(new_n23508), .B(new_n23501), .Y(new_n23509));
  and_5  g21161(.A(new_n23509), .B(new_n22373), .Y(new_n23510));
  or_5   g21162(.A(new_n23510), .B(new_n23507), .Y(n20935));
  xnor_4 g21163(.A(new_n21791), .B(new_n21777), .Y(n20936));
  xnor_4 g21164(.A(new_n16763), .B(new_n16762), .Y(n21008));
  xnor_4 g21165(.A(new_n19301), .B(new_n19263), .Y(n21017));
  and_5  g21166(.A(new_n22883), .B(new_n21226_1), .Y(new_n23515));
  nor_5  g21167(.A(new_n22883), .B(new_n21226_1), .Y(new_n23516));
  nor_5  g21168(.A(new_n22888), .B(new_n23516), .Y(new_n23517));
  or_5   g21169(.A(new_n23517), .B(new_n22882), .Y(new_n23518));
  nor_5  g21170(.A(new_n23518), .B(new_n23515), .Y(n21034));
  xor_4  g21171(.A(new_n21932), .B(new_n21931), .Y(n21046));
  xnor_4 g21172(.A(new_n8564), .B(new_n8545), .Y(n21062));
  xor_4  g21173(.A(new_n22624), .B(new_n22616), .Y(new_n23522));
  xnor_4 g21174(.A(new_n23522), .B(new_n22531), .Y(n21093));
  xnor_4 g21175(.A(new_n9725), .B(new_n7884_1), .Y(n21094));
  xnor_4 g21176(.A(new_n14622), .B(new_n14599), .Y(n21123));
  xnor_4 g21177(.A(new_n18686), .B(new_n17923), .Y(n21154));
  xnor_4 g21178(.A(new_n15453), .B(new_n15431), .Y(n21157));
  xnor_4 g21179(.A(new_n20923_1), .B(new_n20915_1), .Y(n21168));
  xnor_4 g21180(.A(new_n7400), .B(new_n7398), .Y(n21173));
  xnor_4 g21181(.A(new_n4596), .B(new_n4571), .Y(n21176));
  xnor_4 g21182(.A(new_n14279), .B(new_n14272), .Y(n21182));
  nor_5  g21183(.A(new_n21762), .B(new_n20949), .Y(new_n23532));
  nor_5  g21184(.A(new_n21800_1), .B(new_n20950), .Y(new_n23533));
  nor_5  g21185(.A(new_n23533), .B(new_n23532), .Y(new_n23534));
  nor_5  g21186(.A(new_n21799), .B(new_n20960), .Y(new_n23535));
  nor_5  g21187(.A(new_n23535), .B(new_n21765_1), .Y(new_n23536));
  and_5  g21188(.A(new_n23536), .B(new_n23534), .Y(n21193));
  xnor_4 g21189(.A(new_n9469), .B(new_n9468), .Y(n21203));
  xnor_4 g21190(.A(new_n16346), .B(new_n2544), .Y(n21225));
  xnor_4 g21191(.A(new_n19661), .B(new_n19614), .Y(n21238));
  xnor_4 g21192(.A(new_n13773), .B(new_n13754_1), .Y(n21254));
  xnor_4 g21193(.A(new_n19873_1), .B(new_n19845), .Y(n21298));
  xnor_4 g21194(.A(new_n19641_1), .B(new_n9376), .Y(n21302));
  xnor_4 g21195(.A(new_n19722), .B(new_n19719), .Y(n21349));
  xnor_4 g21196(.A(new_n15962), .B(new_n15961), .Y(n21365));
  xnor_4 g21197(.A(new_n15117), .B(new_n15104), .Y(n21367));
  xnor_4 g21198(.A(new_n11783), .B(new_n11755), .Y(n21396));
  xnor_4 g21199(.A(new_n7602), .B(new_n7556), .Y(n21399));
  xnor_4 g21200(.A(new_n3401), .B(new_n3396), .Y(n21404));
  xnor_4 g21201(.A(new_n8465), .B(new_n8454), .Y(n21446));
  xnor_4 g21202(.A(new_n11626), .B(new_n11618), .Y(n21472));
  xnor_4 g21203(.A(new_n7421_1), .B(new_n7375), .Y(n21525));
  xnor_4 g21204(.A(new_n17126), .B(new_n17102), .Y(n21549));
  xnor_4 g21205(.A(new_n19556), .B(new_n19553), .Y(n21615));
  nor_5  g21206(.A(new_n22164), .B(new_n7835), .Y(new_n23555));
  xnor_4 g21207(.A(new_n22164), .B(new_n13394), .Y(new_n23556));
  nor_5  g21208(.A(new_n17427), .B(new_n13394), .Y(new_n23557));
  and_5  g21209(.A(new_n17457), .B(new_n17429), .Y(new_n23558));
  or_5   g21210(.A(new_n23558), .B(new_n23557), .Y(new_n23559));
  and_5  g21211(.A(new_n23559), .B(new_n23556), .Y(new_n23560));
  nor_5  g21212(.A(new_n23560), .B(new_n23555), .Y(n21628));
  nor_5  g21213(.A(new_n21433), .B(new_n20955), .Y(new_n23562));
  xnor_4 g21214(.A(new_n21433), .B(new_n20957), .Y(new_n23563));
  nor_5  g21215(.A(new_n21437), .B(new_n20957), .Y(new_n23564));
  nor_5  g21216(.A(new_n22745), .B(new_n22742), .Y(new_n23565));
  or_5   g21217(.A(new_n23565), .B(new_n23564), .Y(new_n23566));
  and_5  g21218(.A(new_n23566), .B(new_n23563), .Y(new_n23567));
  nor_5  g21219(.A(new_n23567), .B(new_n23562), .Y(n21637));
  xnor_4 g21220(.A(new_n21374), .B(new_n21367_1), .Y(n21645));
  xnor_4 g21221(.A(new_n12032), .B(new_n22664), .Y(n21665));
  xnor_4 g21222(.A(new_n14844), .B(new_n14821), .Y(n21680));
  xnor_4 g21223(.A(new_n21863), .B(new_n21830), .Y(n21685));
  xnor_4 g21224(.A(new_n18438), .B(new_n18414_1), .Y(n21717));
  xnor_4 g21225(.A(new_n16751), .B(new_n16746), .Y(n21719));
  xnor_4 g21226(.A(new_n18430), .B(new_n18427), .Y(n21750));
  xnor_4 g21227(.A(new_n21626), .B(new_n21625), .Y(n21765));
  xnor_4 g21228(.A(new_n23498), .B(new_n23497), .Y(n21800));
  xnor_4 g21229(.A(new_n4299), .B(new_n4296), .Y(new_n23578));
  xnor_4 g21230(.A(new_n23578), .B(new_n4304), .Y(n21820));
  xnor_4 g21231(.A(new_n19295), .B(new_n19273), .Y(n21874));
  xnor_4 g21232(.A(new_n13294), .B(new_n13282), .Y(n21943));
  xnor_4 g21233(.A(new_n15966), .B(new_n15945), .Y(n21960));
  xnor_4 g21234(.A(new_n7159), .B(new_n7157), .Y(n21976));
  xnor_4 g21235(.A(new_n11263), .B(new_n11235), .Y(n21986));
  xnor_4 g21236(.A(new_n11081), .B(new_n11041), .Y(n22016));
  xnor_4 g21237(.A(new_n18432), .B(new_n18423), .Y(n22027));
  xnor_4 g21238(.A(new_n13089), .B(new_n13080), .Y(n22050));
  xnor_4 g21239(.A(new_n4158), .B(new_n4157), .Y(n22063));
  xnor_4 g21240(.A(new_n20921), .B(new_n20918), .Y(n22076));
  nor_5  g21241(.A(new_n20086_1), .B(new_n13736), .Y(new_n23590));
  and_5  g21242(.A(new_n20433), .B(new_n20414), .Y(new_n23591));
  nor_5  g21243(.A(new_n23591), .B(new_n23590), .Y(n22090));
  xnor_4 g21244(.A(new_n22351), .B(new_n22344), .Y(n22107));
  xnor_4 g21245(.A(new_n17619), .B(new_n17593), .Y(n22113));
  nor_5  g21246(.A(new_n13735), .B(new_n13673), .Y(new_n23595));
  nor_5  g21247(.A(new_n13781_1), .B(new_n23595), .Y(new_n23596));
  nor_5  g21248(.A(new_n13736), .B(new_n13674), .Y(new_n23597));
  nor_5  g21249(.A(new_n13780), .B(new_n23597), .Y(new_n23598));
  nor_5  g21250(.A(new_n23598), .B(new_n23596), .Y(n22124));
  nor_5  g21251(.A(new_n22984), .B(new_n19162), .Y(new_n23600));
  and_5  g21252(.A(new_n22988), .B(new_n22985), .Y(new_n23601));
  nor_5  g21253(.A(new_n23601), .B(new_n23600), .Y(n22126));
  nor_5  g21254(.A(new_n23509), .B(new_n23506), .Y(new_n23603));
  xnor_4 g21255(.A(new_n23603), .B(new_n22373), .Y(n22130));
  xor_4  g21256(.A(new_n17799), .B(new_n17798), .Y(n22144));
  xnor_4 g21257(.A(new_n22736), .B(new_n22732), .Y(n22150));
  xnor_4 g21258(.A(new_n19490), .B(new_n19484), .Y(n22157));
  xnor_4 g21259(.A(new_n23306), .B(new_n23303), .Y(n22213));
  xnor_4 g21260(.A(new_n10389), .B(new_n10388_1), .Y(n22283));
  xor_4  g21261(.A(new_n20123), .B(new_n20122), .Y(n22311));
  xnor_4 g21262(.A(new_n8907), .B(new_n8858), .Y(n22317));
  xnor_4 g21263(.A(new_n17384), .B(new_n17371), .Y(n22341));
  nor_5  g21264(.A(new_n7194), .B(new_n7182), .Y(new_n23613));
  and_5  g21265(.A(new_n23613), .B(new_n7178), .Y(new_n23614));
  nand_5 g21266(.A(new_n7194), .B(new_n7182), .Y(new_n23615));
  nor_5  g21267(.A(new_n23615), .B(new_n7178), .Y(new_n23616));
  nor_5  g21268(.A(new_n23616), .B(new_n23614), .Y(new_n23617));
  xnor_4 g21269(.A(new_n23617), .B(new_n18081), .Y(n22353));
  xnor_4 g21270(.A(new_n17382), .B(new_n17374), .Y(n22444));
  xnor_4 g21271(.A(new_n10143), .B(new_n10141), .Y(n22467));
  xnor_4 g21272(.A(new_n20132), .B(new_n8885), .Y(n22484));
  xnor_4 g21273(.A(new_n4606), .B(new_n4546), .Y(n22489));
  xnor_4 g21274(.A(new_n8389), .B(new_n8344), .Y(n22494));
  xnor_4 g21275(.A(new_n10395), .B(new_n10373), .Y(n22533));
  xnor_4 g21276(.A(new_n22319), .B(new_n22317_1), .Y(n22584));
  nor_5  g21277(.A(new_n17805), .B(new_n17783), .Y(new_n23626));
  nor_5  g21278(.A(new_n23626), .B(new_n17744), .Y(n22589));
  xnor_4 g21279(.A(new_n23347), .B(new_n23344), .Y(n22620));
  xnor_4 g21280(.A(new_n8460), .B(new_n8459), .Y(n22623));
  xnor_4 g21281(.A(new_n16874), .B(new_n16860), .Y(n22697));
  xnor_4 g21282(.A(new_n8897), .B(new_n8879), .Y(n22714));
  xnor_4 g21283(.A(new_n11904), .B(new_n11854), .Y(n22761));
  xnor_4 g21284(.A(new_n18852), .B(new_n18836), .Y(n22779));
  xnor_4 g21285(.A(new_n22329), .B(new_n22299), .Y(n22787));
  xnor_4 g21286(.A(new_n2538), .B(new_n2506), .Y(n22819));
  xnor_4 g21287(.A(new_n9203), .B(new_n4586), .Y(n22858));
  xnor_4 g21288(.A(new_n20987), .B(new_n11592), .Y(new_n23637_1));
  xnor_4 g21289(.A(new_n23637_1), .B(new_n22797), .Y(n22870));
  xor_4  g21290(.A(new_n9693), .B(new_n9676), .Y(n22891));
  xor_4  g21291(.A(new_n19444), .B(new_n19431), .Y(n22897));
  xnor_4 g21292(.A(new_n10161), .B(new_n10104), .Y(n22903));
  xnor_4 g21293(.A(new_n14293), .B(new_n14251), .Y(n22907));
  xnor_4 g21294(.A(new_n7164), .B(new_n7163), .Y(n22910));
  xnor_4 g21295(.A(new_n12321), .B(new_n12315_1), .Y(n22914));
  xnor_4 g21296(.A(new_n5769), .B(new_n5853), .Y(n22939));
  xnor_4 g21297(.A(new_n18961), .B(new_n4417), .Y(new_n23646));
  xnor_4 g21298(.A(new_n23646), .B(new_n18959), .Y(n22998));
  xnor_4 g21299(.A(new_n8893), .B(new_n8892), .Y(n23006));
  xnor_4 g21300(.A(new_n12748), .B(new_n12739), .Y(n23007));
  xnor_4 g21301(.A(new_n17990), .B(new_n17987), .Y(n23009));
  xnor_4 g21302(.A(new_n16732), .B(new_n16675), .Y(n23014));
  xor_4  g21303(.A(new_n23566), .B(new_n23563), .Y(n23047));
  xnor_4 g21304(.A(new_n17450_1), .B(new_n17438), .Y(n23058));
  and_5  g21305(.A(new_n18451), .B(new_n18446), .Y(n23066));
  and_5  g21306(.A(new_n18339), .B(new_n10209), .Y(new_n23655));
  nor_5  g21307(.A(new_n23655), .B(new_n18341), .Y(new_n23656));
  xor_4  g21308(.A(new_n23656), .B(new_n18336), .Y(n23067));
  xor_4  g21309(.A(new_n15957), .B(new_n15952), .Y(n23238));
  xnor_4 g21310(.A(new_n17202_1), .B(new_n17187), .Y(n23247));
  xor_4  g21311(.A(new_n14966), .B(new_n14958), .Y(n23248));
  xnor_4 g21312(.A(new_n17281), .B(new_n17270), .Y(n23270));
  xnor_4 g21313(.A(new_n22382), .B(new_n22378), .Y(n23289));
  xnor_4 g21314(.A(new_n5449), .B(new_n5406), .Y(n23305));
  xnor_4 g21315(.A(new_n20724), .B(new_n20721), .Y(n23341));
  xnor_4 g21316(.A(new_n9376), .B(new_n4943), .Y(n23342));
  and_5  g21317(.A(new_n21028), .B(new_n23275), .Y(new_n23666));
  nor_5  g21318(.A(new_n21052), .B(new_n23666), .Y(new_n23667));
  nor_5  g21319(.A(new_n21028), .B(new_n23275), .Y(new_n23668));
  nor_5  g21320(.A(new_n21051), .B(new_n23668), .Y(new_n23669_1));
  nor_5  g21321(.A(new_n23669_1), .B(new_n23667), .Y(n23355));
  xnor_4 g21322(.A(new_n19055), .B(new_n19052), .Y(n23371));
  xnor_4 g21323(.A(new_n15323), .B(new_n15284), .Y(n23401));
  xnor_4 g21324(.A(new_n13087), .B(new_n13086), .Y(n23414));
  xnor_4 g21325(.A(new_n17287), .B(new_n17264), .Y(n23429));
  nor_5  g21326(.A(new_n21280), .B(new_n21274), .Y(new_n23675));
  not_8  g21327(.A(new_n21276_1), .Y(new_n23676));
  nor_5  g21328(.A(new_n23676), .B(new_n21274), .Y(new_n23677));
  nor_5  g21329(.A(new_n23677), .B(new_n21279), .Y(new_n23678));
  nor_5  g21330(.A(new_n23678), .B(new_n23675), .Y(n23433));
  xnor_4 g21331(.A(new_n18270), .B(new_n18256), .Y(n23434));
  nor_5  g21332(.A(new_n22984), .B(new_n21402), .Y(new_n23681));
  nor_5  g21333(.A(new_n23681), .B(new_n23001), .Y(new_n23682));
  nor_5  g21334(.A(new_n22983), .B(new_n21401), .Y(new_n23683));
  nor_5  g21335(.A(new_n23683), .B(new_n23000), .Y(new_n23684_1));
  nor_5  g21336(.A(new_n23684_1), .B(new_n23682), .Y(n23450));
  xnor_4 g21337(.A(new_n16730), .B(new_n16679), .Y(n23471));
  xnor_4 g21338(.A(new_n20734), .B(new_n20706), .Y(n23480));
  xor_4  g21339(.A(new_n17651), .B(new_n17646), .Y(n23546));
  xnor_4 g21340(.A(new_n20368), .B(new_n20360), .Y(n23550));
  xnor_4 g21341(.A(new_n7415), .B(new_n7387), .Y(n23585));
  xor_4  g21342(.A(new_n19442), .B(new_n19434), .Y(n23588));
  xor_4  g21343(.A(new_n20612), .B(new_n20611), .Y(n23619));
  xnor_4 g21344(.A(new_n3072), .B(new_n3061), .Y(n23624));
  xnor_4 g21345(.A(new_n11775_1), .B(new_n11768), .Y(n23628));
  xnor_4 g21346(.A(new_n21527), .B(new_n21514), .Y(n23637));
  xnor_4 g21347(.A(new_n22113_1), .B(new_n22110), .Y(n23663));
  xnor_4 g21348(.A(new_n11777), .B(new_n11764), .Y(n23669));
  xnor_4 g21349(.A(new_n12985_1), .B(new_n12958), .Y(n23684));
  xnor_4 g21350(.A(new_n18777), .B(new_n18768), .Y(n23690));
  xnor_4 g21351(.A(new_n21861), .B(new_n21832_1), .Y(n23714));
  nor_5  g21352(.A(new_n23035_1), .B(new_n23032), .Y(n23719));
  xnor_4 g21353(.A(new_n21001), .B(new_n20998), .Y(n23748));
  xnor_4 g21354(.A(new_n10855), .B(new_n7198), .Y(n23856));
  xnor_4 g21355(.A(new_n7413), .B(new_n7412), .Y(n23883));
  xnor_4 g21356(.A(new_n14273), .B(new_n5809), .Y(new_n23705));
  xnor_4 g21357(.A(new_n23705), .B(new_n14276), .Y(n23888));
  xnor_4 g21358(.A(new_n3381), .B(new_n3356), .Y(n23899));
  xnor_4 g21359(.A(new_n14772_1), .B(new_n9461), .Y(n23903));
  xnor_4 g21360(.A(new_n12728), .B(new_n12702_1), .Y(n23924));
  xnor_4 g21361(.A(new_n16410), .B(new_n16409), .Y(n23935));
  xnor_4 g21362(.A(new_n12981), .B(new_n12966), .Y(n23942));
  xnor_4 g21363(.A(new_n17483), .B(new_n17475), .Y(n23954));
  xnor_4 g21364(.A(new_n18516), .B(new_n18496_1), .Y(n23958));
  xor_4  g21365(.A(new_n21992), .B(new_n21991), .Y(n23986));
  xor_4  g21366(.A(new_n16765), .B(new_n16760), .Y(n24002));
  xnor_4 g21367(.A(new_n12876), .B(new_n12868), .Y(n24039));
  xnor_4 g21368(.A(new_n22967), .B(new_n22966), .Y(n24052));
  xnor_4 g21369(.A(new_n20055), .B(new_n20038), .Y(n24092));
  xnor_4 g21370(.A(new_n15449), .B(new_n15448), .Y(n24096));
  xnor_4 g21371(.A(new_n12097), .B(new_n12072_1), .Y(n24097));
  xnor_4 g21372(.A(new_n11781), .B(new_n11758), .Y(n24105));
  xnor_4 g21373(.A(new_n17972), .B(new_n17954_1), .Y(n24119));
  xnor_4 g21374(.A(new_n14842), .B(new_n14824), .Y(n24133));
  xnor_4 g21375(.A(new_n19653), .B(new_n19626), .Y(n24141));
  xnor_4 g21376(.A(new_n20897), .B(new_n20873), .Y(new_n23725));
  xnor_4 g21377(.A(new_n23725), .B(new_n20933), .Y(n24145));
  xnor_4 g21378(.A(new_n21602), .B(new_n21599_1), .Y(n24146));
  xnor_4 g21379(.A(new_n12661), .B(new_n12609), .Y(n24155));
  xnor_4 g21380(.A(new_n23210), .B(new_n23207), .Y(n24160));
  xnor_4 g21381(.A(new_n9217_1), .B(new_n9185), .Y(n24167));
  and_5  g21382(.A(new_n20183), .B(new_n20178), .Y(n24172));
  xnor_4 g21383(.A(new_n14281), .B(new_n14269), .Y(n24177));
  xor_4  g21384(.A(new_n23072), .B(new_n23071), .Y(n24228));
  xnor_4 g21385(.A(new_n17386), .B(new_n17368), .Y(n24258));
  nor_5  g21386(.A(new_n18081), .B(new_n7182), .Y(new_n23735));
  and_5  g21387(.A(new_n23616), .B(new_n18083), .Y(new_n23736));
  nor_5  g21388(.A(new_n23736), .B(new_n23614), .Y(new_n23737));
  nor_5  g21389(.A(new_n23737), .B(new_n23735), .Y(n24260));
  xnor_4 g21390(.A(new_n18856), .B(new_n18830_1), .Y(n24289));
  xnor_4 g21391(.A(new_n4749), .B(new_n4738), .Y(n24297));
  xnor_4 g21392(.A(new_n11773), .B(new_n3909_1), .Y(n24307));
  xnor_4 g21393(.A(new_n2532), .B(new_n2520), .Y(n24342));
  xnor_4 g21394(.A(new_n15964), .B(new_n15947_1), .Y(n24345));
  xnor_4 g21395(.A(new_n9471), .B(new_n9459_1), .Y(n24347));
  xnor_4 g21396(.A(new_n5022), .B(new_n4979), .Y(n24373));
  xnor_4 g21397(.A(new_n17911_1), .B(new_n21267), .Y(n24406));
  xnor_4 g21398(.A(new_n13638), .B(new_n13626_1), .Y(n24415));
  xnor_4 g21399(.A(new_n10758), .B(new_n10756_1), .Y(n24421));
  xnor_4 g21400(.A(new_n13480), .B(new_n13457_1), .Y(n24431));
  xnor_4 g21401(.A(new_n11894), .B(new_n11871), .Y(n24472));
  and_5  g21402(.A(new_n22389), .B(new_n21918), .Y(new_n23751));
  nor_5  g21403(.A(new_n23751), .B(new_n22391), .Y(new_n23752));
  xor_4  g21404(.A(new_n23752), .B(new_n22386), .Y(n24476));
  xnor_4 g21405(.A(new_n10155), .B(new_n10116), .Y(n24483));
  xnor_4 g21406(.A(new_n22896), .B(new_n13376), .Y(n24501));
  xnor_4 g21407(.A(new_n18011), .B(new_n18008), .Y(n24512));
  xnor_4 g21408(.A(new_n4752), .B(new_n4751), .Y(n24558));
  xnor_4 g21409(.A(new_n2829), .B(new_n2826_1), .Y(n24576));
  xnor_4 g21410(.A(new_n2831), .B(new_n2830), .Y(n24579));
  xnor_4 g21411(.A(new_n20127), .B(new_n20115), .Y(n24602));
  xnor_4 g21412(.A(new_n14156), .B(new_n14123), .Y(n24604));
  xnor_4 g21413(.A(new_n22503), .B(new_n22500), .Y(n24626));
  xnor_4 g21414(.A(new_n21612), .B(new_n21610), .Y(n24629));
  xnor_4 g21415(.A(new_n21376), .B(new_n21365_1), .Y(n24636));
  xnor_4 g21416(.A(new_n21126), .B(new_n21123_1), .Y(n24715));
  xnor_4 g21417(.A(new_n20067), .B(new_n20018), .Y(n24723));
  xnor_4 g21418(.A(new_n16666), .B(new_n16627), .Y(new_n23767));
  xnor_4 g21419(.A(new_n23767), .B(new_n16736), .Y(n24749));
  xnor_4 g21420(.A(new_n20057), .B(new_n20035), .Y(n24758));
  xnor_4 g21421(.A(new_n22579), .B(new_n22576), .Y(n24784));
  xnor_4 g21422(.A(new_n16117), .B(new_n16116), .Y(n24807));
  xnor_4 g21423(.A(new_n9720), .B(new_n7889), .Y(n24826));
  xnor_4 g21424(.A(new_n7598_1), .B(new_n7564), .Y(n24840));
  xnor_4 g21425(.A(new_n9968_1), .B(new_n9955), .Y(n24841));
  xnor_4 g21426(.A(new_n5211_1), .B(new_n5199), .Y(n24853));
  xnor_4 g21427(.A(new_n3076_1), .B(new_n3051), .Y(n24857));
  xnor_4 g21428(.A(new_n6407_1), .B(new_n6393), .Y(n24887));
  xor_4  g21429(.A(new_n9207), .B(new_n9200), .Y(n24934));
  xnor_4 g21430(.A(new_n7425), .B(new_n7367), .Y(n24998));
  xnor_4 g21431(.A(new_n11567), .B(new_n11555), .Y(n25006));
  xnor_4 g21432(.A(new_n20429_1), .B(new_n20418), .Y(n25032));
  xnor_4 g21433(.A(new_n16068_1), .B(new_n16050), .Y(n25062));
  xnor_4 g21434(.A(new_n19253), .B(new_n16627), .Y(new_n23783));
  xnor_4 g21435(.A(new_n23783), .B(new_n19307), .Y(n25083));
  xor_4  g21436(.A(new_n12977), .B(new_n12974), .Y(n25097));
  xnor_4 g21437(.A(new_n17644), .B(new_n17641), .Y(n25133));
  xnor_4 g21438(.A(new_n18272), .B(new_n18253), .Y(n25155));
  xnor_4 g21439(.A(new_n23504), .B(new_n22377), .Y(new_n23788));
  xnor_4 g21440(.A(new_n23788), .B(new_n23501), .Y(n25181));
  xnor_4 g21441(.A(new_n20431), .B(new_n20416), .Y(n25200));
  nor_5  g21442(.A(new_n21141), .B(new_n21138_1), .Y(new_n23791));
  xnor_4 g21443(.A(new_n21135), .B(new_n16797), .Y(new_n23792));
  xnor_4 g21444(.A(new_n23792), .B(new_n23791), .Y(n25209));
  xnor_4 g21445(.A(new_n15038), .B(new_n15037), .Y(n25215));
  xor_4  g21446(.A(new_n18087), .B(new_n18084), .Y(n25244));
  xnor_4 g21447(.A(new_n17727), .B(new_n17708), .Y(n25254));
  xor_4  g21448(.A(new_n20617), .B(new_n20590_1), .Y(n25256));
  nor_5  g21449(.A(new_n22929), .B(new_n21220), .Y(new_n23798));
  nor_5  g21450(.A(new_n23798), .B(new_n22935), .Y(new_n23799));
  xnor_4 g21451(.A(new_n22928), .B(new_n22007), .Y(new_n23800));
  xnor_4 g21452(.A(new_n23800), .B(new_n23799), .Y(n25293));
  xor_4  g21453(.A(new_n20607), .B(new_n20600), .Y(n25328));
  xnor_4 g21454(.A(new_n11060), .B(new_n4301), .Y(n25332));
  nor_5  g21455(.A(new_n22564), .B(new_n21291), .Y(new_n23804));
  nor_5  g21456(.A(new_n22587), .B(new_n23804), .Y(new_n23805));
  and_5  g21457(.A(new_n22564), .B(new_n21291), .Y(new_n23806));
  nor_5  g21458(.A(new_n22586), .B(new_n23806), .Y(new_n23807));
  nor_5  g21459(.A(new_n23807), .B(new_n23805), .Y(n25337));
  xnor_4 g21460(.A(new_n11398_1), .B(new_n10840), .Y(new_n23809));
  xnor_4 g21461(.A(new_n23809), .B(new_n11403_1), .Y(n25356));
  xnor_4 g21462(.A(new_n9042_1), .B(new_n9031), .Y(n25362));
  xnor_4 g21463(.A(new_n14399), .B(new_n14382), .Y(n25412));
  xor_4  g21464(.A(new_n15312), .B(new_n15311), .Y(n25460));
  xnor_4 g21465(.A(new_n7417), .B(new_n7383), .Y(n25468));
  xnor_4 g21466(.A(new_n14401), .B(new_n14379), .Y(n25499));
  xnor_4 g21467(.A(new_n19643), .B(new_n19642), .Y(n25513));
  xnor_4 g21468(.A(new_n12095), .B(new_n12074), .Y(n25518));
  xnor_4 g21469(.A(new_n13302), .B(new_n13268), .Y(n25532));
  xnor_4 g21470(.A(new_n19970), .B(new_n19952), .Y(n25539));
  xnor_4 g21471(.A(new_n16872), .B(new_n16864), .Y(n25550));
  xnor_4 g21472(.A(new_n20728), .B(new_n20715), .Y(n25611));
  xnor_4 g21473(.A(new_n5433), .B(new_n5432), .Y(new_n23822));
  xnor_4 g21474(.A(new_n23822), .B(new_n5437), .Y(n25614));
  xnor_4 g21475(.A(new_n12726), .B(new_n12705), .Y(n25619));
  nor_5  g21476(.A(new_n22818), .B(new_n22682), .Y(new_n23825));
  nor_5  g21477(.A(new_n22823), .B(new_n23825), .Y(new_n23826));
  nor_5  g21478(.A(new_n22817), .B(new_n22683), .Y(new_n23827));
  nor_5  g21479(.A(new_n22822), .B(new_n23827), .Y(new_n23828));
  nor_5  g21480(.A(new_n23828), .B(new_n23826), .Y(n25665));
  xnor_4 g21481(.A(new_n9213), .B(new_n9191_1), .Y(n25706));
  xnor_4 g21482(.A(new_n22818), .B(new_n23461), .Y(new_n23831_1));
  xnor_4 g21483(.A(new_n23831_1), .B(new_n23466), .Y(n25719));
  xor_4  g21484(.A(new_n9701), .B(new_n9655_1), .Y(n25756));
  and_5  g21485(.A(new_n23201), .B(new_n12904_1), .Y(new_n23834));
  nor_5  g21486(.A(new_n12989), .B(new_n23834), .Y(new_n23835));
  nor_5  g21487(.A(new_n23201), .B(new_n12904_1), .Y(new_n23836));
  nor_5  g21488(.A(new_n12988), .B(new_n23836), .Y(new_n23837));
  nor_5  g21489(.A(new_n23837), .B(new_n23835), .Y(n25758));
  xnor_4 g21490(.A(new_n14772_1), .B(new_n5771), .Y(n25773));
  xnor_4 g21491(.A(new_n20520), .B(new_n17611), .Y(n25784));
  xnor_4 g21492(.A(new_n8380), .B(new_n8357), .Y(n25792));
  xnor_4 g21493(.A(new_n6958), .B(new_n6925), .Y(n25816));
  xnor_4 g21494(.A(new_n6413), .B(new_n6380), .Y(n25826));
  xnor_4 g21495(.A(new_n12287), .B(new_n12285), .Y(n25839));
  xnor_4 g21496(.A(new_n13984), .B(new_n13944), .Y(n25840));
  xnor_4 g21497(.A(new_n8192), .B(new_n8162), .Y(n25873));
  xor_4  g21498(.A(new_n23559), .B(new_n23556), .Y(n25934));
  xnor_4 g21499(.A(new_n20925), .B(new_n20912), .Y(n25938));
  xnor_4 g21500(.A(new_n21239), .B(new_n21236), .Y(n25985));
  xnor_4 g21501(.A(new_n13799), .B(new_n9033), .Y(n25994));
  nor_5  g21502(.A(new_n18224), .B(new_n18144), .Y(new_n23851));
  nor_5  g21503(.A(new_n18284), .B(new_n18225), .Y(new_n23852));
  or_5   g21504(.A(new_n23852), .B(new_n23851), .Y(n26084));
  xnor_4 g21505(.A(new_n22583), .B(new_n22570), .Y(n26096));
  or_5   g21506(.A(new_n11585), .B(new_n11523), .Y(new_n23855));
  nor_5  g21507(.A(new_n23855), .B(new_n11502), .Y(n26111));
  xnor_4 g21508(.A(new_n11572), .B(new_n11549), .Y(n26113));
  xor_4  g21509(.A(new_n20076), .B(new_n20073), .Y(n26156));
  xnor_4 g21510(.A(new_n17072), .B(new_n17050), .Y(n26159));
  xnor_4 g21511(.A(new_n3719), .B(new_n3674), .Y(n26179));
  xor_4  g21512(.A(new_n13970), .B(new_n13969), .Y(n26220));
  xnor_4 g21513(.A(new_n22622), .B(new_n22619_1), .Y(n26229));
  xnor_4 g21514(.A(new_n12655), .B(new_n12624), .Y(n26237));
  xnor_4 g21515(.A(new_n15707), .B(new_n15693), .Y(n26250));
  xor_4  g21516(.A(new_n20965), .B(new_n20962), .Y(n26274));
  xnor_4 g21517(.A(new_n15711), .B(new_n15685), .Y(n26287));
  xnor_4 g21518(.A(new_n21156), .B(new_n20438), .Y(new_n23867));
  xnor_4 g21519(.A(new_n23867), .B(new_n23387), .Y(n26317));
  nor_5  g21520(.A(new_n18553), .B(new_n18533), .Y(new_n23869));
  nor_5  g21521(.A(new_n23869), .B(new_n18549), .Y(new_n23870));
  nor_5  g21522(.A(new_n18552), .B(new_n18531), .Y(new_n23871));
  nor_5  g21523(.A(new_n23871), .B(new_n18548), .Y(new_n23872));
  nor_5  g21524(.A(new_n23872), .B(new_n23870), .Y(n26353));
  xnor_4 g21525(.A(new_n20125), .B(new_n20117), .Y(n26375));
  nor_5  g21526(.A(new_n22960), .B(new_n21276_1), .Y(new_n23875));
  nor_5  g21527(.A(new_n22969), .B(new_n22961), .Y(new_n23876));
  nor_5  g21528(.A(new_n23876), .B(new_n23875), .Y(n26396));
  xnor_4 g21529(.A(new_n22874), .B(new_n5435), .Y(n26429));
  xnor_4 g21530(.A(new_n14473), .B(new_n14458), .Y(n26431));
  xnor_4 g21531(.A(new_n7176), .B(new_n7120), .Y(n26439));
  xnor_4 g21532(.A(new_n20366_1), .B(new_n20365), .Y(n26492));
  xnor_4 g21533(.A(new_n10148), .B(new_n10147), .Y(n26515));
  xnor_4 g21534(.A(new_n2536), .B(new_n2510), .Y(n26538));
  xnor_4 g21535(.A(new_n14968), .B(new_n14955), .Y(n26590));
  xnor_4 g21536(.A(new_n19286), .B(new_n16714), .Y(n26598));
  xnor_4 g21537(.A(new_n22928), .B(new_n21220), .Y(new_n23886));
  xnor_4 g21538(.A(new_n23886), .B(new_n22933), .Y(n26605));
  xnor_4 g21539(.A(new_n22904), .B(new_n22898), .Y(new_n23888_1));
  xnor_4 g21540(.A(new_n23888_1), .B(new_n22901), .Y(n26656));
  xnor_4 g21541(.A(new_n11562), .B(new_n11561), .Y(n26674));
  xnor_4 g21542(.A(new_n9565), .B(new_n9549), .Y(n26675));
  xnor_4 g21543(.A(new_n20376), .B(new_n20347), .Y(n26681));
  nor_5  g21544(.A(new_n5698), .B(new_n5498), .Y(new_n23893));
  nor_5  g21545(.A(new_n5767), .B(new_n23893), .Y(new_n23894));
  nor_5  g21546(.A(new_n5699), .B(new_n5499), .Y(new_n23895_1));
  nor_5  g21547(.A(new_n5766), .B(new_n23895_1), .Y(new_n23896));
  nor_5  g21548(.A(new_n23896), .B(new_n23894), .Y(n26696));
  xnor_4 g21549(.A(new_n14730), .B(new_n14712), .Y(n26698));
  xnor_4 g21550(.A(new_n15442), .B(new_n5800), .Y(n26707));
  xor_4  g21551(.A(new_n23329), .B(new_n23327), .Y(n26719));
  xnor_4 g21552(.A(new_n9209), .B(new_n9197), .Y(n26727));
  nor_5  g21553(.A(new_n21290), .B(new_n19127), .Y(new_n23902));
  and_5  g21554(.A(new_n21295), .B(new_n21292), .Y(new_n23903_1));
  nor_5  g21555(.A(new_n23903_1), .B(new_n23902), .Y(n26729));
  xor_4  g21556(.A(new_n21315), .B(new_n21312), .Y(n26745));
  xnor_4 g21557(.A(new_n7906), .B(new_n7868), .Y(n26775));
  xnor_4 g21558(.A(new_n10501), .B(new_n10483), .Y(n26780));
  xor_4  g21559(.A(new_n21716), .B(new_n21709), .Y(n26794));
  xnor_4 g21560(.A(new_n3389), .B(new_n3340_1), .Y(n26795));
  xnor_4 g21561(.A(new_n10773), .B(new_n10735), .Y(n26801));
  xnor_4 g21562(.A(new_n11141), .B(new_n11123), .Y(n26815));
  xnor_4 g21563(.A(new_n23021), .B(new_n23018), .Y(n26847));
  xnor_4 g21564(.A(new_n18553), .B(new_n7361), .Y(new_n23913_1));
  xnor_4 g21565(.A(new_n23913_1), .B(new_n23141), .Y(n26900));
  xor_4  g21566(.A(new_n18693_1), .B(new_n18692), .Y(n26902));
  xor_4  g21567(.A(new_n17323), .B(new_n17320_1), .Y(n26905));
  xnor_4 g21568(.A(new_n8194_1), .B(new_n8157), .Y(n26921));
  xnor_4 g21569(.A(new_n22058), .B(new_n22045), .Y(n26923));
  xnor_4 g21570(.A(new_n10857), .B(new_n10856), .Y(n26929));
  xnor_4 g21571(.A(new_n12665_1), .B(new_n12599), .Y(n26930));
  xnor_4 g21572(.A(new_n15709), .B(new_n15689), .Y(n26943));
  xnor_4 g21573(.A(new_n14403), .B(new_n14376), .Y(n26970));
  xnor_4 g21574(.A(new_n20865), .B(new_n20854), .Y(n27004));
  xnor_4 g21575(.A(new_n10407), .B(new_n10353), .Y(n27011));
  xnor_4 g21576(.A(new_n19305), .B(new_n19256), .Y(n27019));
  xnor_4 g21577(.A(new_n5012), .B(new_n5001), .Y(n27031));
  xnor_4 g21578(.A(new_n21761), .B(new_n20960), .Y(new_n23927));
  xnor_4 g21579(.A(new_n23927), .B(new_n21800_1), .Y(n27051));
  xor_4  g21580(.A(new_n17197), .B(new_n17194), .Y(n27072));
  xnor_4 g21581(.A(new_n15327_1), .B(new_n15276), .Y(n27079));
  xnor_4 g21582(.A(new_n4302), .B(new_n4301), .Y(n27096));
  xor_4  g21583(.A(new_n14149), .B(new_n14138), .Y(n27110));
  xnor_4 g21584(.A(new_n13580), .B(new_n13577), .Y(n27112));
  xnor_4 g21585(.A(new_n22064), .B(new_n21612), .Y(n27130));
  xnor_4 g21586(.A(new_n16064), .B(new_n16056), .Y(n27145));
  nor_5  g21587(.A(new_n16501), .B(new_n14513), .Y(new_n23936));
  and_5  g21588(.A(new_n21462), .B(new_n21459), .Y(new_n23937));
  nor_5  g21589(.A(new_n23937), .B(new_n23936), .Y(n27158));
  xnor_4 g21590(.A(new_n21076), .B(new_n21073), .Y(n27163));
  xnor_4 g21591(.A(new_n23163), .B(new_n20872), .Y(new_n23940));
  xnor_4 g21592(.A(new_n23940), .B(new_n23168), .Y(n27194));
endmodule


