// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Sun Jun 23 19:37:07 2024

module top_810026173_826291639_946996917_1246901 ( 
    n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213, n223,
    n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414, n424,
    n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649, n653,
    n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788, n801,
    n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764,
    n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156, n174,
    n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299, n317,
    n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457, n460,
    n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547, n549,
    n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648, n665,
    n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773, n790,
    n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888, n891,
    n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989, n991,
    n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103, n1113,
    n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183, n1191,
    n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255, n1260,
    n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347, n1348,
    n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426, n1440,
    n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502, n1507,
    n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633, n1635,
    n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690, n1721,
    n1727, n1729, n1731, n1737, n1746  );
  input  n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213,
    n223, n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414,
    n424, n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649,
    n653, n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788,
    n801, n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764;
  output n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156,
    n174, n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299,
    n317, n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457,
    n460, n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547,
    n549, n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648,
    n665, n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773,
    n790, n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888,
    n891, n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989,
    n991, n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103,
    n1113, n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183,
    n1191, n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255,
    n1260, n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347,
    n1348, n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426,
    n1440, n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502,
    n1507, n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633,
    n1635, n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690,
    n1721, n1727, n1729, n1731, n1737, n1746;
  wire new_n276_1, new_n277_1, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290_1, new_n291, new_n292_1, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299_1, new_n300, new_n301,
    new_n302, new_n303_1, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317_1, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329_1,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347_1, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353_1, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372_1, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378_1, new_n379_1, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387_1, new_n388, new_n389, new_n390,
    new_n391_1, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401_1, new_n402_1, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414_1, new_n415, new_n416_1,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423_1,
    new_n424_1, new_n425, new_n426_1, new_n427, new_n428, new_n429_1,
    new_n430, new_n431, new_n432_1, new_n433_1, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444_1, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452_1, new_n453, new_n455, new_n456,
    new_n457_1, new_n458, new_n459, new_n460_1, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469_1,
    new_n470, new_n471, new_n472_1, new_n473, new_n474, new_n475,
    new_n476_1, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482_1, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488_1, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498_1, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510_1, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517_1, new_n518, new_n519, new_n520, new_n521, new_n522_1,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532_1, new_n533, new_n534_1, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541_1, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547_1, new_n548,
    new_n549_1, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555_1, new_n556, new_n557_1, new_n558, new_n559_1, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569_1, new_n570, new_n572, new_n573_1, new_n574,
    new_n575, new_n576, new_n577, new_n579, new_n581, new_n582, new_n585_1,
    new_n586, new_n587, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599_1, new_n600_1,
    new_n603, new_n604, new_n605, new_n606, new_n607_1, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627_1, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638_1, new_n639, new_n640, new_n641, new_n642, new_n643_1,
    new_n644, new_n645, new_n646_1, new_n647_1, new_n648_1, new_n649_1,
    new_n650, new_n651, new_n652, new_n653_1, new_n654, new_n655_1,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665_1, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675_1, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682_1,
    new_n683_1, new_n684_1, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693_1, new_n694,
    new_n695_1, new_n696, new_n697, new_n698, new_n699_1, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712_1, new_n713, new_n714,
    new_n715_1, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724_1, new_n725_1, new_n726, new_n727,
    new_n728, new_n729_1, new_n730, new_n731_1, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738_1, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747_1,
    new_n748_1, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759_1, new_n760,
    new_n761_1, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770_1, new_n771, new_n772, new_n773_1,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788_1,
    new_n789, new_n790_1, new_n791, new_n792_1, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801_1,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813_1, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823_1, new_n824_1, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836_1, new_n837, new_n838, new_n839_1, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846_1, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858_1, new_n859, new_n860, new_n862_1,
    new_n863, new_n864, new_n865_1, new_n866, new_n867_1, new_n868,
    new_n869, new_n870_1, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882_1,
    new_n883_1, new_n884, new_n885, new_n886, new_n887, new_n888_1,
    new_n889, new_n890, new_n891_1, new_n892_1, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902_1, new_n903, new_n904, new_n905_1, new_n906_1, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912_1, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927_1, new_n928, new_n929,
    new_n930, new_n931_1, new_n932, new_n933, new_n934, new_n935_1,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942_1,
    new_n943, new_n944_1, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952_1, new_n953_1, new_n954, new_n955,
    new_n957, new_n959, new_n960, new_n961_1, new_n964, new_n966, new_n967,
    new_n968_1, new_n970, new_n971, new_n972, new_n973, new_n974_1,
    new_n975, new_n976, new_n977, new_n978, new_n979_1, new_n980_1,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n991_1, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000_1, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005_1, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012_1, new_n1013, new_n1014,
    new_n1015_1, new_n1016_1, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025_1, new_n1026,
    new_n1028, new_n1029, new_n1030_1, new_n1031, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062_1, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067_1, new_n1068_1, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103_1, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113_1,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119_1,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135_1, new_n1136, new_n1137,
    new_n1138_1, new_n1140_1, new_n1142_1, new_n1144, new_n1145_1,
    new_n1146, new_n1147, new_n1148, new_n1149_1, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161_1, new_n1162_1, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172_1, new_n1173, new_n1174, new_n1175_1,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183_1, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191_1, new_n1192, new_n1193, new_n1194_1,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199_1, new_n1200,
    new_n1201_1, new_n1202_1, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222_1, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234_1, new_n1235_1, new_n1236,
    new_n1237_1, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249_1,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255_1,
    new_n1256, new_n1259, new_n1261, new_n1262, new_n1263_1, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277_1,
    new_n1278_1, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283_1,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296_1, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305_1, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315_1, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321_1, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330_1, new_n1331,
    new_n1332_1, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338_1, new_n1339, new_n1340_1, new_n1341_1, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347_1, new_n1348_1, new_n1349_1,
    new_n1350, new_n1351_1, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363_1, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369_1, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1380, new_n1382,
    new_n1383_1, new_n1384, new_n1385_1, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393_1, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399_1, new_n1400,
    new_n1402, new_n1404, new_n1405, new_n1408, new_n1409, new_n1410,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1423, new_n1424,
    new_n1425_1, new_n1426_1, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1432, new_n1433, new_n1434, new_n1435_1, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440_1, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453_1, new_n1455, new_n1457_1, new_n1460_1,
    new_n1461_1, new_n1462, new_n1463_1, new_n1464, new_n1465, new_n1466,
    new_n1468, new_n1469, new_n1471, new_n1474, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481_1, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495_1,
    new_n1496, new_n1497, new_n1498_1, new_n1499, new_n1500, new_n1501_1,
    new_n1502_1, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507_1,
    new_n1508, new_n1509, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525_1, new_n1526,
    new_n1527_1, new_n1528, new_n1529, new_n1530_1, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535_1, new_n1536, new_n1537_1, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544_1,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1555, new_n1556_1, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595_1,
    new_n1596, new_n1597_1, new_n1598, new_n1599, new_n1600_1, new_n1601_1,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613_1,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622_1, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1629_1, new_n1630, new_n1631,
    new_n1632, new_n1633_1, new_n1634, new_n1635_1, new_n1636, new_n1637,
    new_n1638, new_n1639, new_n1640, new_n1641, new_n1642_1, new_n1643_1,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654_1, new_n1655,
    new_n1656, new_n1657_1, new_n1658, new_n1659, new_n1660_1, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675_1, new_n1676, new_n1677_1, new_n1678_1, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683_1, new_n1684, new_n1685,
    new_n1686_1, new_n1687, new_n1688_1, new_n1689, new_n1690_1, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1703, new_n1706,
    new_n1707_1, new_n1708, new_n1709, new_n1710, new_n1711, new_n1713,
    new_n1717, new_n1719, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727_1, new_n1729_1, new_n1730, new_n1731_1, new_n1732,
    new_n1733, new_n1736, new_n1738, new_n1740, new_n1741, new_n1742,
    new_n1743_1, new_n1744, new_n1745, new_n1746_1, new_n1747_1, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757_1, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763_1, new_n1764_1, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1776, new_n1779, new_n1782, new_n1783,
    new_n1785, new_n1787, new_n1789, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1796, new_n1798, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1807, new_n1809,
    new_n1812, new_n1814, new_n1816, new_n1817, new_n1818, new_n1820,
    new_n1822, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1830, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1854,
    new_n1855, new_n1856, new_n1858, new_n1859, new_n1860, new_n1863,
    new_n1864, new_n1867, new_n1870, new_n1873, new_n1875, new_n1876,
    new_n1877, new_n1878, new_n1880, new_n1882, new_n1883, new_n1885,
    new_n1887, new_n1889, new_n1891, new_n1892, new_n1893, new_n1894,
    new_n1895, new_n1897, new_n1899, new_n1901, new_n1905, new_n1906,
    new_n1907, new_n1908, new_n1910, new_n1911, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1918, new_n1919, new_n1921, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1943, new_n1945,
    new_n1946, new_n1949, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1957, new_n1959, new_n1961, new_n1962, new_n1963, new_n1965,
    new_n1966, new_n1969, new_n1970, new_n1972, new_n1974, new_n1976,
    new_n1978, new_n1980, new_n1982, new_n1983, new_n1984, new_n1986,
    new_n1987, new_n1989, new_n1991, new_n1993, new_n1995, new_n1996,
    new_n1998, new_n2002, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2009, new_n2012, new_n2014, new_n2016, new_n2018, new_n2021,
    new_n2024, new_n2025, new_n2027, new_n2029, new_n2030, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2038, new_n2042, new_n2043,
    new_n2045, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2055, new_n2057, new_n2059, new_n2060, new_n2061, new_n2063,
    new_n2064, new_n2065;
not_13 g0000(n36, new_n276_1);
not_13 g0001(n1643, new_n277_1);
and_7  g0002(new_n277_1, new_n276_1, new_n278);
xor_5  g0003(n1643, n36, new_n279);
or_2   g0004(n788, n555, new_n280);
not_13 g0005(new_n280, new_n281);
and_7  g0006(n788, n555, new_n282);
not_13 g0007(new_n282, new_n283);
and_7  g0008(new_n283, new_n280, new_n284);
not_13 g0009(n353, new_n285);
not_13 g0010(n747, new_n286);
and_7  g0011(new_n286, new_n285, new_n287);
xor_5  g0012(n747, new_n285, new_n288);
or_2   g0013(n952, n329, new_n289);
and_7  g0014(n1145, n931, new_n290_1);
nor_6  g0015(n952, n329, new_n291);
and_7  g0016(n952, n329, new_n292_1);
or_2   g0017(new_n292_1, new_n291, new_n293);
or_2   g0018(new_n293, new_n290_1, new_n294);
and_7  g0019(new_n294, new_n289, new_n295);
nor_6  g0020(new_n295, new_n288, new_n296);
or_2   g0021(new_n296, new_n287, new_n297);
and_7  g0022(new_n297, new_n284, new_n298);
or_2   g0023(new_n298, new_n281, new_n299_1);
and_7  g0024(new_n299_1, new_n279, new_n300);
nor_6  g0025(new_n300, new_n278, new_n301);
and_7  g0026(new_n301, n1501, new_n302);
and_7  g0027(new_n302, n433, new_n303_1);
nor_6  g0028(new_n302, n433, new_n304);
nor_6  g0029(new_n304, new_n303_1, new_n305);
and_7  g0030(n1000, n870, new_n306);
not_13 g0031(n1000, new_n307);
and_7  g0032(new_n307, n66, new_n308);
nor_6  g0033(new_n308, new_n306, new_n309);
and_7  g0034(n1000, n585, new_n310);
and_7  g0035(new_n307, n968, new_n311);
nor_6  g0036(new_n311, new_n310, new_n312);
and_7  g0037(new_n312, new_n309, new_n313);
and_7  g0038(n1000, n155, new_n314);
not_13 g0039(new_n314, new_n315);
not_13 g0040(n1435, new_n316);
or_2   g0041(new_n316, n1000, new_n317_1);
and_7  g0042(new_n317_1, new_n315, new_n318);
and_7  g0043(new_n318, new_n313, new_n319);
or_2   g0044(n1000, n682, new_n320);
or_2   g0045(n1678, new_n307, new_n321);
and_7  g0046(new_n321, new_n320, new_n322);
and_7  g0047(new_n322, new_n319, new_n323);
xor_5  g0048(n1597, n682, new_n324);
nor_6  g0049(new_n324, n1000, new_n325);
xor_5  g0050(n1678, n607, new_n326);
and_7  g0051(new_n326, n1000, new_n327);
nor_6  g0052(new_n327, new_n325, new_n328);
and_7  g0053(new_n328, new_n323, new_n329_1);
not_13 g0054(new_n323, new_n330);
or_2   g0055(new_n327, new_n325, new_n331);
and_7  g0056(new_n331, new_n330, new_n332);
or_2   g0057(new_n332, new_n329_1, new_n333);
not_13 g0058(n682, new_n334);
and_7  g0059(new_n307, new_n334, new_n335);
not_13 g0060(n1678, new_n336);
and_7  g0061(new_n336, n1000, new_n337);
or_2   g0062(new_n337, new_n335, new_n338);
xor_5  g0063(new_n338, new_n319, new_n339);
and_7  g0064(n1435, new_n307, new_n340);
or_2   g0065(new_n340, new_n314, new_n341);
xor_5  g0066(new_n341, new_n313, new_n342);
not_13 g0067(n693, new_n343);
xor_5  g0068(new_n312, new_n309, new_n344);
and_7  g0069(new_n344, new_n343, new_n345);
or_2   g0070(new_n344, new_n343, new_n346);
not_13 g0071(n1763, new_n347_1);
or_2   g0072(new_n311, new_n310, new_n348);
or_2   g0073(new_n348, new_n347_1, new_n349);
and_7  g0074(new_n348, new_n347_1, new_n350);
not_13 g0075(n1530, new_n351);
and_7  g0076(n1461, n1000, new_n352);
and_7  g0077(new_n307, n347, new_n353_1);
nor_6  g0078(new_n353_1, new_n352, new_n354);
or_2   g0079(new_n354, new_n351, new_n355);
or_2   g0080(new_n355, new_n350, new_n356);
and_7  g0081(new_n356, new_n349, new_n357);
and_7  g0082(new_n357, new_n346, new_n358);
nor_6  g0083(new_n358, new_n345, new_n359);
and_7  g0084(new_n359, new_n342, new_n360);
and_7  g0085(new_n360, new_n339, new_n361);
and_7  g0086(new_n361, new_n333, new_n362);
not_13 g0087(n26, new_n363);
and_7  g0088(n1678, n607, new_n364);
not_13 g0089(new_n364, new_n365);
and_7  g0090(new_n365, new_n363, new_n366);
and_7  g0091(n607, n26, new_n367);
and_7  g0092(new_n367, n1678, new_n368);
or_2   g0093(new_n368, new_n366, new_n369);
and_7  g0094(new_n369, n1000, new_n370);
or_2   g0095(n1597, n46, new_n371);
or_2   g0096(new_n371, n682, new_n372_1);
not_13 g0097(n46, new_n373);
not_13 g0098(n1597, new_n374);
and_7  g0099(new_n374, new_n334, new_n375);
or_2   g0100(new_n375, new_n373, new_n376);
and_7  g0101(new_n376, new_n372_1, new_n377);
and_7  g0102(new_n377, new_n307, new_n378_1);
or_2   g0103(new_n378_1, new_n370, new_n379_1);
nor_6  g0104(new_n379_1, new_n329_1, new_n380);
and_7  g0105(new_n379_1, new_n329_1, new_n381);
or_2   g0106(new_n381, new_n380, new_n382);
and_7  g0107(new_n382, new_n362, new_n383);
nor_6  g0108(new_n382, new_n362, new_n384);
nor_6  g0109(new_n384, new_n383, new_n385);
and_7  g0110(new_n385, new_n305, new_n386);
nor_6  g0111(new_n385, new_n305, new_n387_1);
or_2   g0112(new_n387_1, new_n386, new_n388);
nor_6  g0113(new_n361, new_n333, new_n389);
nor_6  g0114(new_n389, new_n362, new_n390);
not_13 g0115(n1501, new_n391_1);
or_2   g0116(new_n300, new_n278, new_n392);
or_2   g0117(new_n392, new_n391_1, new_n393);
or_2   g0118(new_n301, n1501, new_n394);
and_7  g0119(new_n394, new_n393, new_n395);
nor_6  g0120(new_n395, new_n390, new_n396);
and_7  g0121(new_n395, new_n390, new_n397);
nor_6  g0122(new_n397, new_n396, new_n398);
nor_6  g0123(new_n360, new_n339, new_n399);
nor_6  g0124(new_n399, new_n361, new_n400);
nor_6  g0125(new_n299_1, new_n279, new_n401_1);
or_2   g0126(new_n401_1, new_n300, new_n402_1);
and_7  g0127(new_n402_1, new_n400, new_n403);
nor_6  g0128(new_n359, new_n342, new_n404);
nor_6  g0129(new_n404, new_n360, new_n405);
nor_6  g0130(new_n297, new_n284, new_n406);
or_2   g0131(new_n406, new_n298, new_n407);
nor_6  g0132(new_n407, new_n405, new_n408);
and_7  g0133(new_n407, new_n405, new_n409);
nor_6  g0134(new_n409, new_n408, new_n410);
and_7  g0135(new_n295, new_n288, new_n411);
or_2   g0136(new_n411, new_n296, new_n412);
xor_5  g0137(n1145, n931, new_n413);
xor_5  g0138(new_n354, new_n351, new_n414_1);
and_7  g0139(new_n414_1, new_n413, new_n415);
not_13 g0140(new_n292_1, new_n416_1);
and_7  g0141(new_n416_1, new_n289, new_n417);
xor_5  g0142(new_n417, new_n290_1, new_n418);
nor_6  g0143(new_n418, new_n415, new_n419);
not_13 g0144(n1145, new_n420);
xor_5  g0145(new_n420, n931, new_n421);
xor_5  g0146(new_n354, n1530, new_n422);
or_2   g0147(new_n422, new_n421, new_n423_1);
or_2   g0148(new_n423_1, new_n293, new_n424_1);
xor_5  g0149(new_n312, new_n347_1, new_n425);
and_7  g0150(new_n425, new_n355, new_n426_1);
or_2   g0151(new_n353_1, new_n352, new_n427);
and_7  g0152(new_n427, n1530, new_n428);
xor_5  g0153(new_n312, n1763, new_n429_1);
and_7  g0154(new_n429_1, new_n428, new_n430);
or_2   g0155(new_n430, new_n426_1, new_n431);
and_7  g0156(new_n431, new_n424_1, new_n432_1);
nor_6  g0157(new_n432_1, new_n419, new_n433_1);
nor_6  g0158(new_n433_1, new_n412, new_n434);
and_7  g0159(new_n433_1, new_n412, new_n435);
xor_5  g0160(new_n348, new_n309, new_n436);
and_7  g0161(new_n436, n693, new_n437);
nor_6  g0162(new_n437, new_n345, new_n438);
nor_6  g0163(new_n438, new_n357, new_n439);
and_7  g0164(new_n438, new_n357, new_n440);
or_2   g0165(new_n440, new_n439, new_n441);
nor_6  g0166(new_n441, new_n435, new_n442);
or_2   g0167(new_n442, new_n434, new_n443);
and_7  g0168(new_n443, new_n410, new_n444_1);
nor_6  g0169(new_n444_1, new_n408, new_n445);
nor_6  g0170(new_n402_1, new_n400, new_n446);
nor_6  g0171(new_n446, new_n403, new_n447);
and_7  g0172(new_n447, new_n445, new_n448);
nor_6  g0173(new_n448, new_n403, new_n449);
and_7  g0174(new_n449, new_n398, new_n450);
nor_6  g0175(new_n450, new_n396, new_n451);
nor_6  g0176(new_n451, new_n388, new_n452_1);
and_7  g0177(new_n451, new_n388, new_n453);
or_2   g0178(new_n453, new_n452_1, n19);
not_13 g0179(n69, new_n455);
not_13 g0180(n1381, new_n456);
and_7  g0181(new_n456, n402, new_n457_1);
nor_6  g0182(new_n457_1, n870, new_n458);
not_13 g0183(n66, new_n459);
and_7  g0184(new_n457_1, new_n459, new_n460_1);
nor_6  g0185(new_n460_1, new_n458, new_n461);
xor_5  g0186(new_n461, new_n455, new_n462);
nor_6  g0187(new_n457_1, n585, new_n463);
not_13 g0188(n968, new_n464);
and_7  g0189(new_n457_1, new_n464, new_n465);
nor_6  g0190(new_n465, new_n463, new_n466);
and_7  g0191(new_n466, n953, new_n467);
nor_6  g0192(new_n457_1, n1461, new_n468);
not_13 g0193(n347, new_n469_1);
and_7  g0194(new_n457_1, new_n469_1, new_n470);
nor_6  g0195(new_n470, new_n468, new_n471);
and_7  g0196(new_n471, n303, new_n472_1);
xor_5  g0197(new_n466, n953, new_n473);
and_7  g0198(new_n473, new_n472_1, new_n474);
nor_6  g0199(new_n474, new_n467, new_n475);
nor_6  g0200(new_n475, new_n462, new_n476_1);
and_7  g0201(new_n475, new_n462, new_n477);
nor_6  g0202(new_n477, new_n476_1, new_n478);
and_7  g0203(new_n478, new_n412, new_n479);
nor_6  g0204(new_n478, new_n412, new_n480);
or_2   g0205(new_n480, new_n479, new_n481);
xor_5  g0206(new_n471, n303, new_n482_1);
and_7  g0207(new_n482_1, new_n413, new_n483);
nor_6  g0208(new_n483, new_n418, new_n484);
nor_6  g0209(new_n473, new_n472_1, new_n485);
or_2   g0210(new_n485, new_n474, new_n486);
and_7  g0211(new_n483, new_n417, new_n487);
nor_6  g0212(new_n487, new_n484, new_n488_1);
and_7  g0213(new_n488_1, new_n486, new_n489);
nor_6  g0214(new_n489, new_n484, new_n490);
and_7  g0215(new_n490, new_n481, new_n491);
nor_6  g0216(new_n490, new_n481, new_n492);
or_2   g0217(new_n492, new_n491, n33);
not_13 g0218(n1642, new_n494);
or_2   g0219(n607, n26, new_n495);
or_2   g0220(new_n495, n247, new_n496);
xor_5  g0221(new_n496, new_n494, new_n497);
and_7  g0222(new_n497, n1381, new_n498_1);
not_13 g0223(n379, new_n499);
not_13 g0224(n1527, new_n500);
and_7  g0225(new_n500, new_n373, new_n501);
and_7  g0226(new_n501, new_n499, new_n502);
not_13 g0227(n402, new_n503);
or_2   g0228(n1527, n46, new_n504);
and_7  g0229(new_n504, n379, new_n505);
or_2   g0230(new_n505, new_n503, new_n506);
or_2   g0231(new_n506, new_n502, new_n507);
and_7  g0232(n1642, new_n456, new_n508);
or_2   g0233(new_n508, new_n457_1, new_n509);
and_7  g0234(new_n509, new_n507, new_n510_1);
or_2   g0235(new_n510_1, new_n498_1, new_n511);
not_13 g0236(n247, new_n512);
xor_5  g0237(new_n495, new_n512, new_n513);
and_7  g0238(new_n513, n1381, new_n514);
and_7  g0239(n1527, n46, new_n515);
not_13 g0240(new_n515, new_n516);
and_7  g0241(new_n516, n402, new_n517_1);
and_7  g0242(new_n517_1, new_n504, new_n518);
not_13 g0243(new_n518, new_n519);
and_7  g0244(new_n456, n247, new_n520);
or_2   g0245(new_n520, new_n457_1, new_n521);
and_7  g0246(new_n521, new_n519, new_n522_1);
or_2   g0247(new_n522_1, new_n514, new_n523);
or_2   g0248(n1381, new_n503, new_n524);
and_7  g0249(new_n524, new_n336, new_n525);
and_7  g0250(new_n457_1, new_n334, new_n526);
or_2   g0251(new_n526, new_n525, new_n527);
and_7  g0252(new_n527, new_n277_1, new_n528);
xor_5  g0253(new_n527, new_n277_1, new_n529);
nor_6  g0254(new_n457_1, n155, new_n530);
and_7  g0255(new_n457_1, new_n316, new_n531);
or_2   g0256(new_n531, new_n530, new_n532_1);
not_13 g0257(new_n532_1, new_n533);
and_7  g0258(new_n533, n555, new_n534_1);
or_2   g0259(new_n461, n353, new_n535);
xor_5  g0260(new_n461, new_n285, new_n536);
or_2   g0261(new_n466, n952, new_n537);
and_7  g0262(new_n471, n1145, new_n538);
not_13 g0263(n952, new_n539);
xor_5  g0264(new_n466, new_n539, new_n540);
or_2   g0265(new_n540, new_n538, new_n541_1);
and_7  g0266(new_n541_1, new_n537, new_n542);
or_2   g0267(new_n542, new_n536, new_n543);
and_7  g0268(new_n543, new_n535, new_n544);
not_13 g0269(n555, new_n545);
xor_5  g0270(new_n532_1, new_n545, new_n546);
and_7  g0271(new_n546, new_n544, new_n547_1);
nor_6  g0272(new_n547_1, new_n534_1, new_n548);
and_7  g0273(new_n548, new_n529, new_n549_1);
nor_6  g0274(new_n549_1, new_n528, new_n550);
and_7  g0275(n1381, n607, new_n551);
and_7  g0276(new_n374, n402, new_n552);
not_13 g0277(n607, new_n553);
and_7  g0278(new_n553, new_n503, new_n554);
or_2   g0279(new_n554, new_n552, new_n555_1);
and_7  g0280(new_n555_1, new_n456, new_n556);
or_2   g0281(new_n556, new_n551, new_n557_1);
not_13 g0282(new_n557_1, new_n558);
and_7  g0283(new_n558, new_n550, new_n559_1);
and_7  g0284(n402, n46, new_n560);
and_7  g0285(new_n503, new_n363, new_n561);
or_2   g0286(new_n561, new_n560, new_n562);
and_7  g0287(new_n562, new_n456, new_n563);
not_13 g0288(new_n367, new_n564);
and_7  g0289(new_n495, new_n564, new_n565);
and_7  g0290(new_n565, n1381, new_n566);
or_2   g0291(new_n566, new_n563, new_n567);
not_13 g0292(new_n567, new_n568);
and_7  g0293(new_n568, new_n559_1, new_n569_1);
and_7  g0294(new_n569_1, new_n523, new_n570);
xor_5  g0295(new_n570, new_n511, n1731);
nor_6  g0296(new_n522_1, new_n514, new_n572);
or_2   g0297(new_n549_1, new_n528, new_n573_1);
or_2   g0298(new_n557_1, new_n573_1, new_n574);
or_2   g0299(new_n567, new_n574, new_n575);
or_2   g0300(new_n575, new_n572, new_n576);
or_2   g0301(new_n569_1, new_n523, new_n577);
and_7  g0302(new_n577, new_n576, n1138);
or_2   g0303(new_n558, new_n550, new_n579);
and_7  g0304(new_n579, new_n574, n1727);
nor_6  g0305(new_n540, new_n538, new_n581);
and_7  g0306(new_n540, new_n538, new_n582);
or_2   g0307(new_n582, new_n581, n1457);
xor_5  g0308(new_n471, n1145, n1183);
or_2   g0309(n1183, n1457, new_n585_1);
not_13 g0310(new_n537, new_n586);
or_2   g0311(new_n581, new_n586, new_n587);
xor_5  g0312(new_n587, new_n536, n416);
or_2   g0313(n416, new_n585_1, new_n589);
nor_6  g0314(new_n546, new_n544, new_n590);
nor_6  g0315(new_n590, new_n547_1, n1721);
nor_6  g0316(n1721, new_n589, new_n592);
nor_6  g0317(new_n548, new_n529, new_n593);
nor_6  g0318(new_n593, new_n549_1, new_n594);
nor_6  g0319(new_n594, new_n592, new_n595);
and_7  g0320(new_n595, n1727, new_n596);
and_7  g0321(new_n596, new_n568, new_n597);
and_7  g0322(new_n597, n1138, new_n598);
nor_6  g0323(new_n598, n1731, new_n599_1);
and_7  g0324(new_n598, new_n511, new_n600_1);
nor_6  g0325(new_n600_1, new_n599_1, n44);
xor_5  g0326(new_n414_1, new_n413, n55);
not_13 g0327(n1707, new_n603);
and_7  g0328(new_n603, new_n277_1, new_n604);
not_13 g0329(new_n604, new_n605);
xor_5  g0330(n1707, new_n277_1, new_n606);
not_13 g0331(n1140, new_n607_1);
and_7  g0332(new_n607_1, new_n545, new_n608);
xor_5  g0333(n1140, n555, new_n609);
not_13 g0334(n1351, new_n610);
and_7  g0335(new_n610, new_n285, new_n611);
xor_5  g0336(n1351, new_n285, new_n612);
or_2   g0337(n952, n729, new_n613);
and_7  g0338(n1145, n684, new_n614);
not_13 g0339(n729, new_n615);
xor_5  g0340(n952, new_n615, new_n616);
or_2   g0341(new_n616, new_n614, new_n617);
and_7  g0342(new_n617, new_n613, new_n618);
nor_6  g0343(new_n618, new_n612, new_n619);
or_2   g0344(new_n619, new_n611, new_n620);
and_7  g0345(new_n620, new_n609, new_n621);
nor_6  g0346(new_n621, new_n608, new_n622);
or_2   g0347(new_n622, new_n606, new_n623);
and_7  g0348(new_n623, new_n605, new_n624);
and_7  g0349(new_n624, n1332, new_n625);
and_7  g0350(new_n625, n391, new_n626);
and_7  g0351(new_n626, n1544, new_n627_1);
not_13 g0352(n1544, new_n628);
not_13 g0353(n391, new_n629);
not_13 g0354(n1332, new_n630);
and_7  g0355(n1707, n1643, new_n631);
not_13 g0356(new_n631, new_n632);
and_7  g0357(new_n632, new_n605, new_n633);
or_2   g0358(new_n621, new_n608, new_n634);
and_7  g0359(new_n634, new_n633, new_n635);
or_2   g0360(new_n635, new_n604, new_n636);
or_2   g0361(new_n636, new_n630, new_n637);
or_2   g0362(new_n637, new_n629, new_n638_1);
and_7  g0363(new_n638_1, new_n628, new_n639);
nor_6  g0364(new_n639, new_n627_1, new_n640);
and_7  g0365(n266, n155, new_n641);
not_13 g0366(n266, new_n642);
and_7  g0367(n1435, new_n642, new_n643_1);
nor_6  g0368(new_n643_1, new_n641, new_n644);
and_7  g0369(n870, n266, new_n645);
and_7  g0370(new_n642, n66, new_n646_1);
nor_6  g0371(new_n646_1, new_n645, new_n647_1);
and_7  g0372(new_n647_1, new_n644, new_n648_1);
and_7  g0373(n1678, n266, new_n649_1);
not_13 g0374(new_n649_1, new_n650);
or_2   g0375(new_n334, n266, new_n651);
and_7  g0376(new_n651, new_n650, new_n652);
and_7  g0377(new_n652, new_n648_1, new_n653_1);
and_7  g0378(n1597, new_n642, new_n654);
and_7  g0379(new_n553, n266, new_n655_1);
or_2   g0380(new_n655_1, new_n654, new_n656);
and_7  g0381(new_n656, new_n653_1, new_n657);
and_7  g0382(n266, new_n363, new_n658);
not_13 g0383(new_n658, new_n659);
xor_5  g0384(n1597, new_n373, new_n660);
or_2   g0385(new_n660, n266, new_n661);
and_7  g0386(new_n661, new_n659, new_n662);
xor_5  g0387(new_n662, new_n657, new_n663);
or_2   g0388(new_n374, n266, new_n664);
or_2   g0389(n607, new_n642, new_n665_1);
and_7  g0390(new_n665_1, new_n664, new_n666);
xor_5  g0391(new_n666, new_n653_1, new_n667);
and_7  g0392(n682, new_n642, new_n668);
or_2   g0393(new_n668, new_n649_1, new_n669);
xor_5  g0394(new_n669, new_n648_1, new_n670);
or_2   g0395(new_n643_1, new_n641, new_n671);
xor_5  g0396(new_n647_1, new_n671, new_n672);
and_7  g0397(new_n672, n223, new_n673);
not_13 g0398(n223, new_n674);
xor_5  g0399(new_n647_1, new_n644, new_n675_1);
and_7  g0400(new_n675_1, new_n674, new_n676);
or_2   g0401(new_n676, new_n673, new_n677);
and_7  g0402(new_n647_1, n444, new_n678);
and_7  g0403(n585, n266, new_n679);
and_7  g0404(n968, new_n642, new_n680);
or_2   g0405(new_n680, new_n679, new_n681);
or_2   g0406(new_n681, n472, new_n682_1);
and_7  g0407(n1461, n266, new_n683_1);
and_7  g0408(n347, new_n642, new_n684_1);
or_2   g0409(new_n684_1, new_n683_1, new_n685);
and_7  g0410(new_n685, n801, new_n686);
not_13 g0411(new_n679, new_n687);
or_2   g0412(new_n464, n266, new_n688);
and_7  g0413(new_n688, new_n687, new_n689);
xor_5  g0414(new_n689, n472, new_n690);
or_2   g0415(new_n690, new_n686, new_n691);
and_7  g0416(new_n691, new_n682_1, new_n692);
xor_5  g0417(new_n647_1, n444, new_n693_1);
and_7  g0418(new_n693_1, new_n692, new_n694);
nor_6  g0419(new_n694, new_n678, new_n695_1);
nor_6  g0420(new_n695_1, new_n677, new_n696);
or_2   g0421(new_n696, new_n673, new_n697);
and_7  g0422(new_n697, new_n670, new_n698);
and_7  g0423(new_n698, new_n667, new_n699_1);
and_7  g0424(new_n699_1, new_n663, new_n700);
nor_6  g0425(new_n660, n266, new_n701);
or_2   g0426(new_n701, new_n658, new_n702);
and_7  g0427(new_n702, new_n657, new_n703);
or_2   g0428(new_n504, n1597, new_n704);
and_7  g0429(new_n374, new_n373, new_n705);
or_2   g0430(new_n705, new_n500, new_n706);
and_7  g0431(new_n706, new_n704, new_n707);
and_7  g0432(new_n707, new_n642, new_n708);
and_7  g0433(n266, new_n512, new_n709);
nor_6  g0434(new_n709, new_n708, new_n710);
xor_5  g0435(new_n710, new_n703, new_n711);
and_7  g0436(new_n711, new_n700, new_n712_1);
nor_6  g0437(new_n711, new_n700, new_n713);
nor_6  g0438(new_n713, new_n712_1, new_n714);
nor_6  g0439(new_n714, new_n640, new_n715_1);
and_7  g0440(new_n714, new_n640, new_n716);
or_2   g0441(new_n716, new_n715_1, new_n717);
or_2   g0442(new_n625, n391, new_n718);
and_7  g0443(new_n718, new_n638_1, new_n719);
nor_6  g0444(new_n699_1, new_n663, new_n720);
nor_6  g0445(new_n720, new_n700, new_n721);
nor_6  g0446(new_n721, new_n719, new_n722);
xor_5  g0447(new_n656, new_n653_1, new_n723);
xor_5  g0448(new_n652, new_n648_1, new_n724_1);
nor_6  g0449(new_n696, new_n673, new_n725_1);
or_2   g0450(new_n725_1, new_n724_1, new_n726);
and_7  g0451(new_n726, new_n723, new_n727);
nor_6  g0452(new_n727, new_n699_1, new_n728);
and_7  g0453(new_n636, new_n630, new_n729_1);
nor_6  g0454(new_n729_1, new_n625, new_n730);
or_2   g0455(new_n730, new_n728, new_n731_1);
nor_6  g0456(new_n730, new_n728, new_n732);
and_7  g0457(new_n730, new_n728, new_n733);
or_2   g0458(new_n733, new_n732, new_n734);
and_7  g0459(new_n725_1, new_n724_1, new_n735);
nor_6  g0460(new_n735, new_n698, new_n736);
and_7  g0461(new_n622, new_n606, new_n737);
or_2   g0462(new_n737, new_n635, new_n738_1);
nor_6  g0463(new_n738_1, new_n736, new_n739);
and_7  g0464(new_n738_1, new_n736, new_n740);
nor_6  g0465(new_n740, new_n739, new_n741);
and_7  g0466(new_n695_1, new_n677, new_n742);
nor_6  g0467(new_n742, new_n696, new_n743);
nor_6  g0468(new_n620, new_n609, new_n744);
or_2   g0469(new_n744, new_n621, new_n745);
nor_6  g0470(new_n745, new_n743, new_n746);
and_7  g0471(new_n745, new_n743, new_n747_1);
or_2   g0472(new_n747_1, new_n746, new_n748_1);
nor_6  g0473(new_n693_1, new_n692, new_n749);
nor_6  g0474(new_n749, new_n694, new_n750);
and_7  g0475(new_n618, new_n612, new_n751);
or_2   g0476(new_n751, new_n619, new_n752);
nor_6  g0477(new_n752, new_n750, new_n753);
not_13 g0478(new_n614, new_n754);
and_7  g0479(n952, n729, new_n755);
not_13 g0480(new_n755, new_n756);
and_7  g0481(new_n756, new_n613, new_n757);
or_2   g0482(new_n757, new_n754, new_n758);
and_7  g0483(new_n757, new_n754, new_n759_1);
xor_5  g0484(n1145, n684, new_n760);
xor_5  g0485(new_n685, n801, new_n761_1);
and_7  g0486(new_n761_1, new_n760, new_n762);
nor_6  g0487(new_n762, new_n759_1, new_n763);
and_7  g0488(new_n763, new_n758, new_n764);
not_13 g0489(new_n686, new_n765);
xor_5  g0490(new_n681, n472, new_n766);
or_2   g0491(new_n766, new_n765, new_n767);
and_7  g0492(new_n767, new_n691, new_n768);
and_7  g0493(new_n762, new_n757, new_n769);
nor_6  g0494(new_n769, new_n764, new_n770_1);
and_7  g0495(new_n770_1, new_n768, new_n771);
or_2   g0496(new_n771, new_n764, new_n772);
and_7  g0497(new_n752, new_n750, new_n773_1);
nor_6  g0498(new_n773_1, new_n753, new_n774);
and_7  g0499(new_n774, new_n772, new_n775);
nor_6  g0500(new_n775, new_n753, new_n776);
nor_6  g0501(new_n776, new_n748_1, new_n777);
or_2   g0502(new_n777, new_n746, new_n778);
and_7  g0503(new_n778, new_n741, new_n779);
nor_6  g0504(new_n779, new_n739, new_n780);
or_2   g0505(new_n780, new_n734, new_n781);
and_7  g0506(new_n781, new_n731_1, new_n782);
and_7  g0507(new_n721, new_n719, new_n783);
or_2   g0508(new_n783, new_n722, new_n784);
nor_6  g0509(new_n784, new_n782, new_n785);
or_2   g0510(new_n785, new_n722, new_n786);
xor_5  g0511(new_n786, new_n717, n56);
or_2   g0512(new_n709, new_n708, new_n788_1);
and_7  g0513(new_n788_1, new_n703, new_n789);
and_7  g0514(new_n494, n266, new_n790_1);
not_13 g0515(new_n790_1, new_n791);
xor_5  g0516(new_n704, new_n499, new_n792_1);
or_2   g0517(new_n792_1, n266, new_n793);
and_7  g0518(new_n793, new_n791, new_n794);
xor_5  g0519(new_n794, new_n789, new_n795);
and_7  g0520(new_n795, new_n712_1, new_n796);
nor_6  g0521(new_n792_1, n266, new_n797);
or_2   g0522(new_n797, new_n790_1, new_n798);
and_7  g0523(new_n798, new_n789, new_n799);
not_13 g0524(n171, new_n800);
and_7  g0525(n266, new_n800, new_n801_1);
not_13 g0526(new_n801_1, new_n802);
or_2   g0527(new_n704, n379, new_n803);
and_7  g0528(new_n803, n1263, new_n804);
not_13 g0529(n1263, new_n805);
and_7  g0530(new_n501, new_n374, new_n806);
and_7  g0531(new_n806, new_n499, new_n807);
and_7  g0532(new_n807, new_n805, new_n808);
or_2   g0533(new_n808, n266, new_n809);
or_2   g0534(new_n809, new_n804, new_n810);
and_7  g0535(new_n810, new_n802, new_n811);
xor_5  g0536(new_n811, new_n799, new_n812);
and_7  g0537(new_n812, new_n796, new_n813_1);
not_13 g0538(new_n804, new_n814);
or_2   g0539(new_n803, n1263, new_n815);
and_7  g0540(new_n815, new_n642, new_n816);
and_7  g0541(new_n816, new_n814, new_n817);
or_2   g0542(new_n817, new_n801_1, new_n818);
and_7  g0543(new_n818, new_n799, new_n819);
and_7  g0544(n557, n266, new_n820);
not_13 g0545(n1422, new_n821);
and_7  g0546(new_n808, new_n821, new_n822);
and_7  g0547(new_n822, new_n642, new_n823_1);
and_7  g0548(new_n816, n1422, new_n824_1);
or_2   g0549(new_n824_1, new_n823_1, new_n825);
or_2   g0550(new_n825, new_n820, new_n826);
xor_5  g0551(new_n826, new_n819, new_n827);
and_7  g0552(new_n827, new_n813_1, new_n828);
nor_6  g0553(new_n827, new_n813_1, new_n829);
or_2   g0554(new_n829, new_n828, new_n830);
and_7  g0555(new_n627_1, n649, new_n831);
nor_6  g0556(new_n812, new_n796, new_n832);
nor_6  g0557(new_n832, new_n813_1, new_n833);
nor_6  g0558(new_n833, new_n831, new_n834);
and_7  g0559(new_n833, new_n831, new_n835);
or_2   g0560(new_n835, new_n834, new_n836_1);
not_13 g0561(n649, new_n837);
or_2   g0562(new_n638_1, new_n628, new_n838);
or_2   g0563(new_n838, new_n837, new_n839_1);
or_2   g0564(new_n627_1, n649, new_n840);
and_7  g0565(new_n840, new_n839_1, new_n841);
nor_6  g0566(new_n795, new_n712_1, new_n842);
nor_6  g0567(new_n842, new_n796, new_n843);
nor_6  g0568(new_n843, new_n841, new_n844);
and_7  g0569(new_n843, new_n841, new_n845);
or_2   g0570(new_n845, new_n844, new_n846_1);
or_2   g0571(new_n714, new_n640, new_n847);
nor_6  g0572(new_n785, new_n722, new_n848);
or_2   g0573(new_n848, new_n717, new_n849);
and_7  g0574(new_n849, new_n847, new_n850);
nor_6  g0575(new_n850, new_n846_1, new_n851);
nor_6  g0576(new_n851, new_n844, new_n852);
nor_6  g0577(new_n852, new_n836_1, new_n853);
or_2   g0578(new_n853, new_n834, new_n854);
or_2   g0579(new_n854, new_n830, new_n855);
nor_6  g0580(new_n829, new_n828, new_n856);
or_2   g0581(new_n833, new_n831, new_n857);
or_2   g0582(new_n852, new_n836_1, new_n858_1);
and_7  g0583(new_n858_1, new_n857, new_n859);
or_2   g0584(new_n859, new_n856, new_n860);
and_7  g0585(new_n860, new_n855, n67);
not_13 g0586(n469, new_n862_1);
xor_5  g0587(n1643, new_n862_1, new_n863);
not_13 g0588(n927, new_n864);
and_7  g0589(new_n864, new_n545, new_n865_1);
not_13 g0590(new_n865_1, new_n866);
xor_5  g0591(n927, new_n545, new_n867_1);
not_13 g0592(n655, new_n868);
and_7  g0593(new_n868, new_n285, new_n869);
not_13 g0594(new_n869, new_n870_1);
xor_5  g0595(n655, new_n285, new_n871);
or_2   g0596(n952, n653, new_n872);
and_7  g0597(n1764, n1145, new_n873);
not_13 g0598(n653, new_n874);
xor_5  g0599(n952, new_n874, new_n875);
or_2   g0600(new_n875, new_n873, new_n876);
and_7  g0601(new_n876, new_n872, new_n877);
or_2   g0602(new_n877, new_n871, new_n878);
and_7  g0603(new_n878, new_n870_1, new_n879);
or_2   g0604(new_n879, new_n867_1, new_n880);
and_7  g0605(new_n880, new_n866, new_n881);
and_7  g0606(new_n881, new_n863, new_n882_1);
not_13 g0607(new_n863, new_n883_1);
and_7  g0608(n927, n555, new_n884);
not_13 g0609(new_n884, new_n885);
and_7  g0610(new_n885, new_n866, new_n886);
nor_6  g0611(new_n877, new_n871, new_n887);
or_2   g0612(new_n887, new_n869, new_n888_1);
and_7  g0613(new_n888_1, new_n886, new_n889);
or_2   g0614(new_n889, new_n865_1, new_n890);
and_7  g0615(new_n890, new_n883_1, new_n891_1);
or_2   g0616(new_n891_1, new_n882_1, new_n892_1);
and_7  g0617(new_n892_1, new_n400, new_n893);
nor_6  g0618(new_n892_1, new_n400, new_n894);
nor_6  g0619(new_n894, new_n893, new_n895);
and_7  g0620(new_n879, new_n867_1, new_n896);
or_2   g0621(new_n896, new_n889, new_n897);
nor_6  g0622(new_n897, new_n405, new_n898);
and_7  g0623(new_n897, new_n405, new_n899);
nor_6  g0624(new_n899, new_n898, new_n900);
not_13 g0625(new_n873, new_n901);
and_7  g0626(n952, n653, new_n902_1);
not_13 g0627(new_n902_1, new_n903);
and_7  g0628(new_n903, new_n872, new_n904);
or_2   g0629(new_n904, new_n901, new_n905_1);
xor_5  g0630(n1764, new_n420, new_n906_1);
or_2   g0631(new_n906_1, new_n422, new_n907);
and_7  g0632(new_n907, new_n876, new_n908);
and_7  g0633(new_n908, new_n905_1, new_n909);
xor_5  g0634(n1764, n1145, new_n910);
and_7  g0635(new_n910, new_n414_1, new_n911);
and_7  g0636(new_n911, new_n904, new_n912_1);
nor_6  g0637(new_n912_1, new_n909, new_n913);
and_7  g0638(new_n913, new_n431, new_n914);
nor_6  g0639(new_n914, new_n909, new_n915);
and_7  g0640(new_n877, new_n871, new_n916);
or_2   g0641(new_n916, new_n887, new_n917);
and_7  g0642(new_n917, new_n915, new_n918);
nor_6  g0643(new_n917, new_n915, new_n919);
nor_6  g0644(new_n919, new_n918, new_n920);
and_7  g0645(new_n920, new_n441, new_n921);
nor_6  g0646(new_n921, new_n918, new_n922);
and_7  g0647(new_n922, new_n900, new_n923);
nor_6  g0648(new_n923, new_n898, new_n924);
xor_5  g0649(new_n924, new_n895, n74);
and_7  g0650(new_n570, new_n511, new_n926);
or_2   g0651(new_n496, n1642, new_n927_1);
xor_5  g0652(new_n927_1, new_n800, new_n928);
and_7  g0653(new_n928, n1381, new_n929);
and_7  g0654(new_n502, new_n805, new_n930);
not_13 g0655(new_n502, new_n931_1);
and_7  g0656(new_n931_1, n1263, new_n932);
or_2   g0657(new_n932, new_n503, new_n933);
or_2   g0658(new_n933, new_n930, new_n934);
and_7  g0659(new_n456, n171, new_n935_1);
or_2   g0660(new_n935_1, new_n457_1, new_n936);
and_7  g0661(new_n936, new_n934, new_n937);
or_2   g0662(new_n937, new_n929, new_n938);
and_7  g0663(new_n938, new_n926, new_n939);
not_13 g0664(n557, new_n940);
not_13 g0665(new_n927_1, new_n941);
and_7  g0666(new_n941, new_n800, new_n942_1);
or_2   g0667(new_n942_1, new_n940, new_n943);
and_7  g0668(new_n942_1, new_n940, new_n944_1);
not_13 g0669(new_n944_1, new_n945);
and_7  g0670(new_n945, n1381, new_n946);
and_7  g0671(new_n946, new_n943, new_n947);
and_7  g0672(n557, new_n503, new_n948);
xor_5  g0673(new_n930, n1422, new_n949);
and_7  g0674(new_n949, n402, new_n950);
nor_6  g0675(new_n950, new_n948, new_n951);
and_7  g0676(new_n951, new_n456, new_n952_1);
nor_6  g0677(new_n952_1, new_n947, new_n953_1);
and_7  g0678(new_n953_1, new_n939, new_n954);
nor_6  g0679(new_n953_1, new_n939, new_n955);
nor_6  g0680(new_n955, new_n954, n156);
nor_6  g0681(new_n938, new_n926, new_n957);
nor_6  g0682(new_n957, new_n939, n1149);
and_7  g0683(n1149, new_n600_1, new_n959);
nor_6  g0684(new_n959, n156, new_n960);
and_7  g0685(new_n959, new_n953_1, new_n961_1);
nor_6  g0686(new_n961_1, new_n960, n106);
xor_5  g0687(new_n568, new_n559_1, n1385);
nor_6  g0688(n1385, new_n596, new_n964);
nor_6  g0689(new_n964, new_n597, n126);
not_13 g0690(new_n746, new_n966);
or_2   g0691(new_n776, new_n748_1, new_n967);
and_7  g0692(new_n967, new_n966, new_n968_1);
xor_5  g0693(new_n968_1, new_n741, n135);
and_7  g0694(new_n652, new_n277_1, new_n970);
xor_5  g0695(new_n652, n1643, new_n971);
or_2   g0696(new_n671, n555, new_n972);
and_7  g0697(new_n647_1, new_n285, new_n973);
not_13 g0698(new_n973, new_n974_1);
xor_5  g0699(new_n647_1, n353, new_n975);
or_2   g0700(new_n681, n952, new_n976);
and_7  g0701(new_n685, n1145, new_n977);
xor_5  g0702(new_n681, new_n539, new_n978);
or_2   g0703(new_n978, new_n977, new_n979_1);
and_7  g0704(new_n979_1, new_n976, new_n980_1);
or_2   g0705(new_n980_1, new_n975, new_n981);
and_7  g0706(new_n981, new_n974_1, new_n982);
xor_5  g0707(new_n644, n555, new_n983);
or_2   g0708(new_n983, new_n982, new_n984);
and_7  g0709(new_n984, new_n972, new_n985);
nor_6  g0710(new_n985, new_n971, new_n986);
or_2   g0711(new_n986, new_n970, new_n987);
or_2   g0712(new_n987, new_n656, new_n988);
xor_5  g0713(new_n988, new_n702, n145);
xor_5  g0714(new_n413, n347, n174);
and_7  g0715(new_n395, n1597, new_n991_1);
and_7  g0716(new_n392, new_n391_1, new_n992);
or_2   g0717(new_n992, new_n302, new_n993);
and_7  g0718(new_n993, new_n374, new_n994);
or_2   g0719(new_n994, new_n991_1, new_n995);
and_7  g0720(new_n402_1, n682, new_n996);
nor_6  g0721(new_n401_1, new_n300, new_n997);
or_2   g0722(new_n997, new_n334, new_n998);
or_2   g0723(new_n402_1, n682, new_n999);
and_7  g0724(new_n999, new_n998, new_n1000_1);
and_7  g0725(new_n407, n1435, new_n1001);
nor_6  g0726(new_n406, new_n298, new_n1002);
and_7  g0727(new_n1002, new_n316, new_n1003);
or_2   g0728(new_n1003, new_n1001, new_n1004);
and_7  g0729(new_n412, n66, new_n1005_1);
nor_6  g0730(new_n412, n66, new_n1006);
nor_6  g0731(new_n1006, new_n1005_1, new_n1007);
or_2   g0732(new_n418, n968, new_n1008);
and_7  g0733(new_n413, n347, new_n1009);
nor_6  g0734(new_n418, n968, new_n1010);
and_7  g0735(new_n418, n968, new_n1011);
or_2   g0736(new_n1011, new_n1010, new_n1012_1);
or_2   g0737(new_n1012_1, new_n1009, new_n1013);
and_7  g0738(new_n1013, new_n1008, new_n1014);
and_7  g0739(new_n1014, new_n1007, new_n1015_1);
nor_6  g0740(new_n1015_1, new_n1005_1, new_n1016_1);
nor_6  g0741(new_n1016_1, new_n1004, new_n1017);
or_2   g0742(new_n1017, new_n1001, new_n1018);
and_7  g0743(new_n1018, new_n1000_1, new_n1019);
nor_6  g0744(new_n1019, new_n996, new_n1020);
nor_6  g0745(new_n1020, new_n995, new_n1021);
and_7  g0746(new_n1020, new_n995, new_n1022);
nor_6  g0747(new_n1022, new_n1021, new_n1023);
nor_6  g0748(new_n1018, new_n1000_1, new_n1024);
nor_6  g0749(new_n1024, new_n1019, new_n1025_1);
nor_6  g0750(new_n1014, new_n1007, new_n1026);
nor_6  g0751(new_n1026, new_n1015_1, n1426);
and_7  g0752(new_n1016_1, new_n1004, new_n1028);
nor_6  g0753(new_n1028, new_n1017, new_n1029);
or_2   g0754(new_n1029, n1426, new_n1030_1);
nor_6  g0755(new_n1030_1, new_n1025_1, new_n1031);
xor_5  g0756(new_n1031, new_n1023, n181);
xor_5  g0757(new_n433_1, new_n412, new_n1033);
xor_5  g0758(new_n1033, new_n441, n208);
not_13 g0759(n213, new_n1035);
and_7  g0760(new_n647_1, new_n1035, new_n1036);
xor_5  g0761(new_n647_1, n213, new_n1037);
not_13 g0762(n1743, new_n1038);
and_7  g0763(new_n689, new_n1038, new_n1039);
not_13 g0764(n600, new_n1040);
not_13 g0765(new_n683_1, new_n1041);
or_2   g0766(new_n469_1, n266, new_n1042);
and_7  g0767(new_n1042, new_n1041, new_n1043);
or_2   g0768(new_n1043, new_n1040, new_n1044);
xor_5  g0769(new_n681, n1743, new_n1045);
and_7  g0770(new_n1045, new_n1044, new_n1046);
nor_6  g0771(new_n1046, new_n1039, new_n1047);
nor_6  g0772(new_n1047, new_n1037, new_n1048);
or_2   g0773(new_n1048, new_n1036, new_n1049);
or_2   g0774(new_n1049, new_n644, new_n1050);
or_2   g0775(new_n1050, new_n652, new_n1051);
or_2   g0776(new_n1051, new_n656, new_n1052);
nor_6  g0777(new_n1048, new_n1036, new_n1053);
and_7  g0778(new_n1053, new_n671, new_n1054);
and_7  g0779(new_n1054, new_n669, new_n1055);
or_2   g0780(new_n1055, new_n666, new_n1056);
and_7  g0781(new_n1056, new_n1052, new_n1057);
not_13 g0782(n17, new_n1058);
not_13 g0783(n424, new_n1059);
and_7  g0784(new_n277_1, new_n1059, new_n1060);
not_13 g0785(new_n1060, new_n1061);
and_7  g0786(n1643, n424, new_n1062_1);
not_13 g0787(new_n1062_1, new_n1063);
and_7  g0788(new_n1063, new_n1061, new_n1064);
not_13 g0789(n1363, new_n1065);
and_7  g0790(new_n1065, new_n545, new_n1066);
xor_5  g0791(n1363, n555, new_n1067_1);
not_13 g0792(n498, new_n1068_1);
and_7  g0793(new_n1068_1, new_n285, new_n1069);
xor_5  g0794(n498, new_n285, new_n1070);
not_13 g0795(n414, new_n1071);
and_7  g0796(new_n539, new_n1071, new_n1072);
and_7  g0797(n1145, n183, new_n1073);
not_13 g0798(new_n1073, new_n1074);
xor_5  g0799(n952, n414, new_n1075);
and_7  g0800(new_n1075, new_n1074, new_n1076);
nor_6  g0801(new_n1076, new_n1072, new_n1077);
nor_6  g0802(new_n1077, new_n1070, new_n1078);
or_2   g0803(new_n1078, new_n1069, new_n1079);
and_7  g0804(new_n1079, new_n1067_1, new_n1080);
or_2   g0805(new_n1080, new_n1066, new_n1081);
and_7  g0806(new_n1081, new_n1064, new_n1082);
or_2   g0807(new_n1082, new_n1060, new_n1083);
or_2   g0808(new_n1083, new_n1058, new_n1084);
xor_5  g0809(n1643, new_n1059, new_n1085);
nor_6  g0810(new_n1080, new_n1066, new_n1086);
or_2   g0811(new_n1086, new_n1085, new_n1087);
and_7  g0812(new_n1087, new_n1061, new_n1088);
or_2   g0813(new_n1088, n17, new_n1089);
and_7  g0814(new_n1089, new_n1084, new_n1090);
and_7  g0815(new_n1090, new_n1057, new_n1091);
nor_6  g0816(new_n1090, new_n1057, new_n1092);
or_2   g0817(new_n1092, new_n1091, new_n1093);
and_7  g0818(new_n1050, new_n652, new_n1094);
nor_6  g0819(new_n1094, new_n1055, new_n1095);
and_7  g0820(new_n1086, new_n1085, new_n1096);
or_2   g0821(new_n1096, new_n1082, new_n1097);
or_2   g0822(new_n1097, new_n1095, new_n1098);
and_7  g0823(new_n1049, new_n644, new_n1099);
nor_6  g0824(new_n1099, new_n1054, new_n1100);
nor_6  g0825(new_n1079, new_n1067_1, new_n1101);
or_2   g0826(new_n1101, new_n1080, new_n1102);
nor_6  g0827(new_n1102, new_n1100, new_n1103_1);
and_7  g0828(new_n1102, new_n1100, new_n1104);
or_2   g0829(new_n1104, new_n1103_1, new_n1105);
and_7  g0830(new_n1047, new_n1037, new_n1106);
nor_6  g0831(new_n1106, new_n1048, new_n1107);
and_7  g0832(new_n1077, new_n1070, new_n1108);
nor_6  g0833(new_n1108, new_n1078, new_n1109);
and_7  g0834(new_n1109, new_n1107, new_n1110);
or_2   g0835(new_n1075, new_n1074, new_n1111);
xor_5  g0836(n1145, n183, new_n1112);
xor_5  g0837(new_n685, n600, new_n1113_1);
and_7  g0838(new_n1113_1, new_n1112, new_n1114);
nor_6  g0839(new_n1114, new_n1076, new_n1115);
and_7  g0840(new_n1115, new_n1111, new_n1116);
not_13 g0841(new_n1044, new_n1117);
xor_5  g0842(new_n681, new_n1038, new_n1118);
or_2   g0843(new_n1118, new_n1117, new_n1119_1);
or_2   g0844(new_n1045, new_n1044, new_n1120);
and_7  g0845(new_n1120, new_n1119_1, new_n1121);
and_7  g0846(new_n1114, new_n1075, new_n1122);
nor_6  g0847(new_n1122, new_n1116, new_n1123);
and_7  g0848(new_n1123, new_n1121, new_n1124);
or_2   g0849(new_n1124, new_n1116, new_n1125);
nor_6  g0850(new_n1109, new_n1107, new_n1126);
nor_6  g0851(new_n1126, new_n1110, new_n1127);
and_7  g0852(new_n1127, new_n1125, new_n1128);
nor_6  g0853(new_n1128, new_n1110, new_n1129);
nor_6  g0854(new_n1129, new_n1105, new_n1130);
nor_6  g0855(new_n1130, new_n1103_1, new_n1131);
nor_6  g0856(new_n1097, new_n1095, new_n1132);
and_7  g0857(new_n1097, new_n1095, new_n1133);
or_2   g0858(new_n1133, new_n1132, new_n1134);
or_2   g0859(new_n1134, new_n1131, new_n1135_1);
and_7  g0860(new_n1135_1, new_n1098, new_n1136);
nor_6  g0861(new_n1136, new_n1093, new_n1137);
and_7  g0862(new_n1136, new_n1093, new_n1138_1);
or_2   g0863(new_n1138_1, new_n1137, n216);
not_13 g0864(new_n1125, new_n1140_1);
xor_5  g0865(new_n1127, new_n1140_1, n218);
and_7  g0866(new_n852, new_n836_1, new_n1142_1);
or_2   g0867(new_n1142_1, new_n853, n231);
not_13 g0868(n1747, new_n1144);
not_13 g0869(n738, new_n1145_1);
not_13 g0870(n961, new_n1146);
or_2   g0871(new_n1084, new_n1146, new_n1147);
or_2   g0872(new_n1147, new_n1145_1, new_n1148);
or_2   g0873(new_n1148, new_n1144, new_n1149_1);
and_7  g0874(new_n1088, n17, new_n1150);
and_7  g0875(new_n1150, n961, new_n1151);
and_7  g0876(new_n1151, n738, new_n1152);
or_2   g0877(new_n1152, n1747, new_n1153);
and_7  g0878(new_n1153, new_n1149_1, new_n1154);
or_2   g0879(new_n1052, new_n702, new_n1155);
or_2   g0880(new_n1155, new_n788_1, new_n1156);
or_2   g0881(new_n1156, new_n798, new_n1157);
and_7  g0882(new_n1055, new_n666, new_n1158);
and_7  g0883(new_n1158, new_n662, new_n1159);
and_7  g0884(new_n1159, new_n710, new_n1160);
or_2   g0885(new_n1160, new_n794, new_n1161_1);
and_7  g0886(new_n1161_1, new_n1157, new_n1162_1);
and_7  g0887(new_n1162_1, new_n1154, new_n1163);
nor_6  g0888(new_n1162_1, new_n1154, new_n1164);
or_2   g0889(new_n1164, new_n1163, new_n1165);
or_2   g0890(new_n1151, n738, new_n1166);
and_7  g0891(new_n1166, new_n1148, new_n1167);
or_2   g0892(new_n1159, new_n710, new_n1168);
and_7  g0893(new_n1168, new_n1156, new_n1169);
or_2   g0894(new_n1169, new_n1167, new_n1170);
nor_6  g0895(new_n1169, new_n1167, new_n1171);
and_7  g0896(new_n1169, new_n1167, new_n1172_1);
or_2   g0897(new_n1172_1, new_n1171, new_n1173);
or_2   g0898(new_n1150, n961, new_n1174);
and_7  g0899(new_n1174, new_n1147, new_n1175_1);
or_2   g0900(new_n1158, new_n662, new_n1176);
and_7  g0901(new_n1176, new_n1155, new_n1177);
nor_6  g0902(new_n1177, new_n1175_1, new_n1178);
and_7  g0903(new_n1177, new_n1175_1, new_n1179);
nor_6  g0904(new_n1179, new_n1178, new_n1180);
or_2   g0905(new_n1137, new_n1092, new_n1181);
and_7  g0906(new_n1181, new_n1180, new_n1182);
nor_6  g0907(new_n1182, new_n1178, new_n1183_1);
or_2   g0908(new_n1183_1, new_n1173, new_n1184);
and_7  g0909(new_n1184, new_n1170, new_n1185);
nor_6  g0910(new_n1185, new_n1165, new_n1186);
and_7  g0911(new_n1185, new_n1165, new_n1187);
or_2   g0912(new_n1187, new_n1186, n238);
and_7  g0913(new_n303_1, n1537, new_n1189);
and_7  g0914(new_n1189, n675, new_n1190);
xor_5  g0915(new_n1190, n1263, new_n1191_1);
not_13 g0916(n675, new_n1192);
not_13 g0917(n1537, new_n1193);
not_13 g0918(n433, new_n1194_1);
or_2   g0919(new_n393, new_n1194_1, new_n1195);
or_2   g0920(new_n1195, new_n1193, new_n1196);
or_2   g0921(new_n1196, new_n1192, new_n1197);
or_2   g0922(new_n1189, n675, new_n1198);
and_7  g0923(new_n1198, new_n1197, new_n1199_1);
and_7  g0924(new_n1199_1, n379, new_n1200);
nor_6  g0925(new_n1199_1, n379, new_n1201_1);
or_2   g0926(new_n1201_1, new_n1200, new_n1202_1);
and_7  g0927(new_n1195, new_n1193, new_n1203);
nor_6  g0928(new_n1203, new_n1189, new_n1204);
and_7  g0929(new_n1204, n1527, new_n1205);
nor_6  g0930(new_n1204, n1527, new_n1206);
or_2   g0931(new_n1206, new_n1205, new_n1207);
or_2   g0932(new_n304, new_n303_1, new_n1208);
or_2   g0933(new_n1208, new_n373, new_n1209);
nor_6  g0934(new_n1021, new_n991_1, new_n1210);
and_7  g0935(new_n305, n46, new_n1211);
and_7  g0936(new_n1208, new_n373, new_n1212);
or_2   g0937(new_n1212, new_n1211, new_n1213);
or_2   g0938(new_n1213, new_n1210, new_n1214);
and_7  g0939(new_n1214, new_n1209, new_n1215);
nor_6  g0940(new_n1215, new_n1207, new_n1216);
nor_6  g0941(new_n1216, new_n1205, new_n1217);
nor_6  g0942(new_n1217, new_n1202_1, new_n1218);
nor_6  g0943(new_n1218, new_n1200, new_n1219);
and_7  g0944(new_n1219, new_n1191_1, new_n1220);
nor_6  g0945(new_n1219, new_n1191_1, new_n1221);
or_2   g0946(new_n1221, new_n1220, new_n1222_1);
and_7  g0947(new_n1217, new_n1202_1, new_n1223);
nor_6  g0948(new_n1223, new_n1218, new_n1224);
and_7  g0949(new_n1215, new_n1207, new_n1225);
nor_6  g0950(new_n1225, new_n1216, new_n1226);
or_2   g0951(new_n1030_1, new_n1025_1, new_n1227);
or_2   g0952(new_n1227, new_n1023, new_n1228);
or_2   g0953(new_n1021, new_n991_1, new_n1229);
xor_5  g0954(new_n305, n46, new_n1230);
and_7  g0955(new_n1230, new_n1229, new_n1231);
and_7  g0956(new_n1213, new_n1210, new_n1232);
nor_6  g0957(new_n1232, new_n1231, new_n1233);
or_2   g0958(new_n1233, new_n1228, new_n1234_1);
or_2   g0959(new_n1234_1, new_n1226, new_n1235_1);
or_2   g0960(new_n1235_1, new_n1224, new_n1236);
and_7  g0961(new_n1236, new_n1222_1, new_n1237_1);
nor_6  g0962(new_n1221, new_n1220, new_n1238);
nor_6  g0963(new_n1235_1, new_n1224, new_n1239);
and_7  g0964(new_n1239, new_n1238, new_n1240);
or_2   g0965(new_n1240, new_n1237_1, n270);
xor_5  g0966(new_n736, new_n402_1, new_n1242);
and_7  g0967(new_n743, new_n407, new_n1243);
nor_6  g0968(new_n743, new_n407, new_n1244);
and_7  g0969(new_n750, new_n412, new_n1245);
or_2   g0970(new_n750, new_n412, new_n1246);
and_7  g0971(new_n761_1, new_n413, new_n1247);
nor_6  g0972(new_n1247, new_n418, new_n1248);
and_7  g0973(new_n1247, new_n417, new_n1249_1);
nor_6  g0974(new_n1249_1, new_n1248, new_n1250);
and_7  g0975(new_n1250, new_n768, new_n1251);
nor_6  g0976(new_n1251, new_n1248, new_n1252);
and_7  g0977(new_n1252, new_n1246, new_n1253);
nor_6  g0978(new_n1253, new_n1245, new_n1254);
nor_6  g0979(new_n1254, new_n1244, new_n1255_1);
or_2   g0980(new_n1255_1, new_n1243, new_n1256);
xor_5  g0981(new_n1256, new_n1242, n276);
xor_5  g0982(new_n910, new_n414_1, n290);
not_13 g0983(new_n1009, new_n1259);
xor_5  g0984(new_n1012_1, new_n1259, n292);
and_7  g0985(new_n1152, n1747, new_n1261);
or_2   g0986(new_n1157, new_n818, new_n1262);
and_7  g0987(new_n1160, new_n794, new_n1263_1);
or_2   g0988(new_n1263_1, new_n811, new_n1264);
and_7  g0989(new_n1264, new_n1262, new_n1265);
nor_6  g0990(new_n1265, new_n1261, new_n1266);
and_7  g0991(new_n1265, new_n1261, new_n1267);
nor_6  g0992(new_n1267, new_n1266, new_n1268);
or_2   g0993(new_n1186, new_n1164, new_n1269);
and_7  g0994(new_n1269, new_n1268, new_n1270);
or_2   g0995(new_n1270, new_n1266, new_n1271);
and_7  g0996(new_n1262, new_n823_1, new_n1272);
and_7  g0997(new_n1272, new_n1271, n299);
not_13 g0998(n1341, new_n1274);
or_2   g0999(new_n532_1, new_n1274, new_n1275);
xor_5  g1000(new_n532_1, n1341, new_n1276);
and_7  g1001(new_n461, n69, new_n1277_1);
nor_6  g1002(new_n476_1, new_n1277_1, new_n1278_1);
or_2   g1003(new_n1278_1, new_n1276, new_n1279);
and_7  g1004(new_n1279, new_n1275, new_n1280);
nor_6  g1005(new_n1280, new_n527, new_n1281);
and_7  g1006(new_n1281, new_n558, new_n1282);
and_7  g1007(new_n1282, new_n568, new_n1283_1);
or_2   g1008(new_n1280, new_n527, new_n1284);
or_2   g1009(new_n1284, new_n557_1, new_n1285);
and_7  g1010(new_n1285, new_n567, new_n1286);
nor_6  g1011(new_n1286, new_n1283_1, new_n1287);
not_13 g1012(n761, new_n1288);
and_7  g1013(new_n277_1, new_n1288, new_n1289);
not_13 g1014(new_n1289, new_n1290);
xor_5  g1015(n1643, new_n1288, new_n1291);
not_13 g1016(n1172, new_n1292);
and_7  g1017(new_n1292, new_n545, new_n1293);
xor_5  g1018(n1172, n555, new_n1294);
not_13 g1019(n695, new_n1295);
and_7  g1020(new_n1295, new_n285, new_n1296_1);
xor_5  g1021(n695, new_n285, new_n1297);
not_13 g1022(n1296, new_n1298);
and_7  g1023(new_n1298, new_n539, new_n1299);
and_7  g1024(n1145, n1062, new_n1300);
not_13 g1025(new_n1300, new_n1301);
xor_5  g1026(n1296, n952, new_n1302);
and_7  g1027(new_n1302, new_n1301, new_n1303);
nor_6  g1028(new_n1303, new_n1299, new_n1304);
nor_6  g1029(new_n1304, new_n1297, new_n1305_1);
or_2   g1030(new_n1305_1, new_n1296_1, new_n1306);
and_7  g1031(new_n1306, new_n1294, new_n1307);
nor_6  g1032(new_n1307, new_n1293, new_n1308);
or_2   g1033(new_n1308, new_n1291, new_n1309);
and_7  g1034(new_n1309, new_n1290, new_n1310);
and_7  g1035(new_n1310, n862, new_n1311);
and_7  g1036(new_n1311, n1222, new_n1312);
not_13 g1037(n1222, new_n1313);
not_13 g1038(n862, new_n1314);
and_7  g1039(n1643, n761, new_n1315_1);
not_13 g1040(new_n1315_1, new_n1316);
and_7  g1041(new_n1316, new_n1290, new_n1317);
or_2   g1042(new_n1307, new_n1293, new_n1318);
and_7  g1043(new_n1318, new_n1317, new_n1319);
or_2   g1044(new_n1319, new_n1289, new_n1320);
or_2   g1045(new_n1320, new_n1314, new_n1321_1);
and_7  g1046(new_n1321_1, new_n1313, new_n1322);
nor_6  g1047(new_n1322, new_n1312, new_n1323);
and_7  g1048(new_n1323, new_n1287, new_n1324);
nor_6  g1049(new_n1323, new_n1287, new_n1325);
or_2   g1050(new_n1325, new_n1324, new_n1326);
and_7  g1051(new_n1284, new_n557_1, new_n1327);
or_2   g1052(new_n1327, new_n1282, new_n1328);
and_7  g1053(new_n1320, new_n1314, new_n1329);
or_2   g1054(new_n1329, new_n1311, new_n1330_1);
and_7  g1055(new_n1330_1, new_n1328, new_n1331);
or_2   g1056(new_n1281, new_n558, new_n1332_1);
and_7  g1057(new_n1332_1, new_n1285, new_n1333);
or_2   g1058(new_n1310, n862, new_n1334);
and_7  g1059(new_n1334, new_n1321_1, new_n1335);
and_7  g1060(new_n1335, new_n1333, new_n1336);
nor_6  g1061(new_n1336, new_n1331, new_n1337);
and_7  g1062(new_n1280, new_n527, new_n1338_1);
nor_6  g1063(new_n1338_1, new_n1281, new_n1339);
and_7  g1064(new_n1308, new_n1291, new_n1340_1);
or_2   g1065(new_n1340_1, new_n1319, new_n1341_1);
nor_6  g1066(new_n1341_1, new_n1339, new_n1342);
and_7  g1067(new_n1341_1, new_n1339, new_n1343);
or_2   g1068(new_n1343, new_n1342, new_n1344);
xor_5  g1069(new_n532_1, new_n1274, new_n1345);
or_2   g1070(new_n476_1, new_n1277_1, new_n1346);
or_2   g1071(new_n1346, new_n1345, new_n1347_1);
and_7  g1072(new_n1347_1, new_n1279, new_n1348_1);
nor_6  g1073(new_n1306, new_n1294, new_n1349_1);
or_2   g1074(new_n1349_1, new_n1307, new_n1350);
nor_6  g1075(new_n1350, new_n1348_1, new_n1351_1);
and_7  g1076(new_n1350, new_n1348_1, new_n1352);
nor_6  g1077(new_n1352, new_n1351_1, new_n1353);
and_7  g1078(new_n1304, new_n1297, new_n1354);
or_2   g1079(new_n1354, new_n1305_1, new_n1355);
nor_6  g1080(new_n1355, new_n478, new_n1356);
and_7  g1081(new_n1355, new_n478, new_n1357);
or_2   g1082(new_n1357, new_n1356, new_n1358);
or_2   g1083(new_n1302, new_n1301, new_n1359);
xor_5  g1084(n1145, n1062, new_n1360);
and_7  g1085(new_n1360, new_n482_1, new_n1361);
nor_6  g1086(new_n1361, new_n1303, new_n1362);
and_7  g1087(new_n1362, new_n1359, new_n1363_1);
and_7  g1088(new_n1361, new_n1302, new_n1364);
nor_6  g1089(new_n1364, new_n1363_1, new_n1365);
and_7  g1090(new_n1365, new_n486, new_n1366);
nor_6  g1091(new_n1366, new_n1363_1, new_n1367);
nor_6  g1092(new_n1367, new_n1358, new_n1368);
or_2   g1093(new_n1368, new_n1356, new_n1369_1);
and_7  g1094(new_n1369_1, new_n1353, new_n1370);
nor_6  g1095(new_n1370, new_n1351_1, new_n1371);
nor_6  g1096(new_n1371, new_n1344, new_n1372);
or_2   g1097(new_n1372, new_n1342, new_n1373);
and_7  g1098(new_n1373, new_n1337, new_n1374);
nor_6  g1099(new_n1374, new_n1331, new_n1375);
and_7  g1100(new_n1375, new_n1326, new_n1376);
nor_6  g1101(new_n1375, new_n1326, new_n1377);
or_2   g1102(new_n1377, new_n1376, n317);
xor_5  g1103(new_n1360, new_n482_1, n372);
not_13 g1104(new_n922, new_n1380);
xor_5  g1105(new_n1380, new_n900, n378);
not_13 g1106(new_n826, new_n1382);
or_2   g1107(new_n988, new_n702, new_n1383_1);
or_2   g1108(new_n1383_1, new_n788_1, new_n1384);
or_2   g1109(new_n1384, new_n798, new_n1385_1);
or_2   g1110(new_n1385_1, new_n818, new_n1386);
or_2   g1111(new_n1386, new_n1382, new_n1387);
or_2   g1112(new_n1387, new_n823_1, new_n1388);
not_13 g1113(new_n823_1, new_n1389);
not_13 g1114(new_n970, new_n1390);
or_2   g1115(new_n985, new_n971, new_n1391);
and_7  g1116(new_n1391, new_n1390, new_n1392);
and_7  g1117(new_n1392, new_n666, new_n1393_1);
and_7  g1118(new_n1393_1, new_n662, new_n1394);
and_7  g1119(new_n1394, new_n710, new_n1395);
and_7  g1120(new_n1395, new_n794, new_n1396);
and_7  g1121(new_n1396, new_n811, new_n1397);
or_2   g1122(new_n1397, new_n1389, new_n1398);
and_7  g1123(new_n1398, new_n1388, new_n1399_1);
and_7  g1124(new_n1385_1, new_n818, new_n1400);
nor_6  g1125(new_n1400, new_n1397, n1249);
and_7  g1126(new_n1383_1, new_n788_1, new_n1402);
nor_6  g1127(new_n1402, new_n1395, n1119);
not_13 g1128(new_n977, new_n1404);
or_2   g1129(new_n685, n1145, new_n1405);
and_7  g1130(new_n1405, new_n1404, n647);
xor_5  g1131(new_n978, new_n1404, n646);
or_2   g1132(n646, n647, new_n1408);
nor_6  g1133(new_n980_1, new_n975, new_n1409);
and_7  g1134(new_n980_1, new_n975, new_n1410);
or_2   g1135(new_n1410, new_n1409, n1016);
nor_6  g1136(n1016, new_n1408, new_n1412);
or_2   g1137(new_n1409, new_n973, new_n1413);
not_13 g1138(new_n983, new_n1414);
or_2   g1139(new_n1414, new_n1413, new_n1415);
and_7  g1140(new_n1415, new_n984, new_n1416);
or_2   g1141(new_n1416, new_n1412, new_n1417);
and_7  g1142(new_n985, new_n971, new_n1418);
nor_6  g1143(new_n1418, new_n986, new_n1419);
nor_6  g1144(new_n1419, new_n1417, new_n1420);
and_7  g1145(new_n987, new_n656, new_n1421);
nor_6  g1146(new_n1421, new_n1393_1, n773);
and_7  g1147(n773, new_n1420, new_n1423);
and_7  g1148(new_n1423, new_n662, new_n1424);
and_7  g1149(new_n1424, n1119, new_n1425_1);
and_7  g1150(new_n1425_1, new_n794, new_n1426_1);
and_7  g1151(new_n1426_1, n1249, new_n1427);
and_7  g1152(new_n1427, new_n826, new_n1428);
nor_6  g1153(new_n1428, new_n1399_1, new_n1429);
and_7  g1154(new_n1428, new_n1399_1, new_n1430);
or_2   g1155(new_n1430, new_n1429, n387);
or_2   g1156(new_n1283_1, new_n523, new_n1432);
or_2   g1157(new_n1285, new_n567, new_n1433);
or_2   g1158(new_n1433, new_n572, new_n1434);
and_7  g1159(new_n1434, new_n1432, new_n1435_1);
not_13 g1160(n1757, new_n1436);
or_2   g1161(new_n1321_1, new_n1313, new_n1437);
or_2   g1162(new_n1437, new_n1436, new_n1438);
or_2   g1163(new_n1312, n1757, new_n1439);
and_7  g1164(new_n1439, new_n1438, new_n1440_1);
and_7  g1165(new_n1440_1, new_n1435_1, new_n1441);
nor_6  g1166(new_n1440_1, new_n1435_1, new_n1442);
nor_6  g1167(new_n1442, new_n1441, new_n1443);
or_2   g1168(new_n1323, new_n1287, new_n1444);
or_2   g1169(new_n1375, new_n1326, new_n1445);
and_7  g1170(new_n1445, new_n1444, new_n1446);
xor_5  g1171(new_n1446, new_n1443, n401);
xor_5  g1172(new_n920, new_n441, n423);
and_7  g1173(new_n1348_1, new_n407, new_n1449);
nor_6  g1174(new_n1348_1, new_n407, new_n1450);
nor_6  g1175(new_n1450, new_n1449, new_n1451);
not_13 g1176(new_n1451, new_n1452);
or_2   g1177(new_n492, new_n480, new_n1453_1);
xor_5  g1178(new_n1453_1, new_n1452, n426);
or_2   g1179(new_n1397, new_n826, new_n1455);
and_7  g1180(new_n1455, new_n1387, n493);
nor_6  g1181(n493, new_n1427, new_n1457_1);
nor_6  g1182(new_n1457_1, new_n1428, n429);
xor_5  g1183(n773, new_n1420, n432);
and_7  g1184(new_n1339, new_n402_1, new_n1460_1);
nor_6  g1185(new_n1339, new_n402_1, new_n1461_1);
or_2   g1186(new_n1461_1, new_n1460_1, new_n1462);
and_7  g1187(new_n1453_1, new_n1451, new_n1463_1);
nor_6  g1188(new_n1463_1, new_n1450, new_n1464);
nor_6  g1189(new_n1464, new_n1462, new_n1465);
and_7  g1190(new_n1464, new_n1462, new_n1466);
or_2   g1191(new_n1466, new_n1465, n452);
nor_6  g1192(new_n1233, new_n1228, new_n1468);
and_7  g1193(new_n1233, new_n1228, new_n1469);
or_2   g1194(new_n1469, new_n1468, n457);
nor_6  g1195(new_n1269, new_n1268, new_n1471);
or_2   g1196(new_n1471, new_n1270, n460);
xor_5  g1197(new_n761_1, new_n760, n476);
not_13 g1198(new_n443, new_n1474);
xor_5  g1199(new_n1474, new_n410, n482);
and_7  g1200(new_n1283_1, new_n523, new_n1476);
and_7  g1201(new_n1476, new_n511, new_n1477);
and_7  g1202(new_n1477, new_n938, new_n1478);
nor_6  g1203(new_n1477, new_n938, new_n1479);
nor_6  g1204(new_n1479, new_n1478, new_n1480);
and_7  g1205(new_n1480, new_n1190, new_n1481_1);
nor_6  g1206(new_n1480, new_n1190, new_n1482);
nor_6  g1207(new_n1482, new_n1481_1, new_n1483);
nor_6  g1208(new_n1476, new_n511, new_n1484);
nor_6  g1209(new_n1484, new_n1477, new_n1485);
nor_6  g1210(new_n1485, new_n1199_1, new_n1486);
and_7  g1211(new_n1485, new_n1199_1, new_n1487);
or_2   g1212(new_n1487, new_n1486, new_n1488);
nor_6  g1213(new_n1435_1, new_n1204, new_n1489);
and_7  g1214(new_n1435_1, new_n1204, new_n1490);
nor_6  g1215(new_n1490, new_n1489, new_n1491);
and_7  g1216(new_n1287, new_n305, new_n1492);
and_7  g1217(new_n1328, new_n993, new_n1493);
or_2   g1218(new_n1333, new_n395, new_n1494);
or_2   g1219(new_n1328, new_n993, new_n1495_1);
and_7  g1220(new_n1495_1, new_n1494, new_n1496);
or_2   g1221(new_n1465, new_n1461_1, new_n1497);
and_7  g1222(new_n1497, new_n1496, new_n1498_1);
nor_6  g1223(new_n1498_1, new_n1493, new_n1499);
nor_6  g1224(new_n1287, new_n305, new_n1500);
nor_6  g1225(new_n1500, new_n1492, new_n1501_1);
and_7  g1226(new_n1501_1, new_n1499, new_n1502_1);
nor_6  g1227(new_n1502_1, new_n1492, new_n1503);
and_7  g1228(new_n1503, new_n1491, new_n1504);
nor_6  g1229(new_n1504, new_n1489, new_n1505);
nor_6  g1230(new_n1505, new_n1488, new_n1506);
or_2   g1231(new_n1506, new_n1486, new_n1507_1);
and_7  g1232(new_n1507_1, new_n1483, new_n1508);
nor_6  g1233(new_n1507_1, new_n1483, new_n1509);
or_2   g1234(new_n1509, new_n1508, n510);
and_7  g1235(new_n1199_1, new_n1162_1, new_n1511);
nor_6  g1236(new_n1199_1, new_n1162_1, new_n1512);
nor_6  g1237(new_n1512, new_n1511, new_n1513);
nor_6  g1238(new_n1204, new_n1169, new_n1514);
and_7  g1239(new_n1204, new_n1169, new_n1515);
or_2   g1240(new_n1515, new_n1514, new_n1516);
or_2   g1241(new_n1177, new_n305, new_n1517);
nor_6  g1242(new_n1177, new_n305, new_n1518);
and_7  g1243(new_n1177, new_n305, new_n1519);
or_2   g1244(new_n1519, new_n1518, new_n1520);
nor_6  g1245(new_n1057, new_n395, new_n1521);
and_7  g1246(new_n1057, new_n395, new_n1522);
nor_6  g1247(new_n1522, new_n1521, new_n1523);
and_7  g1248(new_n1095, new_n402_1, new_n1524);
nor_6  g1249(new_n1100, new_n407, new_n1525_1);
and_7  g1250(new_n1100, new_n407, new_n1526);
or_2   g1251(new_n1526, new_n1525_1, new_n1527_1);
xor_5  g1252(new_n295, new_n288, new_n1528);
and_7  g1253(new_n1107, new_n1528, new_n1529);
nor_6  g1254(new_n1107, new_n1528, new_n1530_1);
nor_6  g1255(new_n1530_1, new_n1529, new_n1531);
and_7  g1256(new_n1113_1, new_n413, new_n1532);
nor_6  g1257(new_n1532, new_n418, new_n1533);
and_7  g1258(new_n1532, new_n417, new_n1534);
nor_6  g1259(new_n1534, new_n1533, new_n1535_1);
and_7  g1260(new_n1535_1, new_n1121, new_n1536);
or_2   g1261(new_n1536, new_n1533, new_n1537_1);
and_7  g1262(new_n1537_1, new_n1531, new_n1538);
nor_6  g1263(new_n1538, new_n1529, new_n1539);
nor_6  g1264(new_n1539, new_n1527_1, new_n1540);
nor_6  g1265(new_n1540, new_n1525_1, new_n1541);
nor_6  g1266(new_n1095, new_n402_1, new_n1542);
nor_6  g1267(new_n1542, new_n1524, new_n1543);
and_7  g1268(new_n1543, new_n1541, new_n1544_1);
nor_6  g1269(new_n1544_1, new_n1524, new_n1545);
and_7  g1270(new_n1545, new_n1523, new_n1546);
nor_6  g1271(new_n1546, new_n1521, new_n1547);
or_2   g1272(new_n1547, new_n1520, new_n1548);
and_7  g1273(new_n1548, new_n1517, new_n1549);
nor_6  g1274(new_n1549, new_n1516, new_n1550);
or_2   g1275(new_n1550, new_n1514, new_n1551);
and_7  g1276(new_n1551, new_n1513, new_n1552);
nor_6  g1277(new_n1551, new_n1513, new_n1553);
or_2   g1278(new_n1553, new_n1552, n517);
and_7  g1279(new_n1199_1, new_n843, new_n1555);
nor_6  g1280(new_n1199_1, new_n843, new_n1556_1);
or_2   g1281(new_n1556_1, new_n1555, new_n1557);
nor_6  g1282(new_n1204, new_n714, new_n1558);
and_7  g1283(new_n1204, new_n714, new_n1559);
or_2   g1284(new_n1559, new_n1558, new_n1560);
nor_6  g1285(new_n721, new_n305, new_n1561);
nor_6  g1286(new_n728, new_n395, new_n1562);
and_7  g1287(new_n728, new_n395, new_n1563);
nor_6  g1288(new_n1563, new_n1562, new_n1564);
and_7  g1289(new_n736, new_n402_1, new_n1565);
or_2   g1290(new_n736, new_n402_1, new_n1566);
and_7  g1291(new_n1256, new_n1566, new_n1567);
nor_6  g1292(new_n1567, new_n1565, new_n1568);
and_7  g1293(new_n1568, new_n1564, new_n1569);
nor_6  g1294(new_n1569, new_n1562, new_n1570);
and_7  g1295(new_n721, new_n305, new_n1571);
or_2   g1296(new_n1571, new_n1561, new_n1572);
nor_6  g1297(new_n1572, new_n1570, new_n1573);
nor_6  g1298(new_n1573, new_n1561, new_n1574);
nor_6  g1299(new_n1574, new_n1560, new_n1575);
or_2   g1300(new_n1575, new_n1558, new_n1576);
xor_5  g1301(new_n1576, new_n1557, n522);
or_2   g1302(new_n1029, new_n1025_1, new_n1578);
or_2   g1303(new_n1578, new_n1023, new_n1579);
or_2   g1304(new_n1579, new_n1233, new_n1580);
or_2   g1305(new_n1580, new_n1226, new_n1581);
nor_6  g1306(new_n1581, new_n1224, new_n1582);
and_7  g1307(new_n1581, new_n1224, new_n1583);
or_2   g1308(new_n1583, new_n1582, n532);
and_7  g1309(new_n822, new_n335, new_n1585);
and_7  g1310(new_n368, n247, new_n1586);
and_7  g1311(new_n1586, n1642, new_n1587);
and_7  g1312(new_n1587, n171, new_n1588);
and_7  g1313(new_n1588, n557, new_n1589);
and_7  g1314(new_n1589, n1000, new_n1590);
not_13 g1315(new_n1590, new_n1591);
xor_5  g1316(new_n368, new_n512, new_n1592);
and_7  g1317(new_n1592, n1000, new_n1593);
or_2   g1318(new_n704, n682, new_n1594);
and_7  g1319(new_n705, new_n334, new_n1595_1);
or_2   g1320(new_n1595_1, new_n500, new_n1596);
and_7  g1321(new_n1596, new_n1594, new_n1597_1);
and_7  g1322(new_n1597_1, new_n307, new_n1598);
or_2   g1323(new_n1598, new_n1593, new_n1599);
and_7  g1324(new_n1599, new_n381, new_n1600_1);
xor_5  g1325(new_n1594, n379, new_n1601_1);
nor_6  g1326(new_n1601_1, n1000, new_n1602);
xor_5  g1327(new_n1586, n1642, new_n1603);
and_7  g1328(new_n1603, n1000, new_n1604);
nor_6  g1329(new_n1604, new_n1602, new_n1605);
and_7  g1330(new_n1605, new_n1600_1, new_n1606);
or_2   g1331(new_n1594, n379, new_n1607);
and_7  g1332(new_n1607, n1263, new_n1608);
and_7  g1333(new_n930, new_n375, new_n1609);
or_2   g1334(new_n1609, new_n1608, new_n1610);
and_7  g1335(new_n1610, new_n307, new_n1611);
or_2   g1336(new_n1587, n171, new_n1612);
not_13 g1337(new_n1588, new_n1613_1);
and_7  g1338(new_n1613_1, n1000, new_n1614);
and_7  g1339(new_n1614, new_n1612, new_n1615);
nor_6  g1340(new_n1615, new_n1611, new_n1616);
and_7  g1341(new_n1616, new_n1606, new_n1617);
not_13 g1342(new_n1585, new_n1618);
and_7  g1343(new_n1614, new_n940, new_n1619);
or_2   g1344(new_n1609, new_n821, new_n1620);
and_7  g1345(new_n1620, new_n307, new_n1621);
or_2   g1346(new_n1621, new_n1590, new_n1622_1);
or_2   g1347(new_n1622_1, new_n1619, new_n1623);
and_7  g1348(new_n1623, new_n1618, new_n1624);
and_7  g1349(new_n1624, new_n1617, new_n1625);
and_7  g1350(new_n1625, new_n1591, new_n1626);
nor_6  g1351(new_n1626, new_n1585, new_n1627);
nor_6  g1352(new_n1624, new_n1617, new_n1628);
or_2   g1353(new_n1628, new_n1625, new_n1629_1);
nor_6  g1354(new_n1605, new_n1600_1, new_n1630);
or_2   g1355(new_n1630, new_n1606, new_n1631);
nor_6  g1356(new_n1599, new_n381, new_n1632);
or_2   g1357(new_n1632, new_n1600_1, new_n1633_1);
and_7  g1358(new_n1633_1, new_n383, new_n1634);
and_7  g1359(new_n1634, new_n1631, new_n1635_1);
nor_6  g1360(new_n1616, new_n1606, new_n1636);
or_2   g1361(new_n1636, new_n1617, new_n1637);
and_7  g1362(new_n1637, new_n1635_1, new_n1638);
and_7  g1363(new_n1638, new_n1629_1, new_n1639);
or_2   g1364(new_n1639, new_n1627, new_n1640);
nor_6  g1365(new_n1638, new_n1629_1, new_n1641);
nor_6  g1366(new_n1641, new_n1639, new_n1642_1);
and_7  g1367(new_n277_1, new_n862_1, new_n1643_1);
not_13 g1368(new_n1643_1, new_n1644);
or_2   g1369(new_n881, new_n863, new_n1645);
and_7  g1370(new_n1645, new_n1644, new_n1646);
and_7  g1371(new_n1646, n49, new_n1647);
and_7  g1372(new_n1647, n1622, new_n1648);
and_7  g1373(new_n1648, n906, new_n1649);
and_7  g1374(new_n1649, n277, new_n1650);
nor_6  g1375(new_n1637, new_n1635_1, new_n1651);
nor_6  g1376(new_n1651, new_n1638, new_n1652);
nor_6  g1377(new_n1652, new_n1650, new_n1653);
and_7  g1378(new_n1652, new_n1650, new_n1654_1);
or_2   g1379(new_n1654_1, new_n1653, new_n1655);
not_13 g1380(n277, new_n1656);
not_13 g1381(n906, new_n1657_1);
not_13 g1382(n1622, new_n1658);
not_13 g1383(n49, new_n1659);
or_2   g1384(new_n891_1, new_n1643_1, new_n1660_1);
or_2   g1385(new_n1660_1, new_n1659, new_n1661);
or_2   g1386(new_n1661, new_n1658, new_n1662);
or_2   g1387(new_n1662, new_n1657_1, new_n1663);
and_7  g1388(new_n1663, new_n1656, new_n1664);
nor_6  g1389(new_n1664, new_n1650, new_n1665);
nor_6  g1390(new_n1634, new_n1631, new_n1666);
nor_6  g1391(new_n1666, new_n1635_1, new_n1667);
or_2   g1392(new_n1667, new_n1665, new_n1668);
nor_6  g1393(new_n1667, new_n1665, new_n1669);
and_7  g1394(new_n1667, new_n1665, new_n1670);
or_2   g1395(new_n1670, new_n1669, new_n1671);
and_7  g1396(new_n1662, new_n1657_1, new_n1672);
nor_6  g1397(new_n1672, new_n1649, new_n1673);
nor_6  g1398(new_n1633_1, new_n383, new_n1674);
nor_6  g1399(new_n1674, new_n1634, new_n1675_1);
nor_6  g1400(new_n1675_1, new_n1673, new_n1676);
and_7  g1401(new_n1675_1, new_n1673, new_n1677_1);
or_2   g1402(new_n1677_1, new_n1676, new_n1678_1);
or_2   g1403(new_n1647, n1622, new_n1679);
and_7  g1404(new_n1679, new_n1662, new_n1680);
nor_6  g1405(new_n1680, new_n385, new_n1681);
and_7  g1406(new_n1680, new_n385, new_n1682);
nor_6  g1407(new_n1682, new_n1681, new_n1683_1);
and_7  g1408(new_n1660_1, new_n1659, new_n1684);
nor_6  g1409(new_n1684, new_n1647, new_n1685);
and_7  g1410(new_n1685, new_n390, new_n1686_1);
nor_6  g1411(new_n1685, new_n390, new_n1687);
or_2   g1412(new_n1687, new_n1686_1, new_n1688_1);
and_7  g1413(new_n924, new_n895, new_n1689);
nor_6  g1414(new_n1689, new_n893, new_n1690_1);
nor_6  g1415(new_n1690_1, new_n1688_1, new_n1691);
nor_6  g1416(new_n1691, new_n1686_1, new_n1692);
and_7  g1417(new_n1692, new_n1683_1, new_n1693);
nor_6  g1418(new_n1693, new_n1681, new_n1694);
nor_6  g1419(new_n1694, new_n1678_1, new_n1695);
nor_6  g1420(new_n1695, new_n1676, new_n1696);
or_2   g1421(new_n1696, new_n1671, new_n1697);
and_7  g1422(new_n1697, new_n1668, new_n1698);
nor_6  g1423(new_n1698, new_n1655, new_n1699);
nor_6  g1424(new_n1699, new_n1653, new_n1700);
and_7  g1425(new_n1700, new_n1642_1, new_n1701);
nor_6  g1426(new_n1701, new_n1640, n534);
and_7  g1427(n1721, new_n589, new_n1703);
or_2   g1428(new_n1703, new_n592, n541);
or_2   g1429(new_n1026, new_n1015_1, n547);
nor_6  g1430(new_n1265, new_n1190, new_n1706);
and_7  g1431(new_n1265, new_n1190, new_n1707_1);
or_2   g1432(new_n1707_1, new_n1706, new_n1708);
nor_6  g1433(new_n1552, new_n1512, new_n1709);
nor_6  g1434(new_n1709, new_n1708, new_n1710);
or_2   g1435(new_n1710, new_n1706, new_n1711);
and_7  g1436(new_n1711, new_n1272, n549);
and_7  g1437(new_n1572, new_n1570, new_n1713);
or_2   g1438(new_n1713, new_n1573, n559);
not_13 g1439(new_n1419, n569);
xor_5  g1440(new_n1543, new_n1541, n573);
and_7  g1441(new_n1709, new_n1708, new_n1717);
or_2   g1442(new_n1717, new_n1710, n588);
not_13 g1443(new_n585_1, new_n1719);
xor_5  g1444(n416, new_n1719, n599);
nor_6  g1445(new_n1427, new_n1398, n627);
and_7  g1446(new_n1263_1, new_n811, new_n1722);
xor_5  g1447(new_n1722, new_n1382, new_n1723);
or_2   g1448(new_n1723, new_n1271, new_n1724);
nor_6  g1449(new_n1270, new_n1266, new_n1725);
xor_5  g1450(new_n1722, new_n826, new_n1726);
or_2   g1451(new_n1726, new_n1725, new_n1727_1);
and_7  g1452(new_n1727_1, new_n1724, n638);
and_7  g1453(new_n930, new_n821, new_n1729_1);
and_7  g1454(new_n1729_1, new_n457_1, new_n1730);
and_7  g1455(new_n944_1, n1381, new_n1731_1);
or_2   g1456(new_n1731_1, new_n1730, new_n1732);
not_13 g1457(new_n1732, new_n1733);
nor_6  g1458(new_n1733, new_n954, n643);
xor_5  g1459(new_n1690_1, new_n1688_1, n648);
or_2   g1460(new_n779, new_n739, new_n1736);
xor_5  g1461(new_n1736, new_n734, n665);
or_2   g1462(new_n1182, new_n1178, new_n1738);
xor_5  g1463(new_n1738, new_n1173, n683);
or_2   g1464(new_n1642_1, new_n1190, new_n1740);
nor_6  g1465(new_n1642_1, new_n1190, new_n1741);
and_7  g1466(new_n1642_1, new_n1190, new_n1742);
or_2   g1467(new_n1742, new_n1741, new_n1743_1);
or_2   g1468(new_n1652, new_n1190, new_n1744);
nor_6  g1469(new_n1652, new_n1190, new_n1745);
and_7  g1470(new_n1652, new_n1190, new_n1746_1);
or_2   g1471(new_n1746_1, new_n1745, new_n1747_1);
nor_6  g1472(new_n1667, new_n1199_1, new_n1748);
and_7  g1473(new_n1667, new_n1199_1, new_n1749);
nor_6  g1474(new_n1749, new_n1748, new_n1750);
nor_6  g1475(new_n1675_1, new_n1204, new_n1751);
and_7  g1476(new_n1675_1, new_n1204, new_n1752);
or_2   g1477(new_n1752, new_n1751, new_n1753);
nor_6  g1478(new_n452_1, new_n387_1, new_n1754);
nor_6  g1479(new_n1754, new_n1753, new_n1755);
or_2   g1480(new_n1755, new_n1751, new_n1756);
and_7  g1481(new_n1756, new_n1750, new_n1757_1);
nor_6  g1482(new_n1757_1, new_n1748, new_n1758);
or_2   g1483(new_n1758, new_n1747_1, new_n1759);
and_7  g1484(new_n1759, new_n1744, new_n1760);
or_2   g1485(new_n1760, new_n1743_1, new_n1761);
and_7  g1486(new_n1761, new_n1740, new_n1762);
or_2   g1487(new_n1617, new_n1591, new_n1763_1);
and_7  g1488(new_n1763_1, new_n1627, new_n1764_1);
nor_6  g1489(new_n1764_1, new_n1639, new_n1765);
and_7  g1490(new_n1764_1, new_n1639, new_n1766);
nor_6  g1491(new_n1766, new_n1765, new_n1767);
nor_6  g1492(new_n1767, new_n1762, new_n1768);
and_7  g1493(new_n1767, new_n1197, new_n1769);
and_7  g1494(new_n1761, new_n1190, new_n1770);
or_2   g1495(new_n1770, new_n1769, new_n1771);
nor_6  g1496(new_n1771, new_n1768, new_n1772);
nor_6  g1497(new_n1772, new_n1640, new_n1773);
and_7  g1498(new_n1772, new_n1640, new_n1774);
or_2   g1499(new_n1774, new_n1773, n699);
not_13 g1500(new_n431, new_n1776);
xor_5  g1501(new_n913, new_n1776, n712);
not_13 g1502(new_n594, n715);
nor_6  g1503(new_n1423, n145, new_n1779);
nor_6  g1504(new_n1779, new_n1424, n724);
not_13 g1505(n647, n1255);
xor_5  g1506(new_n978, new_n977, new_n1782);
and_7  g1507(new_n1782, n1255, new_n1783);
xor_5  g1508(n1016, new_n1783, n725);
and_7  g1509(new_n1574, new_n1560, new_n1785);
or_2   g1510(new_n1785, new_n1575, n731);
and_7  g1511(new_n1754, new_n1753, new_n1787);
or_2   g1512(new_n1787, new_n1755, n748);
or_2   g1513(new_n1502_1, new_n1492, new_n1789);
xor_5  g1514(new_n1789, new_n1491, n759);
and_7  g1515(new_n1582, new_n1238, new_n1791);
and_7  g1516(new_n1197, new_n805, new_n1792);
nor_6  g1517(new_n1220, new_n1792, new_n1793);
nor_6  g1518(new_n1793, n1422, new_n1794);
and_7  g1519(new_n1794, new_n1791, n770);
or_2   g1520(new_n1544_1, new_n1524, new_n1796);
xor_5  g1521(new_n1796, new_n1523, n790);
and_7  g1522(new_n1190, new_n833, new_n1798);
nor_6  g1523(new_n1190, new_n833, new_n1799);
or_2   g1524(new_n1799, new_n1798, new_n1800);
nor_6  g1525(new_n1556_1, new_n1555, new_n1801);
and_7  g1526(new_n1576, new_n1801, new_n1802);
nor_6  g1527(new_n1802, new_n1556_1, new_n1803);
nor_6  g1528(new_n1803, new_n1800, new_n1804);
and_7  g1529(new_n1803, new_n1800, new_n1805);
or_2   g1530(new_n1805, new_n1804, n792);
not_13 g1531(new_n1131, new_n1807);
xor_5  g1532(new_n1134, new_n1807, n813);
and_7  g1533(new_n1367, new_n1358, new_n1809);
or_2   g1534(new_n1809, new_n1368, n823);
and_7  g1535(new_n1386, new_n823_1, n824);
not_13 g1536(new_n486, new_n1812);
xor_5  g1537(new_n488_1, new_n1812, n836);
or_2   g1538(new_n1749, new_n1748, new_n1814);
xor_5  g1539(new_n1756, new_n1814, n846);
not_13 g1540(new_n1342, new_n1816);
or_2   g1541(new_n1371, new_n1344, new_n1817);
and_7  g1542(new_n1817, new_n1816, new_n1818);
xor_5  g1543(new_n1818, new_n1337, n858);
or_2   g1544(new_n1395, new_n794, new_n1820);
and_7  g1545(new_n1820, new_n1385_1, n865);
and_7  g1546(new_n1549, new_n1516, new_n1822);
or_2   g1547(new_n1822, new_n1550, n867);
or_2   g1548(new_n952_1, new_n947, new_n1824);
xor_5  g1549(new_n1478, new_n1824, new_n1825);
or_2   g1550(new_n1508, new_n1482, new_n1826);
and_7  g1551(new_n1826, new_n1825, new_n1827);
nor_6  g1552(new_n1826, new_n1825, new_n1828);
nor_6  g1553(new_n1828, new_n1827, n883);
and_7  g1554(new_n784, new_n782, new_n1830);
or_2   g1555(new_n1830, new_n785, n888);
xor_5  g1556(new_n1478, new_n953_1, new_n1832);
and_7  g1557(new_n1312, n1757, new_n1833);
and_7  g1558(new_n1833, n839, new_n1834);
or_2   g1559(new_n1834, new_n1480, new_n1835);
nor_6  g1560(new_n1834, new_n1480, new_n1836);
and_7  g1561(new_n1834, new_n1480, new_n1837);
or_2   g1562(new_n1837, new_n1836, new_n1838);
not_13 g1563(n839, new_n1839);
and_7  g1564(new_n1438, new_n1839, new_n1840);
nor_6  g1565(new_n1840, new_n1834, new_n1841);
or_2   g1566(new_n1841, new_n1485, new_n1842);
nor_6  g1567(new_n1841, new_n1485, new_n1843);
and_7  g1568(new_n1841, new_n1485, new_n1844);
or_2   g1569(new_n1844, new_n1843, new_n1845);
or_2   g1570(new_n1377, new_n1325, new_n1846);
and_7  g1571(new_n1846, new_n1443, new_n1847);
nor_6  g1572(new_n1847, new_n1442, new_n1848);
or_2   g1573(new_n1848, new_n1845, new_n1849);
and_7  g1574(new_n1849, new_n1842, new_n1850);
or_2   g1575(new_n1850, new_n1838, new_n1851);
and_7  g1576(new_n1851, new_n1835, new_n1852);
or_2   g1577(new_n1852, new_n1832, new_n1853);
nor_6  g1578(new_n1850, new_n1838, new_n1854);
or_2   g1579(new_n1854, new_n1836, new_n1855);
or_2   g1580(new_n1855, new_n1825, new_n1856);
and_7  g1581(new_n1856, new_n1853, n891);
and_7  g1582(new_n1478, new_n953_1, new_n1858);
and_7  g1583(new_n1852, new_n1832, new_n1859);
nor_6  g1584(new_n1859, new_n1858, new_n1860);
and_7  g1585(new_n1860, new_n1732, n892);
xor_5  g1586(new_n1113_1, new_n1112, n902);
not_13 g1587(new_n1254, new_n1863);
xor_5  g1588(new_n743, new_n407, new_n1864);
xor_5  g1589(new_n1864, new_n1863, n905);
xor_5  g1590(new_n1468, new_n1226, n912);
nor_6  g1591(n1149, new_n600_1, new_n1867);
nor_6  g1592(new_n1867, new_n959, n935);
xor_5  g1593(new_n1424, n1119, n942);
or_2   g1594(new_n1179, new_n1178, new_n1870);
xor_5  g1595(new_n1181, new_n1870, n944);
and_7  g1596(n770, n547, n974);
or_2   g1597(new_n448, new_n403, new_n1873);
xor_5  g1598(new_n1873, new_n398, n979);
and_7  g1599(new_n1382, new_n819, new_n1875);
not_13 g1600(new_n1875, new_n1876);
and_7  g1601(new_n1876, new_n1389, new_n1877);
nor_6  g1602(new_n1877, new_n828, new_n1878);
and_7  g1603(new_n1878, new_n855, n980);
or_2   g1604(new_n1546, new_n1521, new_n1880);
xor_5  g1605(new_n1880, new_n1520, n989);
nor_6  g1606(new_n1758, new_n1747_1, new_n1882);
or_2   g1607(new_n1882, new_n1745, new_n1883);
xor_5  g1608(new_n1883, new_n1743_1, n991);
or_2   g1609(new_n1847, new_n1442, new_n1885);
xor_5  g1610(new_n1885, new_n1845, n1005);
and_7  g1611(new_n1505, new_n1488, new_n1887);
or_2   g1612(new_n1887, new_n1506, n1012);
nor_6  g1613(new_n1029, new_n1025_1, new_n1889);
xor_5  g1614(new_n1889, new_n1023, n1015);
and_7  g1615(new_n859, new_n856, new_n1891);
and_7  g1616(new_n1877, new_n1891, new_n1892);
and_7  g1617(new_n1877, new_n828, new_n1893);
or_2   g1618(new_n1893, new_n1878, new_n1894);
and_7  g1619(new_n1894, new_n855, new_n1895);
or_2   g1620(new_n1895, new_n1892, n1025);
and_7  g1621(new_n1850, new_n1838, new_n1897);
or_2   g1622(new_n1897, new_n1854, n1030);
and_7  g1623(new_n850, new_n846_1, new_n1899);
or_2   g1624(new_n1899, new_n851, n1067);
nor_6  g1625(new_n1860, new_n1732, new_n1901);
or_2   g1626(new_n1901, n892, n1068);
xor_5  g1627(new_n594, new_n592, n1103);
xor_5  g1628(new_n482_1, new_n413, n1113);
or_2   g1629(new_n1581, new_n1224, new_n1905);
or_2   g1630(new_n1905, new_n1222_1, new_n1906);
and_7  g1631(new_n1793, n1422, new_n1907);
and_7  g1632(new_n1907, new_n1906, new_n1908);
or_2   g1633(new_n1908, n770, n1135);
and_7  g1634(new_n1764_1, new_n1701, new_n1910);
nor_6  g1635(new_n1767, new_n1701, new_n1911);
or_2   g1636(new_n1911, new_n1910, n1142);
nor_6  g1637(new_n1767, new_n1197, new_n1913);
nor_6  g1638(new_n1913, new_n1769, new_n1914);
nor_6  g1639(new_n1914, new_n1762, new_n1915);
and_7  g1640(new_n1914, new_n1762, new_n1916);
nor_6  g1641(new_n1916, new_n1915, n1161);
nor_6  g1642(new_n1579, new_n1233, new_n1918);
and_7  g1643(new_n1579, new_n1233, new_n1919);
or_2   g1644(new_n1919, new_n1918, n1162);
nor_6  g1645(n865, new_n1425_1, new_n1921);
nor_6  g1646(new_n1921, new_n1426_1, n1175);
or_2   g1647(new_n1190, new_n833, new_n1923);
or_2   g1648(new_n1803, new_n1800, new_n1924);
and_7  g1649(new_n1924, new_n1923, new_n1925);
and_7  g1650(new_n1190, new_n830, new_n1926);
or_2   g1651(new_n1926, new_n1925, new_n1927);
and_7  g1652(new_n1197, new_n856, new_n1928);
or_2   g1653(new_n1928, new_n1804, new_n1929);
and_7  g1654(new_n1929, new_n1927, new_n1930);
and_7  g1655(new_n1930, new_n1894, new_n1931);
nor_6  g1656(new_n1893, new_n1878, new_n1932);
or_2   g1657(new_n1804, new_n1799, new_n1933);
or_2   g1658(new_n1197, new_n856, new_n1934);
and_7  g1659(new_n1934, new_n1933, new_n1935);
or_2   g1660(new_n1190, new_n830, new_n1936);
and_7  g1661(new_n1936, new_n1924, new_n1937);
or_2   g1662(new_n1937, new_n1935, new_n1938);
and_7  g1663(new_n1938, new_n1932, new_n1939);
nor_6  g1664(new_n1939, new_n1931, n1191);
xor_5  g1665(new_n1918, new_n1226, n1194);
xor_5  g1666(new_n447, new_n445, n1199);
nor_6  g1667(new_n1537_1, new_n1531, new_n1943);
or_2   g1668(new_n1943, new_n1538, n1201);
not_13 g1669(new_n979_1, new_n1945);
and_7  g1670(new_n1405, new_n1945, new_n1946);
or_2   g1671(new_n1946, new_n1783, n1202);
xor_5  g1672(new_n1419, new_n1417, n1234);
and_7  g1673(new_n1905, new_n1222_1, new_n1949);
or_2   g1674(new_n1949, new_n1791, n1235);
not_13 g1675(n1183, n1237);
and_7  g1676(new_n1722, new_n826, new_n1952);
and_7  g1677(new_n1726, new_n1725, new_n1953);
nor_6  g1678(new_n1953, new_n1952, new_n1954);
nor_6  g1679(new_n1954, new_n823_1, new_n1955);
or_2   g1680(new_n1955, n299, n1260);
nor_6  g1681(new_n1426_1, n1249, new_n1957);
nor_6  g1682(new_n1957, new_n1427, n1277);
nor_6  g1683(new_n1828, new_n1858, new_n1959);
and_7  g1684(new_n1959, new_n1732, n1278);
and_7  g1685(new_n431, new_n419, new_n1961);
or_2   g1686(new_n431, new_n424_1, new_n1962);
and_7  g1687(new_n1962, new_n433_1, new_n1963);
nor_6  g1688(new_n1963, new_n1961, n1283);
or_2   g1689(new_n1236, new_n1222_1, new_n1965);
and_7  g1690(new_n1907, new_n1965, new_n1966);
or_2   g1691(new_n1966, n974, n1305);
xor_5  g1692(new_n595, n1727, n1315);
nor_6  g1693(new_n1696, new_n1671, new_n1969);
and_7  g1694(new_n1696, new_n1671, new_n1970);
or_2   g1695(new_n1970, new_n1969, n1330);
nor_6  g1696(new_n1568, new_n1564, new_n1972);
or_2   g1697(new_n1972, new_n1569, n1338);
not_13 g1698(new_n770_1, new_n1974);
xor_5  g1699(new_n1974, new_n768, n1340);
nor_6  g1700(new_n1700, new_n1642_1, new_n1976);
nor_6  g1701(new_n1976, new_n1701, n1347);
and_7  g1702(new_n1733, new_n954, new_n1978);
or_2   g1703(new_n1978, n643, n1348);
and_7  g1704(new_n1371, new_n1344, new_n1980);
or_2   g1705(new_n1980, new_n1372, n1349);
nor_6  g1706(new_n1907, new_n1794, new_n1982);
nor_6  g1707(new_n1982, new_n1791, new_n1983);
and_7  g1708(new_n1982, new_n1791, new_n1984);
nor_6  g1709(new_n1984, new_n1983, n1369);
nor_6  g1710(new_n1982, new_n1240, new_n1986);
and_7  g1711(new_n1982, new_n1240, new_n1987);
nor_6  g1712(new_n1987, new_n1986, n1383);
or_2   g1713(new_n1691, new_n1686_1, new_n1989);
xor_5  g1714(new_n1989, new_n1683_1, n1393);
not_13 g1715(new_n1535_1, new_n1991);
xor_5  g1716(new_n1991, new_n1121, n1399);
xor_5  g1717(new_n750, new_n412, new_n1993);
xor_5  g1718(new_n1993, new_n1252, n1407);
and_7  g1719(new_n1397, new_n826, new_n1995);
and_7  g1720(new_n1995, new_n1389, new_n1996);
or_2   g1721(n824, new_n1996, n1425);
or_2   g1722(new_n1733, new_n954, new_n1998);
nor_6  g1723(new_n1998, new_n961_1, n1440);
or_2   g1724(new_n1028, new_n1017, n1601);
xor_5  g1725(n1601, new_n1025_1, n1453);
not_13 g1726(new_n1250, new_n2002);
xor_5  g1727(new_n2002, new_n768, n1460);
and_7  g1728(new_n1936, new_n1934, new_n2004);
or_2   g1729(new_n2004, new_n1933, new_n2005);
or_2   g1730(new_n1928, new_n1926, new_n2006);
or_2   g1731(new_n2006, new_n1925, new_n2007);
and_7  g1732(new_n2007, new_n2005, n1463);
and_7  g1733(new_n1235_1, new_n1224, new_n2009);
or_2   g1734(new_n2009, new_n1239, n1470);
xor_5  g1735(new_n1113_1, new_n413, n1481);
not_13 g1736(new_n772, new_n2012);
xor_5  g1737(new_n774, new_n2012, n1495);
and_7  g1738(new_n1129, new_n1105, new_n2014);
or_2   g1739(new_n2014, new_n1130, n1498);
and_7  g1740(new_n1694, new_n1678_1, new_n2016);
or_2   g1741(new_n2016, new_n1695, n1502);
not_13 g1742(new_n1353, new_n2018);
xor_5  g1743(new_n1369_1, new_n2018, n1507);
xor_5  g1744(new_n1416, new_n1412, n1525);
and_7  g1745(new_n776, new_n748_1, new_n2021);
or_2   g1746(new_n2021, new_n777, n1535);
xor_5  g1747(new_n1029, n547, n1556);
and_7  g1748(n1348, new_n961_1, new_n2024);
nor_6  g1749(n1348, new_n961_1, new_n2025);
nor_6  g1750(new_n2025, new_n2024, n1595);
and_7  g1751(new_n1539, new_n1527_1, new_n2027);
or_2   g1752(new_n2027, new_n1540, n1600);
or_2   g1753(new_n471, n1145, new_n2029);
and_7  g1754(new_n2029, new_n581, new_n2030);
or_2   g1755(new_n2030, new_n1719, n1613);
xor_5  g1756(new_n1365, new_n1812, n1629);
or_2   g1757(new_n1877, new_n828, new_n2033);
and_7  g1758(new_n1938, new_n2033, new_n2034);
and_7  g1759(new_n1928, new_n1925, new_n2035);
or_2   g1760(new_n2035, new_n1893, new_n2036);
nor_6  g1761(new_n2036, new_n2034, n1633);
and_7  g1762(n1601, n547, new_n2038);
xor_5  g1763(new_n2038, new_n1025_1, n1635);
xor_5  g1764(new_n1501_1, new_n1499, n1654);
xor_5  g1765(new_n597, n1138, n1657);
or_2   g1766(new_n1828, new_n1858, new_n2042);
and_7  g1767(new_n2042, new_n1733, new_n2043);
or_2   g1768(new_n2043, n1278, n1660);
not_13 g1769(new_n1123, new_n2045);
xor_5  g1770(new_n2045, new_n1121, n1675);
not_13 g1771(new_n1416, n1683);
or_2   g1772(new_n1723, new_n1711, new_n2048);
or_2   g1773(new_n1265, new_n1190, new_n2049);
or_2   g1774(new_n1709, new_n1708, new_n2050);
and_7  g1775(new_n2050, new_n2049, new_n2051);
or_2   g1776(new_n1726, new_n2051, new_n2052);
and_7  g1777(new_n2052, new_n2048, n1686);
xor_5  g1778(new_n761_1, new_n413, n1688);
and_7  g1779(new_n1698, new_n1655, new_n2055);
or_2   g1780(new_n2055, new_n1699, n1690);
and_7  g1781(new_n1758, new_n1747_1, new_n2057);
or_2   g1782(new_n2057, new_n1882, n1729);
and_7  g1783(new_n1726, new_n2051, new_n2059);
nor_6  g1784(new_n2059, new_n1952, new_n2060);
nor_6  g1785(new_n2060, new_n823_1, new_n2061);
or_2   g1786(new_n2061, n549, n1737);
not_13 g1787(new_n1461_1, new_n2063);
or_2   g1788(new_n1464, new_n1462, new_n2064);
and_7  g1789(new_n2064, new_n2063, new_n2065);
xor_5  g1790(new_n2065, new_n1496, n1746);
xor_5  g1791(new_n413, n347, n488);
xor_5  g1792(new_n1012_1, new_n1259, n1677);
endmodule


