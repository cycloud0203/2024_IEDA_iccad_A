// Benchmark "top_810026173_826291639_946996917_1246901" written by ABC on Sun Jun 23 19:37:07 2024

module top_810026173_826291639_946996917_1246901 ( 
    n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213, n223,
    n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414, n424,
    n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649, n653,
    n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788, n801,
    n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764,
    n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156, n174,
    n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299, n317,
    n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457, n460,
    n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547, n549,
    n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648, n665,
    n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773, n790,
    n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888, n891,
    n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989, n991,
    n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103, n1113,
    n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183, n1191,
    n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255, n1260,
    n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347, n1348,
    n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426, n1440,
    n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502, n1507,
    n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633, n1635,
    n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690, n1721,
    n1727, n1729, n1731, n1737, n1746  );
  input  n14, n17, n26, n36, n46, n49, n66, n69, n155, n171, n183, n213,
    n223, n247, n266, n277, n303, n329, n347, n353, n379, n391, n402, n414,
    n424, n433, n444, n469, n472, n498, n555, n557, n585, n600, n607, n649,
    n653, n655, n675, n682, n684, n693, n695, n729, n738, n747, n761, n788,
    n801, n839, n862, n870, n882, n906, n927, n931, n952, n953, n961, n968,
    n1000, n1062, n1140, n1145, n1172, n1222, n1263, n1296, n1321, n1332,
    n1341, n1351, n1363, n1381, n1422, n1435, n1461, n1501, n1527, n1530,
    n1537, n1544, n1597, n1622, n1642, n1643, n1678, n1707, n1743, n1747,
    n1757, n1763, n1764;
  output n19, n33, n44, n55, n56, n67, n74, n106, n126, n135, n145, n156,
    n174, n181, n208, n216, n218, n231, n238, n270, n276, n290, n292, n299,
    n317, n372, n378, n387, n401, n416, n423, n426, n429, n432, n452, n457,
    n460, n476, n482, n488, n493, n510, n517, n522, n532, n534, n541, n547,
    n549, n559, n569, n573, n588, n599, n627, n638, n643, n646, n647, n648,
    n665, n683, n699, n712, n715, n724, n725, n731, n748, n759, n770, n773,
    n790, n792, n813, n823, n824, n836, n846, n858, n865, n867, n883, n888,
    n891, n892, n902, n905, n912, n935, n942, n944, n974, n979, n980, n989,
    n991, n1005, n1012, n1015, n1016, n1025, n1030, n1067, n1068, n1103,
    n1113, n1119, n1135, n1138, n1142, n1149, n1161, n1162, n1175, n1183,
    n1191, n1194, n1199, n1201, n1202, n1234, n1235, n1237, n1249, n1255,
    n1260, n1277, n1278, n1283, n1305, n1315, n1330, n1338, n1340, n1347,
    n1348, n1349, n1369, n1383, n1385, n1393, n1399, n1407, n1425, n1426,
    n1440, n1453, n1457, n1460, n1463, n1470, n1481, n1495, n1498, n1502,
    n1507, n1525, n1535, n1556, n1595, n1600, n1601, n1613, n1629, n1633,
    n1635, n1654, n1657, n1660, n1675, n1677, n1683, n1686, n1688, n1690,
    n1721, n1727, n1729, n1731, n1737, n1746;
  wire new_n276_1, new_n277_1, new_n278, new_n279, new_n280, new_n281,
    new_n282, new_n283, new_n284, new_n285, new_n286, new_n287, new_n288,
    new_n289, new_n290_1, new_n291, new_n292_1, new_n293, new_n294,
    new_n295, new_n296, new_n297, new_n298, new_n299_1, new_n300, new_n301,
    new_n302, new_n303_1, new_n304, new_n305, new_n306, new_n307, new_n308,
    new_n309, new_n310, new_n311, new_n312, new_n313, new_n314, new_n315,
    new_n316, new_n317_1, new_n318, new_n319, new_n320, new_n321, new_n322,
    new_n323, new_n324, new_n325, new_n326, new_n327, new_n328, new_n329_1,
    new_n330, new_n331, new_n332, new_n333, new_n334, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347_1, new_n348, new_n349, new_n350,
    new_n351, new_n352, new_n353_1, new_n354, new_n355, new_n356, new_n357,
    new_n358, new_n359, new_n360, new_n361, new_n362, new_n363, new_n364,
    new_n365, new_n366, new_n367, new_n368, new_n369, new_n370, new_n371,
    new_n372_1, new_n373, new_n374, new_n375, new_n376, new_n377,
    new_n378_1, new_n379_1, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387_1, new_n388, new_n389, new_n390,
    new_n391_1, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401_1, new_n402_1, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414_1, new_n415, new_n416_1,
    new_n417, new_n418, new_n419, new_n420, new_n421, new_n422, new_n423_1,
    new_n424_1, new_n425, new_n426_1, new_n427, new_n428, new_n429_1,
    new_n430, new_n431, new_n432_1, new_n433_1, new_n434, new_n435,
    new_n436, new_n437, new_n438, new_n439, new_n440, new_n441, new_n442,
    new_n443, new_n444_1, new_n445, new_n446, new_n447, new_n448, new_n449,
    new_n450, new_n451, new_n452_1, new_n453, new_n455, new_n456,
    new_n457_1, new_n458, new_n459, new_n460_1, new_n461, new_n462,
    new_n463, new_n464, new_n465, new_n466, new_n467, new_n468, new_n469_1,
    new_n470, new_n471, new_n472_1, new_n473, new_n474, new_n475,
    new_n476_1, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482_1, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488_1, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498_1, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510_1, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517_1, new_n518, new_n519, new_n520, new_n521, new_n522_1,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532_1, new_n533, new_n534_1, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541_1, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547_1, new_n548,
    new_n549_1, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555_1, new_n556, new_n557_1, new_n558, new_n559_1, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569_1, new_n570, new_n572, new_n573_1, new_n574,
    new_n575, new_n576, new_n577, new_n579, new_n581, new_n582, new_n585_1,
    new_n586, new_n587, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599_1, new_n600_1,
    new_n603, new_n604, new_n605, new_n606, new_n607_1, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627_1, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638_1, new_n639, new_n640, new_n641, new_n642, new_n643_1,
    new_n644, new_n645, new_n646_1, new_n647_1, new_n648_1, new_n649_1,
    new_n650, new_n651, new_n652, new_n653_1, new_n654, new_n655_1,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665_1, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675_1, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682_1,
    new_n683_1, new_n684_1, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693_1, new_n694,
    new_n695_1, new_n696, new_n697, new_n698, new_n699_1, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712_1, new_n713, new_n714,
    new_n715_1, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724_1, new_n725_1, new_n726, new_n727,
    new_n728, new_n729_1, new_n730, new_n731_1, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738_1, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747_1,
    new_n748_1, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759_1, new_n760,
    new_n761_1, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770_1, new_n771, new_n772, new_n773_1,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788_1,
    new_n789, new_n790_1, new_n791, new_n792_1, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801_1,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813_1, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823_1, new_n824_1, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836_1, new_n837, new_n838, new_n839_1, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846_1, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858_1, new_n859, new_n860, new_n862_1,
    new_n863, new_n864, new_n865_1, new_n866, new_n867_1, new_n868,
    new_n869, new_n870_1, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882_1,
    new_n883_1, new_n884, new_n885, new_n886, new_n887, new_n888_1,
    new_n889, new_n890, new_n891_1, new_n892_1, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902_1, new_n903, new_n904, new_n905_1, new_n906_1, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912_1, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927_1, new_n928, new_n929,
    new_n930, new_n931_1, new_n932, new_n933, new_n934, new_n935_1,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942_1,
    new_n943, new_n944_1, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952_1, new_n953_1, new_n954, new_n955,
    new_n957, new_n959, new_n960, new_n961_1, new_n964, new_n966, new_n967,
    new_n968_1, new_n970, new_n971, new_n972, new_n973, new_n974_1,
    new_n975, new_n976, new_n977, new_n978, new_n979_1, new_n980_1,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n991_1, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000_1, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005_1, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012_1, new_n1013, new_n1014,
    new_n1015_1, new_n1016_1, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025_1, new_n1026,
    new_n1028, new_n1029, new_n1030_1, new_n1031, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062_1, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067_1, new_n1068_1, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103_1, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113_1,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119_1,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135_1, new_n1136, new_n1137,
    new_n1138_1, new_n1140_1, new_n1142_1, new_n1144, new_n1145_1,
    new_n1146, new_n1147, new_n1148, new_n1149_1, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161_1, new_n1162_1, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172_1, new_n1173, new_n1174, new_n1175_1,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183_1, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191_1, new_n1192, new_n1193, new_n1194_1,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199_1, new_n1200,
    new_n1201_1, new_n1202_1, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222_1, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234_1, new_n1235_1, new_n1236,
    new_n1237_1, new_n1238, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249_1,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255_1,
    new_n1256, new_n1259, new_n1261, new_n1262, new_n1263_1, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1274, new_n1275, new_n1276, new_n1277_1,
    new_n1278_1, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283_1,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296_1, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305_1, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315_1, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321_1, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330_1, new_n1331,
    new_n1332_1, new_n1333, new_n1334, new_n1335, new_n1336, new_n1337,
    new_n1338_1, new_n1339, new_n1340_1, new_n1341_1, new_n1342, new_n1343,
    new_n1344, new_n1345, new_n1346, new_n1347_1, new_n1348_1, new_n1349_1,
    new_n1350, new_n1351_1, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363_1, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369_1, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1380, new_n1382,
    new_n1383_1, new_n1384, new_n1385_1, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393_1, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399_1, new_n1400,
    new_n1402, new_n1404, new_n1405, new_n1408, new_n1409, new_n1410,
    new_n1412, new_n1413, new_n1414, new_n1415, new_n1416, new_n1417,
    new_n1418, new_n1419, new_n1420, new_n1421, new_n1423, new_n1424,
    new_n1425_1, new_n1426_1, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1432, new_n1433, new_n1434, new_n1435_1, new_n1436, new_n1437,
    new_n1438, new_n1439, new_n1440_1, new_n1441, new_n1442, new_n1443,
    new_n1444, new_n1445, new_n1446, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453_1, new_n1455, new_n1457_1, new_n1460_1,
    new_n1461_1, new_n1462, new_n1463_1, new_n1464, new_n1465, new_n1466,
    new_n1468, new_n1469, new_n1471, new_n1474, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1481_1, new_n1482, new_n1483,
    new_n1484, new_n1485, new_n1486, new_n1487, new_n1488, new_n1489,
    new_n1490, new_n1491, new_n1492, new_n1493, new_n1494, new_n1495_1,
    new_n1496, new_n1497, new_n1498_1, new_n1499, new_n1500, new_n1501_1,
    new_n1502_1, new_n1503, new_n1504, new_n1505, new_n1506, new_n1507_1,
    new_n1508, new_n1509, new_n1511, new_n1512, new_n1513, new_n1514,
    new_n1515, new_n1516, new_n1517, new_n1518, new_n1519, new_n1520,
    new_n1521, new_n1522, new_n1523, new_n1524, new_n1525_1, new_n1526,
    new_n1527_1, new_n1528, new_n1529, new_n1530_1, new_n1531, new_n1532,
    new_n1533, new_n1534, new_n1535_1, new_n1536, new_n1537_1, new_n1538,
    new_n1539, new_n1540, new_n1541, new_n1542, new_n1543, new_n1544_1,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1555, new_n1556_1, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1562, new_n1563,
    new_n1564, new_n1565, new_n1566, new_n1567, new_n1568, new_n1569,
    new_n1570, new_n1571, new_n1572, new_n1573, new_n1574, new_n1575,
    new_n1576, new_n1578, new_n1579, new_n1580, new_n1581, new_n1582,
    new_n1583, new_n1585, new_n1586, new_n1587, new_n1588, new_n1589,
    new_n1590, new_n1591, new_n1592, new_n1593, new_n1594, new_n1595_1,
    new_n1596, new_n1597_1, new_n1598, new_n1599, new_n1600_1, new_n1601_1,
    new_n1602, new_n1603, new_n1604, new_n1605, new_n1606, new_n1607,
    new_n1608, new_n1609, new_n1610, new_n1611, new_n1612, new_n1613_1,
    new_n1614, new_n1615, new_n1616, new_n1617, new_n1618, new_n1619,
    new_n1620, new_n1621, new_n1622_1, new_n1623, new_n1624, new_n1625,
    new_n1626, new_n1627, new_n1628, new_n1629_1, new_n1630, new_n1631,
    new_n1632, new_n1633_1, new_n1634, new_n1635_1, new_n1636, new_n1637,
    new_n1638, new_n1639, new_n1640, new_n1641, new_n1642_1, new_n1643_1,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1654_1, new_n1655,
    new_n1656, new_n1657_1, new_n1658, new_n1659, new_n1660_1, new_n1661,
    new_n1662, new_n1663, new_n1664, new_n1665, new_n1666, new_n1667,
    new_n1668, new_n1669, new_n1670, new_n1671, new_n1672, new_n1673,
    new_n1674, new_n1675_1, new_n1676, new_n1677_1, new_n1678_1, new_n1679,
    new_n1680, new_n1681, new_n1682, new_n1683_1, new_n1684, new_n1685,
    new_n1686_1, new_n1687, new_n1688_1, new_n1689, new_n1690_1, new_n1691,
    new_n1692, new_n1693, new_n1694, new_n1695, new_n1696, new_n1697,
    new_n1698, new_n1699, new_n1700, new_n1701, new_n1703, new_n1706,
    new_n1707_1, new_n1708, new_n1709, new_n1710, new_n1711, new_n1713,
    new_n1717, new_n1719, new_n1722, new_n1723, new_n1724, new_n1725,
    new_n1726, new_n1727_1, new_n1729_1, new_n1730, new_n1731_1, new_n1732,
    new_n1733, new_n1736, new_n1738, new_n1740, new_n1741, new_n1742,
    new_n1743_1, new_n1744, new_n1745, new_n1746_1, new_n1747_1, new_n1748,
    new_n1749, new_n1750, new_n1751, new_n1752, new_n1753, new_n1754,
    new_n1755, new_n1756, new_n1757_1, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763_1, new_n1764_1, new_n1765, new_n1766,
    new_n1767, new_n1768, new_n1769, new_n1770, new_n1771, new_n1772,
    new_n1773, new_n1774, new_n1776, new_n1779, new_n1782, new_n1783,
    new_n1785, new_n1787, new_n1789, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1796, new_n1798, new_n1799, new_n1800, new_n1801,
    new_n1802, new_n1803, new_n1804, new_n1805, new_n1807, new_n1809,
    new_n1812, new_n1814, new_n1816, new_n1817, new_n1818, new_n1820,
    new_n1822, new_n1824, new_n1825, new_n1826, new_n1827, new_n1828,
    new_n1830, new_n1832, new_n1833, new_n1834, new_n1835, new_n1836,
    new_n1837, new_n1838, new_n1839, new_n1840, new_n1841, new_n1842,
    new_n1843, new_n1844, new_n1845, new_n1846, new_n1847, new_n1848,
    new_n1849, new_n1850, new_n1851, new_n1852, new_n1853, new_n1854,
    new_n1855, new_n1856, new_n1858, new_n1859, new_n1860, new_n1863,
    new_n1864, new_n1867, new_n1870, new_n1873, new_n1875, new_n1876,
    new_n1877, new_n1878, new_n1880, new_n1882, new_n1883, new_n1885,
    new_n1887, new_n1889, new_n1891, new_n1892, new_n1893, new_n1894,
    new_n1895, new_n1897, new_n1899, new_n1901, new_n1905, new_n1906,
    new_n1907, new_n1908, new_n1910, new_n1911, new_n1913, new_n1914,
    new_n1915, new_n1916, new_n1918, new_n1919, new_n1921, new_n1923,
    new_n1924, new_n1925, new_n1926, new_n1927, new_n1928, new_n1929,
    new_n1930, new_n1931, new_n1932, new_n1933, new_n1934, new_n1935,
    new_n1936, new_n1937, new_n1938, new_n1939, new_n1943, new_n1945,
    new_n1946, new_n1949, new_n1952, new_n1953, new_n1954, new_n1955,
    new_n1957, new_n1959, new_n1961, new_n1962, new_n1963, new_n1965,
    new_n1966, new_n1969, new_n1970, new_n1972, new_n1974, new_n1976,
    new_n1978, new_n1980, new_n1982, new_n1983, new_n1984, new_n1986,
    new_n1987, new_n1989, new_n1991, new_n1993, new_n1995, new_n1996,
    new_n1998, new_n2002, new_n2004, new_n2005, new_n2006, new_n2007,
    new_n2009, new_n2012, new_n2014, new_n2016, new_n2018, new_n2021,
    new_n2024, new_n2025, new_n2027, new_n2029, new_n2030, new_n2033,
    new_n2034, new_n2035, new_n2036, new_n2038, new_n2042, new_n2043,
    new_n2045, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2055, new_n2057, new_n2059, new_n2060, new_n2061, new_n2063,
    new_n2064, new_n2065;
  not_13 g0000(.A(n36), .Y(new_n276_1));
  not_13 g0001(.A(n1643), .Y(new_n277_1));
  and_7  g0002(.A(new_n277_1), .B(new_n276_1), .Y(new_n278));
  xor_5  g0003(.A(n1643), .B(n36), .Y(new_n279));
  or_2   g0004(.A(n788), .B(n555), .Y(new_n280));
  not_13 g0005(.A(new_n280), .Y(new_n281));
  and_7  g0006(.A(n788), .B(n555), .Y(new_n282));
  not_13 g0007(.A(new_n282), .Y(new_n283));
  and_7  g0008(.A(new_n283), .B(new_n280), .Y(new_n284));
  not_13 g0009(.A(n353), .Y(new_n285));
  not_13 g0010(.A(n747), .Y(new_n286));
  and_7  g0011(.A(new_n286), .B(new_n285), .Y(new_n287));
  xor_5  g0012(.A(n747), .B(new_n285), .Y(new_n288));
  or_2   g0013(.A(n952), .B(n329), .Y(new_n289));
  and_7  g0014(.A(n1145), .B(n931), .Y(new_n290_1));
  nor_6  g0015(.A(n952), .B(n329), .Y(new_n291));
  and_7  g0016(.A(n952), .B(n329), .Y(new_n292_1));
  or_2   g0017(.A(new_n292_1), .B(new_n291), .Y(new_n293));
  or_2   g0018(.A(new_n293), .B(new_n290_1), .Y(new_n294));
  and_7  g0019(.A(new_n294), .B(new_n289), .Y(new_n295));
  nor_6  g0020(.A(new_n295), .B(new_n288), .Y(new_n296));
  or_2   g0021(.A(new_n296), .B(new_n287), .Y(new_n297));
  and_7  g0022(.A(new_n297), .B(new_n284), .Y(new_n298));
  or_2   g0023(.A(new_n298), .B(new_n281), .Y(new_n299_1));
  and_7  g0024(.A(new_n299_1), .B(new_n279), .Y(new_n300));
  nor_6  g0025(.A(new_n300), .B(new_n278), .Y(new_n301));
  and_7  g0026(.A(new_n301), .B(n1501), .Y(new_n302));
  and_7  g0027(.A(new_n302), .B(n433), .Y(new_n303_1));
  nor_6  g0028(.A(new_n302), .B(n433), .Y(new_n304));
  nor_6  g0029(.A(new_n304), .B(new_n303_1), .Y(new_n305));
  and_7  g0030(.A(n1000), .B(n870), .Y(new_n306));
  not_13 g0031(.A(n1000), .Y(new_n307));
  and_7  g0032(.A(new_n307), .B(n66), .Y(new_n308));
  nor_6  g0033(.A(new_n308), .B(new_n306), .Y(new_n309));
  and_7  g0034(.A(n1000), .B(n585), .Y(new_n310));
  and_7  g0035(.A(new_n307), .B(n968), .Y(new_n311));
  nor_6  g0036(.A(new_n311), .B(new_n310), .Y(new_n312));
  and_7  g0037(.A(new_n312), .B(new_n309), .Y(new_n313));
  and_7  g0038(.A(n1000), .B(n155), .Y(new_n314));
  not_13 g0039(.A(new_n314), .Y(new_n315));
  not_13 g0040(.A(n1435), .Y(new_n316));
  or_2   g0041(.A(new_n316), .B(n1000), .Y(new_n317_1));
  and_7  g0042(.A(new_n317_1), .B(new_n315), .Y(new_n318));
  and_7  g0043(.A(new_n318), .B(new_n313), .Y(new_n319));
  or_2   g0044(.A(n1000), .B(n682), .Y(new_n320));
  or_2   g0045(.A(n1678), .B(new_n307), .Y(new_n321));
  and_7  g0046(.A(new_n321), .B(new_n320), .Y(new_n322));
  and_7  g0047(.A(new_n322), .B(new_n319), .Y(new_n323));
  xor_5  g0048(.A(n1597), .B(n682), .Y(new_n324));
  nor_6  g0049(.A(new_n324), .B(n1000), .Y(new_n325));
  xor_5  g0050(.A(n1678), .B(n607), .Y(new_n326));
  and_7  g0051(.A(new_n326), .B(n1000), .Y(new_n327));
  nor_6  g0052(.A(new_n327), .B(new_n325), .Y(new_n328));
  and_7  g0053(.A(new_n328), .B(new_n323), .Y(new_n329_1));
  not_13 g0054(.A(new_n323), .Y(new_n330));
  or_2   g0055(.A(new_n327), .B(new_n325), .Y(new_n331));
  and_7  g0056(.A(new_n331), .B(new_n330), .Y(new_n332));
  or_2   g0057(.A(new_n332), .B(new_n329_1), .Y(new_n333));
  not_13 g0058(.A(n682), .Y(new_n334));
  and_7  g0059(.A(new_n307), .B(new_n334), .Y(new_n335));
  not_13 g0060(.A(n1678), .Y(new_n336));
  and_7  g0061(.A(new_n336), .B(n1000), .Y(new_n337));
  or_2   g0062(.A(new_n337), .B(new_n335), .Y(new_n338));
  xor_5  g0063(.A(new_n338), .B(new_n319), .Y(new_n339));
  and_7  g0064(.A(n1435), .B(new_n307), .Y(new_n340));
  or_2   g0065(.A(new_n340), .B(new_n314), .Y(new_n341));
  xor_5  g0066(.A(new_n341), .B(new_n313), .Y(new_n342));
  not_13 g0067(.A(n693), .Y(new_n343));
  xor_5  g0068(.A(new_n312), .B(new_n309), .Y(new_n344));
  and_7  g0069(.A(new_n344), .B(new_n343), .Y(new_n345));
  or_2   g0070(.A(new_n344), .B(new_n343), .Y(new_n346));
  not_13 g0071(.A(n1763), .Y(new_n347_1));
  or_2   g0072(.A(new_n311), .B(new_n310), .Y(new_n348));
  or_2   g0073(.A(new_n348), .B(new_n347_1), .Y(new_n349));
  and_7  g0074(.A(new_n348), .B(new_n347_1), .Y(new_n350));
  not_13 g0075(.A(n1530), .Y(new_n351));
  and_7  g0076(.A(n1461), .B(n1000), .Y(new_n352));
  and_7  g0077(.A(new_n307), .B(n347), .Y(new_n353_1));
  nor_6  g0078(.A(new_n353_1), .B(new_n352), .Y(new_n354));
  or_2   g0079(.A(new_n354), .B(new_n351), .Y(new_n355));
  or_2   g0080(.A(new_n355), .B(new_n350), .Y(new_n356));
  and_7  g0081(.A(new_n356), .B(new_n349), .Y(new_n357));
  and_7  g0082(.A(new_n357), .B(new_n346), .Y(new_n358));
  nor_6  g0083(.A(new_n358), .B(new_n345), .Y(new_n359));
  and_7  g0084(.A(new_n359), .B(new_n342), .Y(new_n360));
  and_7  g0085(.A(new_n360), .B(new_n339), .Y(new_n361));
  and_7  g0086(.A(new_n361), .B(new_n333), .Y(new_n362));
  not_13 g0087(.A(n26), .Y(new_n363));
  and_7  g0088(.A(n1678), .B(n607), .Y(new_n364));
  not_13 g0089(.A(new_n364), .Y(new_n365));
  and_7  g0090(.A(new_n365), .B(new_n363), .Y(new_n366));
  and_7  g0091(.A(n607), .B(n26), .Y(new_n367));
  and_7  g0092(.A(new_n367), .B(n1678), .Y(new_n368));
  or_2   g0093(.A(new_n368), .B(new_n366), .Y(new_n369));
  and_7  g0094(.A(new_n369), .B(n1000), .Y(new_n370));
  or_2   g0095(.A(n1597), .B(n46), .Y(new_n371));
  or_2   g0096(.A(new_n371), .B(n682), .Y(new_n372_1));
  not_13 g0097(.A(n46), .Y(new_n373));
  not_13 g0098(.A(n1597), .Y(new_n374));
  and_7  g0099(.A(new_n374), .B(new_n334), .Y(new_n375));
  or_2   g0100(.A(new_n375), .B(new_n373), .Y(new_n376));
  and_7  g0101(.A(new_n376), .B(new_n372_1), .Y(new_n377));
  and_7  g0102(.A(new_n377), .B(new_n307), .Y(new_n378_1));
  or_2   g0103(.A(new_n378_1), .B(new_n370), .Y(new_n379_1));
  nor_6  g0104(.A(new_n379_1), .B(new_n329_1), .Y(new_n380));
  and_7  g0105(.A(new_n379_1), .B(new_n329_1), .Y(new_n381));
  or_2   g0106(.A(new_n381), .B(new_n380), .Y(new_n382));
  and_7  g0107(.A(new_n382), .B(new_n362), .Y(new_n383));
  nor_6  g0108(.A(new_n382), .B(new_n362), .Y(new_n384));
  nor_6  g0109(.A(new_n384), .B(new_n383), .Y(new_n385));
  and_7  g0110(.A(new_n385), .B(new_n305), .Y(new_n386));
  nor_6  g0111(.A(new_n385), .B(new_n305), .Y(new_n387_1));
  or_2   g0112(.A(new_n387_1), .B(new_n386), .Y(new_n388));
  nor_6  g0113(.A(new_n361), .B(new_n333), .Y(new_n389));
  nor_6  g0114(.A(new_n389), .B(new_n362), .Y(new_n390));
  not_13 g0115(.A(n1501), .Y(new_n391_1));
  or_2   g0116(.A(new_n300), .B(new_n278), .Y(new_n392));
  or_2   g0117(.A(new_n392), .B(new_n391_1), .Y(new_n393));
  or_2   g0118(.A(new_n301), .B(n1501), .Y(new_n394));
  and_7  g0119(.A(new_n394), .B(new_n393), .Y(new_n395));
  nor_6  g0120(.A(new_n395), .B(new_n390), .Y(new_n396));
  and_7  g0121(.A(new_n395), .B(new_n390), .Y(new_n397));
  nor_6  g0122(.A(new_n397), .B(new_n396), .Y(new_n398));
  nor_6  g0123(.A(new_n360), .B(new_n339), .Y(new_n399));
  nor_6  g0124(.A(new_n399), .B(new_n361), .Y(new_n400));
  nor_6  g0125(.A(new_n299_1), .B(new_n279), .Y(new_n401_1));
  or_2   g0126(.A(new_n401_1), .B(new_n300), .Y(new_n402_1));
  and_7  g0127(.A(new_n402_1), .B(new_n400), .Y(new_n403));
  nor_6  g0128(.A(new_n359), .B(new_n342), .Y(new_n404));
  nor_6  g0129(.A(new_n404), .B(new_n360), .Y(new_n405));
  nor_6  g0130(.A(new_n297), .B(new_n284), .Y(new_n406));
  or_2   g0131(.A(new_n406), .B(new_n298), .Y(new_n407));
  nor_6  g0132(.A(new_n407), .B(new_n405), .Y(new_n408));
  and_7  g0133(.A(new_n407), .B(new_n405), .Y(new_n409));
  nor_6  g0134(.A(new_n409), .B(new_n408), .Y(new_n410));
  and_7  g0135(.A(new_n295), .B(new_n288), .Y(new_n411));
  or_2   g0136(.A(new_n411), .B(new_n296), .Y(new_n412));
  xor_5  g0137(.A(n1145), .B(n931), .Y(new_n413));
  xor_5  g0138(.A(new_n354), .B(new_n351), .Y(new_n414_1));
  and_7  g0139(.A(new_n414_1), .B(new_n413), .Y(new_n415));
  not_13 g0140(.A(new_n292_1), .Y(new_n416_1));
  and_7  g0141(.A(new_n416_1), .B(new_n289), .Y(new_n417));
  xor_5  g0142(.A(new_n417), .B(new_n290_1), .Y(new_n418));
  nor_6  g0143(.A(new_n418), .B(new_n415), .Y(new_n419));
  not_13 g0144(.A(n1145), .Y(new_n420));
  xor_5  g0145(.A(new_n420), .B(n931), .Y(new_n421));
  xor_5  g0146(.A(new_n354), .B(n1530), .Y(new_n422));
  or_2   g0147(.A(new_n422), .B(new_n421), .Y(new_n423_1));
  or_2   g0148(.A(new_n423_1), .B(new_n293), .Y(new_n424_1));
  xor_5  g0149(.A(new_n312), .B(new_n347_1), .Y(new_n425));
  and_7  g0150(.A(new_n425), .B(new_n355), .Y(new_n426_1));
  or_2   g0151(.A(new_n353_1), .B(new_n352), .Y(new_n427));
  and_7  g0152(.A(new_n427), .B(n1530), .Y(new_n428));
  xor_5  g0153(.A(new_n312), .B(n1763), .Y(new_n429_1));
  and_7  g0154(.A(new_n429_1), .B(new_n428), .Y(new_n430));
  or_2   g0155(.A(new_n430), .B(new_n426_1), .Y(new_n431));
  and_7  g0156(.A(new_n431), .B(new_n424_1), .Y(new_n432_1));
  nor_6  g0157(.A(new_n432_1), .B(new_n419), .Y(new_n433_1));
  nor_6  g0158(.A(new_n433_1), .B(new_n412), .Y(new_n434));
  and_7  g0159(.A(new_n433_1), .B(new_n412), .Y(new_n435));
  xor_5  g0160(.A(new_n348), .B(new_n309), .Y(new_n436));
  and_7  g0161(.A(new_n436), .B(n693), .Y(new_n437));
  nor_6  g0162(.A(new_n437), .B(new_n345), .Y(new_n438));
  nor_6  g0163(.A(new_n438), .B(new_n357), .Y(new_n439));
  and_7  g0164(.A(new_n438), .B(new_n357), .Y(new_n440));
  or_2   g0165(.A(new_n440), .B(new_n439), .Y(new_n441));
  nor_6  g0166(.A(new_n441), .B(new_n435), .Y(new_n442));
  or_2   g0167(.A(new_n442), .B(new_n434), .Y(new_n443));
  and_7  g0168(.A(new_n443), .B(new_n410), .Y(new_n444_1));
  nor_6  g0169(.A(new_n444_1), .B(new_n408), .Y(new_n445));
  nor_6  g0170(.A(new_n402_1), .B(new_n400), .Y(new_n446));
  nor_6  g0171(.A(new_n446), .B(new_n403), .Y(new_n447));
  and_7  g0172(.A(new_n447), .B(new_n445), .Y(new_n448));
  nor_6  g0173(.A(new_n448), .B(new_n403), .Y(new_n449));
  and_7  g0174(.A(new_n449), .B(new_n398), .Y(new_n450));
  nor_6  g0175(.A(new_n450), .B(new_n396), .Y(new_n451));
  nor_6  g0176(.A(new_n451), .B(new_n388), .Y(new_n452_1));
  and_7  g0177(.A(new_n451), .B(new_n388), .Y(new_n453));
  or_2   g0178(.A(new_n453), .B(new_n452_1), .Y(n19));
  not_13 g0179(.A(n69), .Y(new_n455));
  not_13 g0180(.A(n1381), .Y(new_n456));
  and_7  g0181(.A(new_n456), .B(n402), .Y(new_n457_1));
  nor_6  g0182(.A(new_n457_1), .B(n870), .Y(new_n458));
  not_13 g0183(.A(n66), .Y(new_n459));
  and_7  g0184(.A(new_n457_1), .B(new_n459), .Y(new_n460_1));
  nor_6  g0185(.A(new_n460_1), .B(new_n458), .Y(new_n461));
  xor_5  g0186(.A(new_n461), .B(new_n455), .Y(new_n462));
  nor_6  g0187(.A(new_n457_1), .B(n585), .Y(new_n463));
  not_13 g0188(.A(n968), .Y(new_n464));
  and_7  g0189(.A(new_n457_1), .B(new_n464), .Y(new_n465));
  nor_6  g0190(.A(new_n465), .B(new_n463), .Y(new_n466));
  and_7  g0191(.A(new_n466), .B(n953), .Y(new_n467));
  nor_6  g0192(.A(new_n457_1), .B(n1461), .Y(new_n468));
  not_13 g0193(.A(n347), .Y(new_n469_1));
  and_7  g0194(.A(new_n457_1), .B(new_n469_1), .Y(new_n470));
  nor_6  g0195(.A(new_n470), .B(new_n468), .Y(new_n471));
  and_7  g0196(.A(new_n471), .B(n303), .Y(new_n472_1));
  xor_5  g0197(.A(new_n466), .B(n953), .Y(new_n473));
  and_7  g0198(.A(new_n473), .B(new_n472_1), .Y(new_n474));
  nor_6  g0199(.A(new_n474), .B(new_n467), .Y(new_n475));
  nor_6  g0200(.A(new_n475), .B(new_n462), .Y(new_n476_1));
  and_7  g0201(.A(new_n475), .B(new_n462), .Y(new_n477));
  nor_6  g0202(.A(new_n477), .B(new_n476_1), .Y(new_n478));
  and_7  g0203(.A(new_n478), .B(new_n412), .Y(new_n479));
  nor_6  g0204(.A(new_n478), .B(new_n412), .Y(new_n480));
  or_2   g0205(.A(new_n480), .B(new_n479), .Y(new_n481));
  xor_5  g0206(.A(new_n471), .B(n303), .Y(new_n482_1));
  and_7  g0207(.A(new_n482_1), .B(new_n413), .Y(new_n483));
  nor_6  g0208(.A(new_n483), .B(new_n418), .Y(new_n484));
  nor_6  g0209(.A(new_n473), .B(new_n472_1), .Y(new_n485));
  or_2   g0210(.A(new_n485), .B(new_n474), .Y(new_n486));
  and_7  g0211(.A(new_n483), .B(new_n417), .Y(new_n487));
  nor_6  g0212(.A(new_n487), .B(new_n484), .Y(new_n488_1));
  and_7  g0213(.A(new_n488_1), .B(new_n486), .Y(new_n489));
  nor_6  g0214(.A(new_n489), .B(new_n484), .Y(new_n490));
  and_7  g0215(.A(new_n490), .B(new_n481), .Y(new_n491));
  nor_6  g0216(.A(new_n490), .B(new_n481), .Y(new_n492));
  or_2   g0217(.A(new_n492), .B(new_n491), .Y(n33));
  not_13 g0218(.A(n1642), .Y(new_n494));
  or_2   g0219(.A(n607), .B(n26), .Y(new_n495));
  or_2   g0220(.A(new_n495), .B(n247), .Y(new_n496));
  xor_5  g0221(.A(new_n496), .B(new_n494), .Y(new_n497));
  and_7  g0222(.A(new_n497), .B(n1381), .Y(new_n498_1));
  not_13 g0223(.A(n379), .Y(new_n499));
  not_13 g0224(.A(n1527), .Y(new_n500));
  and_7  g0225(.A(new_n500), .B(new_n373), .Y(new_n501));
  and_7  g0226(.A(new_n501), .B(new_n499), .Y(new_n502));
  not_13 g0227(.A(n402), .Y(new_n503));
  or_2   g0228(.A(n1527), .B(n46), .Y(new_n504));
  and_7  g0229(.A(new_n504), .B(n379), .Y(new_n505));
  or_2   g0230(.A(new_n505), .B(new_n503), .Y(new_n506));
  or_2   g0231(.A(new_n506), .B(new_n502), .Y(new_n507));
  and_7  g0232(.A(n1642), .B(new_n456), .Y(new_n508));
  or_2   g0233(.A(new_n508), .B(new_n457_1), .Y(new_n509));
  and_7  g0234(.A(new_n509), .B(new_n507), .Y(new_n510_1));
  or_2   g0235(.A(new_n510_1), .B(new_n498_1), .Y(new_n511));
  not_13 g0236(.A(n247), .Y(new_n512));
  xor_5  g0237(.A(new_n495), .B(new_n512), .Y(new_n513));
  and_7  g0238(.A(new_n513), .B(n1381), .Y(new_n514));
  and_7  g0239(.A(n1527), .B(n46), .Y(new_n515));
  not_13 g0240(.A(new_n515), .Y(new_n516));
  and_7  g0241(.A(new_n516), .B(n402), .Y(new_n517_1));
  and_7  g0242(.A(new_n517_1), .B(new_n504), .Y(new_n518));
  not_13 g0243(.A(new_n518), .Y(new_n519));
  and_7  g0244(.A(new_n456), .B(n247), .Y(new_n520));
  or_2   g0245(.A(new_n520), .B(new_n457_1), .Y(new_n521));
  and_7  g0246(.A(new_n521), .B(new_n519), .Y(new_n522_1));
  or_2   g0247(.A(new_n522_1), .B(new_n514), .Y(new_n523));
  or_2   g0248(.A(n1381), .B(new_n503), .Y(new_n524));
  and_7  g0249(.A(new_n524), .B(new_n336), .Y(new_n525));
  and_7  g0250(.A(new_n457_1), .B(new_n334), .Y(new_n526));
  or_2   g0251(.A(new_n526), .B(new_n525), .Y(new_n527));
  and_7  g0252(.A(new_n527), .B(new_n277_1), .Y(new_n528));
  xor_5  g0253(.A(new_n527), .B(new_n277_1), .Y(new_n529));
  nor_6  g0254(.A(new_n457_1), .B(n155), .Y(new_n530));
  and_7  g0255(.A(new_n457_1), .B(new_n316), .Y(new_n531));
  or_2   g0256(.A(new_n531), .B(new_n530), .Y(new_n532_1));
  not_13 g0257(.A(new_n532_1), .Y(new_n533));
  and_7  g0258(.A(new_n533), .B(n555), .Y(new_n534_1));
  or_2   g0259(.A(new_n461), .B(n353), .Y(new_n535));
  xor_5  g0260(.A(new_n461), .B(new_n285), .Y(new_n536));
  or_2   g0261(.A(new_n466), .B(n952), .Y(new_n537));
  and_7  g0262(.A(new_n471), .B(n1145), .Y(new_n538));
  not_13 g0263(.A(n952), .Y(new_n539));
  xor_5  g0264(.A(new_n466), .B(new_n539), .Y(new_n540));
  or_2   g0265(.A(new_n540), .B(new_n538), .Y(new_n541_1));
  and_7  g0266(.A(new_n541_1), .B(new_n537), .Y(new_n542));
  or_2   g0267(.A(new_n542), .B(new_n536), .Y(new_n543));
  and_7  g0268(.A(new_n543), .B(new_n535), .Y(new_n544));
  not_13 g0269(.A(n555), .Y(new_n545));
  xor_5  g0270(.A(new_n532_1), .B(new_n545), .Y(new_n546));
  and_7  g0271(.A(new_n546), .B(new_n544), .Y(new_n547_1));
  nor_6  g0272(.A(new_n547_1), .B(new_n534_1), .Y(new_n548));
  and_7  g0273(.A(new_n548), .B(new_n529), .Y(new_n549_1));
  nor_6  g0274(.A(new_n549_1), .B(new_n528), .Y(new_n550));
  and_7  g0275(.A(n1381), .B(n607), .Y(new_n551));
  and_7  g0276(.A(new_n374), .B(n402), .Y(new_n552));
  not_13 g0277(.A(n607), .Y(new_n553));
  and_7  g0278(.A(new_n553), .B(new_n503), .Y(new_n554));
  or_2   g0279(.A(new_n554), .B(new_n552), .Y(new_n555_1));
  and_7  g0280(.A(new_n555_1), .B(new_n456), .Y(new_n556));
  or_2   g0281(.A(new_n556), .B(new_n551), .Y(new_n557_1));
  not_13 g0282(.A(new_n557_1), .Y(new_n558));
  and_7  g0283(.A(new_n558), .B(new_n550), .Y(new_n559_1));
  and_7  g0284(.A(n402), .B(n46), .Y(new_n560));
  and_7  g0285(.A(new_n503), .B(new_n363), .Y(new_n561));
  or_2   g0286(.A(new_n561), .B(new_n560), .Y(new_n562));
  and_7  g0287(.A(new_n562), .B(new_n456), .Y(new_n563));
  not_13 g0288(.A(new_n367), .Y(new_n564));
  and_7  g0289(.A(new_n495), .B(new_n564), .Y(new_n565));
  and_7  g0290(.A(new_n565), .B(n1381), .Y(new_n566));
  or_2   g0291(.A(new_n566), .B(new_n563), .Y(new_n567));
  not_13 g0292(.A(new_n567), .Y(new_n568));
  and_7  g0293(.A(new_n568), .B(new_n559_1), .Y(new_n569_1));
  and_7  g0294(.A(new_n569_1), .B(new_n523), .Y(new_n570));
  xor_5  g0295(.A(new_n570), .B(new_n511), .Y(n1731));
  nor_6  g0296(.A(new_n522_1), .B(new_n514), .Y(new_n572));
  or_2   g0297(.A(new_n549_1), .B(new_n528), .Y(new_n573_1));
  or_2   g0298(.A(new_n557_1), .B(new_n573_1), .Y(new_n574));
  or_2   g0299(.A(new_n567), .B(new_n574), .Y(new_n575));
  or_2   g0300(.A(new_n575), .B(new_n572), .Y(new_n576));
  or_2   g0301(.A(new_n569_1), .B(new_n523), .Y(new_n577));
  and_7  g0302(.A(new_n577), .B(new_n576), .Y(n1138));
  or_2   g0303(.A(new_n558), .B(new_n550), .Y(new_n579));
  and_7  g0304(.A(new_n579), .B(new_n574), .Y(n1727));
  nor_6  g0305(.A(new_n540), .B(new_n538), .Y(new_n581));
  and_7  g0306(.A(new_n540), .B(new_n538), .Y(new_n582));
  or_2   g0307(.A(new_n582), .B(new_n581), .Y(n1457));
  xor_5  g0308(.A(new_n471), .B(n1145), .Y(n1183));
  or_2   g0309(.A(n1183), .B(n1457), .Y(new_n585_1));
  not_13 g0310(.A(new_n537), .Y(new_n586));
  or_2   g0311(.A(new_n581), .B(new_n586), .Y(new_n587));
  xor_5  g0312(.A(new_n587), .B(new_n536), .Y(n416));
  or_2   g0313(.A(n416), .B(new_n585_1), .Y(new_n589));
  nor_6  g0314(.A(new_n546), .B(new_n544), .Y(new_n590));
  nor_6  g0315(.A(new_n590), .B(new_n547_1), .Y(n1721));
  nor_6  g0316(.A(n1721), .B(new_n589), .Y(new_n592));
  nor_6  g0317(.A(new_n548), .B(new_n529), .Y(new_n593));
  nor_6  g0318(.A(new_n593), .B(new_n549_1), .Y(new_n594));
  nor_6  g0319(.A(new_n594), .B(new_n592), .Y(new_n595));
  and_7  g0320(.A(new_n595), .B(n1727), .Y(new_n596));
  and_7  g0321(.A(new_n596), .B(new_n568), .Y(new_n597));
  and_7  g0322(.A(new_n597), .B(n1138), .Y(new_n598));
  nor_6  g0323(.A(new_n598), .B(n1731), .Y(new_n599_1));
  and_7  g0324(.A(new_n598), .B(new_n511), .Y(new_n600_1));
  nor_6  g0325(.A(new_n600_1), .B(new_n599_1), .Y(n44));
  xor_5  g0326(.A(new_n414_1), .B(new_n413), .Y(n55));
  not_13 g0327(.A(n1707), .Y(new_n603));
  and_7  g0328(.A(new_n603), .B(new_n277_1), .Y(new_n604));
  not_13 g0329(.A(new_n604), .Y(new_n605));
  xor_5  g0330(.A(n1707), .B(new_n277_1), .Y(new_n606));
  not_13 g0331(.A(n1140), .Y(new_n607_1));
  and_7  g0332(.A(new_n607_1), .B(new_n545), .Y(new_n608));
  xor_5  g0333(.A(n1140), .B(n555), .Y(new_n609));
  not_13 g0334(.A(n1351), .Y(new_n610));
  and_7  g0335(.A(new_n610), .B(new_n285), .Y(new_n611));
  xor_5  g0336(.A(n1351), .B(new_n285), .Y(new_n612));
  or_2   g0337(.A(n952), .B(n729), .Y(new_n613));
  and_7  g0338(.A(n1145), .B(n684), .Y(new_n614));
  not_13 g0339(.A(n729), .Y(new_n615));
  xor_5  g0340(.A(n952), .B(new_n615), .Y(new_n616));
  or_2   g0341(.A(new_n616), .B(new_n614), .Y(new_n617));
  and_7  g0342(.A(new_n617), .B(new_n613), .Y(new_n618));
  nor_6  g0343(.A(new_n618), .B(new_n612), .Y(new_n619));
  or_2   g0344(.A(new_n619), .B(new_n611), .Y(new_n620));
  and_7  g0345(.A(new_n620), .B(new_n609), .Y(new_n621));
  nor_6  g0346(.A(new_n621), .B(new_n608), .Y(new_n622));
  or_2   g0347(.A(new_n622), .B(new_n606), .Y(new_n623));
  and_7  g0348(.A(new_n623), .B(new_n605), .Y(new_n624));
  and_7  g0349(.A(new_n624), .B(n1332), .Y(new_n625));
  and_7  g0350(.A(new_n625), .B(n391), .Y(new_n626));
  and_7  g0351(.A(new_n626), .B(n1544), .Y(new_n627_1));
  not_13 g0352(.A(n1544), .Y(new_n628));
  not_13 g0353(.A(n391), .Y(new_n629));
  not_13 g0354(.A(n1332), .Y(new_n630));
  and_7  g0355(.A(n1707), .B(n1643), .Y(new_n631));
  not_13 g0356(.A(new_n631), .Y(new_n632));
  and_7  g0357(.A(new_n632), .B(new_n605), .Y(new_n633));
  or_2   g0358(.A(new_n621), .B(new_n608), .Y(new_n634));
  and_7  g0359(.A(new_n634), .B(new_n633), .Y(new_n635));
  or_2   g0360(.A(new_n635), .B(new_n604), .Y(new_n636));
  or_2   g0361(.A(new_n636), .B(new_n630), .Y(new_n637));
  or_2   g0362(.A(new_n637), .B(new_n629), .Y(new_n638_1));
  and_7  g0363(.A(new_n638_1), .B(new_n628), .Y(new_n639));
  nor_6  g0364(.A(new_n639), .B(new_n627_1), .Y(new_n640));
  and_7  g0365(.A(n266), .B(n155), .Y(new_n641));
  not_13 g0366(.A(n266), .Y(new_n642));
  and_7  g0367(.A(n1435), .B(new_n642), .Y(new_n643_1));
  nor_6  g0368(.A(new_n643_1), .B(new_n641), .Y(new_n644));
  and_7  g0369(.A(n870), .B(n266), .Y(new_n645));
  and_7  g0370(.A(new_n642), .B(n66), .Y(new_n646_1));
  nor_6  g0371(.A(new_n646_1), .B(new_n645), .Y(new_n647_1));
  and_7  g0372(.A(new_n647_1), .B(new_n644), .Y(new_n648_1));
  and_7  g0373(.A(n1678), .B(n266), .Y(new_n649_1));
  not_13 g0374(.A(new_n649_1), .Y(new_n650));
  or_2   g0375(.A(new_n334), .B(n266), .Y(new_n651));
  and_7  g0376(.A(new_n651), .B(new_n650), .Y(new_n652));
  and_7  g0377(.A(new_n652), .B(new_n648_1), .Y(new_n653_1));
  and_7  g0378(.A(n1597), .B(new_n642), .Y(new_n654));
  and_7  g0379(.A(new_n553), .B(n266), .Y(new_n655_1));
  or_2   g0380(.A(new_n655_1), .B(new_n654), .Y(new_n656));
  and_7  g0381(.A(new_n656), .B(new_n653_1), .Y(new_n657));
  and_7  g0382(.A(n266), .B(new_n363), .Y(new_n658));
  not_13 g0383(.A(new_n658), .Y(new_n659));
  xor_5  g0384(.A(n1597), .B(new_n373), .Y(new_n660));
  or_2   g0385(.A(new_n660), .B(n266), .Y(new_n661));
  and_7  g0386(.A(new_n661), .B(new_n659), .Y(new_n662));
  xor_5  g0387(.A(new_n662), .B(new_n657), .Y(new_n663));
  or_2   g0388(.A(new_n374), .B(n266), .Y(new_n664));
  or_2   g0389(.A(n607), .B(new_n642), .Y(new_n665_1));
  and_7  g0390(.A(new_n665_1), .B(new_n664), .Y(new_n666));
  xor_5  g0391(.A(new_n666), .B(new_n653_1), .Y(new_n667));
  and_7  g0392(.A(n682), .B(new_n642), .Y(new_n668));
  or_2   g0393(.A(new_n668), .B(new_n649_1), .Y(new_n669));
  xor_5  g0394(.A(new_n669), .B(new_n648_1), .Y(new_n670));
  or_2   g0395(.A(new_n643_1), .B(new_n641), .Y(new_n671));
  xor_5  g0396(.A(new_n647_1), .B(new_n671), .Y(new_n672));
  and_7  g0397(.A(new_n672), .B(n223), .Y(new_n673));
  not_13 g0398(.A(n223), .Y(new_n674));
  xor_5  g0399(.A(new_n647_1), .B(new_n644), .Y(new_n675_1));
  and_7  g0400(.A(new_n675_1), .B(new_n674), .Y(new_n676));
  or_2   g0401(.A(new_n676), .B(new_n673), .Y(new_n677));
  and_7  g0402(.A(new_n647_1), .B(n444), .Y(new_n678));
  and_7  g0403(.A(n585), .B(n266), .Y(new_n679));
  and_7  g0404(.A(n968), .B(new_n642), .Y(new_n680));
  or_2   g0405(.A(new_n680), .B(new_n679), .Y(new_n681));
  or_2   g0406(.A(new_n681), .B(n472), .Y(new_n682_1));
  and_7  g0407(.A(n1461), .B(n266), .Y(new_n683_1));
  and_7  g0408(.A(n347), .B(new_n642), .Y(new_n684_1));
  or_2   g0409(.A(new_n684_1), .B(new_n683_1), .Y(new_n685));
  and_7  g0410(.A(new_n685), .B(n801), .Y(new_n686));
  not_13 g0411(.A(new_n679), .Y(new_n687));
  or_2   g0412(.A(new_n464), .B(n266), .Y(new_n688));
  and_7  g0413(.A(new_n688), .B(new_n687), .Y(new_n689));
  xor_5  g0414(.A(new_n689), .B(n472), .Y(new_n690));
  or_2   g0415(.A(new_n690), .B(new_n686), .Y(new_n691));
  and_7  g0416(.A(new_n691), .B(new_n682_1), .Y(new_n692));
  xor_5  g0417(.A(new_n647_1), .B(n444), .Y(new_n693_1));
  and_7  g0418(.A(new_n693_1), .B(new_n692), .Y(new_n694));
  nor_6  g0419(.A(new_n694), .B(new_n678), .Y(new_n695_1));
  nor_6  g0420(.A(new_n695_1), .B(new_n677), .Y(new_n696));
  or_2   g0421(.A(new_n696), .B(new_n673), .Y(new_n697));
  and_7  g0422(.A(new_n697), .B(new_n670), .Y(new_n698));
  and_7  g0423(.A(new_n698), .B(new_n667), .Y(new_n699_1));
  and_7  g0424(.A(new_n699_1), .B(new_n663), .Y(new_n700));
  nor_6  g0425(.A(new_n660), .B(n266), .Y(new_n701));
  or_2   g0426(.A(new_n701), .B(new_n658), .Y(new_n702));
  and_7  g0427(.A(new_n702), .B(new_n657), .Y(new_n703));
  or_2   g0428(.A(new_n504), .B(n1597), .Y(new_n704));
  and_7  g0429(.A(new_n374), .B(new_n373), .Y(new_n705));
  or_2   g0430(.A(new_n705), .B(new_n500), .Y(new_n706));
  and_7  g0431(.A(new_n706), .B(new_n704), .Y(new_n707));
  and_7  g0432(.A(new_n707), .B(new_n642), .Y(new_n708));
  and_7  g0433(.A(n266), .B(new_n512), .Y(new_n709));
  nor_6  g0434(.A(new_n709), .B(new_n708), .Y(new_n710));
  xor_5  g0435(.A(new_n710), .B(new_n703), .Y(new_n711));
  and_7  g0436(.A(new_n711), .B(new_n700), .Y(new_n712_1));
  nor_6  g0437(.A(new_n711), .B(new_n700), .Y(new_n713));
  nor_6  g0438(.A(new_n713), .B(new_n712_1), .Y(new_n714));
  nor_6  g0439(.A(new_n714), .B(new_n640), .Y(new_n715_1));
  and_7  g0440(.A(new_n714), .B(new_n640), .Y(new_n716));
  or_2   g0441(.A(new_n716), .B(new_n715_1), .Y(new_n717));
  or_2   g0442(.A(new_n625), .B(n391), .Y(new_n718));
  and_7  g0443(.A(new_n718), .B(new_n638_1), .Y(new_n719));
  nor_6  g0444(.A(new_n699_1), .B(new_n663), .Y(new_n720));
  nor_6  g0445(.A(new_n720), .B(new_n700), .Y(new_n721));
  nor_6  g0446(.A(new_n721), .B(new_n719), .Y(new_n722));
  xor_5  g0447(.A(new_n656), .B(new_n653_1), .Y(new_n723));
  xor_5  g0448(.A(new_n652), .B(new_n648_1), .Y(new_n724_1));
  nor_6  g0449(.A(new_n696), .B(new_n673), .Y(new_n725_1));
  or_2   g0450(.A(new_n725_1), .B(new_n724_1), .Y(new_n726));
  and_7  g0451(.A(new_n726), .B(new_n723), .Y(new_n727));
  nor_6  g0452(.A(new_n727), .B(new_n699_1), .Y(new_n728));
  and_7  g0453(.A(new_n636), .B(new_n630), .Y(new_n729_1));
  nor_6  g0454(.A(new_n729_1), .B(new_n625), .Y(new_n730));
  or_2   g0455(.A(new_n730), .B(new_n728), .Y(new_n731_1));
  nor_6  g0456(.A(new_n730), .B(new_n728), .Y(new_n732));
  and_7  g0457(.A(new_n730), .B(new_n728), .Y(new_n733));
  or_2   g0458(.A(new_n733), .B(new_n732), .Y(new_n734));
  and_7  g0459(.A(new_n725_1), .B(new_n724_1), .Y(new_n735));
  nor_6  g0460(.A(new_n735), .B(new_n698), .Y(new_n736));
  and_7  g0461(.A(new_n622), .B(new_n606), .Y(new_n737));
  or_2   g0462(.A(new_n737), .B(new_n635), .Y(new_n738_1));
  nor_6  g0463(.A(new_n738_1), .B(new_n736), .Y(new_n739));
  and_7  g0464(.A(new_n738_1), .B(new_n736), .Y(new_n740));
  nor_6  g0465(.A(new_n740), .B(new_n739), .Y(new_n741));
  and_7  g0466(.A(new_n695_1), .B(new_n677), .Y(new_n742));
  nor_6  g0467(.A(new_n742), .B(new_n696), .Y(new_n743));
  nor_6  g0468(.A(new_n620), .B(new_n609), .Y(new_n744));
  or_2   g0469(.A(new_n744), .B(new_n621), .Y(new_n745));
  nor_6  g0470(.A(new_n745), .B(new_n743), .Y(new_n746));
  and_7  g0471(.A(new_n745), .B(new_n743), .Y(new_n747_1));
  or_2   g0472(.A(new_n747_1), .B(new_n746), .Y(new_n748_1));
  nor_6  g0473(.A(new_n693_1), .B(new_n692), .Y(new_n749));
  nor_6  g0474(.A(new_n749), .B(new_n694), .Y(new_n750));
  and_7  g0475(.A(new_n618), .B(new_n612), .Y(new_n751));
  or_2   g0476(.A(new_n751), .B(new_n619), .Y(new_n752));
  nor_6  g0477(.A(new_n752), .B(new_n750), .Y(new_n753));
  not_13 g0478(.A(new_n614), .Y(new_n754));
  and_7  g0479(.A(n952), .B(n729), .Y(new_n755));
  not_13 g0480(.A(new_n755), .Y(new_n756));
  and_7  g0481(.A(new_n756), .B(new_n613), .Y(new_n757));
  or_2   g0482(.A(new_n757), .B(new_n754), .Y(new_n758));
  and_7  g0483(.A(new_n757), .B(new_n754), .Y(new_n759_1));
  xor_5  g0484(.A(n1145), .B(n684), .Y(new_n760));
  xor_5  g0485(.A(new_n685), .B(n801), .Y(new_n761_1));
  and_7  g0486(.A(new_n761_1), .B(new_n760), .Y(new_n762));
  nor_6  g0487(.A(new_n762), .B(new_n759_1), .Y(new_n763));
  and_7  g0488(.A(new_n763), .B(new_n758), .Y(new_n764));
  not_13 g0489(.A(new_n686), .Y(new_n765));
  xor_5  g0490(.A(new_n681), .B(n472), .Y(new_n766));
  or_2   g0491(.A(new_n766), .B(new_n765), .Y(new_n767));
  and_7  g0492(.A(new_n767), .B(new_n691), .Y(new_n768));
  and_7  g0493(.A(new_n762), .B(new_n757), .Y(new_n769));
  nor_6  g0494(.A(new_n769), .B(new_n764), .Y(new_n770_1));
  and_7  g0495(.A(new_n770_1), .B(new_n768), .Y(new_n771));
  or_2   g0496(.A(new_n771), .B(new_n764), .Y(new_n772));
  and_7  g0497(.A(new_n752), .B(new_n750), .Y(new_n773_1));
  nor_6  g0498(.A(new_n773_1), .B(new_n753), .Y(new_n774));
  and_7  g0499(.A(new_n774), .B(new_n772), .Y(new_n775));
  nor_6  g0500(.A(new_n775), .B(new_n753), .Y(new_n776));
  nor_6  g0501(.A(new_n776), .B(new_n748_1), .Y(new_n777));
  or_2   g0502(.A(new_n777), .B(new_n746), .Y(new_n778));
  and_7  g0503(.A(new_n778), .B(new_n741), .Y(new_n779));
  nor_6  g0504(.A(new_n779), .B(new_n739), .Y(new_n780));
  or_2   g0505(.A(new_n780), .B(new_n734), .Y(new_n781));
  and_7  g0506(.A(new_n781), .B(new_n731_1), .Y(new_n782));
  and_7  g0507(.A(new_n721), .B(new_n719), .Y(new_n783));
  or_2   g0508(.A(new_n783), .B(new_n722), .Y(new_n784));
  nor_6  g0509(.A(new_n784), .B(new_n782), .Y(new_n785));
  or_2   g0510(.A(new_n785), .B(new_n722), .Y(new_n786));
  xor_5  g0511(.A(new_n786), .B(new_n717), .Y(n56));
  or_2   g0512(.A(new_n709), .B(new_n708), .Y(new_n788_1));
  and_7  g0513(.A(new_n788_1), .B(new_n703), .Y(new_n789));
  and_7  g0514(.A(new_n494), .B(n266), .Y(new_n790_1));
  not_13 g0515(.A(new_n790_1), .Y(new_n791));
  xor_5  g0516(.A(new_n704), .B(new_n499), .Y(new_n792_1));
  or_2   g0517(.A(new_n792_1), .B(n266), .Y(new_n793));
  and_7  g0518(.A(new_n793), .B(new_n791), .Y(new_n794));
  xor_5  g0519(.A(new_n794), .B(new_n789), .Y(new_n795));
  and_7  g0520(.A(new_n795), .B(new_n712_1), .Y(new_n796));
  nor_6  g0521(.A(new_n792_1), .B(n266), .Y(new_n797));
  or_2   g0522(.A(new_n797), .B(new_n790_1), .Y(new_n798));
  and_7  g0523(.A(new_n798), .B(new_n789), .Y(new_n799));
  not_13 g0524(.A(n171), .Y(new_n800));
  and_7  g0525(.A(n266), .B(new_n800), .Y(new_n801_1));
  not_13 g0526(.A(new_n801_1), .Y(new_n802));
  or_2   g0527(.A(new_n704), .B(n379), .Y(new_n803));
  and_7  g0528(.A(new_n803), .B(n1263), .Y(new_n804));
  not_13 g0529(.A(n1263), .Y(new_n805));
  and_7  g0530(.A(new_n501), .B(new_n374), .Y(new_n806));
  and_7  g0531(.A(new_n806), .B(new_n499), .Y(new_n807));
  and_7  g0532(.A(new_n807), .B(new_n805), .Y(new_n808));
  or_2   g0533(.A(new_n808), .B(n266), .Y(new_n809));
  or_2   g0534(.A(new_n809), .B(new_n804), .Y(new_n810));
  and_7  g0535(.A(new_n810), .B(new_n802), .Y(new_n811));
  xor_5  g0536(.A(new_n811), .B(new_n799), .Y(new_n812));
  and_7  g0537(.A(new_n812), .B(new_n796), .Y(new_n813_1));
  not_13 g0538(.A(new_n804), .Y(new_n814));
  or_2   g0539(.A(new_n803), .B(n1263), .Y(new_n815));
  and_7  g0540(.A(new_n815), .B(new_n642), .Y(new_n816));
  and_7  g0541(.A(new_n816), .B(new_n814), .Y(new_n817));
  or_2   g0542(.A(new_n817), .B(new_n801_1), .Y(new_n818));
  and_7  g0543(.A(new_n818), .B(new_n799), .Y(new_n819));
  and_7  g0544(.A(n557), .B(n266), .Y(new_n820));
  not_13 g0545(.A(n1422), .Y(new_n821));
  and_7  g0546(.A(new_n808), .B(new_n821), .Y(new_n822));
  and_7  g0547(.A(new_n822), .B(new_n642), .Y(new_n823_1));
  and_7  g0548(.A(new_n816), .B(n1422), .Y(new_n824_1));
  or_2   g0549(.A(new_n824_1), .B(new_n823_1), .Y(new_n825));
  or_2   g0550(.A(new_n825), .B(new_n820), .Y(new_n826));
  xor_5  g0551(.A(new_n826), .B(new_n819), .Y(new_n827));
  and_7  g0552(.A(new_n827), .B(new_n813_1), .Y(new_n828));
  nor_6  g0553(.A(new_n827), .B(new_n813_1), .Y(new_n829));
  or_2   g0554(.A(new_n829), .B(new_n828), .Y(new_n830));
  and_7  g0555(.A(new_n627_1), .B(n649), .Y(new_n831));
  nor_6  g0556(.A(new_n812), .B(new_n796), .Y(new_n832));
  nor_6  g0557(.A(new_n832), .B(new_n813_1), .Y(new_n833));
  nor_6  g0558(.A(new_n833), .B(new_n831), .Y(new_n834));
  and_7  g0559(.A(new_n833), .B(new_n831), .Y(new_n835));
  or_2   g0560(.A(new_n835), .B(new_n834), .Y(new_n836_1));
  not_13 g0561(.A(n649), .Y(new_n837));
  or_2   g0562(.A(new_n638_1), .B(new_n628), .Y(new_n838));
  or_2   g0563(.A(new_n838), .B(new_n837), .Y(new_n839_1));
  or_2   g0564(.A(new_n627_1), .B(n649), .Y(new_n840));
  and_7  g0565(.A(new_n840), .B(new_n839_1), .Y(new_n841));
  nor_6  g0566(.A(new_n795), .B(new_n712_1), .Y(new_n842));
  nor_6  g0567(.A(new_n842), .B(new_n796), .Y(new_n843));
  nor_6  g0568(.A(new_n843), .B(new_n841), .Y(new_n844));
  and_7  g0569(.A(new_n843), .B(new_n841), .Y(new_n845));
  or_2   g0570(.A(new_n845), .B(new_n844), .Y(new_n846_1));
  or_2   g0571(.A(new_n714), .B(new_n640), .Y(new_n847));
  nor_6  g0572(.A(new_n785), .B(new_n722), .Y(new_n848));
  or_2   g0573(.A(new_n848), .B(new_n717), .Y(new_n849));
  and_7  g0574(.A(new_n849), .B(new_n847), .Y(new_n850));
  nor_6  g0575(.A(new_n850), .B(new_n846_1), .Y(new_n851));
  nor_6  g0576(.A(new_n851), .B(new_n844), .Y(new_n852));
  nor_6  g0577(.A(new_n852), .B(new_n836_1), .Y(new_n853));
  or_2   g0578(.A(new_n853), .B(new_n834), .Y(new_n854));
  or_2   g0579(.A(new_n854), .B(new_n830), .Y(new_n855));
  nor_6  g0580(.A(new_n829), .B(new_n828), .Y(new_n856));
  or_2   g0581(.A(new_n833), .B(new_n831), .Y(new_n857));
  or_2   g0582(.A(new_n852), .B(new_n836_1), .Y(new_n858_1));
  and_7  g0583(.A(new_n858_1), .B(new_n857), .Y(new_n859));
  or_2   g0584(.A(new_n859), .B(new_n856), .Y(new_n860));
  and_7  g0585(.A(new_n860), .B(new_n855), .Y(n67));
  not_13 g0586(.A(n469), .Y(new_n862_1));
  xor_5  g0587(.A(n1643), .B(new_n862_1), .Y(new_n863));
  not_13 g0588(.A(n927), .Y(new_n864));
  and_7  g0589(.A(new_n864), .B(new_n545), .Y(new_n865_1));
  not_13 g0590(.A(new_n865_1), .Y(new_n866));
  xor_5  g0591(.A(n927), .B(new_n545), .Y(new_n867_1));
  not_13 g0592(.A(n655), .Y(new_n868));
  and_7  g0593(.A(new_n868), .B(new_n285), .Y(new_n869));
  not_13 g0594(.A(new_n869), .Y(new_n870_1));
  xor_5  g0595(.A(n655), .B(new_n285), .Y(new_n871));
  or_2   g0596(.A(n952), .B(n653), .Y(new_n872));
  and_7  g0597(.A(n1764), .B(n1145), .Y(new_n873));
  not_13 g0598(.A(n653), .Y(new_n874));
  xor_5  g0599(.A(n952), .B(new_n874), .Y(new_n875));
  or_2   g0600(.A(new_n875), .B(new_n873), .Y(new_n876));
  and_7  g0601(.A(new_n876), .B(new_n872), .Y(new_n877));
  or_2   g0602(.A(new_n877), .B(new_n871), .Y(new_n878));
  and_7  g0603(.A(new_n878), .B(new_n870_1), .Y(new_n879));
  or_2   g0604(.A(new_n879), .B(new_n867_1), .Y(new_n880));
  and_7  g0605(.A(new_n880), .B(new_n866), .Y(new_n881));
  and_7  g0606(.A(new_n881), .B(new_n863), .Y(new_n882_1));
  not_13 g0607(.A(new_n863), .Y(new_n883_1));
  and_7  g0608(.A(n927), .B(n555), .Y(new_n884));
  not_13 g0609(.A(new_n884), .Y(new_n885));
  and_7  g0610(.A(new_n885), .B(new_n866), .Y(new_n886));
  nor_6  g0611(.A(new_n877), .B(new_n871), .Y(new_n887));
  or_2   g0612(.A(new_n887), .B(new_n869), .Y(new_n888_1));
  and_7  g0613(.A(new_n888_1), .B(new_n886), .Y(new_n889));
  or_2   g0614(.A(new_n889), .B(new_n865_1), .Y(new_n890));
  and_7  g0615(.A(new_n890), .B(new_n883_1), .Y(new_n891_1));
  or_2   g0616(.A(new_n891_1), .B(new_n882_1), .Y(new_n892_1));
  and_7  g0617(.A(new_n892_1), .B(new_n400), .Y(new_n893));
  nor_6  g0618(.A(new_n892_1), .B(new_n400), .Y(new_n894));
  nor_6  g0619(.A(new_n894), .B(new_n893), .Y(new_n895));
  and_7  g0620(.A(new_n879), .B(new_n867_1), .Y(new_n896));
  or_2   g0621(.A(new_n896), .B(new_n889), .Y(new_n897));
  nor_6  g0622(.A(new_n897), .B(new_n405), .Y(new_n898));
  and_7  g0623(.A(new_n897), .B(new_n405), .Y(new_n899));
  nor_6  g0624(.A(new_n899), .B(new_n898), .Y(new_n900));
  not_13 g0625(.A(new_n873), .Y(new_n901));
  and_7  g0626(.A(n952), .B(n653), .Y(new_n902_1));
  not_13 g0627(.A(new_n902_1), .Y(new_n903));
  and_7  g0628(.A(new_n903), .B(new_n872), .Y(new_n904));
  or_2   g0629(.A(new_n904), .B(new_n901), .Y(new_n905_1));
  xor_5  g0630(.A(n1764), .B(new_n420), .Y(new_n906_1));
  or_2   g0631(.A(new_n906_1), .B(new_n422), .Y(new_n907));
  and_7  g0632(.A(new_n907), .B(new_n876), .Y(new_n908));
  and_7  g0633(.A(new_n908), .B(new_n905_1), .Y(new_n909));
  xor_5  g0634(.A(n1764), .B(n1145), .Y(new_n910));
  and_7  g0635(.A(new_n910), .B(new_n414_1), .Y(new_n911));
  and_7  g0636(.A(new_n911), .B(new_n904), .Y(new_n912_1));
  nor_6  g0637(.A(new_n912_1), .B(new_n909), .Y(new_n913));
  and_7  g0638(.A(new_n913), .B(new_n431), .Y(new_n914));
  nor_6  g0639(.A(new_n914), .B(new_n909), .Y(new_n915));
  and_7  g0640(.A(new_n877), .B(new_n871), .Y(new_n916));
  or_2   g0641(.A(new_n916), .B(new_n887), .Y(new_n917));
  and_7  g0642(.A(new_n917), .B(new_n915), .Y(new_n918));
  nor_6  g0643(.A(new_n917), .B(new_n915), .Y(new_n919));
  nor_6  g0644(.A(new_n919), .B(new_n918), .Y(new_n920));
  and_7  g0645(.A(new_n920), .B(new_n441), .Y(new_n921));
  nor_6  g0646(.A(new_n921), .B(new_n918), .Y(new_n922));
  and_7  g0647(.A(new_n922), .B(new_n900), .Y(new_n923));
  nor_6  g0648(.A(new_n923), .B(new_n898), .Y(new_n924));
  xor_5  g0649(.A(new_n924), .B(new_n895), .Y(n74));
  and_7  g0650(.A(new_n570), .B(new_n511), .Y(new_n926));
  or_2   g0651(.A(new_n496), .B(n1642), .Y(new_n927_1));
  xor_5  g0652(.A(new_n927_1), .B(new_n800), .Y(new_n928));
  and_7  g0653(.A(new_n928), .B(n1381), .Y(new_n929));
  and_7  g0654(.A(new_n502), .B(new_n805), .Y(new_n930));
  not_13 g0655(.A(new_n502), .Y(new_n931_1));
  and_7  g0656(.A(new_n931_1), .B(n1263), .Y(new_n932));
  or_2   g0657(.A(new_n932), .B(new_n503), .Y(new_n933));
  or_2   g0658(.A(new_n933), .B(new_n930), .Y(new_n934));
  and_7  g0659(.A(new_n456), .B(n171), .Y(new_n935_1));
  or_2   g0660(.A(new_n935_1), .B(new_n457_1), .Y(new_n936));
  and_7  g0661(.A(new_n936), .B(new_n934), .Y(new_n937));
  or_2   g0662(.A(new_n937), .B(new_n929), .Y(new_n938));
  and_7  g0663(.A(new_n938), .B(new_n926), .Y(new_n939));
  not_13 g0664(.A(n557), .Y(new_n940));
  not_13 g0665(.A(new_n927_1), .Y(new_n941));
  and_7  g0666(.A(new_n941), .B(new_n800), .Y(new_n942_1));
  or_2   g0667(.A(new_n942_1), .B(new_n940), .Y(new_n943));
  and_7  g0668(.A(new_n942_1), .B(new_n940), .Y(new_n944_1));
  not_13 g0669(.A(new_n944_1), .Y(new_n945));
  and_7  g0670(.A(new_n945), .B(n1381), .Y(new_n946));
  and_7  g0671(.A(new_n946), .B(new_n943), .Y(new_n947));
  and_7  g0672(.A(n557), .B(new_n503), .Y(new_n948));
  xor_5  g0673(.A(new_n930), .B(n1422), .Y(new_n949));
  and_7  g0674(.A(new_n949), .B(n402), .Y(new_n950));
  nor_6  g0675(.A(new_n950), .B(new_n948), .Y(new_n951));
  and_7  g0676(.A(new_n951), .B(new_n456), .Y(new_n952_1));
  nor_6  g0677(.A(new_n952_1), .B(new_n947), .Y(new_n953_1));
  and_7  g0678(.A(new_n953_1), .B(new_n939), .Y(new_n954));
  nor_6  g0679(.A(new_n953_1), .B(new_n939), .Y(new_n955));
  nor_6  g0680(.A(new_n955), .B(new_n954), .Y(n156));
  nor_6  g0681(.A(new_n938), .B(new_n926), .Y(new_n957));
  nor_6  g0682(.A(new_n957), .B(new_n939), .Y(n1149));
  and_7  g0683(.A(n1149), .B(new_n600_1), .Y(new_n959));
  nor_6  g0684(.A(new_n959), .B(n156), .Y(new_n960));
  and_7  g0685(.A(new_n959), .B(new_n953_1), .Y(new_n961_1));
  nor_6  g0686(.A(new_n961_1), .B(new_n960), .Y(n106));
  xor_5  g0687(.A(new_n568), .B(new_n559_1), .Y(n1385));
  nor_6  g0688(.A(n1385), .B(new_n596), .Y(new_n964));
  nor_6  g0689(.A(new_n964), .B(new_n597), .Y(n126));
  not_13 g0690(.A(new_n746), .Y(new_n966));
  or_2   g0691(.A(new_n776), .B(new_n748_1), .Y(new_n967));
  and_7  g0692(.A(new_n967), .B(new_n966), .Y(new_n968_1));
  xor_5  g0693(.A(new_n968_1), .B(new_n741), .Y(n135));
  and_7  g0694(.A(new_n652), .B(new_n277_1), .Y(new_n970));
  xor_5  g0695(.A(new_n652), .B(n1643), .Y(new_n971));
  or_2   g0696(.A(new_n671), .B(n555), .Y(new_n972));
  and_7  g0697(.A(new_n647_1), .B(new_n285), .Y(new_n973));
  not_13 g0698(.A(new_n973), .Y(new_n974_1));
  xor_5  g0699(.A(new_n647_1), .B(n353), .Y(new_n975));
  or_2   g0700(.A(new_n681), .B(n952), .Y(new_n976));
  and_7  g0701(.A(new_n685), .B(n1145), .Y(new_n977));
  xor_5  g0702(.A(new_n681), .B(new_n539), .Y(new_n978));
  or_2   g0703(.A(new_n978), .B(new_n977), .Y(new_n979_1));
  and_7  g0704(.A(new_n979_1), .B(new_n976), .Y(new_n980_1));
  or_2   g0705(.A(new_n980_1), .B(new_n975), .Y(new_n981));
  and_7  g0706(.A(new_n981), .B(new_n974_1), .Y(new_n982));
  xor_5  g0707(.A(new_n644), .B(n555), .Y(new_n983));
  or_2   g0708(.A(new_n983), .B(new_n982), .Y(new_n984));
  and_7  g0709(.A(new_n984), .B(new_n972), .Y(new_n985));
  nor_6  g0710(.A(new_n985), .B(new_n971), .Y(new_n986));
  or_2   g0711(.A(new_n986), .B(new_n970), .Y(new_n987));
  or_2   g0712(.A(new_n987), .B(new_n656), .Y(new_n988));
  xor_5  g0713(.A(new_n988), .B(new_n702), .Y(n145));
  xor_5  g0714(.A(new_n413), .B(n347), .Y(n174));
  and_7  g0715(.A(new_n395), .B(n1597), .Y(new_n991_1));
  and_7  g0716(.A(new_n392), .B(new_n391_1), .Y(new_n992));
  or_2   g0717(.A(new_n992), .B(new_n302), .Y(new_n993));
  and_7  g0718(.A(new_n993), .B(new_n374), .Y(new_n994));
  or_2   g0719(.A(new_n994), .B(new_n991_1), .Y(new_n995));
  and_7  g0720(.A(new_n402_1), .B(n682), .Y(new_n996));
  nor_6  g0721(.A(new_n401_1), .B(new_n300), .Y(new_n997));
  or_2   g0722(.A(new_n997), .B(new_n334), .Y(new_n998));
  or_2   g0723(.A(new_n402_1), .B(n682), .Y(new_n999));
  and_7  g0724(.A(new_n999), .B(new_n998), .Y(new_n1000_1));
  and_7  g0725(.A(new_n407), .B(n1435), .Y(new_n1001));
  nor_6  g0726(.A(new_n406), .B(new_n298), .Y(new_n1002));
  and_7  g0727(.A(new_n1002), .B(new_n316), .Y(new_n1003));
  or_2   g0728(.A(new_n1003), .B(new_n1001), .Y(new_n1004));
  and_7  g0729(.A(new_n412), .B(n66), .Y(new_n1005_1));
  nor_6  g0730(.A(new_n412), .B(n66), .Y(new_n1006));
  nor_6  g0731(.A(new_n1006), .B(new_n1005_1), .Y(new_n1007));
  or_2   g0732(.A(new_n418), .B(n968), .Y(new_n1008));
  and_7  g0733(.A(new_n413), .B(n347), .Y(new_n1009));
  nor_6  g0734(.A(new_n418), .B(n968), .Y(new_n1010));
  and_7  g0735(.A(new_n418), .B(n968), .Y(new_n1011));
  or_2   g0736(.A(new_n1011), .B(new_n1010), .Y(new_n1012_1));
  or_2   g0737(.A(new_n1012_1), .B(new_n1009), .Y(new_n1013));
  and_7  g0738(.A(new_n1013), .B(new_n1008), .Y(new_n1014));
  and_7  g0739(.A(new_n1014), .B(new_n1007), .Y(new_n1015_1));
  nor_6  g0740(.A(new_n1015_1), .B(new_n1005_1), .Y(new_n1016_1));
  nor_6  g0741(.A(new_n1016_1), .B(new_n1004), .Y(new_n1017));
  or_2   g0742(.A(new_n1017), .B(new_n1001), .Y(new_n1018));
  and_7  g0743(.A(new_n1018), .B(new_n1000_1), .Y(new_n1019));
  nor_6  g0744(.A(new_n1019), .B(new_n996), .Y(new_n1020));
  nor_6  g0745(.A(new_n1020), .B(new_n995), .Y(new_n1021));
  and_7  g0746(.A(new_n1020), .B(new_n995), .Y(new_n1022));
  nor_6  g0747(.A(new_n1022), .B(new_n1021), .Y(new_n1023));
  nor_6  g0748(.A(new_n1018), .B(new_n1000_1), .Y(new_n1024));
  nor_6  g0749(.A(new_n1024), .B(new_n1019), .Y(new_n1025_1));
  nor_6  g0750(.A(new_n1014), .B(new_n1007), .Y(new_n1026));
  nor_6  g0751(.A(new_n1026), .B(new_n1015_1), .Y(n1426));
  and_7  g0752(.A(new_n1016_1), .B(new_n1004), .Y(new_n1028));
  nor_6  g0753(.A(new_n1028), .B(new_n1017), .Y(new_n1029));
  or_2   g0754(.A(new_n1029), .B(n1426), .Y(new_n1030_1));
  nor_6  g0755(.A(new_n1030_1), .B(new_n1025_1), .Y(new_n1031));
  xor_5  g0756(.A(new_n1031), .B(new_n1023), .Y(n181));
  xor_5  g0757(.A(new_n433_1), .B(new_n412), .Y(new_n1033));
  xor_5  g0758(.A(new_n1033), .B(new_n441), .Y(n208));
  not_13 g0759(.A(n213), .Y(new_n1035));
  and_7  g0760(.A(new_n647_1), .B(new_n1035), .Y(new_n1036));
  xor_5  g0761(.A(new_n647_1), .B(n213), .Y(new_n1037));
  not_13 g0762(.A(n1743), .Y(new_n1038));
  and_7  g0763(.A(new_n689), .B(new_n1038), .Y(new_n1039));
  not_13 g0764(.A(n600), .Y(new_n1040));
  not_13 g0765(.A(new_n683_1), .Y(new_n1041));
  or_2   g0766(.A(new_n469_1), .B(n266), .Y(new_n1042));
  and_7  g0767(.A(new_n1042), .B(new_n1041), .Y(new_n1043));
  or_2   g0768(.A(new_n1043), .B(new_n1040), .Y(new_n1044));
  xor_5  g0769(.A(new_n681), .B(n1743), .Y(new_n1045));
  and_7  g0770(.A(new_n1045), .B(new_n1044), .Y(new_n1046));
  nor_6  g0771(.A(new_n1046), .B(new_n1039), .Y(new_n1047));
  nor_6  g0772(.A(new_n1047), .B(new_n1037), .Y(new_n1048));
  or_2   g0773(.A(new_n1048), .B(new_n1036), .Y(new_n1049));
  or_2   g0774(.A(new_n1049), .B(new_n644), .Y(new_n1050));
  or_2   g0775(.A(new_n1050), .B(new_n652), .Y(new_n1051));
  or_2   g0776(.A(new_n1051), .B(new_n656), .Y(new_n1052));
  nor_6  g0777(.A(new_n1048), .B(new_n1036), .Y(new_n1053));
  and_7  g0778(.A(new_n1053), .B(new_n671), .Y(new_n1054));
  and_7  g0779(.A(new_n1054), .B(new_n669), .Y(new_n1055));
  or_2   g0780(.A(new_n1055), .B(new_n666), .Y(new_n1056));
  and_7  g0781(.A(new_n1056), .B(new_n1052), .Y(new_n1057));
  not_13 g0782(.A(n17), .Y(new_n1058));
  not_13 g0783(.A(n424), .Y(new_n1059));
  and_7  g0784(.A(new_n277_1), .B(new_n1059), .Y(new_n1060));
  not_13 g0785(.A(new_n1060), .Y(new_n1061));
  and_7  g0786(.A(n1643), .B(n424), .Y(new_n1062_1));
  not_13 g0787(.A(new_n1062_1), .Y(new_n1063));
  and_7  g0788(.A(new_n1063), .B(new_n1061), .Y(new_n1064));
  not_13 g0789(.A(n1363), .Y(new_n1065));
  and_7  g0790(.A(new_n1065), .B(new_n545), .Y(new_n1066));
  xor_5  g0791(.A(n1363), .B(n555), .Y(new_n1067_1));
  not_13 g0792(.A(n498), .Y(new_n1068_1));
  and_7  g0793(.A(new_n1068_1), .B(new_n285), .Y(new_n1069));
  xor_5  g0794(.A(n498), .B(new_n285), .Y(new_n1070));
  not_13 g0795(.A(n414), .Y(new_n1071));
  and_7  g0796(.A(new_n539), .B(new_n1071), .Y(new_n1072));
  and_7  g0797(.A(n1145), .B(n183), .Y(new_n1073));
  not_13 g0798(.A(new_n1073), .Y(new_n1074));
  xor_5  g0799(.A(n952), .B(n414), .Y(new_n1075));
  and_7  g0800(.A(new_n1075), .B(new_n1074), .Y(new_n1076));
  nor_6  g0801(.A(new_n1076), .B(new_n1072), .Y(new_n1077));
  nor_6  g0802(.A(new_n1077), .B(new_n1070), .Y(new_n1078));
  or_2   g0803(.A(new_n1078), .B(new_n1069), .Y(new_n1079));
  and_7  g0804(.A(new_n1079), .B(new_n1067_1), .Y(new_n1080));
  or_2   g0805(.A(new_n1080), .B(new_n1066), .Y(new_n1081));
  and_7  g0806(.A(new_n1081), .B(new_n1064), .Y(new_n1082));
  or_2   g0807(.A(new_n1082), .B(new_n1060), .Y(new_n1083));
  or_2   g0808(.A(new_n1083), .B(new_n1058), .Y(new_n1084));
  xor_5  g0809(.A(n1643), .B(new_n1059), .Y(new_n1085));
  nor_6  g0810(.A(new_n1080), .B(new_n1066), .Y(new_n1086));
  or_2   g0811(.A(new_n1086), .B(new_n1085), .Y(new_n1087));
  and_7  g0812(.A(new_n1087), .B(new_n1061), .Y(new_n1088));
  or_2   g0813(.A(new_n1088), .B(n17), .Y(new_n1089));
  and_7  g0814(.A(new_n1089), .B(new_n1084), .Y(new_n1090));
  and_7  g0815(.A(new_n1090), .B(new_n1057), .Y(new_n1091));
  nor_6  g0816(.A(new_n1090), .B(new_n1057), .Y(new_n1092));
  or_2   g0817(.A(new_n1092), .B(new_n1091), .Y(new_n1093));
  and_7  g0818(.A(new_n1050), .B(new_n652), .Y(new_n1094));
  nor_6  g0819(.A(new_n1094), .B(new_n1055), .Y(new_n1095));
  and_7  g0820(.A(new_n1086), .B(new_n1085), .Y(new_n1096));
  or_2   g0821(.A(new_n1096), .B(new_n1082), .Y(new_n1097));
  or_2   g0822(.A(new_n1097), .B(new_n1095), .Y(new_n1098));
  and_7  g0823(.A(new_n1049), .B(new_n644), .Y(new_n1099));
  nor_6  g0824(.A(new_n1099), .B(new_n1054), .Y(new_n1100));
  nor_6  g0825(.A(new_n1079), .B(new_n1067_1), .Y(new_n1101));
  or_2   g0826(.A(new_n1101), .B(new_n1080), .Y(new_n1102));
  nor_6  g0827(.A(new_n1102), .B(new_n1100), .Y(new_n1103_1));
  and_7  g0828(.A(new_n1102), .B(new_n1100), .Y(new_n1104));
  or_2   g0829(.A(new_n1104), .B(new_n1103_1), .Y(new_n1105));
  and_7  g0830(.A(new_n1047), .B(new_n1037), .Y(new_n1106));
  nor_6  g0831(.A(new_n1106), .B(new_n1048), .Y(new_n1107));
  and_7  g0832(.A(new_n1077), .B(new_n1070), .Y(new_n1108));
  nor_6  g0833(.A(new_n1108), .B(new_n1078), .Y(new_n1109));
  and_7  g0834(.A(new_n1109), .B(new_n1107), .Y(new_n1110));
  or_2   g0835(.A(new_n1075), .B(new_n1074), .Y(new_n1111));
  xor_5  g0836(.A(n1145), .B(n183), .Y(new_n1112));
  xor_5  g0837(.A(new_n685), .B(n600), .Y(new_n1113_1));
  and_7  g0838(.A(new_n1113_1), .B(new_n1112), .Y(new_n1114));
  nor_6  g0839(.A(new_n1114), .B(new_n1076), .Y(new_n1115));
  and_7  g0840(.A(new_n1115), .B(new_n1111), .Y(new_n1116));
  not_13 g0841(.A(new_n1044), .Y(new_n1117));
  xor_5  g0842(.A(new_n681), .B(new_n1038), .Y(new_n1118));
  or_2   g0843(.A(new_n1118), .B(new_n1117), .Y(new_n1119_1));
  or_2   g0844(.A(new_n1045), .B(new_n1044), .Y(new_n1120));
  and_7  g0845(.A(new_n1120), .B(new_n1119_1), .Y(new_n1121));
  and_7  g0846(.A(new_n1114), .B(new_n1075), .Y(new_n1122));
  nor_6  g0847(.A(new_n1122), .B(new_n1116), .Y(new_n1123));
  and_7  g0848(.A(new_n1123), .B(new_n1121), .Y(new_n1124));
  or_2   g0849(.A(new_n1124), .B(new_n1116), .Y(new_n1125));
  nor_6  g0850(.A(new_n1109), .B(new_n1107), .Y(new_n1126));
  nor_6  g0851(.A(new_n1126), .B(new_n1110), .Y(new_n1127));
  and_7  g0852(.A(new_n1127), .B(new_n1125), .Y(new_n1128));
  nor_6  g0853(.A(new_n1128), .B(new_n1110), .Y(new_n1129));
  nor_6  g0854(.A(new_n1129), .B(new_n1105), .Y(new_n1130));
  nor_6  g0855(.A(new_n1130), .B(new_n1103_1), .Y(new_n1131));
  nor_6  g0856(.A(new_n1097), .B(new_n1095), .Y(new_n1132));
  and_7  g0857(.A(new_n1097), .B(new_n1095), .Y(new_n1133));
  or_2   g0858(.A(new_n1133), .B(new_n1132), .Y(new_n1134));
  or_2   g0859(.A(new_n1134), .B(new_n1131), .Y(new_n1135_1));
  and_7  g0860(.A(new_n1135_1), .B(new_n1098), .Y(new_n1136));
  nor_6  g0861(.A(new_n1136), .B(new_n1093), .Y(new_n1137));
  and_7  g0862(.A(new_n1136), .B(new_n1093), .Y(new_n1138_1));
  or_2   g0863(.A(new_n1138_1), .B(new_n1137), .Y(n216));
  not_13 g0864(.A(new_n1125), .Y(new_n1140_1));
  xor_5  g0865(.A(new_n1127), .B(new_n1140_1), .Y(n218));
  and_7  g0866(.A(new_n852), .B(new_n836_1), .Y(new_n1142_1));
  or_2   g0867(.A(new_n1142_1), .B(new_n853), .Y(n231));
  not_13 g0868(.A(n1747), .Y(new_n1144));
  not_13 g0869(.A(n738), .Y(new_n1145_1));
  not_13 g0870(.A(n961), .Y(new_n1146));
  or_2   g0871(.A(new_n1084), .B(new_n1146), .Y(new_n1147));
  or_2   g0872(.A(new_n1147), .B(new_n1145_1), .Y(new_n1148));
  or_2   g0873(.A(new_n1148), .B(new_n1144), .Y(new_n1149_1));
  and_7  g0874(.A(new_n1088), .B(n17), .Y(new_n1150));
  and_7  g0875(.A(new_n1150), .B(n961), .Y(new_n1151));
  and_7  g0876(.A(new_n1151), .B(n738), .Y(new_n1152));
  or_2   g0877(.A(new_n1152), .B(n1747), .Y(new_n1153));
  and_7  g0878(.A(new_n1153), .B(new_n1149_1), .Y(new_n1154));
  or_2   g0879(.A(new_n1052), .B(new_n702), .Y(new_n1155));
  or_2   g0880(.A(new_n1155), .B(new_n788_1), .Y(new_n1156));
  or_2   g0881(.A(new_n1156), .B(new_n798), .Y(new_n1157));
  and_7  g0882(.A(new_n1055), .B(new_n666), .Y(new_n1158));
  and_7  g0883(.A(new_n1158), .B(new_n662), .Y(new_n1159));
  and_7  g0884(.A(new_n1159), .B(new_n710), .Y(new_n1160));
  or_2   g0885(.A(new_n1160), .B(new_n794), .Y(new_n1161_1));
  and_7  g0886(.A(new_n1161_1), .B(new_n1157), .Y(new_n1162_1));
  and_7  g0887(.A(new_n1162_1), .B(new_n1154), .Y(new_n1163));
  nor_6  g0888(.A(new_n1162_1), .B(new_n1154), .Y(new_n1164));
  or_2   g0889(.A(new_n1164), .B(new_n1163), .Y(new_n1165));
  or_2   g0890(.A(new_n1151), .B(n738), .Y(new_n1166));
  and_7  g0891(.A(new_n1166), .B(new_n1148), .Y(new_n1167));
  or_2   g0892(.A(new_n1159), .B(new_n710), .Y(new_n1168));
  and_7  g0893(.A(new_n1168), .B(new_n1156), .Y(new_n1169));
  or_2   g0894(.A(new_n1169), .B(new_n1167), .Y(new_n1170));
  nor_6  g0895(.A(new_n1169), .B(new_n1167), .Y(new_n1171));
  and_7  g0896(.A(new_n1169), .B(new_n1167), .Y(new_n1172_1));
  or_2   g0897(.A(new_n1172_1), .B(new_n1171), .Y(new_n1173));
  or_2   g0898(.A(new_n1150), .B(n961), .Y(new_n1174));
  and_7  g0899(.A(new_n1174), .B(new_n1147), .Y(new_n1175_1));
  or_2   g0900(.A(new_n1158), .B(new_n662), .Y(new_n1176));
  and_7  g0901(.A(new_n1176), .B(new_n1155), .Y(new_n1177));
  nor_6  g0902(.A(new_n1177), .B(new_n1175_1), .Y(new_n1178));
  and_7  g0903(.A(new_n1177), .B(new_n1175_1), .Y(new_n1179));
  nor_6  g0904(.A(new_n1179), .B(new_n1178), .Y(new_n1180));
  or_2   g0905(.A(new_n1137), .B(new_n1092), .Y(new_n1181));
  and_7  g0906(.A(new_n1181), .B(new_n1180), .Y(new_n1182));
  nor_6  g0907(.A(new_n1182), .B(new_n1178), .Y(new_n1183_1));
  or_2   g0908(.A(new_n1183_1), .B(new_n1173), .Y(new_n1184));
  and_7  g0909(.A(new_n1184), .B(new_n1170), .Y(new_n1185));
  nor_6  g0910(.A(new_n1185), .B(new_n1165), .Y(new_n1186));
  and_7  g0911(.A(new_n1185), .B(new_n1165), .Y(new_n1187));
  or_2   g0912(.A(new_n1187), .B(new_n1186), .Y(n238));
  and_7  g0913(.A(new_n303_1), .B(n1537), .Y(new_n1189));
  and_7  g0914(.A(new_n1189), .B(n675), .Y(new_n1190));
  xor_5  g0915(.A(new_n1190), .B(n1263), .Y(new_n1191_1));
  not_13 g0916(.A(n675), .Y(new_n1192));
  not_13 g0917(.A(n1537), .Y(new_n1193));
  not_13 g0918(.A(n433), .Y(new_n1194_1));
  or_2   g0919(.A(new_n393), .B(new_n1194_1), .Y(new_n1195));
  or_2   g0920(.A(new_n1195), .B(new_n1193), .Y(new_n1196));
  or_2   g0921(.A(new_n1196), .B(new_n1192), .Y(new_n1197));
  or_2   g0922(.A(new_n1189), .B(n675), .Y(new_n1198));
  and_7  g0923(.A(new_n1198), .B(new_n1197), .Y(new_n1199_1));
  and_7  g0924(.A(new_n1199_1), .B(n379), .Y(new_n1200));
  nor_6  g0925(.A(new_n1199_1), .B(n379), .Y(new_n1201_1));
  or_2   g0926(.A(new_n1201_1), .B(new_n1200), .Y(new_n1202_1));
  and_7  g0927(.A(new_n1195), .B(new_n1193), .Y(new_n1203));
  nor_6  g0928(.A(new_n1203), .B(new_n1189), .Y(new_n1204));
  and_7  g0929(.A(new_n1204), .B(n1527), .Y(new_n1205));
  nor_6  g0930(.A(new_n1204), .B(n1527), .Y(new_n1206));
  or_2   g0931(.A(new_n1206), .B(new_n1205), .Y(new_n1207));
  or_2   g0932(.A(new_n304), .B(new_n303_1), .Y(new_n1208));
  or_2   g0933(.A(new_n1208), .B(new_n373), .Y(new_n1209));
  nor_6  g0934(.A(new_n1021), .B(new_n991_1), .Y(new_n1210));
  and_7  g0935(.A(new_n305), .B(n46), .Y(new_n1211));
  and_7  g0936(.A(new_n1208), .B(new_n373), .Y(new_n1212));
  or_2   g0937(.A(new_n1212), .B(new_n1211), .Y(new_n1213));
  or_2   g0938(.A(new_n1213), .B(new_n1210), .Y(new_n1214));
  and_7  g0939(.A(new_n1214), .B(new_n1209), .Y(new_n1215));
  nor_6  g0940(.A(new_n1215), .B(new_n1207), .Y(new_n1216));
  nor_6  g0941(.A(new_n1216), .B(new_n1205), .Y(new_n1217));
  nor_6  g0942(.A(new_n1217), .B(new_n1202_1), .Y(new_n1218));
  nor_6  g0943(.A(new_n1218), .B(new_n1200), .Y(new_n1219));
  and_7  g0944(.A(new_n1219), .B(new_n1191_1), .Y(new_n1220));
  nor_6  g0945(.A(new_n1219), .B(new_n1191_1), .Y(new_n1221));
  or_2   g0946(.A(new_n1221), .B(new_n1220), .Y(new_n1222_1));
  and_7  g0947(.A(new_n1217), .B(new_n1202_1), .Y(new_n1223));
  nor_6  g0948(.A(new_n1223), .B(new_n1218), .Y(new_n1224));
  and_7  g0949(.A(new_n1215), .B(new_n1207), .Y(new_n1225));
  nor_6  g0950(.A(new_n1225), .B(new_n1216), .Y(new_n1226));
  or_2   g0951(.A(new_n1030_1), .B(new_n1025_1), .Y(new_n1227));
  or_2   g0952(.A(new_n1227), .B(new_n1023), .Y(new_n1228));
  or_2   g0953(.A(new_n1021), .B(new_n991_1), .Y(new_n1229));
  xor_5  g0954(.A(new_n305), .B(n46), .Y(new_n1230));
  and_7  g0955(.A(new_n1230), .B(new_n1229), .Y(new_n1231));
  and_7  g0956(.A(new_n1213), .B(new_n1210), .Y(new_n1232));
  nor_6  g0957(.A(new_n1232), .B(new_n1231), .Y(new_n1233));
  or_2   g0958(.A(new_n1233), .B(new_n1228), .Y(new_n1234_1));
  or_2   g0959(.A(new_n1234_1), .B(new_n1226), .Y(new_n1235_1));
  or_2   g0960(.A(new_n1235_1), .B(new_n1224), .Y(new_n1236));
  and_7  g0961(.A(new_n1236), .B(new_n1222_1), .Y(new_n1237_1));
  nor_6  g0962(.A(new_n1221), .B(new_n1220), .Y(new_n1238));
  nor_6  g0963(.A(new_n1235_1), .B(new_n1224), .Y(new_n1239));
  and_7  g0964(.A(new_n1239), .B(new_n1238), .Y(new_n1240));
  or_2   g0965(.A(new_n1240), .B(new_n1237_1), .Y(n270));
  xor_5  g0966(.A(new_n736), .B(new_n402_1), .Y(new_n1242));
  and_7  g0967(.A(new_n743), .B(new_n407), .Y(new_n1243));
  nor_6  g0968(.A(new_n743), .B(new_n407), .Y(new_n1244));
  and_7  g0969(.A(new_n750), .B(new_n412), .Y(new_n1245));
  or_2   g0970(.A(new_n750), .B(new_n412), .Y(new_n1246));
  and_7  g0971(.A(new_n761_1), .B(new_n413), .Y(new_n1247));
  nor_6  g0972(.A(new_n1247), .B(new_n418), .Y(new_n1248));
  and_7  g0973(.A(new_n1247), .B(new_n417), .Y(new_n1249_1));
  nor_6  g0974(.A(new_n1249_1), .B(new_n1248), .Y(new_n1250));
  and_7  g0975(.A(new_n1250), .B(new_n768), .Y(new_n1251));
  nor_6  g0976(.A(new_n1251), .B(new_n1248), .Y(new_n1252));
  and_7  g0977(.A(new_n1252), .B(new_n1246), .Y(new_n1253));
  nor_6  g0978(.A(new_n1253), .B(new_n1245), .Y(new_n1254));
  nor_6  g0979(.A(new_n1254), .B(new_n1244), .Y(new_n1255_1));
  or_2   g0980(.A(new_n1255_1), .B(new_n1243), .Y(new_n1256));
  xor_5  g0981(.A(new_n1256), .B(new_n1242), .Y(n276));
  xor_5  g0982(.A(new_n910), .B(new_n414_1), .Y(n290));
  not_13 g0983(.A(new_n1009), .Y(new_n1259));
  xor_5  g0984(.A(new_n1012_1), .B(new_n1259), .Y(n292));
  and_7  g0985(.A(new_n1152), .B(n1747), .Y(new_n1261));
  or_2   g0986(.A(new_n1157), .B(new_n818), .Y(new_n1262));
  and_7  g0987(.A(new_n1160), .B(new_n794), .Y(new_n1263_1));
  or_2   g0988(.A(new_n1263_1), .B(new_n811), .Y(new_n1264));
  and_7  g0989(.A(new_n1264), .B(new_n1262), .Y(new_n1265));
  nor_6  g0990(.A(new_n1265), .B(new_n1261), .Y(new_n1266));
  and_7  g0991(.A(new_n1265), .B(new_n1261), .Y(new_n1267));
  nor_6  g0992(.A(new_n1267), .B(new_n1266), .Y(new_n1268));
  or_2   g0993(.A(new_n1186), .B(new_n1164), .Y(new_n1269));
  and_7  g0994(.A(new_n1269), .B(new_n1268), .Y(new_n1270));
  or_2   g0995(.A(new_n1270), .B(new_n1266), .Y(new_n1271));
  and_7  g0996(.A(new_n1262), .B(new_n823_1), .Y(new_n1272));
  and_7  g0997(.A(new_n1272), .B(new_n1271), .Y(n299));
  not_13 g0998(.A(n1341), .Y(new_n1274));
  or_2   g0999(.A(new_n532_1), .B(new_n1274), .Y(new_n1275));
  xor_5  g1000(.A(new_n532_1), .B(n1341), .Y(new_n1276));
  and_7  g1001(.A(new_n461), .B(n69), .Y(new_n1277_1));
  nor_6  g1002(.A(new_n476_1), .B(new_n1277_1), .Y(new_n1278_1));
  or_2   g1003(.A(new_n1278_1), .B(new_n1276), .Y(new_n1279));
  and_7  g1004(.A(new_n1279), .B(new_n1275), .Y(new_n1280));
  nor_6  g1005(.A(new_n1280), .B(new_n527), .Y(new_n1281));
  and_7  g1006(.A(new_n1281), .B(new_n558), .Y(new_n1282));
  and_7  g1007(.A(new_n1282), .B(new_n568), .Y(new_n1283_1));
  or_2   g1008(.A(new_n1280), .B(new_n527), .Y(new_n1284));
  or_2   g1009(.A(new_n1284), .B(new_n557_1), .Y(new_n1285));
  and_7  g1010(.A(new_n1285), .B(new_n567), .Y(new_n1286));
  nor_6  g1011(.A(new_n1286), .B(new_n1283_1), .Y(new_n1287));
  not_13 g1012(.A(n761), .Y(new_n1288));
  and_7  g1013(.A(new_n277_1), .B(new_n1288), .Y(new_n1289));
  not_13 g1014(.A(new_n1289), .Y(new_n1290));
  xor_5  g1015(.A(n1643), .B(new_n1288), .Y(new_n1291));
  not_13 g1016(.A(n1172), .Y(new_n1292));
  and_7  g1017(.A(new_n1292), .B(new_n545), .Y(new_n1293));
  xor_5  g1018(.A(n1172), .B(n555), .Y(new_n1294));
  not_13 g1019(.A(n695), .Y(new_n1295));
  and_7  g1020(.A(new_n1295), .B(new_n285), .Y(new_n1296_1));
  xor_5  g1021(.A(n695), .B(new_n285), .Y(new_n1297));
  not_13 g1022(.A(n1296), .Y(new_n1298));
  and_7  g1023(.A(new_n1298), .B(new_n539), .Y(new_n1299));
  and_7  g1024(.A(n1145), .B(n1062), .Y(new_n1300));
  not_13 g1025(.A(new_n1300), .Y(new_n1301));
  xor_5  g1026(.A(n1296), .B(n952), .Y(new_n1302));
  and_7  g1027(.A(new_n1302), .B(new_n1301), .Y(new_n1303));
  nor_6  g1028(.A(new_n1303), .B(new_n1299), .Y(new_n1304));
  nor_6  g1029(.A(new_n1304), .B(new_n1297), .Y(new_n1305_1));
  or_2   g1030(.A(new_n1305_1), .B(new_n1296_1), .Y(new_n1306));
  and_7  g1031(.A(new_n1306), .B(new_n1294), .Y(new_n1307));
  nor_6  g1032(.A(new_n1307), .B(new_n1293), .Y(new_n1308));
  or_2   g1033(.A(new_n1308), .B(new_n1291), .Y(new_n1309));
  and_7  g1034(.A(new_n1309), .B(new_n1290), .Y(new_n1310));
  and_7  g1035(.A(new_n1310), .B(n862), .Y(new_n1311));
  and_7  g1036(.A(new_n1311), .B(n1222), .Y(new_n1312));
  not_13 g1037(.A(n1222), .Y(new_n1313));
  not_13 g1038(.A(n862), .Y(new_n1314));
  and_7  g1039(.A(n1643), .B(n761), .Y(new_n1315_1));
  not_13 g1040(.A(new_n1315_1), .Y(new_n1316));
  and_7  g1041(.A(new_n1316), .B(new_n1290), .Y(new_n1317));
  or_2   g1042(.A(new_n1307), .B(new_n1293), .Y(new_n1318));
  and_7  g1043(.A(new_n1318), .B(new_n1317), .Y(new_n1319));
  or_2   g1044(.A(new_n1319), .B(new_n1289), .Y(new_n1320));
  or_2   g1045(.A(new_n1320), .B(new_n1314), .Y(new_n1321_1));
  and_7  g1046(.A(new_n1321_1), .B(new_n1313), .Y(new_n1322));
  nor_6  g1047(.A(new_n1322), .B(new_n1312), .Y(new_n1323));
  and_7  g1048(.A(new_n1323), .B(new_n1287), .Y(new_n1324));
  nor_6  g1049(.A(new_n1323), .B(new_n1287), .Y(new_n1325));
  or_2   g1050(.A(new_n1325), .B(new_n1324), .Y(new_n1326));
  and_7  g1051(.A(new_n1284), .B(new_n557_1), .Y(new_n1327));
  or_2   g1052(.A(new_n1327), .B(new_n1282), .Y(new_n1328));
  and_7  g1053(.A(new_n1320), .B(new_n1314), .Y(new_n1329));
  or_2   g1054(.A(new_n1329), .B(new_n1311), .Y(new_n1330_1));
  and_7  g1055(.A(new_n1330_1), .B(new_n1328), .Y(new_n1331));
  or_2   g1056(.A(new_n1281), .B(new_n558), .Y(new_n1332_1));
  and_7  g1057(.A(new_n1332_1), .B(new_n1285), .Y(new_n1333));
  or_2   g1058(.A(new_n1310), .B(n862), .Y(new_n1334));
  and_7  g1059(.A(new_n1334), .B(new_n1321_1), .Y(new_n1335));
  and_7  g1060(.A(new_n1335), .B(new_n1333), .Y(new_n1336));
  nor_6  g1061(.A(new_n1336), .B(new_n1331), .Y(new_n1337));
  and_7  g1062(.A(new_n1280), .B(new_n527), .Y(new_n1338_1));
  nor_6  g1063(.A(new_n1338_1), .B(new_n1281), .Y(new_n1339));
  and_7  g1064(.A(new_n1308), .B(new_n1291), .Y(new_n1340_1));
  or_2   g1065(.A(new_n1340_1), .B(new_n1319), .Y(new_n1341_1));
  nor_6  g1066(.A(new_n1341_1), .B(new_n1339), .Y(new_n1342));
  and_7  g1067(.A(new_n1341_1), .B(new_n1339), .Y(new_n1343));
  or_2   g1068(.A(new_n1343), .B(new_n1342), .Y(new_n1344));
  xor_5  g1069(.A(new_n532_1), .B(new_n1274), .Y(new_n1345));
  or_2   g1070(.A(new_n476_1), .B(new_n1277_1), .Y(new_n1346));
  or_2   g1071(.A(new_n1346), .B(new_n1345), .Y(new_n1347_1));
  and_7  g1072(.A(new_n1347_1), .B(new_n1279), .Y(new_n1348_1));
  nor_6  g1073(.A(new_n1306), .B(new_n1294), .Y(new_n1349_1));
  or_2   g1074(.A(new_n1349_1), .B(new_n1307), .Y(new_n1350));
  nor_6  g1075(.A(new_n1350), .B(new_n1348_1), .Y(new_n1351_1));
  and_7  g1076(.A(new_n1350), .B(new_n1348_1), .Y(new_n1352));
  nor_6  g1077(.A(new_n1352), .B(new_n1351_1), .Y(new_n1353));
  and_7  g1078(.A(new_n1304), .B(new_n1297), .Y(new_n1354));
  or_2   g1079(.A(new_n1354), .B(new_n1305_1), .Y(new_n1355));
  nor_6  g1080(.A(new_n1355), .B(new_n478), .Y(new_n1356));
  and_7  g1081(.A(new_n1355), .B(new_n478), .Y(new_n1357));
  or_2   g1082(.A(new_n1357), .B(new_n1356), .Y(new_n1358));
  or_2   g1083(.A(new_n1302), .B(new_n1301), .Y(new_n1359));
  xor_5  g1084(.A(n1145), .B(n1062), .Y(new_n1360));
  and_7  g1085(.A(new_n1360), .B(new_n482_1), .Y(new_n1361));
  nor_6  g1086(.A(new_n1361), .B(new_n1303), .Y(new_n1362));
  and_7  g1087(.A(new_n1362), .B(new_n1359), .Y(new_n1363_1));
  and_7  g1088(.A(new_n1361), .B(new_n1302), .Y(new_n1364));
  nor_6  g1089(.A(new_n1364), .B(new_n1363_1), .Y(new_n1365));
  and_7  g1090(.A(new_n1365), .B(new_n486), .Y(new_n1366));
  nor_6  g1091(.A(new_n1366), .B(new_n1363_1), .Y(new_n1367));
  nor_6  g1092(.A(new_n1367), .B(new_n1358), .Y(new_n1368));
  or_2   g1093(.A(new_n1368), .B(new_n1356), .Y(new_n1369_1));
  and_7  g1094(.A(new_n1369_1), .B(new_n1353), .Y(new_n1370));
  nor_6  g1095(.A(new_n1370), .B(new_n1351_1), .Y(new_n1371));
  nor_6  g1096(.A(new_n1371), .B(new_n1344), .Y(new_n1372));
  or_2   g1097(.A(new_n1372), .B(new_n1342), .Y(new_n1373));
  and_7  g1098(.A(new_n1373), .B(new_n1337), .Y(new_n1374));
  nor_6  g1099(.A(new_n1374), .B(new_n1331), .Y(new_n1375));
  and_7  g1100(.A(new_n1375), .B(new_n1326), .Y(new_n1376));
  nor_6  g1101(.A(new_n1375), .B(new_n1326), .Y(new_n1377));
  or_2   g1102(.A(new_n1377), .B(new_n1376), .Y(n317));
  xor_5  g1103(.A(new_n1360), .B(new_n482_1), .Y(n372));
  not_13 g1104(.A(new_n922), .Y(new_n1380));
  xor_5  g1105(.A(new_n1380), .B(new_n900), .Y(n378));
  not_13 g1106(.A(new_n826), .Y(new_n1382));
  or_2   g1107(.A(new_n988), .B(new_n702), .Y(new_n1383_1));
  or_2   g1108(.A(new_n1383_1), .B(new_n788_1), .Y(new_n1384));
  or_2   g1109(.A(new_n1384), .B(new_n798), .Y(new_n1385_1));
  or_2   g1110(.A(new_n1385_1), .B(new_n818), .Y(new_n1386));
  or_2   g1111(.A(new_n1386), .B(new_n1382), .Y(new_n1387));
  or_2   g1112(.A(new_n1387), .B(new_n823_1), .Y(new_n1388));
  not_13 g1113(.A(new_n823_1), .Y(new_n1389));
  not_13 g1114(.A(new_n970), .Y(new_n1390));
  or_2   g1115(.A(new_n985), .B(new_n971), .Y(new_n1391));
  and_7  g1116(.A(new_n1391), .B(new_n1390), .Y(new_n1392));
  and_7  g1117(.A(new_n1392), .B(new_n666), .Y(new_n1393_1));
  and_7  g1118(.A(new_n1393_1), .B(new_n662), .Y(new_n1394));
  and_7  g1119(.A(new_n1394), .B(new_n710), .Y(new_n1395));
  and_7  g1120(.A(new_n1395), .B(new_n794), .Y(new_n1396));
  and_7  g1121(.A(new_n1396), .B(new_n811), .Y(new_n1397));
  or_2   g1122(.A(new_n1397), .B(new_n1389), .Y(new_n1398));
  and_7  g1123(.A(new_n1398), .B(new_n1388), .Y(new_n1399_1));
  and_7  g1124(.A(new_n1385_1), .B(new_n818), .Y(new_n1400));
  nor_6  g1125(.A(new_n1400), .B(new_n1397), .Y(n1249));
  and_7  g1126(.A(new_n1383_1), .B(new_n788_1), .Y(new_n1402));
  nor_6  g1127(.A(new_n1402), .B(new_n1395), .Y(n1119));
  not_13 g1128(.A(new_n977), .Y(new_n1404));
  or_2   g1129(.A(new_n685), .B(n1145), .Y(new_n1405));
  and_7  g1130(.A(new_n1405), .B(new_n1404), .Y(n647));
  xor_5  g1131(.A(new_n978), .B(new_n1404), .Y(n646));
  or_2   g1132(.A(n646), .B(n647), .Y(new_n1408));
  nor_6  g1133(.A(new_n980_1), .B(new_n975), .Y(new_n1409));
  and_7  g1134(.A(new_n980_1), .B(new_n975), .Y(new_n1410));
  or_2   g1135(.A(new_n1410), .B(new_n1409), .Y(n1016));
  nor_6  g1136(.A(n1016), .B(new_n1408), .Y(new_n1412));
  or_2   g1137(.A(new_n1409), .B(new_n973), .Y(new_n1413));
  not_13 g1138(.A(new_n983), .Y(new_n1414));
  or_2   g1139(.A(new_n1414), .B(new_n1413), .Y(new_n1415));
  and_7  g1140(.A(new_n1415), .B(new_n984), .Y(new_n1416));
  or_2   g1141(.A(new_n1416), .B(new_n1412), .Y(new_n1417));
  and_7  g1142(.A(new_n985), .B(new_n971), .Y(new_n1418));
  nor_6  g1143(.A(new_n1418), .B(new_n986), .Y(new_n1419));
  nor_6  g1144(.A(new_n1419), .B(new_n1417), .Y(new_n1420));
  and_7  g1145(.A(new_n987), .B(new_n656), .Y(new_n1421));
  nor_6  g1146(.A(new_n1421), .B(new_n1393_1), .Y(n773));
  and_7  g1147(.A(n773), .B(new_n1420), .Y(new_n1423));
  and_7  g1148(.A(new_n1423), .B(new_n662), .Y(new_n1424));
  and_7  g1149(.A(new_n1424), .B(n1119), .Y(new_n1425_1));
  and_7  g1150(.A(new_n1425_1), .B(new_n794), .Y(new_n1426_1));
  and_7  g1151(.A(new_n1426_1), .B(n1249), .Y(new_n1427));
  and_7  g1152(.A(new_n1427), .B(new_n826), .Y(new_n1428));
  nor_6  g1153(.A(new_n1428), .B(new_n1399_1), .Y(new_n1429));
  and_7  g1154(.A(new_n1428), .B(new_n1399_1), .Y(new_n1430));
  or_2   g1155(.A(new_n1430), .B(new_n1429), .Y(n387));
  or_2   g1156(.A(new_n1283_1), .B(new_n523), .Y(new_n1432));
  or_2   g1157(.A(new_n1285), .B(new_n567), .Y(new_n1433));
  or_2   g1158(.A(new_n1433), .B(new_n572), .Y(new_n1434));
  and_7  g1159(.A(new_n1434), .B(new_n1432), .Y(new_n1435_1));
  not_13 g1160(.A(n1757), .Y(new_n1436));
  or_2   g1161(.A(new_n1321_1), .B(new_n1313), .Y(new_n1437));
  or_2   g1162(.A(new_n1437), .B(new_n1436), .Y(new_n1438));
  or_2   g1163(.A(new_n1312), .B(n1757), .Y(new_n1439));
  and_7  g1164(.A(new_n1439), .B(new_n1438), .Y(new_n1440_1));
  and_7  g1165(.A(new_n1440_1), .B(new_n1435_1), .Y(new_n1441));
  nor_6  g1166(.A(new_n1440_1), .B(new_n1435_1), .Y(new_n1442));
  nor_6  g1167(.A(new_n1442), .B(new_n1441), .Y(new_n1443));
  or_2   g1168(.A(new_n1323), .B(new_n1287), .Y(new_n1444));
  or_2   g1169(.A(new_n1375), .B(new_n1326), .Y(new_n1445));
  and_7  g1170(.A(new_n1445), .B(new_n1444), .Y(new_n1446));
  xor_5  g1171(.A(new_n1446), .B(new_n1443), .Y(n401));
  xor_5  g1172(.A(new_n920), .B(new_n441), .Y(n423));
  and_7  g1173(.A(new_n1348_1), .B(new_n407), .Y(new_n1449));
  nor_6  g1174(.A(new_n1348_1), .B(new_n407), .Y(new_n1450));
  nor_6  g1175(.A(new_n1450), .B(new_n1449), .Y(new_n1451));
  not_13 g1176(.A(new_n1451), .Y(new_n1452));
  or_2   g1177(.A(new_n492), .B(new_n480), .Y(new_n1453_1));
  xor_5  g1178(.A(new_n1453_1), .B(new_n1452), .Y(n426));
  or_2   g1179(.A(new_n1397), .B(new_n826), .Y(new_n1455));
  and_7  g1180(.A(new_n1455), .B(new_n1387), .Y(n493));
  nor_6  g1181(.A(n493), .B(new_n1427), .Y(new_n1457_1));
  nor_6  g1182(.A(new_n1457_1), .B(new_n1428), .Y(n429));
  xor_5  g1183(.A(n773), .B(new_n1420), .Y(n432));
  and_7  g1184(.A(new_n1339), .B(new_n402_1), .Y(new_n1460_1));
  nor_6  g1185(.A(new_n1339), .B(new_n402_1), .Y(new_n1461_1));
  or_2   g1186(.A(new_n1461_1), .B(new_n1460_1), .Y(new_n1462));
  and_7  g1187(.A(new_n1453_1), .B(new_n1451), .Y(new_n1463_1));
  nor_6  g1188(.A(new_n1463_1), .B(new_n1450), .Y(new_n1464));
  nor_6  g1189(.A(new_n1464), .B(new_n1462), .Y(new_n1465));
  and_7  g1190(.A(new_n1464), .B(new_n1462), .Y(new_n1466));
  or_2   g1191(.A(new_n1466), .B(new_n1465), .Y(n452));
  nor_6  g1192(.A(new_n1233), .B(new_n1228), .Y(new_n1468));
  and_7  g1193(.A(new_n1233), .B(new_n1228), .Y(new_n1469));
  or_2   g1194(.A(new_n1469), .B(new_n1468), .Y(n457));
  nor_6  g1195(.A(new_n1269), .B(new_n1268), .Y(new_n1471));
  or_2   g1196(.A(new_n1471), .B(new_n1270), .Y(n460));
  xor_5  g1197(.A(new_n761_1), .B(new_n760), .Y(n476));
  not_13 g1198(.A(new_n443), .Y(new_n1474));
  xor_5  g1199(.A(new_n1474), .B(new_n410), .Y(n482));
  and_7  g1200(.A(new_n1283_1), .B(new_n523), .Y(new_n1476));
  and_7  g1201(.A(new_n1476), .B(new_n511), .Y(new_n1477));
  and_7  g1202(.A(new_n1477), .B(new_n938), .Y(new_n1478));
  nor_6  g1203(.A(new_n1477), .B(new_n938), .Y(new_n1479));
  nor_6  g1204(.A(new_n1479), .B(new_n1478), .Y(new_n1480));
  and_7  g1205(.A(new_n1480), .B(new_n1190), .Y(new_n1481_1));
  nor_6  g1206(.A(new_n1480), .B(new_n1190), .Y(new_n1482));
  nor_6  g1207(.A(new_n1482), .B(new_n1481_1), .Y(new_n1483));
  nor_6  g1208(.A(new_n1476), .B(new_n511), .Y(new_n1484));
  nor_6  g1209(.A(new_n1484), .B(new_n1477), .Y(new_n1485));
  nor_6  g1210(.A(new_n1485), .B(new_n1199_1), .Y(new_n1486));
  and_7  g1211(.A(new_n1485), .B(new_n1199_1), .Y(new_n1487));
  or_2   g1212(.A(new_n1487), .B(new_n1486), .Y(new_n1488));
  nor_6  g1213(.A(new_n1435_1), .B(new_n1204), .Y(new_n1489));
  and_7  g1214(.A(new_n1435_1), .B(new_n1204), .Y(new_n1490));
  nor_6  g1215(.A(new_n1490), .B(new_n1489), .Y(new_n1491));
  and_7  g1216(.A(new_n1287), .B(new_n305), .Y(new_n1492));
  and_7  g1217(.A(new_n1328), .B(new_n993), .Y(new_n1493));
  or_2   g1218(.A(new_n1333), .B(new_n395), .Y(new_n1494));
  or_2   g1219(.A(new_n1328), .B(new_n993), .Y(new_n1495_1));
  and_7  g1220(.A(new_n1495_1), .B(new_n1494), .Y(new_n1496));
  or_2   g1221(.A(new_n1465), .B(new_n1461_1), .Y(new_n1497));
  and_7  g1222(.A(new_n1497), .B(new_n1496), .Y(new_n1498_1));
  nor_6  g1223(.A(new_n1498_1), .B(new_n1493), .Y(new_n1499));
  nor_6  g1224(.A(new_n1287), .B(new_n305), .Y(new_n1500));
  nor_6  g1225(.A(new_n1500), .B(new_n1492), .Y(new_n1501_1));
  and_7  g1226(.A(new_n1501_1), .B(new_n1499), .Y(new_n1502_1));
  nor_6  g1227(.A(new_n1502_1), .B(new_n1492), .Y(new_n1503));
  and_7  g1228(.A(new_n1503), .B(new_n1491), .Y(new_n1504));
  nor_6  g1229(.A(new_n1504), .B(new_n1489), .Y(new_n1505));
  nor_6  g1230(.A(new_n1505), .B(new_n1488), .Y(new_n1506));
  or_2   g1231(.A(new_n1506), .B(new_n1486), .Y(new_n1507_1));
  and_7  g1232(.A(new_n1507_1), .B(new_n1483), .Y(new_n1508));
  nor_6  g1233(.A(new_n1507_1), .B(new_n1483), .Y(new_n1509));
  or_2   g1234(.A(new_n1509), .B(new_n1508), .Y(n510));
  and_7  g1235(.A(new_n1199_1), .B(new_n1162_1), .Y(new_n1511));
  nor_6  g1236(.A(new_n1199_1), .B(new_n1162_1), .Y(new_n1512));
  nor_6  g1237(.A(new_n1512), .B(new_n1511), .Y(new_n1513));
  nor_6  g1238(.A(new_n1204), .B(new_n1169), .Y(new_n1514));
  and_7  g1239(.A(new_n1204), .B(new_n1169), .Y(new_n1515));
  or_2   g1240(.A(new_n1515), .B(new_n1514), .Y(new_n1516));
  or_2   g1241(.A(new_n1177), .B(new_n305), .Y(new_n1517));
  nor_6  g1242(.A(new_n1177), .B(new_n305), .Y(new_n1518));
  and_7  g1243(.A(new_n1177), .B(new_n305), .Y(new_n1519));
  or_2   g1244(.A(new_n1519), .B(new_n1518), .Y(new_n1520));
  nor_6  g1245(.A(new_n1057), .B(new_n395), .Y(new_n1521));
  and_7  g1246(.A(new_n1057), .B(new_n395), .Y(new_n1522));
  nor_6  g1247(.A(new_n1522), .B(new_n1521), .Y(new_n1523));
  and_7  g1248(.A(new_n1095), .B(new_n402_1), .Y(new_n1524));
  nor_6  g1249(.A(new_n1100), .B(new_n407), .Y(new_n1525_1));
  and_7  g1250(.A(new_n1100), .B(new_n407), .Y(new_n1526));
  or_2   g1251(.A(new_n1526), .B(new_n1525_1), .Y(new_n1527_1));
  xor_5  g1252(.A(new_n295), .B(new_n288), .Y(new_n1528));
  and_7  g1253(.A(new_n1107), .B(new_n1528), .Y(new_n1529));
  nor_6  g1254(.A(new_n1107), .B(new_n1528), .Y(new_n1530_1));
  nor_6  g1255(.A(new_n1530_1), .B(new_n1529), .Y(new_n1531));
  and_7  g1256(.A(new_n1113_1), .B(new_n413), .Y(new_n1532));
  nor_6  g1257(.A(new_n1532), .B(new_n418), .Y(new_n1533));
  and_7  g1258(.A(new_n1532), .B(new_n417), .Y(new_n1534));
  nor_6  g1259(.A(new_n1534), .B(new_n1533), .Y(new_n1535_1));
  and_7  g1260(.A(new_n1535_1), .B(new_n1121), .Y(new_n1536));
  or_2   g1261(.A(new_n1536), .B(new_n1533), .Y(new_n1537_1));
  and_7  g1262(.A(new_n1537_1), .B(new_n1531), .Y(new_n1538));
  nor_6  g1263(.A(new_n1538), .B(new_n1529), .Y(new_n1539));
  nor_6  g1264(.A(new_n1539), .B(new_n1527_1), .Y(new_n1540));
  nor_6  g1265(.A(new_n1540), .B(new_n1525_1), .Y(new_n1541));
  nor_6  g1266(.A(new_n1095), .B(new_n402_1), .Y(new_n1542));
  nor_6  g1267(.A(new_n1542), .B(new_n1524), .Y(new_n1543));
  and_7  g1268(.A(new_n1543), .B(new_n1541), .Y(new_n1544_1));
  nor_6  g1269(.A(new_n1544_1), .B(new_n1524), .Y(new_n1545));
  and_7  g1270(.A(new_n1545), .B(new_n1523), .Y(new_n1546));
  nor_6  g1271(.A(new_n1546), .B(new_n1521), .Y(new_n1547));
  or_2   g1272(.A(new_n1547), .B(new_n1520), .Y(new_n1548));
  and_7  g1273(.A(new_n1548), .B(new_n1517), .Y(new_n1549));
  nor_6  g1274(.A(new_n1549), .B(new_n1516), .Y(new_n1550));
  or_2   g1275(.A(new_n1550), .B(new_n1514), .Y(new_n1551));
  and_7  g1276(.A(new_n1551), .B(new_n1513), .Y(new_n1552));
  nor_6  g1277(.A(new_n1551), .B(new_n1513), .Y(new_n1553));
  or_2   g1278(.A(new_n1553), .B(new_n1552), .Y(n517));
  and_7  g1279(.A(new_n1199_1), .B(new_n843), .Y(new_n1555));
  nor_6  g1280(.A(new_n1199_1), .B(new_n843), .Y(new_n1556_1));
  or_2   g1281(.A(new_n1556_1), .B(new_n1555), .Y(new_n1557));
  nor_6  g1282(.A(new_n1204), .B(new_n714), .Y(new_n1558));
  and_7  g1283(.A(new_n1204), .B(new_n714), .Y(new_n1559));
  or_2   g1284(.A(new_n1559), .B(new_n1558), .Y(new_n1560));
  nor_6  g1285(.A(new_n721), .B(new_n305), .Y(new_n1561));
  nor_6  g1286(.A(new_n728), .B(new_n395), .Y(new_n1562));
  and_7  g1287(.A(new_n728), .B(new_n395), .Y(new_n1563));
  nor_6  g1288(.A(new_n1563), .B(new_n1562), .Y(new_n1564));
  and_7  g1289(.A(new_n736), .B(new_n402_1), .Y(new_n1565));
  or_2   g1290(.A(new_n736), .B(new_n402_1), .Y(new_n1566));
  and_7  g1291(.A(new_n1256), .B(new_n1566), .Y(new_n1567));
  nor_6  g1292(.A(new_n1567), .B(new_n1565), .Y(new_n1568));
  and_7  g1293(.A(new_n1568), .B(new_n1564), .Y(new_n1569));
  nor_6  g1294(.A(new_n1569), .B(new_n1562), .Y(new_n1570));
  and_7  g1295(.A(new_n721), .B(new_n305), .Y(new_n1571));
  or_2   g1296(.A(new_n1571), .B(new_n1561), .Y(new_n1572));
  nor_6  g1297(.A(new_n1572), .B(new_n1570), .Y(new_n1573));
  nor_6  g1298(.A(new_n1573), .B(new_n1561), .Y(new_n1574));
  nor_6  g1299(.A(new_n1574), .B(new_n1560), .Y(new_n1575));
  or_2   g1300(.A(new_n1575), .B(new_n1558), .Y(new_n1576));
  xor_5  g1301(.A(new_n1576), .B(new_n1557), .Y(n522));
  or_2   g1302(.A(new_n1029), .B(new_n1025_1), .Y(new_n1578));
  or_2   g1303(.A(new_n1578), .B(new_n1023), .Y(new_n1579));
  or_2   g1304(.A(new_n1579), .B(new_n1233), .Y(new_n1580));
  or_2   g1305(.A(new_n1580), .B(new_n1226), .Y(new_n1581));
  nor_6  g1306(.A(new_n1581), .B(new_n1224), .Y(new_n1582));
  and_7  g1307(.A(new_n1581), .B(new_n1224), .Y(new_n1583));
  or_2   g1308(.A(new_n1583), .B(new_n1582), .Y(n532));
  and_7  g1309(.A(new_n822), .B(new_n335), .Y(new_n1585));
  and_7  g1310(.A(new_n368), .B(n247), .Y(new_n1586));
  and_7  g1311(.A(new_n1586), .B(n1642), .Y(new_n1587));
  and_7  g1312(.A(new_n1587), .B(n171), .Y(new_n1588));
  and_7  g1313(.A(new_n1588), .B(n557), .Y(new_n1589));
  and_7  g1314(.A(new_n1589), .B(n1000), .Y(new_n1590));
  not_13 g1315(.A(new_n1590), .Y(new_n1591));
  xor_5  g1316(.A(new_n368), .B(new_n512), .Y(new_n1592));
  and_7  g1317(.A(new_n1592), .B(n1000), .Y(new_n1593));
  or_2   g1318(.A(new_n704), .B(n682), .Y(new_n1594));
  and_7  g1319(.A(new_n705), .B(new_n334), .Y(new_n1595_1));
  or_2   g1320(.A(new_n1595_1), .B(new_n500), .Y(new_n1596));
  and_7  g1321(.A(new_n1596), .B(new_n1594), .Y(new_n1597_1));
  and_7  g1322(.A(new_n1597_1), .B(new_n307), .Y(new_n1598));
  or_2   g1323(.A(new_n1598), .B(new_n1593), .Y(new_n1599));
  and_7  g1324(.A(new_n1599), .B(new_n381), .Y(new_n1600_1));
  xor_5  g1325(.A(new_n1594), .B(n379), .Y(new_n1601_1));
  nor_6  g1326(.A(new_n1601_1), .B(n1000), .Y(new_n1602));
  xor_5  g1327(.A(new_n1586), .B(n1642), .Y(new_n1603));
  and_7  g1328(.A(new_n1603), .B(n1000), .Y(new_n1604));
  nor_6  g1329(.A(new_n1604), .B(new_n1602), .Y(new_n1605));
  and_7  g1330(.A(new_n1605), .B(new_n1600_1), .Y(new_n1606));
  or_2   g1331(.A(new_n1594), .B(n379), .Y(new_n1607));
  and_7  g1332(.A(new_n1607), .B(n1263), .Y(new_n1608));
  and_7  g1333(.A(new_n930), .B(new_n375), .Y(new_n1609));
  or_2   g1334(.A(new_n1609), .B(new_n1608), .Y(new_n1610));
  and_7  g1335(.A(new_n1610), .B(new_n307), .Y(new_n1611));
  or_2   g1336(.A(new_n1587), .B(n171), .Y(new_n1612));
  not_13 g1337(.A(new_n1588), .Y(new_n1613_1));
  and_7  g1338(.A(new_n1613_1), .B(n1000), .Y(new_n1614));
  and_7  g1339(.A(new_n1614), .B(new_n1612), .Y(new_n1615));
  nor_6  g1340(.A(new_n1615), .B(new_n1611), .Y(new_n1616));
  and_7  g1341(.A(new_n1616), .B(new_n1606), .Y(new_n1617));
  not_13 g1342(.A(new_n1585), .Y(new_n1618));
  and_7  g1343(.A(new_n1614), .B(new_n940), .Y(new_n1619));
  or_2   g1344(.A(new_n1609), .B(new_n821), .Y(new_n1620));
  and_7  g1345(.A(new_n1620), .B(new_n307), .Y(new_n1621));
  or_2   g1346(.A(new_n1621), .B(new_n1590), .Y(new_n1622_1));
  or_2   g1347(.A(new_n1622_1), .B(new_n1619), .Y(new_n1623));
  and_7  g1348(.A(new_n1623), .B(new_n1618), .Y(new_n1624));
  and_7  g1349(.A(new_n1624), .B(new_n1617), .Y(new_n1625));
  and_7  g1350(.A(new_n1625), .B(new_n1591), .Y(new_n1626));
  nor_6  g1351(.A(new_n1626), .B(new_n1585), .Y(new_n1627));
  nor_6  g1352(.A(new_n1624), .B(new_n1617), .Y(new_n1628));
  or_2   g1353(.A(new_n1628), .B(new_n1625), .Y(new_n1629_1));
  nor_6  g1354(.A(new_n1605), .B(new_n1600_1), .Y(new_n1630));
  or_2   g1355(.A(new_n1630), .B(new_n1606), .Y(new_n1631));
  nor_6  g1356(.A(new_n1599), .B(new_n381), .Y(new_n1632));
  or_2   g1357(.A(new_n1632), .B(new_n1600_1), .Y(new_n1633_1));
  and_7  g1358(.A(new_n1633_1), .B(new_n383), .Y(new_n1634));
  and_7  g1359(.A(new_n1634), .B(new_n1631), .Y(new_n1635_1));
  nor_6  g1360(.A(new_n1616), .B(new_n1606), .Y(new_n1636));
  or_2   g1361(.A(new_n1636), .B(new_n1617), .Y(new_n1637));
  and_7  g1362(.A(new_n1637), .B(new_n1635_1), .Y(new_n1638));
  and_7  g1363(.A(new_n1638), .B(new_n1629_1), .Y(new_n1639));
  or_2   g1364(.A(new_n1639), .B(new_n1627), .Y(new_n1640));
  nor_6  g1365(.A(new_n1638), .B(new_n1629_1), .Y(new_n1641));
  nor_6  g1366(.A(new_n1641), .B(new_n1639), .Y(new_n1642_1));
  and_7  g1367(.A(new_n277_1), .B(new_n862_1), .Y(new_n1643_1));
  not_13 g1368(.A(new_n1643_1), .Y(new_n1644));
  or_2   g1369(.A(new_n881), .B(new_n863), .Y(new_n1645));
  and_7  g1370(.A(new_n1645), .B(new_n1644), .Y(new_n1646));
  and_7  g1371(.A(new_n1646), .B(n49), .Y(new_n1647));
  and_7  g1372(.A(new_n1647), .B(n1622), .Y(new_n1648));
  and_7  g1373(.A(new_n1648), .B(n906), .Y(new_n1649));
  and_7  g1374(.A(new_n1649), .B(n277), .Y(new_n1650));
  nor_6  g1375(.A(new_n1637), .B(new_n1635_1), .Y(new_n1651));
  nor_6  g1376(.A(new_n1651), .B(new_n1638), .Y(new_n1652));
  nor_6  g1377(.A(new_n1652), .B(new_n1650), .Y(new_n1653));
  and_7  g1378(.A(new_n1652), .B(new_n1650), .Y(new_n1654_1));
  or_2   g1379(.A(new_n1654_1), .B(new_n1653), .Y(new_n1655));
  not_13 g1380(.A(n277), .Y(new_n1656));
  not_13 g1381(.A(n906), .Y(new_n1657_1));
  not_13 g1382(.A(n1622), .Y(new_n1658));
  not_13 g1383(.A(n49), .Y(new_n1659));
  or_2   g1384(.A(new_n891_1), .B(new_n1643_1), .Y(new_n1660_1));
  or_2   g1385(.A(new_n1660_1), .B(new_n1659), .Y(new_n1661));
  or_2   g1386(.A(new_n1661), .B(new_n1658), .Y(new_n1662));
  or_2   g1387(.A(new_n1662), .B(new_n1657_1), .Y(new_n1663));
  and_7  g1388(.A(new_n1663), .B(new_n1656), .Y(new_n1664));
  nor_6  g1389(.A(new_n1664), .B(new_n1650), .Y(new_n1665));
  nor_6  g1390(.A(new_n1634), .B(new_n1631), .Y(new_n1666));
  nor_6  g1391(.A(new_n1666), .B(new_n1635_1), .Y(new_n1667));
  or_2   g1392(.A(new_n1667), .B(new_n1665), .Y(new_n1668));
  nor_6  g1393(.A(new_n1667), .B(new_n1665), .Y(new_n1669));
  and_7  g1394(.A(new_n1667), .B(new_n1665), .Y(new_n1670));
  or_2   g1395(.A(new_n1670), .B(new_n1669), .Y(new_n1671));
  and_7  g1396(.A(new_n1662), .B(new_n1657_1), .Y(new_n1672));
  nor_6  g1397(.A(new_n1672), .B(new_n1649), .Y(new_n1673));
  nor_6  g1398(.A(new_n1633_1), .B(new_n383), .Y(new_n1674));
  nor_6  g1399(.A(new_n1674), .B(new_n1634), .Y(new_n1675_1));
  nor_6  g1400(.A(new_n1675_1), .B(new_n1673), .Y(new_n1676));
  and_7  g1401(.A(new_n1675_1), .B(new_n1673), .Y(new_n1677_1));
  or_2   g1402(.A(new_n1677_1), .B(new_n1676), .Y(new_n1678_1));
  or_2   g1403(.A(new_n1647), .B(n1622), .Y(new_n1679));
  and_7  g1404(.A(new_n1679), .B(new_n1662), .Y(new_n1680));
  nor_6  g1405(.A(new_n1680), .B(new_n385), .Y(new_n1681));
  and_7  g1406(.A(new_n1680), .B(new_n385), .Y(new_n1682));
  nor_6  g1407(.A(new_n1682), .B(new_n1681), .Y(new_n1683_1));
  and_7  g1408(.A(new_n1660_1), .B(new_n1659), .Y(new_n1684));
  nor_6  g1409(.A(new_n1684), .B(new_n1647), .Y(new_n1685));
  and_7  g1410(.A(new_n1685), .B(new_n390), .Y(new_n1686_1));
  nor_6  g1411(.A(new_n1685), .B(new_n390), .Y(new_n1687));
  or_2   g1412(.A(new_n1687), .B(new_n1686_1), .Y(new_n1688_1));
  and_7  g1413(.A(new_n924), .B(new_n895), .Y(new_n1689));
  nor_6  g1414(.A(new_n1689), .B(new_n893), .Y(new_n1690_1));
  nor_6  g1415(.A(new_n1690_1), .B(new_n1688_1), .Y(new_n1691));
  nor_6  g1416(.A(new_n1691), .B(new_n1686_1), .Y(new_n1692));
  and_7  g1417(.A(new_n1692), .B(new_n1683_1), .Y(new_n1693));
  nor_6  g1418(.A(new_n1693), .B(new_n1681), .Y(new_n1694));
  nor_6  g1419(.A(new_n1694), .B(new_n1678_1), .Y(new_n1695));
  nor_6  g1420(.A(new_n1695), .B(new_n1676), .Y(new_n1696));
  or_2   g1421(.A(new_n1696), .B(new_n1671), .Y(new_n1697));
  and_7  g1422(.A(new_n1697), .B(new_n1668), .Y(new_n1698));
  nor_6  g1423(.A(new_n1698), .B(new_n1655), .Y(new_n1699));
  nor_6  g1424(.A(new_n1699), .B(new_n1653), .Y(new_n1700));
  and_7  g1425(.A(new_n1700), .B(new_n1642_1), .Y(new_n1701));
  nor_6  g1426(.A(new_n1701), .B(new_n1640), .Y(n534));
  and_7  g1427(.A(n1721), .B(new_n589), .Y(new_n1703));
  or_2   g1428(.A(new_n1703), .B(new_n592), .Y(n541));
  or_2   g1429(.A(new_n1026), .B(new_n1015_1), .Y(n547));
  nor_6  g1430(.A(new_n1265), .B(new_n1190), .Y(new_n1706));
  and_7  g1431(.A(new_n1265), .B(new_n1190), .Y(new_n1707_1));
  or_2   g1432(.A(new_n1707_1), .B(new_n1706), .Y(new_n1708));
  nor_6  g1433(.A(new_n1552), .B(new_n1512), .Y(new_n1709));
  nor_6  g1434(.A(new_n1709), .B(new_n1708), .Y(new_n1710));
  or_2   g1435(.A(new_n1710), .B(new_n1706), .Y(new_n1711));
  and_7  g1436(.A(new_n1711), .B(new_n1272), .Y(n549));
  and_7  g1437(.A(new_n1572), .B(new_n1570), .Y(new_n1713));
  or_2   g1438(.A(new_n1713), .B(new_n1573), .Y(n559));
  not_13 g1439(.A(new_n1419), .Y(n569));
  xor_5  g1440(.A(new_n1543), .B(new_n1541), .Y(n573));
  and_7  g1441(.A(new_n1709), .B(new_n1708), .Y(new_n1717));
  or_2   g1442(.A(new_n1717), .B(new_n1710), .Y(n588));
  not_13 g1443(.A(new_n585_1), .Y(new_n1719));
  xor_5  g1444(.A(n416), .B(new_n1719), .Y(n599));
  nor_6  g1445(.A(new_n1427), .B(new_n1398), .Y(n627));
  and_7  g1446(.A(new_n1263_1), .B(new_n811), .Y(new_n1722));
  xor_5  g1447(.A(new_n1722), .B(new_n1382), .Y(new_n1723));
  or_2   g1448(.A(new_n1723), .B(new_n1271), .Y(new_n1724));
  nor_6  g1449(.A(new_n1270), .B(new_n1266), .Y(new_n1725));
  xor_5  g1450(.A(new_n1722), .B(new_n826), .Y(new_n1726));
  or_2   g1451(.A(new_n1726), .B(new_n1725), .Y(new_n1727_1));
  and_7  g1452(.A(new_n1727_1), .B(new_n1724), .Y(n638));
  and_7  g1453(.A(new_n930), .B(new_n821), .Y(new_n1729_1));
  and_7  g1454(.A(new_n1729_1), .B(new_n457_1), .Y(new_n1730));
  and_7  g1455(.A(new_n944_1), .B(n1381), .Y(new_n1731_1));
  or_2   g1456(.A(new_n1731_1), .B(new_n1730), .Y(new_n1732));
  not_13 g1457(.A(new_n1732), .Y(new_n1733));
  nor_6  g1458(.A(new_n1733), .B(new_n954), .Y(n643));
  xor_5  g1459(.A(new_n1690_1), .B(new_n1688_1), .Y(n648));
  or_2   g1460(.A(new_n779), .B(new_n739), .Y(new_n1736));
  xor_5  g1461(.A(new_n1736), .B(new_n734), .Y(n665));
  or_2   g1462(.A(new_n1182), .B(new_n1178), .Y(new_n1738));
  xor_5  g1463(.A(new_n1738), .B(new_n1173), .Y(n683));
  or_2   g1464(.A(new_n1642_1), .B(new_n1190), .Y(new_n1740));
  nor_6  g1465(.A(new_n1642_1), .B(new_n1190), .Y(new_n1741));
  and_7  g1466(.A(new_n1642_1), .B(new_n1190), .Y(new_n1742));
  or_2   g1467(.A(new_n1742), .B(new_n1741), .Y(new_n1743_1));
  or_2   g1468(.A(new_n1652), .B(new_n1190), .Y(new_n1744));
  nor_6  g1469(.A(new_n1652), .B(new_n1190), .Y(new_n1745));
  and_7  g1470(.A(new_n1652), .B(new_n1190), .Y(new_n1746_1));
  or_2   g1471(.A(new_n1746_1), .B(new_n1745), .Y(new_n1747_1));
  nor_6  g1472(.A(new_n1667), .B(new_n1199_1), .Y(new_n1748));
  and_7  g1473(.A(new_n1667), .B(new_n1199_1), .Y(new_n1749));
  nor_6  g1474(.A(new_n1749), .B(new_n1748), .Y(new_n1750));
  nor_6  g1475(.A(new_n1675_1), .B(new_n1204), .Y(new_n1751));
  and_7  g1476(.A(new_n1675_1), .B(new_n1204), .Y(new_n1752));
  or_2   g1477(.A(new_n1752), .B(new_n1751), .Y(new_n1753));
  nor_6  g1478(.A(new_n452_1), .B(new_n387_1), .Y(new_n1754));
  nor_6  g1479(.A(new_n1754), .B(new_n1753), .Y(new_n1755));
  or_2   g1480(.A(new_n1755), .B(new_n1751), .Y(new_n1756));
  and_7  g1481(.A(new_n1756), .B(new_n1750), .Y(new_n1757_1));
  nor_6  g1482(.A(new_n1757_1), .B(new_n1748), .Y(new_n1758));
  or_2   g1483(.A(new_n1758), .B(new_n1747_1), .Y(new_n1759));
  and_7  g1484(.A(new_n1759), .B(new_n1744), .Y(new_n1760));
  or_2   g1485(.A(new_n1760), .B(new_n1743_1), .Y(new_n1761));
  and_7  g1486(.A(new_n1761), .B(new_n1740), .Y(new_n1762));
  or_2   g1487(.A(new_n1617), .B(new_n1591), .Y(new_n1763_1));
  and_7  g1488(.A(new_n1763_1), .B(new_n1627), .Y(new_n1764_1));
  nor_6  g1489(.A(new_n1764_1), .B(new_n1639), .Y(new_n1765));
  and_7  g1490(.A(new_n1764_1), .B(new_n1639), .Y(new_n1766));
  nor_6  g1491(.A(new_n1766), .B(new_n1765), .Y(new_n1767));
  nor_6  g1492(.A(new_n1767), .B(new_n1762), .Y(new_n1768));
  and_7  g1493(.A(new_n1767), .B(new_n1197), .Y(new_n1769));
  and_7  g1494(.A(new_n1761), .B(new_n1190), .Y(new_n1770));
  or_2   g1495(.A(new_n1770), .B(new_n1769), .Y(new_n1771));
  nor_6  g1496(.A(new_n1771), .B(new_n1768), .Y(new_n1772));
  nor_6  g1497(.A(new_n1772), .B(new_n1640), .Y(new_n1773));
  and_7  g1498(.A(new_n1772), .B(new_n1640), .Y(new_n1774));
  or_2   g1499(.A(new_n1774), .B(new_n1773), .Y(n699));
  not_13 g1500(.A(new_n431), .Y(new_n1776));
  xor_5  g1501(.A(new_n913), .B(new_n1776), .Y(n712));
  not_13 g1502(.A(new_n594), .Y(n715));
  nor_6  g1503(.A(new_n1423), .B(n145), .Y(new_n1779));
  nor_6  g1504(.A(new_n1779), .B(new_n1424), .Y(n724));
  not_13 g1505(.A(n647), .Y(n1255));
  xor_5  g1506(.A(new_n978), .B(new_n977), .Y(new_n1782));
  and_7  g1507(.A(new_n1782), .B(n1255), .Y(new_n1783));
  xor_5  g1508(.A(n1016), .B(new_n1783), .Y(n725));
  and_7  g1509(.A(new_n1574), .B(new_n1560), .Y(new_n1785));
  or_2   g1510(.A(new_n1785), .B(new_n1575), .Y(n731));
  and_7  g1511(.A(new_n1754), .B(new_n1753), .Y(new_n1787));
  or_2   g1512(.A(new_n1787), .B(new_n1755), .Y(n748));
  or_2   g1513(.A(new_n1502_1), .B(new_n1492), .Y(new_n1789));
  xor_5  g1514(.A(new_n1789), .B(new_n1491), .Y(n759));
  and_7  g1515(.A(new_n1582), .B(new_n1238), .Y(new_n1791));
  and_7  g1516(.A(new_n1197), .B(new_n805), .Y(new_n1792));
  nor_6  g1517(.A(new_n1220), .B(new_n1792), .Y(new_n1793));
  nor_6  g1518(.A(new_n1793), .B(n1422), .Y(new_n1794));
  and_7  g1519(.A(new_n1794), .B(new_n1791), .Y(n770));
  or_2   g1520(.A(new_n1544_1), .B(new_n1524), .Y(new_n1796));
  xor_5  g1521(.A(new_n1796), .B(new_n1523), .Y(n790));
  and_7  g1522(.A(new_n1190), .B(new_n833), .Y(new_n1798));
  nor_6  g1523(.A(new_n1190), .B(new_n833), .Y(new_n1799));
  or_2   g1524(.A(new_n1799), .B(new_n1798), .Y(new_n1800));
  nor_6  g1525(.A(new_n1556_1), .B(new_n1555), .Y(new_n1801));
  and_7  g1526(.A(new_n1576), .B(new_n1801), .Y(new_n1802));
  nor_6  g1527(.A(new_n1802), .B(new_n1556_1), .Y(new_n1803));
  nor_6  g1528(.A(new_n1803), .B(new_n1800), .Y(new_n1804));
  and_7  g1529(.A(new_n1803), .B(new_n1800), .Y(new_n1805));
  or_2   g1530(.A(new_n1805), .B(new_n1804), .Y(n792));
  not_13 g1531(.A(new_n1131), .Y(new_n1807));
  xor_5  g1532(.A(new_n1134), .B(new_n1807), .Y(n813));
  and_7  g1533(.A(new_n1367), .B(new_n1358), .Y(new_n1809));
  or_2   g1534(.A(new_n1809), .B(new_n1368), .Y(n823));
  and_7  g1535(.A(new_n1386), .B(new_n823_1), .Y(n824));
  not_13 g1536(.A(new_n486), .Y(new_n1812));
  xor_5  g1537(.A(new_n488_1), .B(new_n1812), .Y(n836));
  or_2   g1538(.A(new_n1749), .B(new_n1748), .Y(new_n1814));
  xor_5  g1539(.A(new_n1756), .B(new_n1814), .Y(n846));
  not_13 g1540(.A(new_n1342), .Y(new_n1816));
  or_2   g1541(.A(new_n1371), .B(new_n1344), .Y(new_n1817));
  and_7  g1542(.A(new_n1817), .B(new_n1816), .Y(new_n1818));
  xor_5  g1543(.A(new_n1818), .B(new_n1337), .Y(n858));
  or_2   g1544(.A(new_n1395), .B(new_n794), .Y(new_n1820));
  and_7  g1545(.A(new_n1820), .B(new_n1385_1), .Y(n865));
  and_7  g1546(.A(new_n1549), .B(new_n1516), .Y(new_n1822));
  or_2   g1547(.A(new_n1822), .B(new_n1550), .Y(n867));
  or_2   g1548(.A(new_n952_1), .B(new_n947), .Y(new_n1824));
  xor_5  g1549(.A(new_n1478), .B(new_n1824), .Y(new_n1825));
  or_2   g1550(.A(new_n1508), .B(new_n1482), .Y(new_n1826));
  and_7  g1551(.A(new_n1826), .B(new_n1825), .Y(new_n1827));
  nor_6  g1552(.A(new_n1826), .B(new_n1825), .Y(new_n1828));
  nor_6  g1553(.A(new_n1828), .B(new_n1827), .Y(n883));
  and_7  g1554(.A(new_n784), .B(new_n782), .Y(new_n1830));
  or_2   g1555(.A(new_n1830), .B(new_n785), .Y(n888));
  xor_5  g1556(.A(new_n1478), .B(new_n953_1), .Y(new_n1832));
  and_7  g1557(.A(new_n1312), .B(n1757), .Y(new_n1833));
  and_7  g1558(.A(new_n1833), .B(n839), .Y(new_n1834));
  or_2   g1559(.A(new_n1834), .B(new_n1480), .Y(new_n1835));
  nor_6  g1560(.A(new_n1834), .B(new_n1480), .Y(new_n1836));
  and_7  g1561(.A(new_n1834), .B(new_n1480), .Y(new_n1837));
  or_2   g1562(.A(new_n1837), .B(new_n1836), .Y(new_n1838));
  not_13 g1563(.A(n839), .Y(new_n1839));
  and_7  g1564(.A(new_n1438), .B(new_n1839), .Y(new_n1840));
  nor_6  g1565(.A(new_n1840), .B(new_n1834), .Y(new_n1841));
  or_2   g1566(.A(new_n1841), .B(new_n1485), .Y(new_n1842));
  nor_6  g1567(.A(new_n1841), .B(new_n1485), .Y(new_n1843));
  and_7  g1568(.A(new_n1841), .B(new_n1485), .Y(new_n1844));
  or_2   g1569(.A(new_n1844), .B(new_n1843), .Y(new_n1845));
  or_2   g1570(.A(new_n1377), .B(new_n1325), .Y(new_n1846));
  and_7  g1571(.A(new_n1846), .B(new_n1443), .Y(new_n1847));
  nor_6  g1572(.A(new_n1847), .B(new_n1442), .Y(new_n1848));
  or_2   g1573(.A(new_n1848), .B(new_n1845), .Y(new_n1849));
  and_7  g1574(.A(new_n1849), .B(new_n1842), .Y(new_n1850));
  or_2   g1575(.A(new_n1850), .B(new_n1838), .Y(new_n1851));
  and_7  g1576(.A(new_n1851), .B(new_n1835), .Y(new_n1852));
  or_2   g1577(.A(new_n1852), .B(new_n1832), .Y(new_n1853));
  nor_6  g1578(.A(new_n1850), .B(new_n1838), .Y(new_n1854));
  or_2   g1579(.A(new_n1854), .B(new_n1836), .Y(new_n1855));
  or_2   g1580(.A(new_n1855), .B(new_n1825), .Y(new_n1856));
  and_7  g1581(.A(new_n1856), .B(new_n1853), .Y(n891));
  and_7  g1582(.A(new_n1478), .B(new_n953_1), .Y(new_n1858));
  and_7  g1583(.A(new_n1852), .B(new_n1832), .Y(new_n1859));
  nor_6  g1584(.A(new_n1859), .B(new_n1858), .Y(new_n1860));
  and_7  g1585(.A(new_n1860), .B(new_n1732), .Y(n892));
  xor_5  g1586(.A(new_n1113_1), .B(new_n1112), .Y(n902));
  not_13 g1587(.A(new_n1254), .Y(new_n1863));
  xor_5  g1588(.A(new_n743), .B(new_n407), .Y(new_n1864));
  xor_5  g1589(.A(new_n1864), .B(new_n1863), .Y(n905));
  xor_5  g1590(.A(new_n1468), .B(new_n1226), .Y(n912));
  nor_6  g1591(.A(n1149), .B(new_n600_1), .Y(new_n1867));
  nor_6  g1592(.A(new_n1867), .B(new_n959), .Y(n935));
  xor_5  g1593(.A(new_n1424), .B(n1119), .Y(n942));
  or_2   g1594(.A(new_n1179), .B(new_n1178), .Y(new_n1870));
  xor_5  g1595(.A(new_n1181), .B(new_n1870), .Y(n944));
  and_7  g1596(.A(n770), .B(n547), .Y(n974));
  or_2   g1597(.A(new_n448), .B(new_n403), .Y(new_n1873));
  xor_5  g1598(.A(new_n1873), .B(new_n398), .Y(n979));
  and_7  g1599(.A(new_n1382), .B(new_n819), .Y(new_n1875));
  not_13 g1600(.A(new_n1875), .Y(new_n1876));
  and_7  g1601(.A(new_n1876), .B(new_n1389), .Y(new_n1877));
  nor_6  g1602(.A(new_n1877), .B(new_n828), .Y(new_n1878));
  and_7  g1603(.A(new_n1878), .B(new_n855), .Y(n980));
  or_2   g1604(.A(new_n1546), .B(new_n1521), .Y(new_n1880));
  xor_5  g1605(.A(new_n1880), .B(new_n1520), .Y(n989));
  nor_6  g1606(.A(new_n1758), .B(new_n1747_1), .Y(new_n1882));
  or_2   g1607(.A(new_n1882), .B(new_n1745), .Y(new_n1883));
  xor_5  g1608(.A(new_n1883), .B(new_n1743_1), .Y(n991));
  or_2   g1609(.A(new_n1847), .B(new_n1442), .Y(new_n1885));
  xor_5  g1610(.A(new_n1885), .B(new_n1845), .Y(n1005));
  and_7  g1611(.A(new_n1505), .B(new_n1488), .Y(new_n1887));
  or_2   g1612(.A(new_n1887), .B(new_n1506), .Y(n1012));
  nor_6  g1613(.A(new_n1029), .B(new_n1025_1), .Y(new_n1889));
  xor_5  g1614(.A(new_n1889), .B(new_n1023), .Y(n1015));
  and_7  g1615(.A(new_n859), .B(new_n856), .Y(new_n1891));
  and_7  g1616(.A(new_n1877), .B(new_n1891), .Y(new_n1892));
  and_7  g1617(.A(new_n1877), .B(new_n828), .Y(new_n1893));
  or_2   g1618(.A(new_n1893), .B(new_n1878), .Y(new_n1894));
  and_7  g1619(.A(new_n1894), .B(new_n855), .Y(new_n1895));
  or_2   g1620(.A(new_n1895), .B(new_n1892), .Y(n1025));
  and_7  g1621(.A(new_n1850), .B(new_n1838), .Y(new_n1897));
  or_2   g1622(.A(new_n1897), .B(new_n1854), .Y(n1030));
  and_7  g1623(.A(new_n850), .B(new_n846_1), .Y(new_n1899));
  or_2   g1624(.A(new_n1899), .B(new_n851), .Y(n1067));
  nor_6  g1625(.A(new_n1860), .B(new_n1732), .Y(new_n1901));
  or_2   g1626(.A(new_n1901), .B(n892), .Y(n1068));
  xor_5  g1627(.A(new_n594), .B(new_n592), .Y(n1103));
  xor_5  g1628(.A(new_n482_1), .B(new_n413), .Y(n1113));
  or_2   g1629(.A(new_n1581), .B(new_n1224), .Y(new_n1905));
  or_2   g1630(.A(new_n1905), .B(new_n1222_1), .Y(new_n1906));
  and_7  g1631(.A(new_n1793), .B(n1422), .Y(new_n1907));
  and_7  g1632(.A(new_n1907), .B(new_n1906), .Y(new_n1908));
  or_2   g1633(.A(new_n1908), .B(n770), .Y(n1135));
  and_7  g1634(.A(new_n1764_1), .B(new_n1701), .Y(new_n1910));
  nor_6  g1635(.A(new_n1767), .B(new_n1701), .Y(new_n1911));
  or_2   g1636(.A(new_n1911), .B(new_n1910), .Y(n1142));
  nor_6  g1637(.A(new_n1767), .B(new_n1197), .Y(new_n1913));
  nor_6  g1638(.A(new_n1913), .B(new_n1769), .Y(new_n1914));
  nor_6  g1639(.A(new_n1914), .B(new_n1762), .Y(new_n1915));
  and_7  g1640(.A(new_n1914), .B(new_n1762), .Y(new_n1916));
  nor_6  g1641(.A(new_n1916), .B(new_n1915), .Y(n1161));
  nor_6  g1642(.A(new_n1579), .B(new_n1233), .Y(new_n1918));
  and_7  g1643(.A(new_n1579), .B(new_n1233), .Y(new_n1919));
  or_2   g1644(.A(new_n1919), .B(new_n1918), .Y(n1162));
  nor_6  g1645(.A(n865), .B(new_n1425_1), .Y(new_n1921));
  nor_6  g1646(.A(new_n1921), .B(new_n1426_1), .Y(n1175));
  or_2   g1647(.A(new_n1190), .B(new_n833), .Y(new_n1923));
  or_2   g1648(.A(new_n1803), .B(new_n1800), .Y(new_n1924));
  and_7  g1649(.A(new_n1924), .B(new_n1923), .Y(new_n1925));
  and_7  g1650(.A(new_n1190), .B(new_n830), .Y(new_n1926));
  or_2   g1651(.A(new_n1926), .B(new_n1925), .Y(new_n1927));
  and_7  g1652(.A(new_n1197), .B(new_n856), .Y(new_n1928));
  or_2   g1653(.A(new_n1928), .B(new_n1804), .Y(new_n1929));
  and_7  g1654(.A(new_n1929), .B(new_n1927), .Y(new_n1930));
  and_7  g1655(.A(new_n1930), .B(new_n1894), .Y(new_n1931));
  nor_6  g1656(.A(new_n1893), .B(new_n1878), .Y(new_n1932));
  or_2   g1657(.A(new_n1804), .B(new_n1799), .Y(new_n1933));
  or_2   g1658(.A(new_n1197), .B(new_n856), .Y(new_n1934));
  and_7  g1659(.A(new_n1934), .B(new_n1933), .Y(new_n1935));
  or_2   g1660(.A(new_n1190), .B(new_n830), .Y(new_n1936));
  and_7  g1661(.A(new_n1936), .B(new_n1924), .Y(new_n1937));
  or_2   g1662(.A(new_n1937), .B(new_n1935), .Y(new_n1938));
  and_7  g1663(.A(new_n1938), .B(new_n1932), .Y(new_n1939));
  nor_6  g1664(.A(new_n1939), .B(new_n1931), .Y(n1191));
  xor_5  g1665(.A(new_n1918), .B(new_n1226), .Y(n1194));
  xor_5  g1666(.A(new_n447), .B(new_n445), .Y(n1199));
  nor_6  g1667(.A(new_n1537_1), .B(new_n1531), .Y(new_n1943));
  or_2   g1668(.A(new_n1943), .B(new_n1538), .Y(n1201));
  not_13 g1669(.A(new_n979_1), .Y(new_n1945));
  and_7  g1670(.A(new_n1405), .B(new_n1945), .Y(new_n1946));
  or_2   g1671(.A(new_n1946), .B(new_n1783), .Y(n1202));
  xor_5  g1672(.A(new_n1419), .B(new_n1417), .Y(n1234));
  and_7  g1673(.A(new_n1905), .B(new_n1222_1), .Y(new_n1949));
  or_2   g1674(.A(new_n1949), .B(new_n1791), .Y(n1235));
  not_13 g1675(.A(n1183), .Y(n1237));
  and_7  g1676(.A(new_n1722), .B(new_n826), .Y(new_n1952));
  and_7  g1677(.A(new_n1726), .B(new_n1725), .Y(new_n1953));
  nor_6  g1678(.A(new_n1953), .B(new_n1952), .Y(new_n1954));
  nor_6  g1679(.A(new_n1954), .B(new_n823_1), .Y(new_n1955));
  or_2   g1680(.A(new_n1955), .B(n299), .Y(n1260));
  nor_6  g1681(.A(new_n1426_1), .B(n1249), .Y(new_n1957));
  nor_6  g1682(.A(new_n1957), .B(new_n1427), .Y(n1277));
  nor_6  g1683(.A(new_n1828), .B(new_n1858), .Y(new_n1959));
  and_7  g1684(.A(new_n1959), .B(new_n1732), .Y(n1278));
  and_7  g1685(.A(new_n431), .B(new_n419), .Y(new_n1961));
  or_2   g1686(.A(new_n431), .B(new_n424_1), .Y(new_n1962));
  and_7  g1687(.A(new_n1962), .B(new_n433_1), .Y(new_n1963));
  nor_6  g1688(.A(new_n1963), .B(new_n1961), .Y(n1283));
  or_2   g1689(.A(new_n1236), .B(new_n1222_1), .Y(new_n1965));
  and_7  g1690(.A(new_n1907), .B(new_n1965), .Y(new_n1966));
  or_2   g1691(.A(new_n1966), .B(n974), .Y(n1305));
  xor_5  g1692(.A(new_n595), .B(n1727), .Y(n1315));
  nor_6  g1693(.A(new_n1696), .B(new_n1671), .Y(new_n1969));
  and_7  g1694(.A(new_n1696), .B(new_n1671), .Y(new_n1970));
  or_2   g1695(.A(new_n1970), .B(new_n1969), .Y(n1330));
  nor_6  g1696(.A(new_n1568), .B(new_n1564), .Y(new_n1972));
  or_2   g1697(.A(new_n1972), .B(new_n1569), .Y(n1338));
  not_13 g1698(.A(new_n770_1), .Y(new_n1974));
  xor_5  g1699(.A(new_n1974), .B(new_n768), .Y(n1340));
  nor_6  g1700(.A(new_n1700), .B(new_n1642_1), .Y(new_n1976));
  nor_6  g1701(.A(new_n1976), .B(new_n1701), .Y(n1347));
  and_7  g1702(.A(new_n1733), .B(new_n954), .Y(new_n1978));
  or_2   g1703(.A(new_n1978), .B(n643), .Y(n1348));
  and_7  g1704(.A(new_n1371), .B(new_n1344), .Y(new_n1980));
  or_2   g1705(.A(new_n1980), .B(new_n1372), .Y(n1349));
  nor_6  g1706(.A(new_n1907), .B(new_n1794), .Y(new_n1982));
  nor_6  g1707(.A(new_n1982), .B(new_n1791), .Y(new_n1983));
  and_7  g1708(.A(new_n1982), .B(new_n1791), .Y(new_n1984));
  nor_6  g1709(.A(new_n1984), .B(new_n1983), .Y(n1369));
  nor_6  g1710(.A(new_n1982), .B(new_n1240), .Y(new_n1986));
  and_7  g1711(.A(new_n1982), .B(new_n1240), .Y(new_n1987));
  nor_6  g1712(.A(new_n1987), .B(new_n1986), .Y(n1383));
  or_2   g1713(.A(new_n1691), .B(new_n1686_1), .Y(new_n1989));
  xor_5  g1714(.A(new_n1989), .B(new_n1683_1), .Y(n1393));
  not_13 g1715(.A(new_n1535_1), .Y(new_n1991));
  xor_5  g1716(.A(new_n1991), .B(new_n1121), .Y(n1399));
  xor_5  g1717(.A(new_n750), .B(new_n412), .Y(new_n1993));
  xor_5  g1718(.A(new_n1993), .B(new_n1252), .Y(n1407));
  and_7  g1719(.A(new_n1397), .B(new_n826), .Y(new_n1995));
  and_7  g1720(.A(new_n1995), .B(new_n1389), .Y(new_n1996));
  or_2   g1721(.A(n824), .B(new_n1996), .Y(n1425));
  or_2   g1722(.A(new_n1733), .B(new_n954), .Y(new_n1998));
  nor_6  g1723(.A(new_n1998), .B(new_n961_1), .Y(n1440));
  or_2   g1724(.A(new_n1028), .B(new_n1017), .Y(n1601));
  xor_5  g1725(.A(n1601), .B(new_n1025_1), .Y(n1453));
  not_13 g1726(.A(new_n1250), .Y(new_n2002));
  xor_5  g1727(.A(new_n2002), .B(new_n768), .Y(n1460));
  and_7  g1728(.A(new_n1936), .B(new_n1934), .Y(new_n2004));
  or_2   g1729(.A(new_n2004), .B(new_n1933), .Y(new_n2005));
  or_2   g1730(.A(new_n1928), .B(new_n1926), .Y(new_n2006));
  or_2   g1731(.A(new_n2006), .B(new_n1925), .Y(new_n2007));
  and_7  g1732(.A(new_n2007), .B(new_n2005), .Y(n1463));
  and_7  g1733(.A(new_n1235_1), .B(new_n1224), .Y(new_n2009));
  or_2   g1734(.A(new_n2009), .B(new_n1239), .Y(n1470));
  xor_5  g1735(.A(new_n1113_1), .B(new_n413), .Y(n1481));
  not_13 g1736(.A(new_n772), .Y(new_n2012));
  xor_5  g1737(.A(new_n774), .B(new_n2012), .Y(n1495));
  and_7  g1738(.A(new_n1129), .B(new_n1105), .Y(new_n2014));
  or_2   g1739(.A(new_n2014), .B(new_n1130), .Y(n1498));
  and_7  g1740(.A(new_n1694), .B(new_n1678_1), .Y(new_n2016));
  or_2   g1741(.A(new_n2016), .B(new_n1695), .Y(n1502));
  not_13 g1742(.A(new_n1353), .Y(new_n2018));
  xor_5  g1743(.A(new_n1369_1), .B(new_n2018), .Y(n1507));
  xor_5  g1744(.A(new_n1416), .B(new_n1412), .Y(n1525));
  and_7  g1745(.A(new_n776), .B(new_n748_1), .Y(new_n2021));
  or_2   g1746(.A(new_n2021), .B(new_n777), .Y(n1535));
  xor_5  g1747(.A(new_n1029), .B(n547), .Y(n1556));
  and_7  g1748(.A(n1348), .B(new_n961_1), .Y(new_n2024));
  nor_6  g1749(.A(n1348), .B(new_n961_1), .Y(new_n2025));
  nor_6  g1750(.A(new_n2025), .B(new_n2024), .Y(n1595));
  and_7  g1751(.A(new_n1539), .B(new_n1527_1), .Y(new_n2027));
  or_2   g1752(.A(new_n2027), .B(new_n1540), .Y(n1600));
  or_2   g1753(.A(new_n471), .B(n1145), .Y(new_n2029));
  and_7  g1754(.A(new_n2029), .B(new_n581), .Y(new_n2030));
  or_2   g1755(.A(new_n2030), .B(new_n1719), .Y(n1613));
  xor_5  g1756(.A(new_n1365), .B(new_n1812), .Y(n1629));
  or_2   g1757(.A(new_n1877), .B(new_n828), .Y(new_n2033));
  and_7  g1758(.A(new_n1938), .B(new_n2033), .Y(new_n2034));
  and_7  g1759(.A(new_n1928), .B(new_n1925), .Y(new_n2035));
  or_2   g1760(.A(new_n2035), .B(new_n1893), .Y(new_n2036));
  nor_6  g1761(.A(new_n2036), .B(new_n2034), .Y(n1633));
  and_7  g1762(.A(n1601), .B(n547), .Y(new_n2038));
  xor_5  g1763(.A(new_n2038), .B(new_n1025_1), .Y(n1635));
  xor_5  g1764(.A(new_n1501_1), .B(new_n1499), .Y(n1654));
  xor_5  g1765(.A(new_n597), .B(n1138), .Y(n1657));
  or_2   g1766(.A(new_n1828), .B(new_n1858), .Y(new_n2042));
  and_7  g1767(.A(new_n2042), .B(new_n1733), .Y(new_n2043));
  or_2   g1768(.A(new_n2043), .B(n1278), .Y(n1660));
  not_13 g1769(.A(new_n1123), .Y(new_n2045));
  xor_5  g1770(.A(new_n2045), .B(new_n1121), .Y(n1675));
  not_13 g1771(.A(new_n1416), .Y(n1683));
  or_2   g1772(.A(new_n1723), .B(new_n1711), .Y(new_n2048));
  or_2   g1773(.A(new_n1265), .B(new_n1190), .Y(new_n2049));
  or_2   g1774(.A(new_n1709), .B(new_n1708), .Y(new_n2050));
  and_7  g1775(.A(new_n2050), .B(new_n2049), .Y(new_n2051));
  or_2   g1776(.A(new_n1726), .B(new_n2051), .Y(new_n2052));
  and_7  g1777(.A(new_n2052), .B(new_n2048), .Y(n1686));
  xor_5  g1778(.A(new_n761_1), .B(new_n413), .Y(n1688));
  and_7  g1779(.A(new_n1698), .B(new_n1655), .Y(new_n2055));
  or_2   g1780(.A(new_n2055), .B(new_n1699), .Y(n1690));
  and_7  g1781(.A(new_n1758), .B(new_n1747_1), .Y(new_n2057));
  or_2   g1782(.A(new_n2057), .B(new_n1882), .Y(n1729));
  and_7  g1783(.A(new_n1726), .B(new_n2051), .Y(new_n2059));
  nor_6  g1784(.A(new_n2059), .B(new_n1952), .Y(new_n2060));
  nor_6  g1785(.A(new_n2060), .B(new_n823_1), .Y(new_n2061));
  or_2   g1786(.A(new_n2061), .B(n549), .Y(n1737));
  not_13 g1787(.A(new_n1461_1), .Y(new_n2063));
  or_2   g1788(.A(new_n1464), .B(new_n1462), .Y(new_n2064));
  and_7  g1789(.A(new_n2064), .B(new_n2063), .Y(new_n2065));
  xor_5  g1790(.A(new_n2065), .B(new_n1496), .Y(n1746));
  xor_5  g1791(.A(new_n413), .B(n347), .Y(n488));
  xor_5  g1792(.A(new_n1012_1), .B(new_n1259), .Y(n1677));
endmodule


